//
// Conformal-LEC Version 15.10-d154 ( 22-Jul-2015) ( 64 bit executable)
//
module test ( 
    n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 , 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 );
input 
    n0 , 
    n1 , 
    n2 , 
    n3 , 
    n4 , 
    n5 , 
    n6 , 
    n7 , 
    n8 , 
    n9 , 
    n10 , 
    n11 , 
    n12 , 
    n13 , 
    n14 , 
    n15 , 
    n16 , 
    n17 , 
    n18 , 
    n19 , 
    n20 , 
    n21 , 
    n22 , 
    n23 , 
    n24 , 
    n25 , 
    n26 , 
    n27 , 
    n28 , 
    n29 , 
    n30 , 
    n31 , 
    n32 , 
    n33 , 
    n34 , 
    n35 , 
    n36 , 
    n37 , 
    n38 , 
    n39 , 
    n40 , 
    n41 , 
    n42 , 
    n43 , 
    n44 , 
    n45 , 
    n46 , 
    n47 , 
    n48 , 
    n49 , 
    n50 , 
    n51 , 
    n52 , 
    n53 , 
    n54 , 
    n55 , 
    n56 , 
    n57 , 
    n58 , 
    n59 , 
    n60 , 
    n61 , 
    n62 , 
    n63 , 
    n64 , 
    n65 , 
    n66 , 
    n67 , 
    n68 , 
    n69 , 
    n70 , 
    n71 , 
    n72 , 
    n73 , 
    n74 , 
    n75 , 
    n76 , 
    n77 , 
    n78 , 
    n79 , 
    n80 , 
    n81 , 
    n82 , 
    n83 , 
    n84 , 
    n85 , 
    n86 , 
    n87 , 
    n88 , 
    n89 , 
    n90 , 
    n91 , 
    n92 , 
    n93 , 
    n94 , 
    n95 , 
    n96 , 
    n97 , 
    n98 , 
    n99 , 
    n100 , 
    n101 , 
    n102 , 
    n103 , 
    n104 , 
    n105 , 
    n106 , 
    n107 , 
    n108 , 
    n109 , 
    n110 , 
    n111 , 
    n112 , 
    n113 , 
    n114 , 
    n115 , 
    n116 , 
    n117 , 
    n118 , 
    n119 , 
    n120 , 
    n121 , 
    n122 , 
    n123 , 
    n124 , 
    n125 , 
    n126 , 
    n127 , 
    n128 , 
    n129 , 
    n130 , 
    n131 , 
    n132 , 
    n133 , 
    n134 , 
    n135 , 
    n136 , 
    n137 , 
    n138 , 
    n139 , 
    n140 , 
    n141 , 
    n142 , 
    n143 , 
    n144 , 
    n145 , 
    n146 , 
    n147 , 
    n148 , 
    n149 , 
    n150 , 
    n151 , 
    n152 , 
    n153 , 
    n154 , 
    n155 , 
    n156 , 
    n157 , 
    n158 , 
    n159 ;
output 
    n160 , 
    n161 , 
    n162 , 
    n163 , 
    n164 , 
    n165 , 
    n166 , 
    n167 , 
    n168 , 
    n169 , 
    n170 , 
    n171 , 
    n172 , 
    n173 , 
    n174 , 
    n175 , 
    n176 , 
    n177 , 
    n178 , 
    n179 , 
    n180 , 
    n181 , 
    n182 , 
    n183 , 
    n184 , 
    n185 , 
    n186 , 
    n187 , 
    n188 , 
    n189 , 
    n190 , 
    n191 , 
    n192 , 
    n193 , 
    n194 , 
    n195 , 
    n196 , 
    n197 , 
    n198 , 
    n199 , 
    n200 , 
    n201 , 
    n202 , 
    n203 , 
    n204 , 
    n205 , 
    n206 , 
    n207 , 
    n208 , 
    n209 , 
    n210 , 
    n211 , 
    n212 , 
    n213 , 
    n214 , 
    n215 , 
    n216 , 
    n217 , 
    n218 , 
    n219 , 
    n220 , 
    n221 , 
    n222 , 
    n223 , 
    n224 , 
    n225 , 
    n226 , 
    n227 , 
    n228 , 
    n229 , 
    n230 , 
    n231 , 
    n232 , 
    n233 , 
    n234 , 
    n235 , 
    n236 , 
    n237 , 
    n238 , 
    n239 , 
    n240 , 
    n241 , 
    n242 , 
    n243 , 
    n244 , 
    n245 , 
    n246 , 
    n247 , 
    n248 , 
    n249 , 
    n250 , 
    n251 , 
    n252 , 
    n253 , 
    n254 , 
    n255 , 
    n256 , 
    n257 , 
    n258 , 
    n259 , 
    n260 , 
    n261 , 
    n262 , 
    n263 , 
    n264 , 
    n265 , 
    n266 , 
    n267 , 
    n268 , 
    n269 , 
    n270 , 
    n271 , 
    n272 , 
    n273 , 
    n274 , 
    n275 , 
    n276 , 
    n277 , 
    n278 , 
    n279 , 
    n280 , 
    n281 , 
    n282 , 
    n283 , 
    n284 , 
    n285 , 
    n286 , 
    n287 , 
    n288 , 
    n289 , 
    n290 , 
    n291 , 
    n292 , 
    n293 , 
    n294 , 
    n295 , 
    n296 , 
    n297 , 
    n298 , 
    n299 , 
    n300 , 
    n301 , 
    n302 , 
    n303 , 
    n304 , 
    n305 , 
    n306 , 
    n307 , 
    n308 , 
    n309 , 
    n310 , 
    n311 , 
    n312 , 
    n313 , 
    n314 , 
    n315 , 
    n316 , 
    n317 , 
    n318 , 
    n319 , 
    n320 , 
    n321 , 
    n322 , 
    n323 , 
    n324 , 
    n325 , 
    n326 , 
    n327 , 
    n328 , 
    n329 , 
    n330 , 
    n331 , 
    n332 , 
    n333 , 
    n334 , 
    n335 , 
    n336 , 
    n337 , 
    n338 , 
    n339 , 
    n340 , 
    n341 , 
    n342 , 
    n343 , 
    n344 , 
    n345 , 
    n346 , 
    n347 , 
    n348 , 
    n349 , 
    n350 , 
    n351 , 
    n352 , 
    n353 , 
    n354 , 
    n355 , 
    n356 , 
    n357 , 
    n358 , 
    n359 , 
    n360 , 
    n361 , 
    n362 , 
    n363 , 
    n364 , 
    n365 , 
    n366 , 
    n367 , 
    n368 , 
    n369 , 
    n370 , 
    n371 , 
    n372 , 
    n373 , 
    n374 , 
    n375 , 
    n376 , 
    n377 , 
    n378 , 
    n379 , 
    n380 , 
    n381 , 
    n382 , 
    n383 , 
    n384 , 
    n385 , 
    n386 , 
    n387 , 
    n388 , 
    n389 , 
    n390 , 
    n391 , 
    n392 , 
    n393 , 
    n394 , 
    n395 , 
    n396 , 
    n397 , 
    n398 , 
    n399 , 
    n400 , 
    n401 , 
    n402 , 
    n403 , 
    n404 , 
    n405 , 
    n406 , 
    n407 , 
    n408 , 
    n409 , 
    n410 , 
    n411 , 
    n412 , 
    n413 , 
    n414 , 
    n415 , 
    n416 , 
    n417 , 
    n418 , 
    n419 , 
    n420 , 
    n421 , 
    n422 , 
    n423 , 
    n424 , 
    n425 , 
    n426 , 
    n427 , 
    n428 , 
    n429 , 
    n430 , 
    n431 , 
    n432 , 
    n433 , 
    n434 , 
    n435 , 
    n436 , 
    n437 , 
    n438 , 
    n439 , 
    n440 , 
    n441 , 
    n442 , 
    n443 , 
    n444 , 
    n445 , 
    n446 , 
    n447 , 
    n448 , 
    n449 , 
    n450 , 
    n451 , 
    n452 , 
    n453 , 
    n454 , 
    n455 , 
    n456 , 
    n457 , 
    n458 , 
    n459 , 
    n460 , 
    n461 , 
    n462 , 
    n463 , 
    n464 , 
    n465 , 
    n466 , 
    n467 , 
    n468 , 
    n469 , 
    n470 , 
    n471 , 
    n472 , 
    n473 , 
    n474 , 
    n475 , 
    n476 , 
    n477 , 
    n478 , 
    n479 , 
    n480 , 
    n481 , 
    n482 , 
    n483 , 
    n484 , 
    n485 , 
    n486 , 
    n487 , 
    n488 , 
    n489 , 
    n490 , 
    n491 , 
    n492 , 
    n493 , 
    n494 , 
    n495 , 
    n496 , 
    n497 , 
    n498 , 
    n499 , 
    n500 , 
    n501 , 
    n502 , 
    n503 , 
    n504 , 
    n505 , 
    n506 , 
    n507 , 
    n508 , 
    n509 , 
    n510 , 
    n511 , 
    n512 , 
    n513 , 
    n514 , 
    n515 , 
    n516 , 
    n517 , 
    n518 , 
    n519 , 
    n520 , 
    n521 , 
    n522 , 
    n523 , 
    n524 , 
    n525 , 
    n526 , 
    n527 , 
    n528 , 
    n529 , 
    n530 , 
    n531 , 
    n532 , 
    n533 , 
    n534 , 
    n535 , 
    n536 , 
    n537 , 
    n538 , 
    n539 , 
    n540 , 
    n541 , 
    n542 , 
    n543 , 
    n544 ;

wire 
    n1090 , 
    n1091 , 
    n1092 , 
    n1093 , 
    n1094 , 
    n1095 , 
    n1096 , 
    n1097 , 
    n1098 , 
    n1099 , 
    n1100 , 
    n1101 , 
    n1102 , 
    n1103 , 
    n1104 , 
    n1105 , 
    n1106 , 
    n1107 , 
    n1108 , 
    n1109 , 
    n1110 , 
    n1111 , 
    n1112 , 
    n1113 , 
    n1114 , 
    n1115 , 
    n1116 , 
    n1117 , 
    n1118 , 
    n1119 , 
    n1120 , 
    n1121 , 
    n1122 , 
    n1123 , 
    n1124 , 
    n1125 , 
    n1126 , 
    n1127 , 
    n1128 , 
    n1129 , 
    n1130 , 
    n1131 , 
    n1132 , 
    n1133 , 
    n1134 , 
    n1135 , 
    n1136 , 
    n1137 , 
    n1138 , 
    n1139 , 
    n1140 , 
    n1141 , 
    n1142 , 
    n1143 , 
    n1144 , 
    n1145 , 
    n1146 , 
    n1147 , 
    n1148 , 
    n1149 , 
    n1150 , 
    n1151 , 
    n1152 , 
    n1153 , 
    n1154 , 
    n1155 , 
    n1156 , 
    n1157 , 
    n1158 , 
    n1159 , 
    n1160 , 
    n1161 , 
    n1162 , 
    n1163 , 
    n1164 , 
    n1165 , 
    n1166 , 
    n1167 , 
    n1168 , 
    n1169 , 
    n1170 , 
    n1171 , 
    n1172 , 
    n1173 , 
    n1174 , 
    n1175 , 
    n1176 , 
    n1177 , 
    n1178 , 
    n1179 , 
    n1180 , 
    n1181 , 
    n1182 , 
    n1183 , 
    n1184 , 
    n1185 , 
    n1186 , 
    n1187 , 
    n1188 , 
    n1189 , 
    n1190 , 
    n1191 , 
    n1192 , 
    n1193 , 
    n1194 , 
    n1195 , 
    n1196 , 
    n1197 , 
    n1198 , 
    n1199 , 
    n1200 , 
    n1201 , 
    n1202 , 
    n1203 , 
    n1204 , 
    n1205 , 
    n1206 , 
    n1207 , 
    n1208 , 
    n1209 , 
    n1210 , 
    n1211 , 
    n1212 , 
    n1213 , 
    n1214 , 
    n1215 , 
    n1216 , 
    n1217 , 
    n1218 , 
    n1219 , 
    n1220 , 
    n1221 , 
    n1222 , 
    n1223 , 
    n1224 , 
    n1225 , 
    n1226 , 
    n1227 , 
    n1228 , 
    n1229 , 
    n1230 , 
    n1231 , 
    n1232 , 
    n1233 , 
    n1234 , 
    n1235 , 
    n1236 , 
    n1237 , 
    n1238 , 
    n1239 , 
    n1240 , 
    n1241 , 
    n1242 , 
    n1243 , 
    n1244 , 
    n1245 , 
    n1246 , 
    n1247 , 
    n1248 , 
    n1249 , 
    n1250 , 
    n1251 , 
    n1252 , 
    n1253 , 
    n1254 , 
    n1255 , 
    n1256 , 
    n1257 , 
    n1258 , 
    n1259 , 
    n1260 , 
    n1261 , 
    n1262 , 
    n1263 , 
    n1264 , 
    n1265 , 
    n1266 , 
    n1267 , 
    n1268 , 
    n1269 , 
    n1270 , 
    n1271 , 
    n1272 , 
    n1273 , 
    n1274 , 
    n1275 , 
    n1276 , 
    n1277 , 
    n1278 , 
    n1279 , 
    n1280 , 
    n1281 , 
    n1282 , 
    n1283 , 
    n1284 , 
    n1285 , 
    n1286 , 
    n1287 , 
    n1288 , 
    n1289 , 
    n1290 , 
    n1291 , 
    n1292 , 
    n1293 , 
    n1294 , 
    n1295 , 
    n1296 , 
    n1297 , 
    n1298 , 
    n1299 , 
    n1300 , 
    n1301 , 
    n1302 , 
    n1303 , 
    n1304 , 
    n1305 , 
    n1306 , 
    n1307 , 
    n1308 , 
    n1309 , 
    n1310 , 
    n1311 , 
    n1312 , 
    n1313 , 
    n1314 , 
    n1315 , 
    n1316 , 
    n1317 , 
    n1318 , 
    n1319 , 
    n1320 , 
    n1321 , 
    n1322 , 
    n1323 , 
    n1324 , 
    n1325 , 
    n1326 , 
    n1327 , 
    n1328 , 
    n1329 , 
    n1330 , 
    n1331 , 
    n1332 , 
    n1333 , 
    n1334 , 
    n1335 , 
    n1336 , 
    n1337 , 
    n1338 , 
    n1339 , 
    n1340 , 
    n1341 , 
    n1342 , 
    n1343 , 
    n1344 , 
    n1345 , 
    n1346 , 
    n1347 , 
    n1348 , 
    n1349 , 
    n1350 , 
    n1351 , 
    n1352 , 
    n1353 , 
    n1354 , 
    n1355 , 
    n1356 , 
    n1357 , 
    n1358 , 
    n1359 , 
    n1360 , 
    n1361 , 
    n1362 , 
    n1363 , 
    n1364 , 
    n1365 , 
    n1366 , 
    n1367 , 
    n1368 , 
    n1369 , 
    n1370 , 
    n1371 , 
    n1372 , 
    n1373 , 
    n1374 , 
    n1375 , 
    n1376 , 
    n1377 , 
    n1378 , 
    n1379 , 
    n1380 , 
    n1381 , 
    n1382 , 
    n1383 , 
    n1384 , 
    n1385 , 
    n1386 , 
    n1387 , 
    n1388 , 
    n1389 , 
    n1390 , 
    n1391 , 
    n1392 , 
    n1393 , 
    n1394 , 
    n1395 , 
    n1396 , 
    n1397 , 
    n1398 , 
    n1399 , 
    n1400 , 
    n1401 , 
    n1402 , 
    n1403 , 
    n1404 , 
    n1405 , 
    n1406 , 
    n1407 , 
    n1408 , 
    n1409 , 
    n1410 , 
    n1411 , 
    n1412 , 
    n1413 , 
    n1414 , 
    n1415 , 
    n1416 , 
    n1417 , 
    n1418 , 
    n1419 , 
    n1420 , 
    n1421 , 
    n1422 , 
    n1423 , 
    n1424 , 
    n1425 , 
    n1426 , 
    n1427 , 
    n1428 , 
    n1429 , 
    n1430 , 
    n1431 , 
    n1432 , 
    n1433 , 
    n1434 , 
    n1435 , 
    n1436 , 
    n1437 , 
    n1438 , 
    n1439 , 
    n1440 , 
    n1441 , 
    n1442 , 
    n1443 , 
    n1444 , 
    n1445 , 
    n1446 , 
    n1447 , 
    n1448 , 
    n1449 , 
    n1450 , 
    n1451 , 
    n1452 , 
    n1453 , 
    n1454 , 
    n1455 , 
    n1456 , 
    n1457 , 
    n1458 , 
    n1459 , 
    n1460 , 
    n1461 , 
    n1462 , 
    n1463 , 
    n1464 , 
    n1465 , 
    n1466 , 
    n1467 , 
    n1468 , 
    n1469 , 
    n1470 , 
    n1471 , 
    n1472 , 
    n1473 , 
    n1474 , 
    n1475 , 
    n1476 , 
    n1477 , 
    n1478 , 
    n1479 , 
    n1480 , 
    n1481 , 
    n1482 , 
    n1483 , 
    n1484 , 
    n1485 , 
    n1486 , 
    n1487 , 
    n1488 , 
    n1489 , 
    n1490 , 
    n1491 , 
    n1492 , 
    n1493 , 
    n1494 , 
    n1495 , 
    n1496 , 
    n1497 , 
    n1498 , 
    n1499 , 
    n1500 , 
    n1501 , 
    n1502 , 
    n1503 , 
    n1504 , 
    n1505 , 
    n1506 , 
    n1507 , 
    n1508 , 
    n1509 , 
    n1510 , 
    n1511 , 
    n1512 , 
    n1513 , 
    n1514 , 
    n1515 , 
    n1516 , 
    n1517 , 
    n1518 , 
    n1519 , 
    n1520 , 
    n1521 , 
    n1522 , 
    n1523 , 
    n1524 , 
    n1525 , 
    n1526 , 
    n1527 , 
    n1528 , 
    n1529 , 
    n1530 , 
    n1531 , 
    n1532 , 
    n1533 , 
    n1534 , 
    n1535 , 
    n1536 , 
    n1537 , 
    n1538 , 
    n1539 , 
    n1540 , 
    n1541 , 
    n1542 , 
    n1543 , 
    n1544 , 
    n1545 , 
    n1546 , 
    n1547 , 
    n1548 , 
    n1549 , 
    n1550 , 
    n1551 , 
    n1552 , 
    n1553 , 
    n1554 , 
    n1555 , 
    n1556 , 
    n1557 , 
    n1558 , 
    n1559 , 
    n1560 , 
    n1561 , 
    n1562 , 
    n1563 , 
    n1564 , 
    n1565 , 
    n1566 , 
    n1567 , 
    n1568 , 
    n1569 , 
    n1570 , 
    n1571 , 
    n1572 , 
    n1573 , 
    n1574 , 
    n1575 , 
    n1576 , 
    n1577 , 
    n1578 , 
    n1579 , 
    n1580 , 
    n1581 , 
    n1582 , 
    n1583 , 
    n1584 , 
    n1585 , 
    n1586 , 
    n1587 , 
    n1588 , 
    n1589 , 
    n1590 , 
    n1591 , 
    n1592 , 
    n1593 , 
    n1594 , 
    n1595 , 
    n1596 , 
    n1597 , 
    n1598 , 
    n1599 , 
    n1600 , 
    n1601 , 
    n1602 , 
    n1603 , 
    n1604 , 
    n1605 , 
    n1606 , 
    n1607 , 
    n1608 , 
    n1609 , 
    n1610 , 
    n1611 , 
    n1612 , 
    n1613 , 
    n1614 , 
    n1615 , 
    n1616 , 
    n1617 , 
    n1618 , 
    n1619 , 
    n1620 , 
    n1621 , 
    n1622 , 
    n1623 , 
    n1624 , 
    n1625 , 
    n1626 , 
    n1627 , 
    n1628 , 
    n1629 , 
    n1630 , 
    n1631 , 
    n1632 , 
    n1633 , 
    n1634 ;
wire n528834 , n528835 , n528836 , n528837 , n528838 , n528839 , n528840 , n528841 , n528842 , 
     n528843 , n528844 , n528845 , n528846 , n528847 , n528848 , n528849 , n528850 , n528851 , n528852 , 
     n528853 , n528854 , n528855 , n528856 , n528857 , n528858 , n528859 , n528860 , n528861 , n528862 , 
     n528863 , n528864 , n528865 , n528866 , n528867 , n528868 , n528869 , n528870 , n528871 , n528872 , 
     n528873 , n528874 , n528875 , n528876 , n528877 , n528878 , n528879 , n528880 , n528881 , n528882 , 
     n528883 , n528884 , n528885 , n528886 , n528887 , n528888 , n528889 , n528890 , n528891 , n528892 , 
     n528893 , n528894 , n528895 , n528896 , n528897 , n528898 , n528899 , n528900 , n528901 , n528902 , 
     n528903 , n528904 , n528905 , n528906 , n528907 , n528908 , n528909 , n528910 , n528911 , n528912 , 
     n528913 , n528914 , n528915 , n528916 , n528917 , n528918 , n528919 , n528920 , n528921 , n528922 , 
     n528923 , n528924 , n528925 , n528926 , n528927 , n528928 , n528929 , n528930 , n528931 , n528932 , 
     n528933 , n528934 , n528935 , n528936 , n528937 , n528938 , n528939 , n528940 , n528941 , n528942 , 
     n528943 , n528944 , n528945 , n528946 , n528947 , n528948 , n528949 , n528950 , n528951 , n528952 , 
     n528953 , n528954 , n528955 , n528956 , n528957 , n528958 , n528959 , n528960 , n528961 , n528962 , 
     n528963 , n528964 , n528965 , n528966 , n528967 , n528968 , n528969 , n528970 , n528971 , n528972 , 
     n528973 , n528974 , n528975 , n528976 , n528977 , n528978 , n528979 , n528980 , n528981 , n528982 , 
     n528983 , n528984 , n528985 , n528986 , n528987 , n528988 , n528989 , n528990 , n528991 , n528992 , 
     n528993 , n528994 , n528995 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , 
     n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , 
     n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , 
     n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , 
     n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , 
     n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , 
     n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , 
     n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , 
     n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , 
     n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , 
     n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , 
     n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , 
     n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , 
     n529123 , n529124 , n529125 , n529126 , n529127 , n529128 , n529129 , n529130 , n529131 , n1874 , 
     n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n529140 , n1883 , n529142 , 
     n1885 , n529144 , n1887 , n1888 , n529147 , n1890 , n1891 , n1892 , n1893 , n1894 , 
     n529153 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n529161 , n1904 , 
     n529163 , n1906 , n529165 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n529172 , 
     n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n529181 , n1924 , 
     n529183 , n1926 , n1927 , n1928 , n1929 , n1930 , n529189 , n1932 , n529191 , n1934 , 
     n529193 , n1936 , n1937 , n1938 , n1939 , n1940 , n529199 , n1942 , n529201 , n1944 , 
     n529203 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n529210 , n1953 , n1954 , 
     n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n529219 , n1962 , n529221 , n1964 , 
     n529223 , n1966 , n1967 , n529226 , n1969 , n1970 , n1971 , n1972 , n1973 , n529232 , 
     n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , 
     n1985 , n529244 , n1987 , n529246 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , 
     n529253 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n529261 , n2004 , 
     n529263 , n2006 , n529265 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n529272 , 
     n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n529281 , n2024 , 
     n529283 , n2026 , n529285 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n529292 , 
     n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , 
     n2045 , n2046 , n2047 , n529306 , n2049 , n529308 , n2050 , n2051 , n2052 , n2053 , 
     n2054 , n2055 , n529315 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , 
     n529323 , n2065 , n529325 , n2067 , n529327 , n2069 , n2070 , n2071 , n2072 , n2073 , 
     n2074 , n529334 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , 
     n529343 , n2085 , n529345 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n529352 , 
     n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , 
     n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , 
     n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , 
     n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , 
     n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , 
     n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , 
     n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , 
     n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , 
     n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , 
     n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , 
     n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , 
     n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , 
     n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , 
     n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , 
     n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , 
     n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , 
     n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , 
     n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , 
     n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , 
     n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , 
     n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , 
     n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , 
     n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , 
     n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , 
     n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , 
     n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , 
     n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , 
     n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , 
     n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , 
     n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , 
     n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n529659 , n2401 , n2402 , n2403 , 
     n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , 
     n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , 
     n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , 
     n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , 
     n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , 
     n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , 
     n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , 
     n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , 
     n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , 
     n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , 
     n2504 , n2505 , n2506 , n2507 , n2508 , n529768 , n2510 , n529770 , n2512 , n2513 , 
     n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , 
     n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , 
     n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , 
     n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , 
     n2554 , n529814 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , 
     n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , 
     n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , 
     n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , 
     n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , 
     n529863 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , 
     n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , 
     n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , 
     n2633 , n2634 , n2635 , n2636 , n2637 , n529898 , n2639 , n2640 , n2641 , n2642 , 
     n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , 
     n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , 
     n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , 
     n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , 
     n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , 
     n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , 
     n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , 
     n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n529980 , n2721 , n529982 , 
     n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , 
     n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , 
     n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , 
     n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , 
     n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , 
     n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , 
     n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , 
     n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , 
     n2803 , n2804 , n530065 , n2806 , n530067 , n2808 , n2809 , n2810 , n2811 , n2812 , 
     n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , 
     n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , 
     n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , 
     n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , 
     n2853 , n2854 , n2855 , n2856 , n530117 , n2858 , n530119 , n2860 , n2861 , n2862 , 
     n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , 
     n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , 
     n2883 , n2884 , n530145 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , 
     n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , 
     n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , 
     n2913 , n2914 , n2915 , n2916 , n2917 , n530178 , n2919 , n2920 , n2921 , n2922 , 
     n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , 
     n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , 
     n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , 
     n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , 
     n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n530232 , 
     n2973 , n530234 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , 
     n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , 
     n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , 
     n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , 
     n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , 
     n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , 
     n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , 
     n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , 
     n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n530320 , n3061 , n3062 , 
     n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , 
     n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , 
     n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , 
     n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , 
     n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , 
     n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , 
     n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , 
     n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , 
     n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , 
     n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , 
     n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , 
     n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , 
     n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , 
     n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , 
     n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , 
     n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n530481 , n3222 , 
     n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , 
     n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , 
     n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , 
     n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , 
     n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , 
     n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n530540 , n3281 , n3282 , 
     n3283 , n3284 , n3285 , n530546 , n3287 , n530548 , n3289 , n3290 , n3291 , n3292 , 
     n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , 
     n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , 
     n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , 
     n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n530592 , 
     n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , 
     n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , 
     n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , 
     n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , 
     n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , 
     n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , 
     n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , 
     n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , 
     n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , 
     n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , 
     n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , 
     n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , 
     n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , 
     n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , 
     n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , 
     n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , 
     n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , 
     n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , 
     n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n530781 , n3522 , 
     n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , 
     n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , 
     n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , 
     n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , 
     n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , 
     n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , 
     n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , 
     n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , 
     n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , 
     n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , 
     n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , 
     n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , 
     n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , 
     n3653 , n3654 , n3655 , n3656 , n3657 , n530918 , n3659 , n3660 , n3661 , n3662 , 
     n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , 
     n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , 
     n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , 
     n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , 
     n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , 
     n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , 
     n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , 
     n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , 
     n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , 
     n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , 
     n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , 
     n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , 
     n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , 
     n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n531059 , n3800 , n3801 , n3802 , 
     n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n531072 , 
     n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , 
     n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , 
     n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , 
     n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , 
     n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , 
     n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , 
     n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , 
     n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , 
     n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , 
     n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , 
     n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , 
     n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , 
     n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , 
     n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , 
     n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , 
     n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , 
     n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , 
     n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , 
     n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , 
     n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , 
     n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , 
     n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , 
     n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , 
     n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , 
     n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , 
     n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , 
     n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , 
     n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , 
     n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , 
     n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , 
     n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , 
     n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , 
     n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , 
     n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , 
     n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , 
     n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , 
     n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , 
     n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , 
     n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , 
     n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , 
     n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , 
     n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , 
     n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , 
     n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , 
     n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , 
     n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , 
     n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , 
     n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , 
     n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , 
     n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , 
     n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , 
     n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , 
     n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , 
     n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , 
     n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , 
     n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , 
     n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , 
     n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , 
     n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , 
     n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , 
     n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , 
     n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , 
     n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , 
     n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , 
     n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , 
     n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , 
     n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , 
     n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , 
     n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , 
     n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , 
     n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , 
     n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , 
     n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , 
     n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , 
     n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , 
     n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , 
     n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , 
     n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , 
     n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , 
     n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , 
     n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , 
     n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , 
     n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , 
     n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , 
     n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , 
     n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , 
     n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , 
     n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , 
     n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , 
     n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , 
     n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , 
     n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , 
     n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , 
     n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , 
     n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , 
     n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , 
     n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , 
     n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , 
     n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , 
     n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , 
     n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , 
     n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , 
     n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , 
     n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , 
     n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , 
     n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , 
     n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , 
     n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , 
     n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , 
     n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , 
     n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , 
     n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , 
     n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , 
     n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , 
     n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , 
     n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , 
     n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , 
     n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , 
     n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , 
     n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , 
     n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , 
     n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , 
     n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , 
     n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , 
     n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , 
     n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , 
     n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , 
     n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , 
     n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , 
     n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , 
     n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , 
     n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , 
     n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , 
     n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , 
     n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , 
     n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , 
     n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , 
     n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , 
     n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , 
     n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , 
     n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , 
     n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , 
     n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , 
     n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , 
     n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , 
     n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , 
     n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , 
     n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , 
     n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , 
     n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , 
     n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , 
     n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , 
     n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , 
     n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , 
     n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , 
     n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , 
     n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , 
     n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , 
     n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , 
     n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , 
     n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , 
     n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , 
     n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , 
     n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , 
     n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , 
     n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , 
     n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , 
     n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , 
     n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , 
     n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , 
     n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , 
     n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , 
     n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , 
     n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , 
     n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , 
     n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , 
     n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , 
     n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , 
     n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , 
     n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , 
     n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , 
     n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , 
     n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , 
     n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , 
     n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , 
     n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , 
     n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , 
     n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , 
     n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , 
     n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , 
     n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , 
     n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , 
     n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , 
     n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , 
     n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , 
     n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , 
     n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , 
     n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , 
     n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , 
     n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , 
     n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , 
     n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , 
     n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , 
     n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , 
     n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , 
     n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , 
     n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , 
     n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , 
     n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , 
     n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , 
     n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , 
     n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , 
     n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , 
     n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , 
     n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , 
     n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , 
     n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , 
     n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , 
     n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , 
     n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , 
     n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , 
     n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , 
     n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , 
     n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , 
     n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , 
     n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , 
     n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , 
     n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , 
     n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , 
     n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , 
     n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , 
     n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , 
     n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , 
     n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , 
     n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , 
     n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , 
     n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , 
     n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , 
     n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , 
     n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , 
     n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , 
     n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , 
     n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , 
     n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , 
     n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , 
     n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , 
     n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , 
     n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , 
     n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , 
     n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , 
     n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , 
     n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , 
     n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , 
     n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , 
     n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , 
     n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , 
     n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , 
     n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , 
     n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , 
     n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , 
     n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , 
     n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , 
     n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , 
     n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , 
     n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , 
     n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , 
     n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , 
     n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , 
     n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , 
     n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , 
     n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , 
     n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , 
     n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , 
     n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , 
     n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , 
     n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , 
     n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , 
     n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , 
     n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , 
     n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n533872 , 
     n533873 , n6614 , n533875 , n533876 , n6617 , n533878 , n533879 , n6620 , n533881 , n533882 , 
     n6623 , n533884 , n533885 , n6626 , n533887 , n533888 , n6629 , n533890 , n533891 , n6632 , 
     n533893 , n533894 , n6635 , n533896 , n533897 , n6638 , n533899 , n533900 , n6641 , n533902 , 
     n533903 , n6644 , n533905 , n533906 , n6647 , n533908 , n533909 , n6650 , n533911 , n533912 , 
     n6653 , n533914 , n533915 , n6656 , n533917 , n533918 , n6659 , n533920 , n533921 , n6662 , 
     n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , 
     n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , 
     n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , 
     n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , 
     n6703 , n6704 , n6705 , n533966 , n533967 , n6708 , n6709 , n6710 , n533971 , n533972 , 
     n6713 , n6714 , n6715 , n6716 , n533977 , n533978 , n6719 , n6720 , n6721 , n6722 , 
     n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , 
     n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , 
     n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , 
     n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , 
     n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , 
     n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , 
     n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , 
     n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , 
     n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , 
     n6813 , n534074 , n534075 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , 
     n6823 , n534084 , n534085 , n6826 , n534087 , n534088 , n6829 , n534090 , n534091 , n6832 , 
     n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n534101 , n534102 , 
     n6843 , n6844 , n6845 , n534106 , n534107 , n6848 , n6849 , n6850 , n6851 , n6852 , 
     n6853 , n6854 , n534115 , n534116 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , 
     n6863 , n6864 , n6865 , n534126 , n534127 , n6868 , n534129 , n534130 , n6871 , n534132 , 
     n534133 , n6874 , n534135 , n534136 , n6877 , n534138 , n534139 , n6880 , n534141 , n534142 , 
     n6883 , n534144 , n534145 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , 
     n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , 
     n6903 , n6904 , n6905 , n6906 , n534167 , n534168 , n6909 , n6910 , n6911 , n534172 , 
     n534173 , n6914 , n6915 , n6916 , n6917 , n534178 , n534179 , n6920 , n6921 , n6922 , 
     n6923 , n6924 , n6925 , n534186 , n534187 , n6928 , n6929 , n6930 , n6931 , n6932 , 
     n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , 
     n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , 
     n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , 
     n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , 
     n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , 
     n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , 
     n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , 
     n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , 
     n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n534280 , n534281 , n7022 , 
     n7023 , n7024 , n534285 , n534286 , n7027 , n7028 , n7029 , n7030 , n534291 , n534292 , 
     n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , 
     n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , 
     n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , 
     n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , 
     n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , 
     n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , 
     n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , 
     n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , 
     n7113 , n7114 , n7115 , n7116 , n7117 , n534378 , n534379 , n7120 , n7121 , n7122 , 
     n7123 , n7124 , n7125 , n7126 , n7127 , n534388 , n534389 , n7130 , n7131 , n7132 , 
     n534393 , n534394 , n7135 , n7136 , n7137 , n7138 , n534399 , n534400 , n7141 , n7142 , 
     n7143 , n7144 , n7145 , n7146 , n534407 , n534408 , n7149 , n7150 , n7151 , n7152 , 
     n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , 
     n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , 
     n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , 
     n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , 
     n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , 
     n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , 
     n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , 
     n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , 
     n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , 
     n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , 
     n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , 
     n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , 
     n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , 
     n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , 
     n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , 
     n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , 
     n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , 
     n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , 
     n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , 
     n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , 
     n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , 
     n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , 
     n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , 
     n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , 
     n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , 
     n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , 
     n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , 
     n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , 
     n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , 
     n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , 
     n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , 
     n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , 
     n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , 
     n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , 
     n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , 
     n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , 
     n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , 
     n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , 
     n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , 
     n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , 
     n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , 
     n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , 
     n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , 
     n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , 
     n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , 
     n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , 
     n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , 
     n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , 
     n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , 
     n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , 
     n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , 
     n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n534929 , n534930 , n7671 , n7672 , 
     n7673 , n534934 , n534935 , n7676 , n7677 , n534938 , n534939 , n7680 , n7681 , n7682 , 
     n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , 
     n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , 
     n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n534969 , n534970 , n7711 , n7712 , 
     n7713 , n7714 , n7715 , n534976 , n534977 , n7718 , n7719 , n7720 , n534981 , n534982 , 
     n7723 , n7724 , n7725 , n534986 , n534987 , n7728 , n7729 , n7730 , n7731 , n7732 , 
     n7733 , n7734 , n534995 , n534996 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , 
     n7743 , n7744 , n7745 , n535006 , n535007 , n7748 , n7749 , n7750 , n535011 , n535012 , 
     n7753 , n7754 , n7755 , n535016 , n535017 , n7758 , n7759 , n7760 , n7761 , n7762 , 
     n7763 , n7764 , n535025 , n535026 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , 
     n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n535041 , n535042 , 
     n7783 , n7784 , n7785 , n535046 , n535047 , n7788 , n7789 , n7790 , n535051 , n535052 , 
     n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n535060 , n535061 , n7802 , 
     n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n535070 , n535071 , n7812 , 
     n7813 , n7814 , n535075 , n535076 , n7817 , n7818 , n7819 , n535080 , n535081 , n7822 , 
     n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n535089 , n535090 , n7831 , n7832 , 
     n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n535101 , n535102 , 
     n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n535110 , n535111 , n7852 , 
     n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , 
     n7863 , n7864 , n7865 , n7866 , n7867 , n535128 , n535129 , n7870 , n7871 , n7872 , 
     n7873 , n7874 , n7875 , n7876 , n535137 , n535138 , n7879 , n7880 , n7881 , n7882 , 
     n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , 
     n7893 , n7894 , n7895 , n535156 , n535157 , n7898 , n535159 , n535160 , n7901 , n535162 , 
     n535163 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , 
     n535173 , n535174 , n7915 , n7916 , n7917 , n535178 , n535179 , n7920 , n7921 , n7922 , 
     n7923 , n7924 , n7925 , n7926 , n535187 , n535188 , n7929 , n7930 , n7931 , n7932 , 
     n7933 , n7934 , n7935 , n7936 , n535197 , n535198 , n7939 , n535200 , n535201 , n535202 , 
     n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n535212 , 
     n535213 , n7954 , n7955 , n7956 , n535217 , n535218 , n7959 , n7960 , n7961 , n7962 , 
     n7963 , n7964 , n7965 , n535226 , n535227 , n7968 , n7969 , n7970 , n7971 , n7972 , 
     n7973 , n7974 , n7975 , n7976 , n535237 , n535238 , n7979 , n535240 , n535241 , n7982 , 
     n7983 , n7984 , n535245 , n535246 , n7987 , n7988 , n535249 , n535250 , n7991 , n7992 , 
     n7993 , n7994 , n7995 , n7996 , n7997 , n535258 , n535259 , n8000 , n8001 , n8002 , 
     n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , 
     n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n535279 , n535280 , n8021 , n8022 , 
     n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , 
     n8033 , n8034 , n8035 , n8036 , n535297 , n535298 , n8039 , n8040 , n8041 , n8042 , 
     n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , 
     n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , 
     n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n535329 , n535330 , n8071 , n8072 , 
     n8073 , n535334 , n535335 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , 
     n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n535349 , n535350 , n8091 , n535352 , 
     n535353 , n8094 , n8095 , n8096 , n535357 , n535358 , n8099 , n8100 , n535361 , n535362 , 
     n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n535369 , n535370 , n8111 , n8112 , 
     n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , 
     n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , 
     n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , 
     n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , 
     n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , 
     n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , 
     n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , 
     n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , 
     n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , 
     n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , 
     n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , 
     n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , 
     n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , 
     n535503 , n535504 , n8245 , n8246 , n535507 , n535508 , n8249 , n8250 , n8251 , n8252 , 
     n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , 
     n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , 
     n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , 
     n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , 
     n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , 
     n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , 
     n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , 
     n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n535592 , 
     n535593 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , 
     n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , 
     n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , 
     n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , 
     n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , 
     n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , 
     n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , 
     n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , 
     n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , 
     n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , 
     n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , 
     n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , 
     n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , 
     n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , 
     n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , 
     n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , 
     n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , 
     n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , 
     n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , 
     n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , 
     n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , 
     n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , 
     n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , 
     n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , 
     n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , 
     n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , 
     n535853 , n535854 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n535862 , 
     n535863 , n8604 , n8605 , n8606 , n535867 , n535868 , n8609 , n8610 , n8611 , n8612 , 
     n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , 
     n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , 
     n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , 
     n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , 
     n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , 
     n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , 
     n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , 
     n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , 
     n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , 
     n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , 
     n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , 
     n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , 
     n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , 
     n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , 
     n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , 
     n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , 
     n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , 
     n536043 , n536044 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , 
     n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , 
     n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , 
     n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , 
     n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , 
     n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , 
     n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , 
     n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , 
     n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , 
     n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , 
     n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , 
     n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , 
     n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , 
     n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , 
     n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , 
     n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , 
     n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , 
     n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , 
     n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , 
     n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , 
     n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , 
     n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , 
     n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , 
     n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , 
     n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , 
     n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , 
     n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , 
     n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , 
     n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , 
     n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n536342 , 
     n536343 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , 
     n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , 
     n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , 
     n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , 
     n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , 
     n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , 
     n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , 
     n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n536420 , n536421 , n9162 , 
     n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , 
     n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , 
     n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , 
     n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , 
     n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , 
     n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , 
     n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , 
     n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , 
     n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , 
     n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , 
     n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , 
     n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , 
     n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , 
     n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , 
     n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , 
     n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , 
     n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , 
     n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , 
     n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , 
     n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , 
     n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , 
     n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , 
     n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , 
     n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , 
     n9403 , n9404 , n9405 , n9406 , n9407 , n536668 , n536669 , n9410 , n9411 , n9412 , 
     n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , 
     n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , 
     n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , 
     n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , 
     n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , 
     n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , 
     n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n536740 , n536741 , n9482 , 
     n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , 
     n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , 
     n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , 
     n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , 
     n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , 
     n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , 
     n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , 
     n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , 
     n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , 
     n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , 
     n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , 
     n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , 
     n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , 
     n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , 
     n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , 
     n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , 
     n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , 
     n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , 
     n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , 
     n9673 , n536934 , n536935 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , 
     n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , 
     n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , 
     n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , 
     n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , 
     n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , 
     n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , 
     n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , 
     n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , 
     n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , 
     n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , 
     n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , 
     n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , 
     n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n537071 , n9812 , 
     n537073 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , 
     n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , 
     n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , 
     n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , 
     n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , 
     n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , 
     n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , 
     n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , 
     n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , 
     n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , 
     n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , 
     n537183 , n537184 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , 
     n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , 
     n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , 
     n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , 
     n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , 
     n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , 
     n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , 
     n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , 
     n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , 
     n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , 
     n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , 
     n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , 
     n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , 
     n537313 , n537314 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , 
     n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , 
     n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , 
     n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , 
     n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , 
     n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , 
     n10113 , n10114 , n10115 , n10116 , n10117 , n537378 , n537379 , n10120 , n10121 , n10122 , 
     n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , 
     n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , 
     n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , 
     n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , 
     n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , 
     n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , 
     n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , 
     n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , 
     n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , 
     n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , 
     n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , 
     n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , 
     n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , 
     n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , 
     n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , 
     n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , 
     n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , 
     n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , 
     n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , 
     n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , 
     n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , 
     n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , 
     n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , 
     n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , 
     n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , 
     n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , 
     n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , 
     n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , 
     n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , 
     n10413 , n10414 , n10415 , n10416 , n537677 , n537678 , n10419 , n10420 , n10421 , n10422 , 
     n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , 
     n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , 
     n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , 
     n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , 
     n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , 
     n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , 
     n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , 
     n10493 , n10494 , n10495 , n10496 , n537757 , n537758 , n10499 , n10500 , n10501 , n10502 , 
     n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , 
     n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , 
     n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , 
     n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , 
     n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , 
     n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , 
     n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , 
     n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , 
     n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , 
     n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , 
     n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , 
     n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , 
     n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , 
     n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , 
     n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , 
     n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , 
     n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , 
     n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , 
     n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , 
     n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , 
     n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , 
     n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , 
     n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , 
     n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , 
     n10743 , n10744 , n538005 , n538006 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , 
     n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , 
     n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , 
     n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , 
     n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , 
     n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , 
     n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , 
     n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , 
     n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , 
     n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n538100 , n538101 , n10842 , 
     n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , 
     n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , 
     n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , 
     n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , 
     n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , 
     n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , 
     n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , 
     n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , 
     n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , 
     n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , 
     n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , 
     n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , 
     n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , 
     n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , 
     n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , 
     n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , 
     n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , 
     n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , 
     n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , 
     n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , 
     n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , 
     n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , 
     n11063 , n11064 , n11065 , n538326 , n538327 , n11068 , n11069 , n11070 , n11071 , n11072 , 
     n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , 
     n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , 
     n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , 
     n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , 
     n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , 
     n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , 
     n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , 
     n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , 
     n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , 
     n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , 
     n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , 
     n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , 
     n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , 
     n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , 
     n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , 
     n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , 
     n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , 
     n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , 
     n11253 , n11254 , n11255 , n11256 , n11257 , n538518 , n538519 , n11260 , n11261 , n11262 , 
     n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , 
     n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , 
     n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , 
     n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , 
     n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , 
     n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , 
     n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , 
     n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , 
     n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , 
     n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , 
     n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , 
     n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , 
     n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , 
     n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , 
     n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n538671 , n538672 , 
     n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , 
     n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , 
     n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , 
     n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , 
     n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , 
     n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , 
     n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , 
     n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , 
     n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , 
     n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , 
     n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , 
     n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , 
     n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , 
     n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , 
     n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , 
     n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , 
     n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n538839 , n538840 , n11581 , n11582 , 
     n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , 
     n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , 
     n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , 
     n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , 
     n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , 
     n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , 
     n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , 
     n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , 
     n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , 
     n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , 
     n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , 
     n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , 
     n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , 
     n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , 
     n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , 
     n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , 
     n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , 
     n11753 , n11754 , n539015 , n539016 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , 
     n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , 
     n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , 
     n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , 
     n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , 
     n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , 
     n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , 
     n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , 
     n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , 
     n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , 
     n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n539120 , n539121 , n11862 , 
     n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , 
     n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , 
     n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , 
     n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , 
     n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , 
     n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , 
     n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , 
     n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , 
     n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , 
     n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , 
     n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , 
     n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , 
     n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , 
     n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , 
     n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , 
     n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , 
     n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , 
     n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , 
     n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , 
     n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , 
     n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , 
     n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , 
     n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , 
     n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n539359 , n539360 , n12101 , n12102 , 
     n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , 
     n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , 
     n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , 
     n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , 
     n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , 
     n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , 
     n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , 
     n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , 
     n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , 
     n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , 
     n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , 
     n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , 
     n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , 
     n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , 
     n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n539512 , 
     n539513 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , 
     n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , 
     n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , 
     n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , 
     n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , 
     n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , 
     n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , 
     n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , 
     n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , 
     n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , 
     n12353 , n12354 , n12355 , n12356 , n539617 , n539618 , n12359 , n12360 , n12361 , n12362 , 
     n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , 
     n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , 
     n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , 
     n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , 
     n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , 
     n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , 
     n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , 
     n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , 
     n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , 
     n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , 
     n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , 
     n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , 
     n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , 
     n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , 
     n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , 
     n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n539780 , n539781 , n12522 , 
     n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , 
     n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , 
     n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , 
     n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , 
     n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , 
     n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , 
     n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , 
     n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , 
     n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , 
     n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , 
     n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , 
     n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , 
     n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , 
     n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , 
     n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , 
     n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , 
     n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , 
     n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , 
     n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , 
     n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , 
     n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , 
     n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , 
     n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , 
     n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , 
     n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , 
     n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n540041 , n540042 , 
     n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , 
     n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , 
     n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , 
     n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , 
     n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , 
     n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , 
     n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , 
     n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , 
     n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , 
     n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , 
     n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , 
     n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , 
     n12903 , n12904 , n540165 , n540166 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , 
     n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , 
     n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , 
     n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , 
     n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , 
     n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , 
     n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , 
     n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , 
     n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , 
     n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , 
     n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , 
     n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , 
     n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , 
     n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , 
     n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , 
     n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , 
     n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , 
     n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , 
     n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , 
     n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , 
     n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , 
     n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , 
     n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , 
     n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , 
     n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , 
     n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , 
     n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , 
     n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , 
     n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , 
     n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , 
     n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , 
     n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , 
     n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , 
     n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , 
     n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , 
     n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , 
     n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , 
     n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , 
     n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , 
     n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , 
     n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , 
     n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , 
     n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , 
     n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , 
     n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , 
     n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , 
     n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , 
     n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , 
     n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , 
     n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , 
     n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , 
     n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , 
     n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , 
     n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , 
     n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , 
     n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , 
     n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , 
     n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , 
     n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , 
     n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , 
     n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , 
     n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , 
     n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , 
     n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , 
     n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , 
     n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , 
     n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , 
     n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , 
     n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , 
     n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , 
     n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , 
     n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , 
     n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , 
     n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , 
     n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , 
     n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , 
     n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , 
     n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , 
     n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , 
     n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , 
     n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , 
     n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , 
     n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , 
     n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , 
     n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , 
     n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , 
     n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , 
     n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , 
     n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , 
     n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , 
     n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , 
     n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , 
     n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , 
     n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , 
     n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , 
     n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , 
     n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , 
     n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , 
     n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , 
     n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , 
     n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , 
     n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , 
     n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , 
     n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , 
     n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , 
     n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , 
     n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , 
     n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , 
     n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , 
     n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , 
     n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , 
     n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , 
     n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , 
     n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , 
     n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , 
     n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , 
     n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , 
     n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , 
     n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , 
     n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , 
     n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , 
     n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , 
     n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , 
     n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , 
     n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , 
     n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , 
     n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , 
     n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , 
     n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , 
     n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , 
     n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , 
     n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , 
     n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , 
     n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , 
     n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , 
     n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , 
     n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , 
     n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , 
     n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , 
     n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , 
     n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , 
     n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , 
     n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , 
     n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , 
     n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , 
     n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , 
     n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , 
     n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , 
     n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , 
     n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , 
     n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , 
     n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , 
     n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , 
     n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , 
     n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , 
     n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , 
     n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , 
     n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , 
     n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , 
     n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , 
     n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , 
     n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , 
     n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , 
     n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , 
     n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , 
     n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , 
     n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , 
     n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , 
     n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , 
     n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , 
     n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , 
     n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , 
     n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , 
     n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , 
     n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , 
     n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , 
     n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , 
     n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , 
     n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , 
     n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , 
     n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , 
     n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , 
     n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , 
     n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , 
     n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , 
     n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , 
     n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , 
     n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , 
     n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , 
     n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , 
     n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , 
     n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , 
     n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , 
     n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , 
     n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , 
     n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , 
     n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , 
     n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , 
     n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , 
     n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , 
     n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , 
     n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , 
     n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , 
     n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , 
     n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , 
     n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , 
     n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , 
     n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , 
     n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , 
     n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , 
     n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , 
     n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , 
     n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , 
     n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , 
     n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , 
     n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , 
     n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , 
     n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , 
     n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , 
     n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , 
     n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , 
     n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , 
     n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , 
     n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , 
     n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , 
     n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , 
     n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , 
     n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , 
     n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , 
     n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , 
     n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , 
     n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , 
     n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , 
     n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , 
     n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , 
     n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , 
     n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , 
     n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , 
     n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , 
     n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , 
     n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , 
     n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , 
     n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , 
     n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , 
     n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , 
     n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , 
     n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , 
     n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , 
     n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , 
     n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , 
     n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , 
     n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , 
     n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , 
     n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , 
     n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , 
     n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , 
     n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , 
     n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , 
     n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , 
     n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , 
     n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , 
     n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , 
     n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , 
     n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , 
     n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , 
     n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , 
     n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , 
     n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , 
     n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , 
     n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , 
     n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , 
     n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , 
     n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , 
     n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , 
     n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , 
     n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , 
     n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , 
     n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , 
     n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , 
     n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , 
     n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , 
     n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , 
     n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , 
     n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , 
     n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , 
     n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , 
     n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , 
     n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , 
     n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , 
     n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , 
     n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , 
     n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , 
     n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , 
     n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , 
     n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , 
     n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , 
     n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , 
     n15873 , n543134 , n543135 , n15876 , n543137 , n543138 , n15879 , n543140 , n543141 , n15882 , 
     n543143 , n543144 , n15885 , n543146 , n543147 , n15888 , n543149 , n543150 , n15891 , n543152 , 
     n543153 , n15894 , n543155 , n543156 , n15897 , n543158 , n543159 , n15900 , n543161 , n543162 , 
     n15903 , n543164 , n543165 , n15906 , n543167 , n543168 , n15909 , n543170 , n543171 , n15912 , 
     n543173 , n543174 , n15915 , n543176 , n543177 , n15918 , n543179 , n543180 , n15921 , n543182 , 
     n543183 , n15924 , n543185 , n543186 , n15927 , n543188 , n543189 , n15930 , n543191 , n543192 , 
     n15933 , n543194 , n543195 , n15936 , n543197 , n543198 , n15939 , n543200 , n543201 , n15942 , 
     n543203 , n543204 , n15945 , n543206 , n543207 , n15948 , n543209 , n543210 , n15951 , n543212 , 
     n543213 , n15954 , n543215 , n543216 , n15957 , n543218 , n543219 , n15960 , n543221 , n543222 , 
     n15963 , n543224 , n543225 , n15966 , n543227 , n543228 , n15969 , n543230 , n543231 , n15972 , 
     n543233 , n543234 , n15975 , n543236 , n543237 , n15978 , n543239 , n543240 , n15981 , n543242 , 
     n543243 , n15984 , n543245 , n543246 , n15987 , n543248 , n543249 , n15990 , n543251 , n543252 , 
     n15993 , n543254 , n543255 , n15996 , n543257 , n543258 , n15999 , n543260 , n543261 , n16002 , 
     n543263 , n543264 , n16005 , n543266 , n543267 , n16008 , n543269 , n543270 , n16011 , n543272 , 
     n543273 , n16014 , n543275 , n543276 , n16017 , n543278 , n543279 , n16020 , n543281 , n543282 , 
     n16023 , n543284 , n543285 , n16026 , n543287 , n543288 , n16029 , n543290 , n543291 , n16032 , 
     n543293 , n543294 , n16035 , n543296 , n543297 , n16038 , n543299 , n543300 , n16041 , n543302 , 
     n543303 , n16044 , n543305 , n543306 , n16047 , n543308 , n543309 , n16050 , n543311 , n543312 , 
     n16053 , n543314 , n543315 , n16056 , n543317 , n543318 , n16059 , n543320 , n543321 , n16062 , 
     n543323 , n543324 , n543325 , n16066 , n543327 , n16068 , n543329 , n16070 , n16071 , n543332 , 
     n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , 
     n16083 , n543344 , n16085 , n543346 , n16087 , n543348 , n16089 , n16090 , n16091 , n16092 , 
     n16093 , n16094 , n543355 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , 
     n16103 , n543364 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , 
     n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n543381 , n16122 , 
     n543383 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , 
     n16133 , n543394 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , 
     n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n543409 , n16150 , n16151 , n16152 , 
     n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , 
     n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , 
     n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n543440 , n16181 , n543442 , 
     n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , 
     n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , 
     n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , 
     n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , 
     n16223 , n16224 , n16225 , n16226 , n16227 , n543488 , n16229 , n16230 , n16231 , n16232 , 
     n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , 
     n16243 , n16244 , n16245 , n543506 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , 
     n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , 
     n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , 
     n16273 , n16274 , n16275 , n16276 , n16277 , n543538 , n16279 , n16280 , n16281 , n16282 , 
     n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , 
     n543553 , n16294 , n543555 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , 
     n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , 
     n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , 
     n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , 
     n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , 
     n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , 
     n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , 
     n16363 , n543624 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , 
     n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , 
     n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n543649 , n16390 , n543651 , n16392 , 
     n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , 
     n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , 
     n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , 
     n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , 
     n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , 
     n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , 
     n16453 , n16454 , n16455 , n543716 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , 
     n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n543731 , n16472 , 
     n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , 
     n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , 
     n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , 
     n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n543769 , n16510 , n16511 , n16512 , 
     n16513 , n16514 , n543775 , n16516 , n543777 , n16518 , n16519 , n16520 , n16521 , n16522 , 
     n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , 
     n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , 
     n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , 
     n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , 
     n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , 
     n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , 
     n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , 
     n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , 
     n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n543870 , n16611 , n16612 , 
     n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , 
     n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , 
     n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n543901 , n16642 , 
     n543903 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , 
     n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , 
     n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , 
     n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , 
     n16683 , n16684 , n16685 , n16686 , n543947 , n16688 , n16689 , n16690 , n16691 , n16692 , 
     n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , 
     n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , 
     n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , 
     n16723 , n543984 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , 
     n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , 
     n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , 
     n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , 
     n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , 
     n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , 
     n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , 
     n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , 
     n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , 
     n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n544079 , n16820 , n16821 , n16822 , 
     n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , 
     n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n544102 , 
     n16843 , n544104 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , 
     n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , 
     n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , 
     n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , 
     n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , 
     n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , 
     n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , 
     n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , 
     n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , 
     n16933 , n16934 , n544195 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , 
     n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , 
     n16953 , n16954 , n16955 , n544216 , n544217 , n16958 , n544219 , n16960 , n16961 , n16962 , 
     n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , 
     n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , 
     n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , 
     n16993 , n544254 , n16995 , n544256 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , 
     n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , 
     n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , 
     n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , 
     n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , 
     n17043 , n544304 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , 
     n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , 
     n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , 
     n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , 
     n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , 
     n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , 
     n17103 , n17104 , n17105 , n544366 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , 
     n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , 
     n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , 
     n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , 
     n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , 
     n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , 
     n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , 
     n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , 
     n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , 
     n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , 
     n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n544469 , n17210 , n544471 , n17212 , 
     n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , 
     n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , 
     n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n544499 , n17240 , n17241 , n17242 , 
     n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , 
     n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , 
     n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , 
     n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , 
     n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , 
     n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , 
     n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , 
     n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , 
     n17323 , n17324 , n17325 , n544586 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , 
     n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , 
     n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , 
     n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , 
     n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , 
     n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , 
     n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , 
     n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , 
     n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , 
     n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , 
     n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , 
     n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , 
     n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n544711 , n17452 , 
     n544713 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , 
     n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , 
     n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n544741 , n17482 , 
     n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , 
     n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , 
     n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , 
     n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , 
     n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n544789 , n17530 , n17531 , n17532 , 
     n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , 
     n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , 
     n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , 
     n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , 
     n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , 
     n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , 
     n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , 
     n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , 
     n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , 
     n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , 
     n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , 
     n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , 
     n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , 
     n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , 
     n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , 
     n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , 
     n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , 
     n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , 
     n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n544980 , n17721 , n544982 , 
     n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , 
     n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , 
     n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , 
     n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , 
     n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , 
     n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , 
     n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , 
     n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , 
     n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , 
     n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , 
     n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , 
     n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , 
     n545103 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , 
     n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , 
     n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , 
     n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , 
     n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , 
     n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , 
     n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , 
     n545173 , n17914 , n545175 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , 
     n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , 
     n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , 
     n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , 
     n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , 
     n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , 
     n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , 
     n17983 , n545244 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , 
     n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , 
     n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , 
     n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , 
     n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , 
     n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , 
     n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , 
     n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , 
     n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , 
     n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , 
     n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , 
     n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , 
     n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , 
     n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , 
     n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , 
     n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , 
     n18143 , n545404 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , 
     n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , 
     n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , 
     n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , 
     n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , 
     n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n545462 , 
     n18203 , n18204 , n18205 , n18206 , n18207 , n545468 , n18209 , n545470 , n18211 , n18212 , 
     n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , 
     n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , 
     n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , 
     n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , 
     n18253 , n545514 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , 
     n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , 
     n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , 
     n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , 
     n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , 
     n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , 
     n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , 
     n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , 
     n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , 
     n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , 
     n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , 
     n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , 
     n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , 
     n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , 
     n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , 
     n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , 
     n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , 
     n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , 
     n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , 
     n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , 
     n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , 
     n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , 
     n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , 
     n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , 
     n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , 
     n18503 , n18504 , n545765 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , 
     n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , 
     n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , 
     n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , 
     n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , 
     n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , 
     n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , 
     n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , 
     n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , 
     n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , 
     n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , 
     n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , 
     n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , 
     n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , 
     n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , 
     n545913 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , 
     n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , 
     n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , 
     n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , 
     n18693 , n545954 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , 
     n18703 , n18704 , n18705 , n18706 , n545967 , n18708 , n18709 , n18710 , n18711 , n18712 , 
     n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , 
     n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , 
     n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , 
     n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , 
     n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , 
     n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , 
     n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , 
     n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , 
     n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , 
     n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , 
     n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , 
     n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , 
     n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , 
     n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , 
     n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , 
     n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , 
     n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , 
     n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , 
     n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , 
     n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , 
     n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , 
     n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , 
     n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , 
     n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , 
     n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , 
     n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , 
     n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , 
     n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , 
     n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , 
     n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , 
     n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , 
     n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , 
     n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , 
     n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , 
     n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , 
     n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , 
     n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , 
     n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , 
     n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , 
     n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , 
     n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , 
     n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , 
     n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , 
     n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , 
     n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , 
     n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , 
     n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , 
     n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , 
     n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , 
     n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , 
     n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , 
     n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , 
     n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , 
     n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , 
     n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , 
     n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , 
     n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , 
     n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , 
     n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , 
     n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , 
     n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , 
     n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , 
     n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , 
     n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , 
     n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , 
     n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , 
     n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , 
     n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , 
     n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , 
     n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , 
     n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , 
     n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , 
     n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , 
     n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , 
     n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , 
     n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , 
     n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , 
     n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , 
     n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , 
     n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , 
     n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , 
     n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , 
     n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , 
     n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , 
     n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , 
     n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , 
     n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , 
     n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , 
     n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , 
     n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , 
     n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , 
     n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , 
     n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , 
     n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , 
     n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , 
     n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , 
     n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , 
     n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , 
     n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , 
     n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , 
     n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , 
     n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , 
     n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , 
     n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , 
     n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , 
     n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , 
     n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , 
     n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , 
     n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , 
     n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , 
     n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , 
     n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , 
     n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , 
     n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , 
     n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , 
     n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , 
     n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , 
     n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , 
     n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , 
     n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , 
     n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , 
     n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , 
     n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , 
     n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , 
     n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , 
     n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , 
     n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , 
     n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , 
     n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , 
     n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , 
     n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , 
     n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , 
     n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , 
     n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , 
     n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , 
     n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , 
     n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , 
     n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , 
     n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , 
     n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , 
     n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , 
     n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , 
     n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , 
     n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , 
     n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , 
     n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , 
     n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , 
     n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , 
     n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , 
     n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , 
     n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , 
     n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , 
     n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , 
     n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , 
     n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , 
     n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , 
     n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , 
     n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , 
     n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , 
     n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , 
     n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , 
     n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , 
     n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , 
     n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , 
     n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , 
     n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , 
     n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , 
     n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , 
     n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , 
     n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , 
     n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , 
     n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , 
     n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , 
     n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , 
     n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , 
     n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , 
     n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , 
     n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , 
     n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , 
     n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , 
     n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , 
     n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , 
     n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , 
     n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , 
     n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , 
     n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , 
     n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , 
     n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , 
     n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , 
     n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , 
     n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , 
     n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , 
     n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , 
     n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , 
     n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , 
     n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , 
     n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , 
     n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , 
     n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , 
     n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , 
     n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , 
     n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , 
     n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , 
     n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , 
     n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , 
     n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , 
     n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , 
     n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , 
     n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , 
     n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , 
     n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , 
     n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , 
     n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , 
     n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , 
     n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , 
     n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , 
     n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , 
     n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , 
     n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , 
     n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , 
     n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , 
     n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , 
     n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , 
     n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , 
     n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , 
     n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , 
     n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , 
     n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , 
     n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , 
     n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , 
     n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , 
     n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , 
     n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , 
     n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , 
     n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , 
     n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , 
     n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , 
     n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , 
     n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , 
     n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , 
     n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , 
     n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , 
     n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , 
     n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , 
     n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , 
     n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , 
     n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , 
     n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , 
     n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , 
     n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , 
     n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , 
     n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , 
     n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , 
     n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , 
     n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , 
     n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , 
     n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , 
     n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , 
     n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , 
     n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , 
     n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , 
     n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , 
     n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , 
     n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , 
     n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , 
     n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , 
     n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , 
     n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , 
     n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , 
     n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , 
     n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , 
     n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , 
     n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , 
     n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , 
     n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , 
     n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , 
     n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , 
     n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , 
     n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , 
     n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , 
     n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , 
     n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , 
     n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , 
     n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , 
     n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , 
     n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , 
     n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , 
     n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , 
     n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , 
     n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , 
     n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , 
     n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , 
     n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , 
     n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , 
     n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , 
     n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , 
     n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , 
     n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , 
     n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , 
     n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , 
     n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , 
     n21723 , n21724 , n21725 , n548986 , n548987 , n21728 , n548989 , n21730 , n548991 , n21732 , 
     n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , 
     n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , 
     n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n549020 , n549021 , n21762 , 
     n21763 , n21764 , n21765 , n21766 , n549027 , n549028 , n21769 , n549030 , n21771 , n549032 , 
     n21773 , n21774 , n549035 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n549042 , 
     n549043 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n549052 , 
     n549053 , n21794 , n549055 , n21796 , n549057 , n21798 , n21799 , n549060 , n21801 , n21802 , 
     n21803 , n21804 , n21805 , n21806 , n549067 , n549068 , n21809 , n21810 , n21811 , n21812 , 
     n21813 , n21814 , n21815 , n21816 , n21817 , n549078 , n549079 , n21820 , n549081 , n21822 , 
     n549083 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n549091 , n549092 , 
     n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , 
     n21843 , n549104 , n549105 , n21846 , n549107 , n21848 , n21849 , n549110 , n21851 , n21852 , 
     n21853 , n21854 , n21855 , n21856 , n549117 , n549118 , n21859 , n21860 , n21861 , n21862 , 
     n21863 , n21864 , n21865 , n21866 , n21867 , n549128 , n549129 , n21870 , n549131 , n21872 , 
     n549133 , n21874 , n21875 , n549136 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , 
     n549143 , n549144 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , 
     n549153 , n549154 , n21895 , n549156 , n21897 , n549158 , n21899 , n21900 , n21901 , n21902 , 
     n21903 , n21904 , n21905 , n549166 , n549167 , n21908 , n21909 , n21910 , n21911 , n21912 , 
     n21913 , n21914 , n21915 , n21916 , n549177 , n549178 , n21919 , n549180 , n21921 , n549182 , 
     n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n549190 , n549191 , n21932 , 
     n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , 
     n21943 , n21944 , n549205 , n549206 , n21947 , n549208 , n21949 , n549210 , n21951 , n21952 , 
     n549213 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n549220 , n549221 , n21962 , 
     n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n549230 , n549231 , n21972 , 
     n549233 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n549241 , n549242 , 
     n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , 
     n549253 , n549254 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , 
     n22003 , n549264 , n549265 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n549272 , 
     n549273 , n22014 , n549275 , n22016 , n549277 , n22018 , n22019 , n22020 , n22021 , n22022 , 
     n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n549291 , n549292 , 
     n22033 , n549294 , n22035 , n22036 , n22037 , n22038 , n549299 , n549300 , n22041 , n22042 , 
     n22043 , n22044 , n22045 , n22046 , n549307 , n549308 , n22049 , n22050 , n22051 , n22052 , 
     n22053 , n549314 , n549315 , n22056 , n549317 , n22058 , n22059 , n22060 , n22061 , n22062 , 
     n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , 
     n22073 , n22074 , n22075 , n22076 , n22077 , n549338 , n549339 , n22080 , n22081 , n22082 , 
     n22083 , n549344 , n549345 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n549352 , 
     n549353 , n22094 , n22095 , n22096 , n22097 , n22098 , n549359 , n549360 , n22101 , n22102 , 
     n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , 
     n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n549382 , 
     n549383 , n22124 , n22125 , n22126 , n549387 , n549388 , n22129 , n22130 , n22131 , n22132 , 
     n22133 , n22134 , n549395 , n549396 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , 
     n22143 , n22144 , n22145 , n549406 , n549407 , n22148 , n22149 , n22150 , n22151 , n22152 , 
     n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , 
     n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , 
     n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , 
     n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n549449 , n22190 , n22191 , n22192 , 
     n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , 
     n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , 
     n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , 
     n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , 
     n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n549502 , 
     n549503 , n22244 , n549505 , n22246 , n549507 , n22248 , n22249 , n22250 , n22251 , n22252 , 
     n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , 
     n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n549531 , n549532 , 
     n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , 
     n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , 
     n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n549560 , n22301 , n22302 , 
     n22303 , n22304 , n22305 , n22306 , n22307 , n549568 , n549569 , n22310 , n22311 , n22312 , 
     n22313 , n22314 , n22315 , n22316 , n22317 , n549578 , n22319 , n22320 , n22321 , n22322 , 
     n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , 
     n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , 
     n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , 
     n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , 
     n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , 
     n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , 
     n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , 
     n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , 
     n22403 , n22404 , n22405 , n22406 , n549667 , n549668 , n22409 , n22410 , n22411 , n22412 , 
     n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , 
     n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , 
     n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , 
     n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , 
     n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , 
     n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , 
     n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , 
     n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , 
     n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , 
     n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , 
     n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , 
     n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , 
     n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , 
     n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , 
     n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , 
     n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , 
     n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , 
     n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , 
     n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , 
     n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , 
     n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , 
     n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , 
     n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , 
     n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , 
     n22653 , n22654 , n22655 , n22656 , n549917 , n549918 , n22659 , n22660 , n22661 , n549922 , 
     n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , 
     n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , 
     n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , 
     n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , 
     n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , 
     n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , 
     n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , 
     n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , 
     n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , 
     n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , 
     n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , 
     n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , 
     n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , 
     n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , 
     n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , 
     n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n550081 , n550082 , 
     n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , 
     n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , 
     n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , 
     n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , 
     n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , 
     n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , 
     n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , 
     n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , 
     n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , 
     n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , 
     n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , 
     n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , 
     n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , 
     n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , 
     n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , 
     n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , 
     n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , 
     n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , 
     n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , 
     n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , 
     n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , 
     n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , 
     n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , 
     n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , 
     n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , 
     n550333 , n550334 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , 
     n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , 
     n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , 
     n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , 
     n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , 
     n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , 
     n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , 
     n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , 
     n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , 
     n23162 , n550424 , n550425 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , 
     n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , 
     n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , 
     n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , 
     n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , 
     n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , 
     n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , 
     n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , 
     n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , 
     n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n550521 , n23261 , 
     n550523 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , 
     n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , 
     n550543 , n550544 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , 
     n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , 
     n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , 
     n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , 
     n23322 , n550584 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , 
     n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , 
     n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , 
     n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , 
     n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , 
     n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , 
     n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , 
     n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , 
     n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , 
     n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , 
     n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , 
     n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , 
     n23441 , n23442 , n23443 , n550706 , n550707 , n23446 , n23447 , n23448 , n23449 , n23450 , 
     n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , 
     n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , 
     n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , 
     n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , 
     n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , 
     n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , 
     n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , 
     n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , 
     n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , 
     n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , 
     n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , 
     n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , 
     n23571 , n23572 , n550835 , n550836 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , 
     n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , 
     n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , 
     n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , 
     n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , 
     n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , 
     n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , 
     n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , 
     n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , 
     n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , 
     n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , 
     n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , 
     n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , 
     n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , 
     n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , 
     n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , 
     n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , 
     n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , 
     n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , 
     n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , 
     n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , 
     n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , 
     n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , 
     n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , 
     n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , 
     n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , 
     n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , 
     n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , 
     n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , 
     n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , 
     n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , 
     n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , 
     n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , 
     n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , 
     n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , 
     n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , 
     n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , 
     n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , 
     n23951 , n551214 , n551215 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , 
     n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , 
     n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , 
     n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , 
     n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , 
     n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n551271 , n551272 , 
     n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , 
     n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , 
     n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , 
     n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , 
     n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , 
     n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , 
     n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , 
     n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , 
     n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , 
     n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , 
     n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , 
     n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , 
     n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , 
     n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , 
     n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , 
     n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , 
     n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , 
     n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , 
     n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , 
     n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , 
     n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , 
     n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , 
     n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , 
     n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , 
     n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , 
     n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , 
     n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , 
     n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , 
     n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , 
     n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , 
     n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , 
     n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , 
     n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , 
     n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , 
     n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , 
     n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , 
     n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , 
     n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , 
     n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , 
     n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , 
     n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , 
     n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , 
     n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , 
     n24441 , n24442 , n24443 , n551706 , n551707 , n24446 , n24447 , n24448 , n24449 , n24450 , 
     n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , 
     n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , 
     n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , 
     n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , 
     n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , 
     n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , 
     n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , 
     n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , 
     n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , 
     n24541 , n551804 , n551805 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , 
     n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , 
     n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , 
     n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , 
     n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , 
     n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , 
     n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , 
     n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , 
     n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , 
     n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , 
     n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , 
     n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , 
     n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , 
     n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , 
     n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , 
     n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , 
     n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , 
     n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , 
     n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , 
     n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , 
     n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , 
     n552013 , n552014 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , 
     n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , 
     n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , 
     n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , 
     n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , 
     n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , 
     n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , 
     n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , 
     n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , 
     n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , 
     n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , 
     n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , 
     n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , 
     n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , 
     n24891 , n24892 , n24893 , n552156 , n552157 , n24896 , n24897 , n24898 , n24899 , n24900 , 
     n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , 
     n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , 
     n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , 
     n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , 
     n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , 
     n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , 
     n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , 
     n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , 
     n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , 
     n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , 
     n25001 , n552264 , n552265 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , 
     n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , 
     n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , 
     n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , 
     n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , 
     n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , 
     n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , 
     n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n552341 , n552342 , 
     n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , 
     n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , 
     n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , 
     n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , 
     n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , 
     n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , 
     n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , 
     n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , 
     n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , 
     n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , 
     n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , 
     n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , 
     n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , 
     n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , 
     n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , 
     n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , 
     n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , 
     n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , 
     n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , 
     n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , 
     n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , 
     n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , 
     n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , 
     n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , 
     n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , 
     n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n552599 , n552600 , n25337 , n25338 , 
     n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n552609 , n552610 , n25347 , n25348 , 
     n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , 
     n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , 
     n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , 
     n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , 
     n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , 
     n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , 
     n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , 
     n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n552689 , n552690 , n25427 , n25428 , 
     n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , 
     n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , 
     n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , 
     n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , 
     n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , 
     n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , 
     n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , 
     n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , 
     n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , 
     n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , 
     n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , 
     n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , 
     n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , 
     n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , 
     n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , 
     n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , 
     n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , 
     n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , 
     n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , 
     n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , 
     n25629 , n25630 , n552895 , n552896 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , 
     n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , 
     n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , 
     n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , 
     n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , 
     n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , 
     n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , 
     n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , 
     n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , 
     n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , 
     n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , 
     n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , 
     n25749 , n25750 , n553015 , n553016 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , 
     n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , 
     n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , 
     n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , 
     n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , 
     n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , 
     n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , 
     n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , 
     n25829 , n25830 , n553095 , n553096 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , 
     n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , 
     n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , 
     n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , 
     n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , 
     n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , 
     n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , 
     n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , 
     n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , 
     n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , 
     n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , 
     n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , 
     n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , 
     n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , 
     n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , 
     n25979 , n25980 , n25981 , n25982 , n25983 , n553248 , n553249 , n25986 , n25987 , n25988 , 
     n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , 
     n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , 
     n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , 
     n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , 
     n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , 
     n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , 
     n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , 
     n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , 
     n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , 
     n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , 
     n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , 
     n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n553369 , n553370 , n26107 , n26108 , 
     n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , 
     n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , 
     n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , 
     n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , 
     n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , 
     n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , 
     n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , 
     n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , 
     n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , 
     n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , 
     n26209 , n26210 , n26211 , n553476 , n553477 , n26214 , n26215 , n26216 , n26217 , n26218 , 
     n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , 
     n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , 
     n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , 
     n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , 
     n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , 
     n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , 
     n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , 
     n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , 
     n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , 
     n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , 
     n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , 
     n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , 
     n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , 
     n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n553622 , 
     n553623 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n553630 , n553631 , n26368 , 
     n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , 
     n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , 
     n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , 
     n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , 
     n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , 
     n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , 
     n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , 
     n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , 
     n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , 
     n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , 
     n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , 
     n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , 
     n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , 
     n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , 
     n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , 
     n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , 
     n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , 
     n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , 
     n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , 
     n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , 
     n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , 
     n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , 
     n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , 
     n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , 
     n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , 
     n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , 
     n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , 
     n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , 
     n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , 
     n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , 
     n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , 
     n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , 
     n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , 
     n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , 
     n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , 
     n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , 
     n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , 
     n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , 
     n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , 
     n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , 
     n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , 
     n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , 
     n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , 
     n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , 
     n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , 
     n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , 
     n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , 
     n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , 
     n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , 
     n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , 
     n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , 
     n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , 
     n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , 
     n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , 
     n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , 
     n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , 
     n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , 
     n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , 
     n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , 
     n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , 
     n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , 
     n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , 
     n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , 
     n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , 
     n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , 
     n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , 
     n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , 
     n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , 
     n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , 
     n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , 
     n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , 
     n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , 
     n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , 
     n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , 
     n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , 
     n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , 
     n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , 
     n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , 
     n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , 
     n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , 
     n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , 
     n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , 
     n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , 
     n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , 
     n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , 
     n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , 
     n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , 
     n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , 
     n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , 
     n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , 
     n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , 
     n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , 
     n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , 
     n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , 
     n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , 
     n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , 
     n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , 
     n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , 
     n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , 
     n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , 
     n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , 
     n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , 
     n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , 
     n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , 
     n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , 
     n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , 
     n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , 
     n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , 
     n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , 
     n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , 
     n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , 
     n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , 
     n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , 
     n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , 
     n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , 
     n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , 
     n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , 
     n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , 
     n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , 
     n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , 
     n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , 
     n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , 
     n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , 
     n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , 
     n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , 
     n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , 
     n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , 
     n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , 
     n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , 
     n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , 
     n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , 
     n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , 
     n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , 
     n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , 
     n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , 
     n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , 
     n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , 
     n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , 
     n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , 
     n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , 
     n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , 
     n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , 
     n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , 
     n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , 
     n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , 
     n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , 
     n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , 
     n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , 
     n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , 
     n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , 
     n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , 
     n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , 
     n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , 
     n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , 
     n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , 
     n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , 
     n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , 
     n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , 
     n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , 
     n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , 
     n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , 
     n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , 
     n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , 
     n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , 
     n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , 
     n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , 
     n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , 
     n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , 
     n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , 
     n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , 
     n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , 
     n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , 
     n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , 
     n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , 
     n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , 
     n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , 
     n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , 
     n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , 
     n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , 
     n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , 
     n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , 
     n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , 
     n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , 
     n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , 
     n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , 
     n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , 
     n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , 
     n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , 
     n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , 
     n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , 
     n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , 
     n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , 
     n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , 
     n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , 
     n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , 
     n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , 
     n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , 
     n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , 
     n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , 
     n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , 
     n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , 
     n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , 
     n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , 
     n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , 
     n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , 
     n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , 
     n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , 
     n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , 
     n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , 
     n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , 
     n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , 
     n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , 
     n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , 
     n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , 
     n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , 
     n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , 
     n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , 
     n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , 
     n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , 
     n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , 
     n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , 
     n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , 
     n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , 
     n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , 
     n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , 
     n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , 
     n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , 
     n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , 
     n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , 
     n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , 
     n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , 
     n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , 
     n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , 
     n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , 
     n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , 
     n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , 
     n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , 
     n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , 
     n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , 
     n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , 
     n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , 
     n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , 
     n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , 
     n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , 
     n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , 
     n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , 
     n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , 
     n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , 
     n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , 
     n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , 
     n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , 
     n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , 
     n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , 
     n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , 
     n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , 
     n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , 
     n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , 
     n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , 
     n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , 
     n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , 
     n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , 
     n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , 
     n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , 
     n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , 
     n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , 
     n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , 
     n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , 
     n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , 
     n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , 
     n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , 
     n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , 
     n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , 
     n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , 
     n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , 
     n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , 
     n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , 
     n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , 
     n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , 
     n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , 
     n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , 
     n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , 
     n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , 
     n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , 
     n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , 
     n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , 
     n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , 
     n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , 
     n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , 
     n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , 
     n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , 
     n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , 
     n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , 
     n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , 
     n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , 
     n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , 
     n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , 
     n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , 
     n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , 
     n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , 
     n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , 
     n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , 
     n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , 
     n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , 
     n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , 
     n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , 
     n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , 
     n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , 
     n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , 
     n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , 
     n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , 
     n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , 
     n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , 
     n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , 
     n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , 
     n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , 
     n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , 
     n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , 
     n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , 
     n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , 
     n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , 
     n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , 
     n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , 
     n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , 
     n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , 
     n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , 
     n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , 
     n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , 
     n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , 
     n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , 
     n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , 
     n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , 
     n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , 
     n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , 
     n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , 
     n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , 
     n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , 
     n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , 
     n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , 
     n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , 
     n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , 
     n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , 
     n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , 
     n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , 
     n29799 , n29800 , n29801 , n29802 , n557067 , n557068 , n29805 , n557070 , n557071 , n29808 , 
     n557073 , n557074 , n29811 , n557076 , n557077 , n29814 , n557079 , n557080 , n29817 , n557082 , 
     n557083 , n29820 , n557085 , n557086 , n29823 , n557088 , n557089 , n29826 , n557091 , n557092 , 
     n29829 , n557094 , n557095 , n29832 , n557097 , n557098 , n29835 , n557100 , n557101 , n29838 , 
     n557103 , n557104 , n29841 , n557106 , n557107 , n29844 , n557109 , n557110 , n29847 , n557112 , 
     n557113 , n29850 , n557115 , n557116 , n29853 , n557118 , n557119 , n29856 , n557121 , n557122 , 
     n29859 , n557124 , n557125 , n29862 , n557127 , n557128 , n29865 , n557130 , n557131 , n29868 , 
     n557133 , n557134 , n29871 , n557136 , n557137 , n29874 , n557139 , n557140 , n29877 , n557142 , 
     n557143 , n29880 , n557145 , n557146 , n29883 , n557148 , n557149 , n29886 , n557151 , n557152 , 
     n29889 , n557154 , n557155 , n29892 , n557157 , n557158 , n29895 , n557160 , n557161 , n29898 , 
     n557163 , n557164 , n29901 , n557166 , n557167 , n29904 , n557169 , n557170 , n29907 , n557172 , 
     n557173 , n29910 , n557175 , n557176 , n29913 , n557178 , n557179 , n29916 , n557181 , n557182 , 
     n29919 , n557184 , n557185 , n29922 , n557187 , n557188 , n29925 , n557190 , n557191 , n29928 , 
     n557193 , n557194 , n29931 , n557196 , n557197 , n29934 , n557199 , n557200 , n29937 , n557202 , 
     n557203 , n29940 , n557205 , n557206 , n29943 , n557208 , n557209 , n29946 , n557211 , n557212 , 
     n29949 , n557214 , n557215 , n29952 , n557217 , n557218 , n29955 , n557220 , n557221 , n29958 , 
     n557223 , n557224 , n29961 , n557226 , n557227 , n29964 , n557229 , n557230 , n29967 , n557232 , 
     n557233 , n29970 , n557235 , n557236 , n29973 , n557238 , n557239 , n29976 , n557241 , n557242 , 
     n29979 , n557244 , n557245 , n29982 , n557247 , n557248 , n29985 , n557250 , n557251 , n29988 , 
     n557253 , n557254 , n29991 , n557256 , n557257 , n29994 , n29995 , n29996 , n29997 , n29998 , 
     n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , 
     n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , 
     n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , 
     n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , 
     n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , 
     n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , 
     n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , 
     n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , 
     n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , 
     n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , 
     n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , 
     n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , 
     n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , 
     n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , 
     n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , 
     n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , 
     n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , 
     n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , 
     n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , 
     n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , 
     n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , 
     n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , 
     n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , 
     n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , 
     n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , 
     n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , 
     n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , 
     n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , 
     n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , 
     n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , 
     n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , 
     n30309 , n30310 , n30311 , n557576 , n30313 , n30314 , n557579 , n30316 , n30317 , n557582 , 
     n30319 , n30320 , n557585 , n30322 , n30323 , n557588 , n30325 , n30326 , n557591 , n30328 , 
     n30329 , n557594 , n30331 , n30332 , n557597 , n30334 , n30335 , n557600 , n30337 , n30338 , 
     n557603 , n30340 , n30341 , n557606 , n30343 , n30344 , n557609 , n30346 , n30347 , n557612 , 
     n30349 , n30350 , n557615 , n30352 , n30353 , n557618 , n30355 , n30356 , n557621 , n30358 , 
     n30359 , n557624 , n30361 , n30362 , n557627 , n30364 , n30365 , n557630 , n30367 , n30368 , 
     n557633 , n30370 , n30371 , n557636 , n30373 , n30374 , n557639 , n30376 , n30377 , n557642 , 
     n30379 , n30380 , n557645 , n30382 , n30383 , n557648 , n30385 , n30386 , n557651 , n30388 , 
     n30389 , n557654 , n30391 , n30392 , n557657 , n30394 , n30395 , n557660 , n30397 , n30398 , 
     n557663 , n30400 , n30401 , n557666 , n30403 , n30404 , n557669 , n30406 , n30407 , n557672 , 
     n30409 , n30410 , n557675 , n30412 , n30413 , n557678 , n30415 , n30416 , n557681 , n30418 , 
     n30419 , n557684 , n30421 , n30422 , n557687 , n30424 , n30425 , n557690 , n30427 , n30428 , 
     n557693 , n30430 , n30431 , n557696 , n30433 , n30434 , n557699 , n30436 , n30437 , n557702 , 
     n30439 , n30440 , n557705 , n30442 , n30443 , n557708 , n30445 , n30446 , n557711 , n30448 , 
     n30449 , n557714 , n30451 , n30452 , n557717 , n30454 , n30455 , n557720 , n30457 , n30458 , 
     n557723 , n30460 , n30461 , n557726 , n30463 , n30464 , n557729 , n30466 , n30467 , n557732 , 
     n30469 , n30470 , n557735 , n30472 , n30473 , n557738 , n30475 , n30476 , n557741 , n30478 , 
     n30479 , n557744 , n30481 , n30482 , n557747 , n30484 , n30485 , n557750 , n30487 , n30488 , 
     n557753 , n30490 , n30491 , n557756 , n30493 , n30494 , n557759 , n30496 , n30497 , n557762 , 
     n30499 , n30500 , n557765 , n30502 , n557767 , n557768 , n557769 , n557770 , n557771 , n557772 , 
     n557773 , n557774 , n557775 , n557776 , n557777 , n557778 , n557779 , n557780 , n557781 , n557782 , 
     n557783 , n557784 , n557785 , n557786 , n557787 , n557788 , n557789 , n557790 , n557791 , n557792 , 
     n557793 , n557794 , n557795 , n557796 , n557797 , n557798 , n557799 , n557800 , n557801 , n557802 , 
     n557803 , n557804 , n557805 , n557806 , n557807 , n557808 , n557809 , n557810 , n557811 , n557812 , 
     n557813 , n557814 , n557815 , n557816 , n557817 , n557818 , n557819 , n557820 , n557821 , n557822 , 
     n557823 , n557824 , n557825 , n557826 , n557827 , n557828 , n557829 , n557830 , n557831 , n557832 , 
     n557833 , n30570 , n557835 , n30572 , n30573 , n557838 , n30575 , n30576 , n557841 , n30578 , 
     n557843 , n30580 , n30581 , n557846 , n30583 , n30584 , n30585 , n557850 , n30587 , n30588 , 
     n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n557861 , n30598 , 
     n30599 , n557864 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n557872 , 
     n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , 
     n557883 , n30620 , n30621 , n557886 , n30623 , n30624 , n30625 , n557890 , n30627 , n30628 , 
     n30629 , n30630 , n557895 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , 
     n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , 
     n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n557921 , n30658 , 
     n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , 
     n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , 
     n557943 , n30680 , n30681 , n30682 , n30683 , n557948 , n30685 , n30686 , n30687 , n30688 , 
     n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , 
     n30699 , n30700 , n557965 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , 
     n30709 , n557974 , n30711 , n30712 , n30713 , n30714 , n557979 , n30716 , n30717 , n30718 , 
     n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , 
     n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , 
     n30739 , n30740 , n30741 , n30742 , n30743 , n558008 , n30745 , n30746 , n558011 , n30748 , 
     n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n558022 , 
     n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , 
     n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , 
     n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , 
     n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , 
     n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , 
     n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , 
     n30819 , n30820 , n30821 , n30822 , n558087 , n30824 , n30825 , n30826 , n30827 , n30828 , 
     n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , 
     n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , 
     n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , 
     n558123 , n30860 , n30861 , n558126 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , 
     n30869 , n30870 , n558135 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , 
     n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , 
     n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , 
     n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , 
     n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , 
     n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n558189 , n30926 , n30927 , n30928 , 
     n30929 , n30930 , n558195 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , 
     n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n558210 , n30947 , n30948 , 
     n558213 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n558221 , n30958 , 
     n30959 , n30960 , n558225 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , 
     n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , 
     n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , 
     n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , 
     n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , 
     n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , 
     n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , 
     n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , 
     n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , 
     n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n558320 , n31057 , n31058 , 
     n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n558329 , n31066 , n31067 , n31068 , 
     n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , 
     n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , 
     n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , 
     n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , 
     n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , 
     n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , 
     n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n558402 , 
     n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , 
     n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , 
     n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n558431 , n31168 , 
     n31169 , n558434 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , 
     n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , 
     n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , 
     n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , 
     n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , 
     n31219 , n31220 , n31221 , n31222 , n558487 , n31224 , n31225 , n31226 , n31227 , n31228 , 
     n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , 
     n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , 
     n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , 
     n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n558532 , 
     n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n558541 , n31278 , 
     n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , 
     n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , 
     n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , 
     n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n558579 , n31316 , n31317 , n31318 , 
     n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , 
     n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , 
     n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , 
     n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , 
     n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , 
     n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , 
     n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , 
     n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , 
     n31399 , n31400 , n31401 , n31402 , n31403 , n558668 , n31405 , n31406 , n31407 , n31408 , 
     n31409 , n31410 , n31411 , n31412 , n558677 , n31414 , n31415 , n31416 , n31417 , n31418 , 
     n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , 
     n558693 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , 
     n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , 
     n31449 , n31450 , n31451 , n558716 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , 
     n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , 
     n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , 
     n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , 
     n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , 
     n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , 
     n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n558780 , n31517 , n31518 , 
     n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , 
     n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , 
     n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n558809 , n31546 , n31547 , n31548 , 
     n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , 
     n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , 
     n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , 
     n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , 
     n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n558860 , n31597 , n31598 , 
     n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , 
     n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n558882 , 
     n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , 
     n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , 
     n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , 
     n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , 
     n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , 
     n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , 
     n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , 
     n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , 
     n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , 
     n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , 
     n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , 
     n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , 
     n31739 , n559004 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , 
     n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , 
     n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n559029 , n31766 , n31767 , n31768 , 
     n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , 
     n31779 , n31780 , n31781 , n559046 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , 
     n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , 
     n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , 
     n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , 
     n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , 
     n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , 
     n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , 
     n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , 
     n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , 
     n31869 , n559134 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , 
     n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n559151 , n31888 , 
     n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , 
     n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , 
     n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , 
     n31919 , n31920 , n31921 , n559186 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , 
     n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , 
     n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , 
     n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , 
     n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , 
     n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , 
     n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , 
     n31989 , n31990 , n31991 , n31992 , n559257 , n31993 , n31994 , n31995 , n559261 , n31997 , 
     n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , 
     n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , 
     n559283 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , 
     n32028 , n32029 , n559295 , n559296 , n559297 , n559298 , n559299 , n559300 , n32030 , n32031 , 
     n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n559311 , n559312 , 
     n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , 
     n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , 
     n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , 
     n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , 
     n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , 
     n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , 
     n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , 
     n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , 
     n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , 
     n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , 
     n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , 
     n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , 
     n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , 
     n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , 
     n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , 
     n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , 
     n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , 
     n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , 
     n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n559499 , n32227 , n32228 , n32229 , 
     n32230 , n32231 , n32232 , n32233 , n559507 , n32235 , n32236 , n32237 , n32238 , n32239 , 
     n32240 , n32241 , n32242 , n559516 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , 
     n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , 
     n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , 
     n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , 
     n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , 
     n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n559569 , n32296 , n32297 , n32298 , 
     n32299 , n32300 , n559575 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , 
     n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , 
     n559593 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , 
     n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , 
     n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , 
     n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , 
     n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , 
     n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , 
     n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , 
     n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , 
     n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , 
     n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , 
     n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , 
     n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , 
     n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , 
     n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , 
     n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , 
     n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , 
     n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n559761 , n32488 , 
     n32489 , n32490 , n32491 , n32492 , n559767 , n32494 , n32495 , n32496 , n32497 , n32498 , 
     n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n559781 , n32508 , 
     n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , 
     n32519 , n32520 , n32521 , n32522 , n32523 , n559798 , n32525 , n32526 , n32527 , n32528 , 
     n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , 
     n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , 
     n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , 
     n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , 
     n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , 
     n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , 
     n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , 
     n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , 
     n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , 
     n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , 
     n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , 
     n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , 
     n32649 , n32650 , n32651 , n32652 , n32653 , n559928 , n32655 , n32656 , n32657 , n32658 , 
     n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , 
     n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , 
     n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , 
     n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , 
     n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , 
     n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , 
     n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , 
     n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , 
     n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , 
     n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , 
     n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , 
     n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , 
     n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , 
     n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , 
     n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , 
     n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , 
     n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , 
     n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , 
     n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , 
     n560123 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , 
     n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n560141 , n32868 , 
     n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , 
     n32879 , n32880 , n560155 , n32882 , n32883 , n32884 , n32885 , n32886 , n560161 , n32888 , 
     n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , 
     n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , 
     n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , 
     n32919 , n32920 , n560195 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , 
     n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , 
     n560213 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , 
     n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , 
     n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , 
     n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , 
     n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , 
     n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , 
     n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , 
     n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , 
     n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , 
     n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , 
     n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , 
     n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , 
     n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , 
     n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , 
     n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , 
     n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , 
     n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , 
     n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , 
     n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , 
     n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , 
     n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , 
     n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , 
     n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , 
     n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , 
     n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , 
     n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , 
     n33199 , n33200 , n33201 , n33202 , n560477 , n33204 , n33205 , n33206 , n33207 , n33208 , 
     n33209 , n33210 , n33211 , n560486 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , 
     n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , 
     n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , 
     n560513 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , 
     n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , 
     n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , 
     n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , 
     n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , 
     n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , 
     n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , 
     n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , 
     n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , 
     n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , 
     n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , 
     n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , 
     n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , 
     n33369 , n33370 , n33371 , n33372 , n560647 , n33374 , n33375 , n33376 , n33377 , n33378 , 
     n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , 
     n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , 
     n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , 
     n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , 
     n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , 
     n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , 
     n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , 
     n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , 
     n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , 
     n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , 
     n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , 
     n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , 
     n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , 
     n33509 , n33510 , n33511 , n560786 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , 
     n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , 
     n33529 , n33530 , n560805 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , 
     n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , 
     n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n560829 , n33556 , n33557 , n33558 , 
     n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , 
     n33569 , n33570 , n33571 , n33572 , n33573 , n560848 , n33575 , n33576 , n33577 , n33578 , 
     n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , 
     n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , 
     n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , 
     n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , 
     n33619 , n33620 , n33621 , n33622 , n560897 , n33624 , n33625 , n33626 , n33627 , n33628 , 
     n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , 
     n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , 
     n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , 
     n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , 
     n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , 
     n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , 
     n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , 
     n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , 
     n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , 
     n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , 
     n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , 
     n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , 
     n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , 
     n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , 
     n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , 
     n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , 
     n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , 
     n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , 
     n33809 , n33810 , n33811 , n33812 , n33813 , n561088 , n33815 , n33816 , n33817 , n33818 , 
     n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , 
     n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , 
     n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , 
     n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , 
     n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , 
     n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , 
     n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , 
     n33889 , n33890 , n33891 , n33892 , n561167 , n33894 , n33895 , n33896 , n33897 , n33898 , 
     n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , 
     n33909 , n33910 , n33911 , n33912 , n561187 , n33914 , n33915 , n33916 , n33917 , n33918 , 
     n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , 
     n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , 
     n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , 
     n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , 
     n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , 
     n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , 
     n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , 
     n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , 
     n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , 
     n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , 
     n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , 
     n34029 , n34030 , n561305 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , 
     n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n561322 , 
     n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , 
     n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , 
     n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , 
     n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , 
     n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , 
     n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , 
     n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , 
     n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , 
     n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , 
     n34139 , n34140 , n34141 , n561416 , n34143 , n34144 , n34145 , n34146 , n34147 , n561422 , 
     n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , 
     n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , 
     n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , 
     n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , 
     n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , 
     n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , 
     n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , 
     n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , 
     n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , 
     n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , 
     n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , 
     n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , 
     n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , 
     n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , 
     n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n561571 , n34298 , 
     n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , 
     n34309 , n34310 , n34311 , n34312 , n34313 , n561588 , n34315 , n34316 , n34317 , n34318 , 
     n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , 
     n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , 
     n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , 
     n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , 
     n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , 
     n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , 
     n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , 
     n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , 
     n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , 
     n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , 
     n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , 
     n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , 
     n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , 
     n34449 , n34450 , n34451 , n561726 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , 
     n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , 
     n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , 
     n561753 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , 
     n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , 
     n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , 
     n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , 
     n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , 
     n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , 
     n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , 
     n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , 
     n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , 
     n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , 
     n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , 
     n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , 
     n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , 
     n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , 
     n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , 
     n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , 
     n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , 
     n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , 
     n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , 
     n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , 
     n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , 
     n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , 
     n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , 
     n34709 , n34710 , n561985 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , 
     n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , 
     n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , 
     n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , 
     n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , 
     n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , 
     n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , 
     n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , 
     n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , 
     n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , 
     n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , 
     n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , 
     n34829 , n34830 , n34831 , n562106 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , 
     n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , 
     n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , 
     n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , 
     n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , 
     n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , 
     n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , 
     n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , 
     n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , 
     n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , 
     n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , 
     n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , 
     n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , 
     n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , 
     n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , 
     n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , 
     n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , 
     n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , 
     n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , 
     n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , 
     n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , 
     n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , 
     n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , 
     n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , 
     n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , 
     n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , 
     n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , 
     n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , 
     n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , 
     n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , 
     n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , 
     n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , 
     n35149 , n35150 , n562425 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , 
     n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , 
     n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , 
     n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , 
     n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , 
     n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , 
     n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , 
     n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , 
     n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , 
     n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , 
     n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , 
     n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , 
     n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , 
     n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , 
     n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , 
     n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , 
     n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , 
     n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , 
     n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , 
     n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , 
     n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , 
     n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , 
     n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , 
     n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , 
     n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , 
     n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , 
     n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , 
     n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , 
     n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , 
     n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , 
     n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , 
     n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , 
     n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , 
     n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , 
     n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , 
     n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , 
     n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , 
     n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , 
     n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , 
     n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , 
     n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n562832 , 
     n35559 , n35560 , n562835 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , 
     n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , 
     n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , 
     n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , 
     n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , 
     n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , 
     n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , 
     n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , 
     n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , 
     n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , 
     n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , 
     n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , 
     n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , 
     n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , 
     n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , 
     n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , 
     n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , 
     n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , 
     n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , 
     n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , 
     n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , 
     n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , 
     n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , 
     n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , 
     n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , 
     n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , 
     n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n563099 , n35825 , n35826 , n35827 , 
     n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , 
     n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , 
     n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , 
     n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , 
     n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , 
     n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , 
     n563163 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , 
     n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , 
     n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , 
     n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , 
     n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , 
     n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , 
     n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , 
     n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , 
     n35968 , n35969 , n35970 , n563246 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , 
     n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , 
     n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , 
     n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , 
     n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , 
     n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , 
     n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , 
     n36037 , n36038 , n563315 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , 
     n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n563329 , n36053 , n36054 , n36055 , 
     n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , 
     n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , 
     n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , 
     n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , 
     n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , 
     n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , 
     n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , 
     n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , 
     n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , 
     n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , 
     n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , 
     n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , 
     n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , 
     n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n563472 , 
     n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , 
     n563483 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , 
     n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , 
     n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , 
     n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , 
     n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , 
     n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , 
     n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , 
     n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , 
     n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , 
     n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , 
     n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , 
     n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , 
     n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , 
     n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , 
     n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , 
     n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , 
     n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , 
     n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , 
     n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , 
     n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , 
     n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , 
     n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , 
     n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , 
     n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , 
     n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , 
     n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , 
     n36465 , n36466 , n36467 , n36468 , n563747 , n36469 , n563749 , n563750 , n36470 , n36471 , 
     n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , 
     n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , 
     n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , 
     n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , 
     n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , 
     n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , 
     n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , 
     n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , 
     n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , 
     n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , 
     n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , 
     n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n563870 , n36589 , n36590 , 
     n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , 
     n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , 
     n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , 
     n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , 
     n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , 
     n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , 
     n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , 
     n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , 
     n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , 
     n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , 
     n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , 
     n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , 
     n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , 
     n36721 , n36722 , n36723 , n36724 , n36725 , n564008 , n36727 , n36728 , n36729 , n36730 , 
     n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , 
     n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , 
     n36751 , n36752 , n564035 , n36754 , n36755 , n36756 , n564039 , n36758 , n36759 , n36760 , 
     n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , 
     n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , 
     n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , 
     n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , 
     n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , 
     n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , 
     n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , 
     n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , 
     n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , 
     n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , 
     n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , 
     n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , 
     n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , 
     n36891 , n36892 , n36893 , n36894 , n36895 , n564178 , n36896 , n564180 , n36897 , n36898 , 
     n36899 , n36900 , n36901 , n564186 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , 
     n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , 
     n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , 
     n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , 
     n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , 
     n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , 
     n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , 
     n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , 
     n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , 
     n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , 
     n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , 
     n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , 
     n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , 
     n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , 
     n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , 
     n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , 
     n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , 
     n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , 
     n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , 
     n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , 
     n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , 
     n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , 
     n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , 
     n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , 
     n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , 
     n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , 
     n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , 
     n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , 
     n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , 
     n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , 
     n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , 
     n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , 
     n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , 
     n37228 , n37229 , n37230 , n564516 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , 
     n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , 
     n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , 
     n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , 
     n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , 
     n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , 
     n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , 
     n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , 
     n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , 
     n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , 
     n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , 
     n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , 
     n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , 
     n564643 , n564644 , n564645 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , 
     n37365 , n37366 , n37367 , n564656 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , 
     n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , 
     n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n564679 , n37392 , n37393 , n37394 , 
     n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , 
     n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , 
     n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , 
     n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , 
     n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , 
     n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , 
     n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , 
     n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , 
     n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , 
     n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , 
     n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , 
     n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , 
     n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , 
     n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , 
     n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , 
     n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , 
     n37555 , n37556 , n564845 , n564846 , n564847 , n37557 , n37558 , n37559 , n37560 , n37561 , 
     n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , 
     n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , 
     n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , 
     n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , 
     n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , 
     n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n564910 , n564911 , n564912 , 
     n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n564921 , n37628 , 
     n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , 
     n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , 
     n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , 
     n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , 
     n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , 
     n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , 
     n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , 
     n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , 
     n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , 
     n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , 
     n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , 
     n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n565042 , 
     n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , 
     n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , 
     n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , 
     n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , 
     n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , 
     n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , 
     n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , 
     n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , 
     n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , 
     n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , 
     n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , 
     n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , 
     n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n565170 , n37877 , n37878 , 
     n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , 
     n37889 , n37890 , n37891 , n37892 , n37893 , n565188 , n565189 , n565190 , n37894 , n37895 , 
     n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , 
     n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , 
     n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , 
     n37926 , n37927 , n37928 , n37929 , n565227 , n565228 , n565229 , n37930 , n37931 , n37932 , 
     n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , 
     n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , 
     n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , 
     n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , 
     n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , 
     n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , 
     n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , 
     n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , 
     n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , 
     n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n565330 , n38031 , n38032 , 
     n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , 
     n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , 
     n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , 
     n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , 
     n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , 
     n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , 
     n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , 
     n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n565412 , 
     n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , 
     n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , 
     n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , 
     n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , 
     n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , 
     n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , 
     n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , 
     n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , 
     n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , 
     n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , 
     n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , 
     n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , 
     n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , 
     n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , 
     n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , 
     n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , 
     n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , 
     n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , 
     n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , 
     n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , 
     n38312 , n38313 , n38314 , n38315 , n38316 , n565618 , n38318 , n38319 , n38320 , n38321 , 
     n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , 
     n38332 , n565634 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , 
     n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , 
     n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , 
     n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , 
     n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , 
     n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , 
     n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , 
     n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , 
     n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , 
     n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , 
     n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , 
     n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n565749 , n38449 , n38450 , n38451 , 
     n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , 
     n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , 
     n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , 
     n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , 
     n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , 
     n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , 
     n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , 
     n38522 , n38523 , n38524 , n38525 , n38526 , n565828 , n38528 , n38529 , n38530 , n38531 , 
     n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , 
     n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , 
     n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , 
     n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , 
     n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , 
     n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , 
     n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , 
     n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , 
     n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , 
     n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , 
     n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , 
     n38642 , n38643 , n38644 , n565946 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , 
     n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , 
     n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , 
     n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , 
     n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , 
     n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , 
     n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , 
     n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , 
     n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , 
     n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , 
     n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , 
     n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , 
     n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n566071 , n38771 , 
     n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , 
     n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , 
     n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , 
     n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , 
     n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , 
     n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , 
     n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n566142 , 
     n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , 
     n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , 
     n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , 
     n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , 
     n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n566189 , n38889 , n38890 , n38891 , 
     n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , 
     n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , 
     n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , 
     n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , 
     n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , 
     n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , 
     n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , 
     n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , 
     n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , 
     n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , 
     n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , 
     n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , 
     n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n566320 , n39020 , n39021 , 
     n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , 
     n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , 
     n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , 
     n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , 
     n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , 
     n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n566379 , n39079 , n39080 , n39081 , 
     n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , 
     n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , 
     n39102 , n39103 , n39104 , n566406 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , 
     n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , 
     n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , 
     n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , 
     n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , 
     n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , 
     n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , 
     n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , 
     n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , 
     n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n566500 , n39200 , n39201 , 
     n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , 
     n39212 , n566514 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , 
     n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , 
     n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , 
     n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , 
     n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , 
     n39262 , n566564 , n39264 , n39265 , n39266 , n39267 , n39268 , n566570 , n39270 , n39271 , 
     n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , 
     n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , 
     n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , 
     n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , 
     n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , 
     n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , 
     n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , 
     n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , 
     n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , 
     n39362 , n566664 , n566665 , n39365 , n566667 , n39367 , n566669 , n39369 , n39370 , n566672 , 
     n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , 
     n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n566690 , n39390 , n39391 , 
     n566693 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , 
     n39402 , n39403 , n39404 , n39405 , n39406 , n566708 , n566709 , n39409 , n39410 , n39411 , 
     n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , 
     n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n566731 , n566732 , 
     n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n566740 , n566741 , n39441 , 
     n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , 
     n39452 , n39453 , n39454 , n39455 , n566757 , n39457 , n566759 , n39459 , n39460 , n39461 , 
     n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n566771 , n566772 , 
     n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , 
     n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n566792 , 
     n566793 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , 
     n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , 
     n39512 , n39513 , n39514 , n39515 , n566817 , n39517 , n566819 , n39519 , n39520 , n39521 , 
     n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , 
     n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , 
     n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n566851 , n566852 , 
     n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , 
     n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , 
     n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , 
     n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , 
     n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , 
     n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , 
     n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n566919 , n566920 , n39620 , n39621 , 
     n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , 
     n39632 , n39633 , n39634 , n39635 , n39636 , n566938 , n39638 , n566940 , n39640 , n39641 , 
     n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n566952 , 
     n566953 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , 
     n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n566969 , n566970 , n39670 , n39671 , 
     n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , 
     n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , 
     n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , 
     n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , 
     n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , 
     n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , 
     n39732 , n39733 , n39734 , n39735 , n567037 , n39737 , n567039 , n39739 , n39740 , n39741 , 
     n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n567051 , n567052 , 
     n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , 
     n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , 
     n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , 
     n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , 
     n39792 , n567094 , n567095 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , 
     n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , 
     n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , 
     n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , 
     n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , 
     n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n567152 , 
     n39852 , n567154 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , 
     n39862 , n39863 , n39864 , n567166 , n567167 , n39867 , n39868 , n39869 , n39870 , n39871 , 
     n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , 
     n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , 
     n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , 
     n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , 
     n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , 
     n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , 
     n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , 
     n39942 , n39943 , n39944 , n39945 , n567247 , n567248 , n39948 , n39949 , n39950 , n39951 , 
     n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , 
     n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , 
     n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , 
     n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , 
     n39992 , n567294 , n39994 , n567296 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , 
     n40002 , n40003 , n40004 , n40005 , n40006 , n567308 , n567309 , n40009 , n40010 , n40011 , 
     n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , 
     n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , 
     n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , 
     n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , 
     n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , 
     n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , 
     n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , 
     n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , 
     n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , 
     n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , 
     n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , 
     n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , 
     n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , 
     n40142 , n40143 , n40144 , n40145 , n567447 , n567448 , n40148 , n40149 , n40150 , n40151 , 
     n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , 
     n40162 , n567464 , n40164 , n567466 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , 
     n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , 
     n40182 , n40183 , n567485 , n567486 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , 
     n40192 , n40193 , n40194 , n567496 , n567497 , n40197 , n40198 , n40199 , n40200 , n40201 , 
     n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , 
     n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , 
     n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , 
     n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , 
     n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , 
     n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , 
     n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , 
     n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , 
     n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , 
     n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , 
     n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , 
     n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , 
     n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , 
     n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , 
     n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , 
     n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , 
     n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n567672 , 
     n567673 , n40373 , n40374 , n40375 , n567677 , n40377 , n567679 , n40379 , n40380 , n40381 , 
     n40382 , n40383 , n40384 , n40385 , n567687 , n567688 , n40388 , n40389 , n40390 , n40391 , 
     n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , 
     n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , 
     n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , 
     n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , 
     n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , 
     n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , 
     n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , 
     n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , 
     n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , 
     n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n567791 , n567792 , 
     n40492 , n40493 , n40494 , n567796 , n40496 , n567798 , n40498 , n40499 , n40500 , n40501 , 
     n40502 , n40503 , n40504 , n567806 , n567807 , n40507 , n40508 , n40509 , n40510 , n40511 , 
     n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , 
     n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , 
     n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , 
     n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , 
     n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , 
     n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , 
     n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , 
     n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , 
     n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , 
     n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , 
     n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , 
     n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , 
     n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , 
     n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , 
     n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , 
     n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , 
     n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , 
     n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , 
     n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , 
     n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , 
     n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , 
     n568023 , n40723 , n568025 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , 
     n40732 , n40733 , n40734 , n40735 , n568037 , n568038 , n40738 , n40739 , n40740 , n40741 , 
     n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , 
     n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , 
     n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , 
     n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , 
     n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , 
     n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , 
     n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , 
     n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , 
     n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , 
     n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , 
     n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , 
     n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , 
     n40862 , n40863 , n40864 , n40865 , n40866 , n568168 , n568169 , n40869 , n40870 , n40871 , 
     n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , 
     n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , 
     n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , 
     n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , 
     n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , 
     n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , 
     n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , 
     n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , 
     n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , 
     n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , 
     n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , 
     n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , 
     n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , 
     n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , 
     n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , 
     n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n568331 , n568332 , 
     n41032 , n41033 , n41034 , n568336 , n41036 , n568338 , n41038 , n41039 , n41040 , n41041 , 
     n41042 , n41043 , n41044 , n568346 , n568347 , n41047 , n41048 , n41049 , n41050 , n41051 , 
     n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , 
     n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , 
     n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , 
     n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , 
     n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , 
     n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , 
     n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , 
     n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , 
     n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , 
     n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , 
     n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , 
     n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , 
     n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n568481 , n568482 , 
     n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n568489 , n41189 , n568491 , n41191 , 
     n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , 
     n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , 
     n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , 
     n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , 
     n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , 
     n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , 
     n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , 
     n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , 
     n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , 
     n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , 
     n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , 
     n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , 
     n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , 
     n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , 
     n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , 
     n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , 
     n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , 
     n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , 
     n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , 
     n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , 
     n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , 
     n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , 
     n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , 
     n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , 
     n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , 
     n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , 
     n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , 
     n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , 
     n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , 
     n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , 
     n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , 
     n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , 
     n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , 
     n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , 
     n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , 
     n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , 
     n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , 
     n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , 
     n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , 
     n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , 
     n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , 
     n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , 
     n41612 , n568914 , n568915 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , 
     n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , 
     n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , 
     n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , 
     n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , 
     n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , 
     n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n568982 , 
     n41682 , n568984 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n568991 , n568992 , 
     n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , 
     n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , 
     n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , 
     n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , 
     n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , 
     n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , 
     n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , 
     n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , 
     n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , 
     n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , 
     n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , 
     n41802 , n41803 , n41804 , n569106 , n569107 , n41807 , n41808 , n41809 , n41810 , n41811 , 
     n41812 , n41813 , n569115 , n569116 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , 
     n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , 
     n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , 
     n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , 
     n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , 
     n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , 
     n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , 
     n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , 
     n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , 
     n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , 
     n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , 
     n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , 
     n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , 
     n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , 
     n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , 
     n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , 
     n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , 
     n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , 
     n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , 
     n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , 
     n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , 
     n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , 
     n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , 
     n42042 , n42043 , n42044 , n42045 , n569347 , n569348 , n42048 , n42049 , n42050 , n42051 , 
     n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n569360 , n569361 , n42061 , 
     n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , 
     n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , 
     n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , 
     n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , 
     n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , 
     n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , 
     n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , 
     n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , 
     n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , 
     n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , 
     n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , 
     n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , 
     n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , 
     n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , 
     n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , 
     n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , 
     n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , 
     n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , 
     n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , 
     n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , 
     n42262 , n42263 , n42264 , n569566 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , 
     n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , 
     n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , 
     n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , 
     n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , 
     n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , 
     n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , 
     n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , 
     n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , 
     n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , 
     n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , 
     n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , 
     n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , 
     n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , 
     n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , 
     n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , 
     n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , 
     n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , 
     n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , 
     n42452 , n42453 , n569755 , n569756 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , 
     n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , 
     n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , 
     n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , 
     n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , 
     n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , 
     n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , 
     n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , 
     n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , 
     n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , 
     n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , 
     n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , 
     n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , 
     n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , 
     n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , 
     n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , 
     n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , 
     n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , 
     n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , 
     n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , 
     n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , 
     n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , 
     n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , 
     n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , 
     n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , 
     n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , 
     n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , 
     n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , 
     n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , 
     n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , 
     n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , 
     n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , 
     n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , 
     n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , 
     n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , 
     n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n570110 , n570111 , n42811 , 
     n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , 
     n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , 
     n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , 
     n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , 
     n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , 
     n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , 
     n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , 
     n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , 
     n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , 
     n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , 
     n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , 
     n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , 
     n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , 
     n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , 
     n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , 
     n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , 
     n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , 
     n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , 
     n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , 
     n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , 
     n43012 , n43013 , n43014 , n43015 , n43016 , n570318 , n570319 , n43019 , n43020 , n43021 , 
     n43022 , n43023 , n43024 , n570326 , n570327 , n43027 , n43028 , n43029 , n43030 , n43031 , 
     n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , 
     n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , 
     n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , 
     n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n570372 , 
     n570373 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , 
     n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , 
     n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , 
     n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , 
     n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , 
     n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , 
     n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , 
     n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , 
     n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , 
     n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , 
     n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , 
     n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n570491 , n570492 , 
     n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n570499 , n570500 , n43200 , n43201 , 
     n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , 
     n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , 
     n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , 
     n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , 
     n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , 
     n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , 
     n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , 
     n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , 
     n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , 
     n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , 
     n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , 
     n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , 
     n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , 
     n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , 
     n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , 
     n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , 
     n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , 
     n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , 
     n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , 
     n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , 
     n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , 
     n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , 
     n43422 , n43423 , n43424 , n43425 , n570727 , n570728 , n43428 , n43429 , n43430 , n570732 , 
     n43431 , n43432 , n43433 , n43434 , n570737 , n570738 , n43437 , n43438 , n43439 , n43440 , 
     n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , 
     n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , 
     n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , 
     n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , 
     n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , 
     n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , 
     n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , 
     n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , 
     n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , 
     n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , 
     n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , 
     n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , 
     n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , 
     n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , 
     n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , 
     n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , 
     n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , 
     n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , 
     n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , 
     n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , 
     n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , 
     n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , 
     n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , 
     n570973 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , 
     n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , 
     n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , 
     n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , 
     n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , 
     n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , 
     n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , 
     n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , 
     n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , 
     n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , 
     n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , 
     n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , 
     n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , 
     n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , 
     n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , 
     n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , 
     n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , 
     n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , 
     n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , 
     n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , 
     n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , 
     n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , 
     n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , 
     n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , 
     n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , 
     n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , 
     n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , 
     n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , 
     n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , 
     n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , 
     n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , 
     n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , 
     n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , 
     n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , 
     n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , 
     n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , 
     n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , 
     n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , 
     n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , 
     n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , 
     n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , 
     n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , 
     n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , 
     n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , 
     n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , 
     n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , 
     n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , 
     n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , 
     n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , 
     n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , 
     n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , 
     n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , 
     n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , 
     n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , 
     n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , 
     n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , 
     n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , 
     n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , 
     n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , 
     n44260 , n44261 , n571565 , n571566 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , 
     n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , 
     n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , 
     n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , 
     n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , 
     n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , 
     n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , 
     n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , 
     n44340 , n44341 , n44342 , n44343 , n44344 , n571648 , n571649 , n44347 , n44348 , n44349 , 
     n44350 , n44351 , n44352 , n44353 , n44354 , n571658 , n571659 , n44357 , n44358 , n44359 , 
     n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , 
     n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , 
     n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , 
     n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , 
     n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , 
     n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , 
     n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , 
     n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , 
     n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , 
     n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n571759 , n571760 , n44458 , n44459 , 
     n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , 
     n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , 
     n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , 
     n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , 
     n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , 
     n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n571821 , n571822 , 
     n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , 
     n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , 
     n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , 
     n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , 
     n44560 , n44561 , n44562 , n571866 , n571867 , n44565 , n44566 , n44567 , n44568 , n44569 , 
     n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , 
     n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , 
     n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , 
     n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , 
     n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , 
     n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , 
     n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , 
     n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , 
     n44650 , n44651 , n44652 , n44653 , n571957 , n571958 , n44656 , n44657 , n44658 , n44659 , 
     n44660 , n44661 , n44662 , n571966 , n571967 , n44665 , n44666 , n44667 , n44668 , n44669 , 
     n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , 
     n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , 
     n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , 
     n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , 
     n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , 
     n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , 
     n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , 
     n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , 
     n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , 
     n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , 
     n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , 
     n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , 
     n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , 
     n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , 
     n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , 
     n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , 
     n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , 
     n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , 
     n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , 
     n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , 
     n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , 
     n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , 
     n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , 
     n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , 
     n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , 
     n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , 
     n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , 
     n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , 
     n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , 
     n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , 
     n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , 
     n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n572292 , 
     n572293 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n572300 , n572301 , n44999 , 
     n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n572309 , n572310 , n45008 , n45009 , 
     n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n572322 , 
     n572323 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , 
     n45030 , n45031 , n572335 , n572336 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , 
     n45040 , n45041 , n45042 , n45043 , n45044 , n572348 , n572349 , n45047 , n45048 , n45049 , 
     n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n572361 , n572362 , 
     n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , 
     n45070 , n572374 , n572375 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , 
     n45080 , n45081 , n45082 , n45083 , n572387 , n572388 , n45086 , n45087 , n45088 , n45089 , 
     n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n572400 , n572401 , n45099 , 
     n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , 
     n572413 , n572414 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , 
     n45120 , n45121 , n45122 , n572426 , n572427 , n45125 , n45126 , n45127 , n45128 , n45129 , 
     n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n572439 , n572440 , n45138 , n45139 , 
     n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n572452 , 
     n572453 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , 
     n45160 , n45161 , n572465 , n572466 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , 
     n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , 
     n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , 
     n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , 
     n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , 
     n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , 
     n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , 
     n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , 
     n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , 
     n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , 
     n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , 
     n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , 
     n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , 
     n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , 
     n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , 
     n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , 
     n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , 
     n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , 
     n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , 
     n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , 
     n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , 
     n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , 
     n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , 
     n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , 
     n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , 
     n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , 
     n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , 
     n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , 
     n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , 
     n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , 
     n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , 
     n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , 
     n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , 
     n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , 
     n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , 
     n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , 
     n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , 
     n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , 
     n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , 
     n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , 
     n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , 
     n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , 
     n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , 
     n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , 
     n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , 
     n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , 
     n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , 
     n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , 
     n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , 
     n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , 
     n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , 
     n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , 
     n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , 
     n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , 
     n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , 
     n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , 
     n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , 
     n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , 
     n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , 
     n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , 
     n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , 
     n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , 
     n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , 
     n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , 
     n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , 
     n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , 
     n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , 
     n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , 
     n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , 
     n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , 
     n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , 
     n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , 
     n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , 
     n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , 
     n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , 
     n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , 
     n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , 
     n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , 
     n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , 
     n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , 
     n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , 
     n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , 
     n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , 
     n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , 
     n46000 , n46001 , n46002 , n46003 , n46004 , n573308 , n573309 , n573310 , n46005 , n46006 , 
     n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , 
     n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , 
     n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , 
     n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , 
     n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , 
     n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , 
     n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , 
     n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , 
     n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , 
     n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , 
     n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , 
     n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , 
     n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , 
     n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , 
     n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , 
     n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , 
     n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , 
     n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , 
     n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , 
     n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , 
     n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , 
     n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , 
     n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , 
     n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , 
     n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , 
     n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , 
     n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , 
     n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , 
     n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , 
     n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , 
     n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , 
     n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , 
     n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , 
     n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , 
     n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , 
     n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , 
     n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , 
     n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , 
     n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , 
     n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , 
     n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , 
     n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , 
     n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , 
     n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n573752 , 
     n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , 
     n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , 
     n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , 
     n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , 
     n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , 
     n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , 
     n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , 
     n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , 
     n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , 
     n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , 
     n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , 
     n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , 
     n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , 
     n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , 
     n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , 
     n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , 
     n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , 
     n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , 
     n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , 
     n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , 
     n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , 
     n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , 
     n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , 
     n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , 
     n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , 
     n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , 
     n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , 
     n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , 
     n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , 
     n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , 
     n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , 
     n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , 
     n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , 
     n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , 
     n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , 
     n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , 
     n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , 
     n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , 
     n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , 
     n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , 
     n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , 
     n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , 
     n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , 
     n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , 
     n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , 
     n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , 
     n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , 
     n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , 
     n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , 
     n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , 
     n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , 
     n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , 
     n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , 
     n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , 
     n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , 
     n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , 
     n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , 
     n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , 
     n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , 
     n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , 
     n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , 
     n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , 
     n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , 
     n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , 
     n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , 
     n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , 
     n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , 
     n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , 
     n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , 
     n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , 
     n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , 
     n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , 
     n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , 
     n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , 
     n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , 
     n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , 
     n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , 
     n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , 
     n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , 
     n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , 
     n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , 
     n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , 
     n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , 
     n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , 
     n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , 
     n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , 
     n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , 
     n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , 
     n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , 
     n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , 
     n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , 
     n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , 
     n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , 
     n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , 
     n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , 
     n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , 
     n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , 
     n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , 
     n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , 
     n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , 
     n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , 
     n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , 
     n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , 
     n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , 
     n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , 
     n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , 
     n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , 
     n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , 
     n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , 
     n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , 
     n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , 
     n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , 
     n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , 
     n574883 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , 
     n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , 
     n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , 
     n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , 
     n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , 
     n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , 
     n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , 
     n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , 
     n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , 
     n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , 
     n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , 
     n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , 
     n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , 
     n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , 
     n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , 
     n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , 
     n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , 
     n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , 
     n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , 
     n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , 
     n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , 
     n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , 
     n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , 
     n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , 
     n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , 
     n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , 
     n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , 
     n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , 
     n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , 
     n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , 
     n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , 
     n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , 
     n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , 
     n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , 
     n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , 
     n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , 
     n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , 
     n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , 
     n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , 
     n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , 
     n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , 
     n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , 
     n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , 
     n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , 
     n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , 
     n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , 
     n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , 
     n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , 
     n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , 
     n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , 
     n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , 
     n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , 
     n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , 
     n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , 
     n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , 
     n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , 
     n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , 
     n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , 
     n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , 
     n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , 
     n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , 
     n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , 
     n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , 
     n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , 
     n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , 
     n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , 
     n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , 
     n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , 
     n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , 
     n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , 
     n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , 
     n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , 
     n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , 
     n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , 
     n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , 
     n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , 
     n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , 
     n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , 
     n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , 
     n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , 
     n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , 
     n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , 
     n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , 
     n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , 
     n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , 
     n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , 
     n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , 
     n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , 
     n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , 
     n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , 
     n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , 
     n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , 
     n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , 
     n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , 
     n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , 
     n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , 
     n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , 
     n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , 
     n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , 
     n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , 
     n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , 
     n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , 
     n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , 
     n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , 
     n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , 
     n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , 
     n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , 
     n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , 
     n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , 
     n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , 
     n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , 
     n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , 
     n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , 
     n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , 
     n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , 
     n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , 
     n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , 
     n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , 
     n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , 
     n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , 
     n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , 
     n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , 
     n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , 
     n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , 
     n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , 
     n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , 
     n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , 
     n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , 
     n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , 
     n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , 
     n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , 
     n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , 
     n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , 
     n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , 
     n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , 
     n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , 
     n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , 
     n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , 
     n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , 
     n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , 
     n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , 
     n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , 
     n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , 
     n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , 
     n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , 
     n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , 
     n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , 
     n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , 
     n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , 
     n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , 
     n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , 
     n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , 
     n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , 
     n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , 
     n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , 
     n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , 
     n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , 
     n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , 
     n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , 
     n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , 
     n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , 
     n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , 
     n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , 
     n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , 
     n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , 
     n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , 
     n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , 
     n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , 
     n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , 
     n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , 
     n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , 
     n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , 
     n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , 
     n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , 
     n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , 
     n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , 
     n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , 
     n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , 
     n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , 
     n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , 
     n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , 
     n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , 
     n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , 
     n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , 
     n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , 
     n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , 
     n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , 
     n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , 
     n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , 
     n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , 
     n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , 
     n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , 
     n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , 
     n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , 
     n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , 
     n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , 
     n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , 
     n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , 
     n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , 
     n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , 
     n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , 
     n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , 
     n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , 
     n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , 
     n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , 
     n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , 
     n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , 
     n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , 
     n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , 
     n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , 
     n49675 , n49676 , n49677 , n49678 , n49679 , n576988 , n49680 , n49681 , n49682 , n49683 , 
     n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , 
     n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , 
     n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , 
     n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , 
     n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , 
     n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , 
     n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , 
     n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , 
     n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , 
     n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , 
     n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , 
     n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , 
     n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , 
     n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , 
     n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , 
     n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , 
     n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , 
     n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , 
     n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , 
     n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , 
     n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , 
     n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , 
     n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , 
     n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , 
     n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , 
     n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , 
     n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , 
     n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , 
     n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , 
     n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , 
     n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , 
     n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , 
     n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , 
     n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , 
     n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , 
     n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , 
     n50044 , n50045 , n50046 , n50047 , n50048 , n577358 , n577359 , n577360 , n50049 , n50050 , 
     n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , 
     n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , 
     n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , 
     n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , 
     n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , 
     n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , 
     n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , 
     n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , 
     n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , 
     n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , 
     n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , 
     n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , 
     n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , 
     n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , 
     n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , 
     n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , 
     n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , 
     n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , 
     n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , 
     n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , 
     n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , 
     n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , 
     n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , 
     n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , 
     n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , 
     n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , 
     n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , 
     n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , 
     n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , 
     n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , 
     n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , 
     n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , 
     n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , 
     n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , 
     n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , 
     n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , 
     n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , 
     n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , 
     n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , 
     n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , 
     n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , 
     n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , 
     n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , 
     n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , 
     n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , 
     n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , 
     n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , 
     n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n577840 , n50528 , n50529 , 
     n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , 
     n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , 
     n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , 
     n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , 
     n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , 
     n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , 
     n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , 
     n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , 
     n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , 
     n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , 
     n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , 
     n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , 
     n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , 
     n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , 
     n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , 
     n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , 
     n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , 
     n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , 
     n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , 
     n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , 
     n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , 
     n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , 
     n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , 
     n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , 
     n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , 
     n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , 
     n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , 
     n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , 
     n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , 
     n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , 
     n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , 
     n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , 
     n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , 
     n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , 
     n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , 
     n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , 
     n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , 
     n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , 
     n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , 
     n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , 
     n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , 
     n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , 
     n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , 
     n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , 
     n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , 
     n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , 
     n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , 
     n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , 
     n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , 
     n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , 
     n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , 
     n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , 
     n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , 
     n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , 
     n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , 
     n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , 
     n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , 
     n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , 
     n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , 
     n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , 
     n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , 
     n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , 
     n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , 
     n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , 
     n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , 
     n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , 
     n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , 
     n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , 
     n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , 
     n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , 
     n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , 
     n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , 
     n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , 
     n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n578582 , 
     n51270 , n578584 , n51272 , n578586 , n51274 , n578588 , n51276 , n578590 , n51278 , n578592 , 
     n51280 , n578594 , n51282 , n578596 , n51284 , n578598 , n51286 , n578600 , n51288 , n578602 , 
     n51290 , n578604 , n51292 , n578606 , n51294 , n578608 , n51296 , n578610 , n51298 , n578612 , 
     n51300 , n578614 , n51302 , n578616 , n51304 , n578618 , n51306 , n578620 , n51308 , n578622 , 
     n51310 , n578624 , n51312 , n578626 , n51314 , n578628 , n51316 , n578630 , n51318 , n578632 , 
     n51320 , n578634 , n51322 , n578636 , n51324 , n578638 , n578639 , n51327 , n578641 , n51329 , 
     n578643 , n51331 , n578645 , n51333 , n578647 , n51335 , n578649 , n51337 , n578651 , n51339 , 
     n578653 , n51341 , n578655 , n51343 , n578657 , n51345 , n578659 , n51347 , n578661 , n51349 , 
     n578663 , n51351 , n578665 , n51353 , n578667 , n51355 , n578669 , n51357 , n578671 , n51359 , 
     n578673 , n51361 , n578675 , n51363 , n578677 , n51365 , n578679 , n578680 , n578681 , n578682 , 
     n578683 , n51368 , n578685 , n51370 , n578687 , n51372 , n578689 , n51374 , n578691 , n51376 , 
     n578693 , n51378 , n578695 , n51380 , n578697 , n51382 , n578699 , n51384 , n578701 , n51386 , 
     n578703 , n51388 , n578705 , n51390 , n578707 , n51392 , n578709 , n51394 , n578711 , n51396 , 
     n578713 , n51398 , n578715 , n51400 , n578717 , n51402 , n578719 , n51404 , n578721 , n51406 , 
     n578723 , n51408 , n578725 , n51410 , n578727 , n51412 , n578729 , n51414 , n578731 , n51416 , 
     n578733 , n51418 , n578735 , n51420 , n578737 , n51422 , n578739 , n51424 , n578741 , n51426 , 
     n578743 , n51428 , n578745 , n51430 , n578747 , n51432 , n578749 , n51434 , n578751 , n51436 , 
     n578753 , n51438 , n578755 , n51440 , n578757 , n51442 , n578759 , n51444 , n578761 , n51446 , 
     n578763 , n51448 , n578765 , n51450 , n578767 , n51452 , n578769 , n51454 , n578771 , n51456 , 
     n578773 , n51458 , n578775 , n51460 , n578777 , n51462 , n578779 , n51464 , n578781 , n51466 , 
     n578783 , n51468 , n578785 , n51470 , n578787 , n51472 , n578789 , n51474 , n578791 , n51476 , 
     n578793 , n51478 , n578795 , n51480 , n578797 , n51482 , n51483 , n578800 , n51485 , n51486 , 
     n578803 , n51488 , n51489 , n578806 , n51491 , n51492 , n578809 , n51494 , n51495 , n578812 , 
     n51497 , n51498 , n578815 , n51500 , n51501 , n578818 , n51503 , n51504 , n578821 , n51506 , 
     n51507 , n578824 , n51509 , n51510 , n578827 , n51512 , n51513 , n578830 , n51515 , n51516 , 
     n578833 , n51518 , n51519 , n578836 , n51521 , n51522 , n578839 , n51524 , n51525 , n578842 , 
     n51527 , n51528 , n578845 , n51530 , n51531 , n578848 , n51533 , n51534 , n578851 , n51536 , 
     n51537 , n578854 , n51539 , n578856 , n578857 , n578858 , n578859 , n578860 , n578861 , n578862 , 
     n578863 , n578864 , n578865 , n578866 , n578867 , n578868 , n578869 , n578870 , n578871 , n578872 , 
     n578873 , n578874 , n578875 , n578876 , n578877 , n578878 , n578879 , n578880 , n578881 , n578882 , 
     n578883 , n578884 , n578885 , n578886 , n578887 , n578888 , n578889 , n578890 , n578891 , n578892 , 
     n578893 , n578894 , n578895 , n578896 , n578897 , n578898 , n578899 , n578900 , n578901 , n578902 , 
     n578903 , n578904 , n578905 , n578906 , n578907 , n578908 , n578909 , n578910 , n578911 , n578912 , 
     n578913 , n578914 , n578915 , n578916 , n578917 , n578918 , n578919 , n578920 , n578921 , n578922 , 
     n578923 , n51608 , n578925 , n578926 , n51611 , n578928 , n578929 , n51614 , n578931 , n578932 , 
     n51617 , n578934 , n578935 , n51620 , n578937 , n578938 , n51623 , n578940 , n578941 , n51626 , 
     n578943 , n578944 , n51629 , n578946 , n578947 , n51632 , n578949 , n578950 , n51635 , n578952 , 
     n578953 , n51638 , n578955 , n578956 , n51641 , n578958 , n578959 , n51644 , n578961 , n578962 , 
     n51647 , n578964 , n578965 , n51650 , n578967 , n578968 , n51653 , n578970 , n578971 , n51656 , 
     n578973 , n578974 , n51659 , n578976 , n578977 , n51662 , n578979 , n578980 , n51665 , n578982 , 
     n578983 , n51668 , n578985 , n578986 , n51671 , n578988 , n578989 , n51674 , n578991 , n578992 , 
     n51677 , n578994 , n578995 , n51680 , n578997 , n578998 , n51683 , n579000 , n579001 , n51686 , 
     n579003 , n579004 , n51689 , n579006 , n579007 , n51692 , n579009 , n579010 , n51695 , n579012 , 
     n579013 , n51698 , n579015 , n579016 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , 
     n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , 
     n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , 
     n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , 
     n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , 
     n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , 
     n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , 
     n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , 
     n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , 
     n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n579111 , n579112 , 
     n51797 , n51798 , n579115 , n579116 , n51801 , n51802 , n579119 , n579120 , n51805 , n51806 , 
     n579123 , n579124 , n51809 , n51810 , n579127 , n579128 , n51813 , n51814 , n579131 , n579132 , 
     n51817 , n51818 , n579135 , n579136 , n51821 , n51822 , n579139 , n579140 , n51825 , n51826 , 
     n579143 , n579144 , n51829 , n51830 , n579147 , n579148 , n51833 , n51834 , n579151 , n579152 , 
     n51837 , n51838 , n579155 , n579156 , n51841 , n51842 , n579159 , n579160 , n51845 , n51846 , 
     n579163 , n579164 , n51849 , n51850 , n579167 , n579168 , n51853 , n51854 , n579171 , n579172 , 
     n51857 , n51858 , n579175 , n579176 , n51861 , n51862 , n579179 , n579180 , n51865 , n51866 , 
     n579183 , n579184 , n51869 , n51870 , n579187 , n579188 , n51873 , n51874 , n579191 , n579192 , 
     n51877 , n51878 , n579195 , n579196 , n51881 , n51882 , n579199 , n579200 , n51885 , n51886 , 
     n579203 , n579204 , n51889 , n51890 , n579207 , n579208 , n51893 , n51894 , n579211 , n579212 , 
     n51897 , n51898 , n579215 , n579216 , n51901 , n51902 , n579219 , n579220 , n51905 , n51906 , 
     n579223 , n579224 , n51909 , n51910 , n579227 , n579228 , n51913 , n51914 , n579231 , n579232 , 
     n51917 , n51918 , n579235 , n579236 , n51921 , n579238 , n579239 , n51924 , n51925 , n51926 , 
     n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , 
     n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , 
     n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , 
     n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n579281 , n51965 , 
     n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , 
     n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , 
     n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , 
     n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , 
     n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , 
     n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , 
     n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , 
     n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , 
     n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , 
     n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , 
     n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , 
     n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , 
     n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , 
     n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , 
     n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , 
     n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , 
     n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , 
     n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , 
     n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , 
     n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , 
     n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , 
     n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , 
     n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , 
     n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , 
     n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , 
     n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , 
     n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , 
     n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , 
     n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , 
     n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , 
     n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , 
     n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , 
     n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , 
     n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , 
     n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , 
     n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , 
     n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , 
     n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , 
     n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , 
     n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , 
     n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , 
     n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , 
     n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , 
     n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , 
     n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , 
     n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , 
     n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , 
     n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , 
     n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , 
     n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , 
     n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , 
     n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , 
     n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , 
     n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , 
     n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , 
     n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , 
     n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , 
     n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , 
     n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , 
     n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , 
     n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , 
     n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , 
     n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , 
     n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , 
     n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , 
     n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , 
     n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , 
     n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , 
     n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , 
     n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , 
     n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , 
     n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , 
     n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , 
     n52696 , n580014 , n580015 , n580016 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , 
     n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , 
     n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , 
     n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , 
     n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , 
     n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , 
     n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , 
     n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , 
     n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , 
     n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , 
     n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , 
     n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , 
     n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , 
     n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , 
     n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , 
     n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , 
     n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , 
     n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , 
     n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , 
     n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , 
     n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , 
     n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , 
     n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , 
     n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , 
     n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , 
     n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , 
     n52953 , n52954 , n580275 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , 
     n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , 
     n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , 
     n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , 
     n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , 
     n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , 
     n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , 
     n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , 
     n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , 
     n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , 
     n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , 
     n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , 
     n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , 
     n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , 
     n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , 
     n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , 
     n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , 
     n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , 
     n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , 
     n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , 
     n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , 
     n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , 
     n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , 
     n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , 
     n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , 
     n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , 
     n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , 
     n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , 
     n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , 
     n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , 
     n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , 
     n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , 
     n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n580602 , 
     n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , 
     n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , 
     n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , 
     n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , 
     n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , 
     n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , 
     n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , 
     n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , 
     n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , 
     n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , 
     n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , 
     n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , 
     n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , 
     n53411 , n53412 , n580735 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , 
     n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , 
     n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , 
     n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , 
     n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , 
     n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , 
     n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , 
     n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , 
     n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , 
     n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , 
     n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , 
     n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , 
     n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , 
     n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , 
     n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , 
     n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , 
     n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , 
     n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , 
     n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , 
     n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , 
     n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , 
     n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , 
     n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , 
     n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , 
     n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , 
     n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , 
     n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , 
     n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , 
     n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , 
     n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , 
     n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , 
     n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , 
     n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , 
     n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , 
     n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , 
     n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , 
     n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , 
     n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , 
     n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , 
     n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , 
     n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , 
     n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , 
     n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , 
     n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , 
     n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , 
     n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , 
     n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , 
     n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , 
     n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , 
     n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , 
     n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , 
     n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , 
     n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , 
     n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , 
     n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , 
     n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , 
     n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , 
     n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , 
     n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , 
     n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , 
     n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , 
     n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , 
     n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , 
     n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , 
     n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , 
     n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , 
     n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , 
     n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , 
     n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , 
     n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , 
     n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , 
     n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , 
     n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , 
     n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , 
     n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , 
     n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , 
     n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , 
     n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , 
     n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , 
     n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , 
     n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , 
     n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , 
     n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , 
     n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , 
     n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , 
     n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , 
     n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , 
     n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , 
     n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , 
     n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , 
     n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , 
     n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , 
     n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , 
     n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , 
     n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , 
     n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , 
     n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , 
     n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , 
     n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , 
     n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , 
     n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , 
     n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , 
     n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , 
     n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , 
     n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , 
     n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , 
     n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , 
     n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , 
     n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , 
     n54500 , n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , n54509 , 
     n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , 
     n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , 
     n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , 
     n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , 
     n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , 
     n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , 
     n54570 , n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , n54579 , 
     n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , 
     n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , 
     n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , 
     n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , 
     n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , 
     n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , 
     n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , 
     n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , 
     n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , 
     n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , 
     n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , 
     n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , 
     n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , 
     n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , 
     n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , 
     n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , 
     n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , 
     n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , 
     n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , 
     n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , 
     n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , 
     n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , 
     n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , 
     n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , 
     n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , 
     n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , 
     n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , 
     n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , 
     n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , 
     n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , 
     n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , 
     n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , 
     n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , 
     n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , 
     n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , 
     n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , 
     n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , 
     n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , 
     n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , 
     n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , 
     n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , 
     n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , 
     n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , 
     n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , 
     n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , 
     n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , 
     n55040 , n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , n55049 , 
     n55050 , n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , n55059 , 
     n55060 , n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , n55069 , 
     n55070 , n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , n55079 , 
     n55080 , n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , n55089 , 
     n55090 , n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , n55099 , 
     n55100 , n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , n55109 , 
     n55110 , n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , n55119 , 
     n55120 , n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , n55127 , n55128 , n55129 , 
     n55130 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , n55139 , 
     n55140 , n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , n55149 , 
     n55150 , n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , 
     n55160 , n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , n55169 , 
     n55170 , n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , n55177 , n55178 , n55179 , 
     n55180 , n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , n55189 , 
     n55190 , n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , n55199 , 
     n55200 , n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , n55209 , 
     n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , n55219 , 
     n55220 , n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , n55229 , 
     n55230 , n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , n55239 , 
     n55240 , n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , n55249 , 
     n55250 , n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , n55259 , 
     n55260 , n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , n55269 , 
     n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , n55279 , 
     n55280 , n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , n55289 , 
     n55290 , n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , n55299 , 
     n55300 , n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , n55309 , 
     n55310 , n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , n55319 , 
     n55320 , n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , n55329 , 
     n55330 , n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , n55339 , 
     n55340 , n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , n55349 , 
     n55350 , n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , n55359 , 
     n55360 , n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , n55367 , n55368 , n55369 , 
     n55370 , n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , n55379 , 
     n55380 , n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , n55387 , n55388 , n55389 , 
     n55390 , n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , n55397 , n55398 , n55399 , 
     n55400 , n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , n55407 , n55408 , n55409 , 
     n55410 , n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , n55417 , n55418 , n55419 , 
     n55420 , n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , n55427 , n55428 , n55429 , 
     n55430 , n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , n55437 , n55438 , n55439 , 
     n55440 , n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , n55447 , n55448 , n55449 , 
     n55450 , n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , n55457 , n55458 , n55459 , 
     n55460 , n55461 , n582785 , n582786 , n55464 , n582788 , n582789 , n582790 , n55468 , n582792 , 
     n55470 , n582794 , n582795 , n55473 , n582797 , n55475 , n582799 , n582800 , n55478 , n582802 , 
     n582803 , n582804 , n582805 , n55483 , n582807 , n582808 , n55486 , n582810 , n582811 , n55489 , 
     n582813 , n582814 , n55492 , n582816 , n582817 , n582818 , n55496 , n582820 , n582821 , n582822 , 
     n55500 , n582824 , n55502 , n582826 , n582827 , n55505 , n582829 , n55507 , n55508 , n55509 , 
     n55510 , n582834 , n582835 , n582836 , n55514 , n582838 , n582839 , n582840 , n582841 , n55519 , 
     n582843 , n582844 , n55522 , n582846 , n582847 , n55525 , n582849 , n582850 , n55528 , n582852 , 
     n582853 , n582854 , n582855 , n55533 , n582857 , n582858 , n582859 , n582860 , n55538 , n582862 , 
     n582863 , n55541 , n582865 , n582866 , n55544 , n582868 , n582869 , n55547 , n55548 , n55549 , 
     n582873 , n582874 , n55552 , n582876 , n55554 , n55555 , n55556 , n55557 , n55558 , n55559 , 
     n582883 , n582884 , n55562 , n582886 , n582887 , n55565 , n582889 , n582890 , n55568 , n582892 , 
     n582893 , n55571 , n582895 , n55573 , n582897 , n55575 , n55576 , n55577 , n55578 , n582902 , 
     n582903 , n55581 , n582905 , n55583 , n582907 , n55585 , n582909 , n582910 , n55588 , n582912 , 
     n582913 , n582914 , n582915 , n55593 , n582917 , n582918 , n55596 , n582920 , n582921 , n55599 , 
     n582923 , n582924 , n55602 , n55603 , n55604 , n582928 , n582929 , n582930 , n55608 , n582932 , 
     n55610 , n55611 , n582935 , n582936 , n55614 , n582938 , n55616 , n55617 , n55618 , n55619 , 
     n55620 , n55621 , n582945 , n55623 , n582947 , n55625 , n582949 , n582950 , n55628 , n582952 , 
     n582953 , n582954 , n582955 , n55633 , n582957 , n582958 , n55636 , n582960 , n582961 , n55639 , 
     n582963 , n582964 , n55642 , n55643 , n55644 , n582968 , n582969 , n582970 , n582971 , n55649 , 
     n582973 , n582974 , n582975 , n55653 , n582977 , n582978 , n55656 , n582980 , n55658 , n582982 , 
     n582983 , n55661 , n582985 , n55663 , n582987 , n55665 , n55666 , n582990 , n582991 , n55669 , 
     n582993 , n582994 , n55672 , n582996 , n582997 , n55675 , n582999 , n583000 , n55678 , n583002 , 
     n583003 , n55681 , n583005 , n583006 , n583007 , n583008 , n55686 , n583010 , n583011 , n55689 , 
     n583013 , n583014 , n55692 , n583016 , n583017 , n55695 , n55696 , n55697 , n583021 , n583022 , 
     n55700 , n55701 , n55702 , n583026 , n583027 , n55705 , n583029 , n55707 , n55708 , n55709 , 
     n55710 , n55711 , n583035 , n55713 , n583037 , n583038 , n55716 , n583040 , n55718 , n583042 , 
     n583043 , n55721 , n55722 , n55723 , n55724 , n583048 , n55726 , n583050 , n55728 , n55729 , 
     n583053 , n55731 , n583055 , n583056 , n55734 , n583058 , n55736 , n55737 , n583061 , n55739 , 
     n55740 , n55741 , n583065 , n55743 , n55744 , n583068 , n55746 , n55747 , n55748 , n583072 , 
     n583073 , n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , n55757 , n55758 , n583082 , 
     n583083 , n583084 , n55762 , n583086 , n583087 , n583088 , n55766 , n583090 , n583091 , n583092 , 
     n55770 , n583094 , n583095 , n55773 , n583097 , n583098 , n55776 , n583100 , n583101 , n583102 , 
     n583103 , n55781 , n583105 , n583106 , n583107 , n583108 , n55786 , n583110 , n583111 , n55789 , 
     n583113 , n583114 , n55792 , n583116 , n583117 , n55795 , n583119 , n583120 , n583121 , n583122 , 
     n55800 , n583124 , n583125 , n583126 , n583127 , n55805 , n583129 , n583130 , n55808 , n583132 , 
     n583133 , n55811 , n583135 , n583136 , n55814 , n583138 , n583139 , n55817 , n583141 , n583142 , 
     n55820 , n55821 , n583145 , n55823 , n583147 , n583148 , n55826 , n55827 , n583151 , n55829 , 
     n583153 , n55831 , n583155 , n55833 , n583157 , n583158 , n55836 , n583160 , n55838 , n583162 , 
     n55840 , n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , n55847 , n55848 , n583172 , 
     n583173 , n55851 , n583175 , n583176 , n583177 , n55855 , n583179 , n583180 , n583181 , n55859 , 
     n583183 , n583184 , n55862 , n583186 , n55864 , n583188 , n583189 , n55867 , n583191 , n55869 , 
     n583193 , n55871 , n55872 , n583196 , n583197 , n55875 , n583199 , n583200 , n55878 , n583202 , 
     n583203 , n55881 , n583205 , n583206 , n583207 , n55885 , n583209 , n583210 , n55888 , n583212 , 
     n55890 , n583214 , n583215 , n583216 , n583217 , n55895 , n583219 , n583220 , n55898 , n583222 , 
     n55900 , n583224 , n55902 , n55903 , n583227 , n583228 , n55906 , n583230 , n583231 , n55909 , 
     n583233 , n583234 , n55912 , n583236 , n583237 , n55915 , n583239 , n583240 , n55918 , n583242 , 
     n583243 , n583244 , n55922 , n583246 , n55924 , n583248 , n583249 , n55927 , n583251 , n55929 , 
     n55930 , n55931 , n583255 , n55933 , n55934 , n55935 , n583259 , n583260 , n55938 , n583262 , 
     n55940 , n55941 , n583265 , n55943 , n583267 , n583268 , n55946 , n55947 , n55948 , n583272 , 
     n583273 , n55951 , n583275 , n583276 , n55954 , n583278 , n583279 , n583280 , n583281 , n55959 , 
     n583283 , n583284 , n55962 , n583286 , n583287 , n55965 , n583289 , n583290 , n55968 , n55969 , 
     n55970 , n583294 , n583295 , n55973 , n55974 , n583298 , n583299 , n55977 , n55978 , n55979 , 
     n583303 , n583304 , n55982 , n583306 , n583307 , n55985 , n583309 , n583310 , n55988 , n55989 , 
     n583313 , n583314 , n55992 , n583316 , n55994 , n55995 , n55996 , n55997 , n55998 , n55999 , 
     n56000 , n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , n56007 , n56008 , n56009 , 
     n56010 , n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , n56017 , n56018 , n56019 , 
     n56020 , n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , n56027 , n56028 , n56029 , 
     n56030 , n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , n56037 , n56038 , n583362 , 
     n583363 , n583364 , n56042 , n583366 , n583367 , n583368 , n583369 , n56047 , n583371 , n583372 , 
     n56050 , n583374 , n583375 , n56053 , n583377 , n583378 , n56056 , n583380 , n583381 , n583382 , 
     n56060 , n583384 , n583385 , n583386 , n56064 , n583388 , n56066 , n583390 , n583391 , n56069 , 
     n583393 , n56071 , n56072 , n583396 , n583397 , n56075 , n583399 , n583400 , n583401 , n583402 , 
     n56080 , n583404 , n583405 , n56083 , n583407 , n583408 , n56086 , n583410 , n583411 , n56089 , 
     n583413 , n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , n56097 , n56098 , n56099 , 
     n583423 , n583424 , n56102 , n56103 , n56104 , n56105 , n583429 , n583430 , n56108 , n583432 , 
     n583433 , n56111 , n583435 , n583436 , n583437 , n583438 , n56116 , n583440 , n583441 , n56119 , 
     n583443 , n583444 , n56122 , n583446 , n583447 , n56125 , n583449 , n583450 , n56128 , n583452 , 
     n56130 , n56131 , n56132 , n56133 , n56134 , n56135 , n583459 , n56137 , n56138 , n56139 , 
     n56140 , n583464 , n583465 , n56143 , n583467 , n56145 , n56146 , n56147 , n56148 , n56149 , 
     n56150 , n56151 , n56152 , n56153 , n56154 , n56155 , n56156 , n56157 , n56158 , n56159 , 
     n583483 , n56161 , n583485 , n583486 , n56164 , n583488 , n56166 , n583490 , n583491 , n56169 , 
     n56170 , n56171 , n583495 , n583496 , n56174 , n56175 , n56176 , n583500 , n583501 , n56179 , 
     n56180 , n56181 , n56182 , n56183 , n56184 , n56185 , n583509 , n583510 , n56188 , n583512 , 
     n56190 , n583514 , n56192 , n583516 , n56194 , n583518 , n56196 , n56197 , n56198 , n56199 , 
     n56200 , n56201 , n56202 , n56203 , n56204 , n56205 , n56206 , n56207 , n56208 , n56209 , 
     n56210 , n56211 , n56212 , n56213 , n56214 , n56215 , n56216 , n56217 , n56218 , n56219 , 
     n56220 , n56221 , n56222 , n56223 , n56224 , n56225 , n56226 , n56227 , n56228 , n56229 , 
     n56230 , n56231 , n56232 , n56233 , n56234 , n56235 , n56236 , n56237 , n56238 , n56239 , 
     n583563 , n56241 , n583565 , n56243 , n56244 , n56245 , n56246 , n56247 , n56248 , n56249 , 
     n56250 , n56251 , n583575 , n583576 , n56254 , n56255 , n56256 , n56257 , n583581 , n56259 , 
     n583583 , n583584 , n56262 , n56263 , n56264 , n56265 , n583589 , n583590 , n56268 , n583592 , 
     n583593 , n56271 , n56272 , n56273 , n56274 , n583598 , n583599 , n56277 , n56278 , n56279 , 
     n56280 , n583604 , n56282 , n583606 , n583607 , n56285 , n583609 , n583610 , n583611 , n583612 , 
     n56290 , n583614 , n583615 , n56293 , n583617 , n583618 , n56296 , n583620 , n583621 , n56299 , 
     n583623 , n583624 , n56302 , n583626 , n583627 , n56305 , n583629 , n583630 , n56308 , n583632 , 
     n583633 , n56311 , n56312 , n583636 , n583637 , n56315 , n56316 , n56317 , n583641 , n56319 , 
     n583643 , n583644 , n56322 , n583646 , n583647 , n56325 , n583649 , n56327 , n56328 , n583652 , 
     n56330 , n583654 , n583655 , n56333 , n56334 , n56335 , n56336 , n583660 , n583661 , n56339 , 
     n583663 , n583664 , n56342 , n583666 , n56344 , n56345 , n583669 , n56347 , n583671 , n583672 , 
     n56350 , n583674 , n583675 , n583676 , n56354 , n583678 , n56356 , n583680 , n583681 , n56359 , 
     n583683 , n56361 , n56362 , n56363 , n56364 , n56365 , n583689 , n583690 , n583691 , n56369 , 
     n583693 , n583694 , n583695 , n583696 , n56374 , n583698 , n583699 , n56377 , n583701 , n583702 , 
     n56380 , n583704 , n583705 , n56383 , n583707 , n56385 , n56386 , n583710 , n56388 , n56389 , 
     n56390 , n56391 , n583715 , n583716 , n56394 , n583718 , n583719 , n583720 , n56398 , n583722 , 
     n583723 , n583724 , n583725 , n56403 , n583727 , n583728 , n56406 , n583730 , n583731 , n56409 , 
     n583733 , n583734 , n56412 , n583736 , n583737 , n583738 , n56416 , n583740 , n583741 , n583742 , 
     n583743 , n56421 , n583745 , n583746 , n56424 , n583748 , n583749 , n56427 , n583751 , n583752 , 
     n56430 , n583754 , n56432 , n56433 , n56434 , n56435 , n56436 , n56437 , n56438 , n56439 , 
     n583763 , n56441 , n583765 , n56443 , n56444 , n583768 , n56446 , n583770 , n56448 , n56449 , 
     n56450 , n56451 , n56452 , n56453 , n583777 , n56455 , n583779 , n583780 , n56458 , n56459 , 
     n583783 , n583784 , n56462 , n56463 , n583787 , n583788 , n56466 , n583790 , n583791 , n56469 , 
     n56470 , n583794 , n583795 , n56473 , n583797 , n583798 , n56476 , n583800 , n583801 , n56479 , 
     n56480 , n56481 , n56482 , n56483 , n56484 , n56485 , n56486 , n583810 , n56488 , n56489 , 
     n56490 , n56491 , n583815 , n56493 , n56494 , n56495 , n56496 , n56497 , n56498 , n56499 , 
     n56500 , n56501 , n56502 , n56503 , n56504 , n583828 , n583829 , n583830 , n56508 , n583832 , 
     n583833 , n56511 , n56512 , n583836 , n56514 , n56515 , n583839 , n583840 , n56518 , n583842 , 
     n583843 , n56521 , n583845 , n583846 , n56524 , n583848 , n583849 , n56527 , n583851 , n583852 , 
     n583853 , n56531 , n583855 , n56533 , n56534 , n56535 , n56536 , n56537 , n56538 , n56539 , 
     n56540 , n56541 , n56542 , n56543 , n56544 , n56545 , n56546 , n56547 , n583871 , n56549 , 
     n583873 , n583874 , n56552 , n583876 , n56554 , n56555 , n56556 , n56557 , n56558 , n56559 , 
     n56560 , n56561 , n56562 , n56563 , n56564 , n583888 , n56566 , n583890 , n583891 , n56569 , 
     n583893 , n583894 , n56572 , n583896 , n583897 , n56575 , n583899 , n56577 , n56578 , n56579 , 
     n56580 , n56581 , n583905 , n56583 , n56584 , n583908 , n56586 , n56587 , n56588 , n56589 , 
     n583913 , n583914 , n583915 , n56593 , n583917 , n583918 , n583919 , n56597 , n583921 , n56599 , 
     n583923 , n583924 , n56602 , n583926 , n56604 , n583928 , n583929 , n583930 , n56608 , n583932 , 
     n583933 , n583934 , n583935 , n56613 , n583937 , n583938 , n56616 , n583940 , n583941 , n56619 , 
     n583943 , n583944 , n56622 , n583946 , n583947 , n56625 , n583949 , n583950 , n56628 , n583952 , 
     n583953 , n583954 , n583955 , n56633 , n583957 , n583958 , n56636 , n583960 , n583961 , n56639 , 
     n583963 , n583964 , n56642 , n583966 , n583967 , n56645 , n56646 , n56647 , n583971 , n583972 , 
     n56650 , n583974 , n583975 , n583976 , n583977 , n56655 , n583979 , n56657 , n583981 , n583982 , 
     n56660 , n583984 , n583985 , n583986 , n583987 , n56665 , n583989 , n583990 , n56668 , n583992 , 
     n56670 , n56671 , n56672 , n56673 , n583997 , n583998 , n56676 , n584000 , n56678 , n584002 , 
     n584003 , n56681 , n584005 , n584006 , n584007 , n56685 , n584009 , n584010 , n584011 , n56689 , 
     n584013 , n584014 , n56692 , n584016 , n56694 , n56695 , n56696 , n56697 , n56698 , n56699 , 
     n584023 , n584024 , n56702 , n584026 , n584027 , n56705 , n584029 , n584030 , n584031 , n56709 , 
     n584033 , n584034 , n56712 , n584036 , n56714 , n56715 , n584039 , n584040 , n56718 , n584042 , 
     n56720 , n56721 , n56722 , n56723 , n56724 , n56725 , n56726 , n56727 , n56728 , n56729 , 
     n56730 , n56731 , n56732 , n56733 , n584057 , n56735 , n56736 , n584060 , n56738 , n56739 , 
     n584063 , n584064 , n56742 , n56743 , n584067 , n584068 , n56746 , n584070 , n584071 , n56749 , 
     n56750 , n584074 , n56752 , n584076 , n584077 , n56755 , n584079 , n584080 , n56758 , n584082 , 
     n584083 , n56761 , n584085 , n584086 , n584087 , n584088 , n56766 , n584090 , n584091 , n56769 , 
     n584093 , n584094 , n56772 , n584096 , n584097 , n56775 , n584099 , n584100 , n584101 , n56779 , 
     n584103 , n584104 , n584105 , n56783 , n584107 , n56785 , n584109 , n584110 , n56788 , n584112 , 
     n56790 , n56791 , n56792 , n56793 , n584117 , n584118 , n56796 , n584120 , n584121 , n584122 , 
     n56800 , n584124 , n56802 , n584126 , n584127 , n56805 , n584129 , n56807 , n56808 , n56809 , 
     n56810 , n56811 , n56812 , n56813 , n56814 , n56815 , n56816 , n56817 , n56818 , n56819 , 
     n56820 , n584144 , n584145 , n56823 , n584147 , n584148 , n584149 , n56827 , n584151 , n56829 , 
     n584153 , n584154 , n56832 , n584156 , n56834 , n584158 , n584159 , n56837 , n584161 , n584162 , 
     n584163 , n56841 , n584165 , n56843 , n584167 , n584168 , n56846 , n584170 , n56848 , n56849 , 
     n56850 , n584174 , n584175 , n56853 , n584177 , n584178 , n584179 , n584180 , n56858 , n584182 , 
     n584183 , n56861 , n584185 , n584186 , n56864 , n56865 , n584189 , n56867 , n56868 , n584192 , 
     n584193 , n56871 , n584195 , n584196 , n56874 , n584198 , n56876 , n56877 , n56878 , n56879 , 
     n56880 , n56881 , n56882 , n56883 , n584207 , n56885 , n584209 , n584210 , n56888 , n56889 , 
     n584213 , n584214 , n56892 , n56893 , n584217 , n56895 , n56896 , n584220 , n56898 , n584222 , 
     n584223 , n56901 , n584225 , n584226 , n584227 , n584228 , n56906 , n584230 , n584231 , n56909 , 
     n584233 , n584234 , n56912 , n584236 , n584237 , n56915 , n56916 , n56917 , n584241 , n584242 , 
     n584243 , n56921 , n584245 , n584246 , n56924 , n584248 , n584249 , n56927 , n584251 , n584252 , 
     n56930 , n56931 , n584255 , n584256 , n56934 , n584258 , n584259 , n56937 , n584261 , n584262 , 
     n56940 , n584264 , n584265 , n56943 , n584267 , n56945 , n56946 , n56947 , n56948 , n56949 , 
     n56950 , n56951 , n56952 , n584276 , n584277 , n56955 , n584279 , n584280 , n584281 , n584282 , 
     n56960 , n584284 , n584285 , n56963 , n584287 , n584288 , n56966 , n584290 , n584291 , n56969 , 
     n56970 , n56971 , n584295 , n584296 , n584297 , n584298 , n56976 , n584300 , n584301 , n584302 , 
     n584303 , n56981 , n584305 , n584306 , n56984 , n584308 , n584309 , n56987 , n584311 , n584312 , 
     n56990 , n56991 , n56992 , n584316 , n584317 , n56995 , n584319 , n584320 , n56998 , n584322 , 
     n584323 , n584324 , n584325 , n57003 , n584327 , n584328 , n57006 , n584330 , n584331 , n57009 , 
     n584333 , n584334 , n57012 , n57013 , n57014 , n584338 , n584339 , n57017 , n584341 , n57019 , 
     n57020 , n57021 , n57022 , n57023 , n57024 , n57025 , n57026 , n57027 , n584351 , n57029 , 
     n57030 , n57031 , n57032 , n57033 , n57034 , n584358 , n584359 , n57037 , n57038 , n57039 , 
     n57040 , n584364 , n57042 , n57043 , n57044 , n57045 , n584369 , n584370 , n57048 , n57049 , 
     n57050 , n57051 , n57052 , n584376 , n57054 , n584378 , n584379 , n57057 , n57058 , n57059 , 
     n57060 , n57061 , n584385 , n584386 , n57064 , n584388 , n57066 , n57067 , n57068 , n57069 , 
     n57070 , n57071 , n57072 , n584396 , n57074 , n584398 , n584399 , n57077 , n584401 , n57079 , 
     n57080 , n57081 , n584405 , n57083 , n584407 , n584408 , n57086 , n57087 , n584411 , n57089 , 
     n584413 , n57091 , n584415 , n584416 , n57094 , n584418 , n584419 , n584420 , n584421 , n57099 , 
     n584423 , n57101 , n584425 , n57103 , n57104 , n584428 , n57106 , n584430 , n584431 , n57109 , 
     n584433 , n584434 , n57112 , n57113 , n57114 , n57115 , n584439 , n584440 , n57118 , n584442 , 
     n584443 , n57121 , n584445 , n57123 , n584447 , n57125 , n57126 , n584450 , n57128 , n584452 , 
     n584453 , n57131 , n584455 , n584456 , n57134 , n584458 , n584459 , n57137 , n584461 , n57139 , 
     n57140 , n57141 , n57142 , n584466 , n584467 , n57145 , n584469 , n57147 , n57148 , n57149 , 
     n57150 , n57151 , n57152 , n57153 , n57154 , n57155 , n57156 , n584480 , n57158 , n57159 , 
     n57160 , n57161 , n57162 , n57163 , n57164 , n57165 , n57166 , n57167 , n57168 , n57169 , 
     n57170 , n57171 , n57172 , n57173 , n57174 , n57175 , n57176 , n57177 , n57178 , n57179 , 
     n57180 , n57181 , n57182 , n57183 , n584507 , n57185 , n57186 , n584510 , n584511 , n57189 , 
     n584513 , n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , n57197 , n57198 , n57199 , 
     n57200 , n57201 , n57202 , n57203 , n57204 , n57205 , n584529 , n584530 , n57208 , n584532 , 
     n57210 , n57211 , n57212 , n57213 , n57214 , n57215 , n57216 , n584540 , n57218 , n57219 , 
     n57220 , n584544 , n57222 , n57223 , n57224 , n57225 , n584549 , n584550 , n57228 , n584552 , 
     n584553 , n57231 , n584555 , n584556 , n57234 , n57235 , n584559 , n584560 , n57238 , n57239 , 
     n584563 , n57241 , n57242 , n584566 , n57244 , n584568 , n584569 , n57247 , n57248 , n57249 , 
     n57250 , n57251 , n57252 , n57253 , n57254 , n57255 , n57256 , n57257 , n57258 , n57259 , 
     n57260 , n584584 , n584585 , n57263 , n584587 , n584588 , n57266 , n584590 , n584591 , n57269 , 
     n57270 , n584594 , n584595 , n57273 , n57274 , n584598 , n57276 , n57277 , n57278 , n57279 , 
     n57280 , n57281 , n57282 , n57283 , n57284 , n57285 , n57286 , n57287 , n57288 , n57289 , 
     n57290 , n57291 , n57292 , n57293 , n57294 , n57295 , n57296 , n57297 , n57298 , n57299 , 
     n57300 , n57301 , n584625 , n584626 , n57304 , n584628 , n57306 , n57307 , n57308 , n584632 , 
     n584633 , n57311 , n584635 , n57313 , n57314 , n57315 , n584639 , n57317 , n584641 , n584642 , 
     n57320 , n584644 , n584645 , n57323 , n57324 , n584648 , n584649 , n57327 , n57328 , n584652 , 
     n584653 , n57331 , n57332 , n57333 , n584657 , n57335 , n584659 , n57337 , n584661 , n57339 , 
     n584663 , n57341 , n57342 , n57343 , n584667 , n57345 , n584669 , n57347 , n584671 , n57349 , 
     n584673 , n57351 , n584675 , n57353 , n57354 , n57355 , n57356 , n584680 , n57358 , n584682 , 
     n57360 , n584684 , n57362 , n57363 , n57364 , n57365 , n584689 , n57367 , n57368 , n584692 , 
     n57370 , n57371 , n57372 , n57373 , n584697 , n584698 , n584699 , n57377 , n584701 , n57379 , 
     n584703 , n584704 , n584705 , n584706 , n57384 , n584708 , n57386 , n57387 , n584711 , n57389 , 
     n57390 , n57391 , n57392 , n584716 , n57394 , n584718 , n584719 , n57397 , n57398 , n57399 , 
     n57400 , n57401 , n57402 , n57403 , n57404 , n57405 , n584729 , n57407 , n57408 , n584732 , 
     n584733 , n57411 , n584735 , n584736 , n57414 , n584738 , n584739 , n57417 , n57418 , n584742 , 
     n584743 , n57421 , n57422 , n57423 , n57424 , n57425 , n584749 , n584750 , n57428 , n584752 , 
     n57430 , n57431 , n57432 , n57433 , n584757 , n57435 , n584759 , n584760 , n57438 , n584762 , 
     n584763 , n57441 , n57442 , n584766 , n584767 , n57445 , n57446 , n584770 , n57448 , n584772 , 
     n584773 , n57451 , n584775 , n57453 , n584777 , n57455 , n57456 , n57457 , n584781 , n584782 , 
     n57460 , n57461 , n584785 , n584786 , n57464 , n57465 , n584789 , n57467 , n57468 , n57469 , 
     n57470 , n584794 , n57472 , n584796 , n584797 , n57475 , n584799 , n57477 , n57478 , n584802 , 
     n57480 , n584804 , n57482 , n584806 , n57484 , n57485 , n584809 , n57487 , n584811 , n57489 , 
     n584813 , n57491 , n57492 , n584816 , n584817 , n57495 , n584819 , n57497 , n57498 , n584822 , 
     n584823 , n584824 , n57502 , n584826 , n584827 , n57505 , n57506 , n57507 , n57508 , n57509 , 
     n57510 , n57511 , n584835 , n57513 , n57514 , n584838 , n584839 , n57517 , n584841 , n584842 , 
     n57520 , n584844 , n584845 , n57523 , n584847 , n57525 , n57526 , n57527 , n57528 , n57529 , 
     n57530 , n57531 , n57532 , n584856 , n584857 , n584858 , n57536 , n584860 , n584861 , n584862 , 
     n584863 , n57541 , n584865 , n584866 , n57544 , n584868 , n584869 , n57547 , n584871 , n584872 , 
     n57550 , n584874 , n584875 , n584876 , n57554 , n584878 , n584879 , n584880 , n584881 , n57559 , 
     n584883 , n584884 , n57562 , n584886 , n584887 , n57565 , n584889 , n584890 , n57568 , n584892 , 
     n57570 , n584894 , n584895 , n57573 , n584897 , n584898 , n584899 , n584900 , n57578 , n584902 , 
     n584903 , n57581 , n57582 , n57583 , n57584 , n57585 , n584909 , n584910 , n57588 , n584912 , 
     n57590 , n584914 , n57592 , n584916 , n584917 , n57595 , n584919 , n584920 , n584921 , n57599 , 
     n584923 , n57601 , n584925 , n584926 , n57604 , n584928 , n57606 , n584930 , n57608 , n57609 , 
     n57610 , n57611 , n584935 , n57613 , n57614 , n57615 , n57616 , n57617 , n57618 , n57619 , 
     n57620 , n57621 , n57622 , n57623 , n584947 , n57625 , n584949 , n584950 , n57628 , n584952 , 
     n57630 , n57631 , n57632 , n57633 , n57634 , n57635 , n57636 , n57637 , n57638 , n57639 , 
     n57640 , n584964 , n57642 , n584966 , n57644 , n57645 , n57646 , n57647 , n57648 , n57649 , 
     n57650 , n57651 , n57652 , n57653 , n57654 , n57655 , n57656 , n57657 , n57658 , n57659 , 
     n57660 , n57661 , n584985 , n57663 , n57664 , n57665 , n57666 , n57667 , n584991 , n57669 , 
     n57670 , n57671 , n57672 , n57673 , n57674 , n57675 , n57676 , n57677 , n57678 , n57679 , 
     n57680 , n57681 , n57682 , n57683 , n57684 , n57685 , n57686 , n57687 , n57688 , n57689 , 
     n57690 , n57691 , n57692 , n57693 , n57694 , n57695 , n57696 , n57697 , n585021 , n585022 , 
     n585023 , n57701 , n585025 , n585026 , n57704 , n57705 , n57706 , n57707 , n585031 , n57709 , 
     n585033 , n57711 , n585035 , n57713 , n585037 , n585038 , n57716 , n585040 , n585041 , n585042 , 
     n57720 , n585044 , n585045 , n57723 , n585047 , n57725 , n57726 , n57727 , n585051 , n57729 , 
     n585053 , n585054 , n57732 , n57733 , n57734 , n57735 , n585059 , n585060 , n57738 , n585062 , 
     n57740 , n57741 , n57742 , n57743 , n57744 , n57745 , n57746 , n57747 , n57748 , n57749 , 
     n57750 , n57751 , n57752 , n57753 , n57754 , n57755 , n57756 , n57757 , n57758 , n57759 , 
     n57760 , n57761 , n57762 , n585086 , n57764 , n57765 , n57766 , n57767 , n57768 , n585092 , 
     n57770 , n57771 , n585095 , n57773 , n57774 , n57775 , n57776 , n585100 , n585101 , n57779 , 
     n57780 , n57781 , n57782 , n57783 , n57784 , n585108 , n57786 , n57787 , n585111 , n57789 , 
     n57790 , n57791 , n57792 , n57793 , n585117 , n57795 , n57796 , n585120 , n585121 , n57799 , 
     n57800 , n585124 , n57802 , n57803 , n57804 , n57805 , n57806 , n585130 , n57808 , n57809 , 
     n57810 , n57811 , n57812 , n57813 , n585137 , n585138 , n585139 , n57817 , n585141 , n585142 , 
     n57820 , n585144 , n585145 , n57823 , n585147 , n585148 , n57826 , n57827 , n585151 , n585152 , 
     n57830 , n585154 , n585155 , n57833 , n585157 , n585158 , n57836 , n585160 , n585161 , n57839 , 
     n585163 , n585164 , n585165 , n585166 , n57844 , n585168 , n585169 , n585170 , n585171 , n57849 , 
     n585173 , n585174 , n57852 , n585176 , n585177 , n57855 , n585179 , n57857 , n585181 , n57859 , 
     n57860 , n585184 , n585185 , n57863 , n585187 , n585188 , n57866 , n585190 , n585191 , n57869 , 
     n585193 , n585194 , n57872 , n585196 , n585197 , n57875 , n585199 , n585200 , n585201 , n57879 , 
     n585203 , n585204 , n57882 , n585206 , n57884 , n585208 , n585209 , n57887 , n57888 , n585212 , 
     n585213 , n57891 , n585215 , n585216 , n57894 , n585218 , n585219 , n57897 , n585221 , n585222 , 
     n57900 , n585224 , n585225 , n585226 , n57904 , n585228 , n585229 , n57907 , n585231 , n585232 , 
     n57910 , n57911 , n585235 , n57913 , n585237 , n585238 , n57916 , n57917 , n585241 , n585242 , 
     n57920 , n57921 , n57922 , n585246 , n585247 , n57925 , n57926 , n57927 , n57928 , n57929 , 
     n585253 , n57931 , n57932 , n57933 , n585257 , n57935 , n585259 , n585260 , n57938 , n585262 , 
     n57940 , n57941 , n57942 , n585266 , n57944 , n585268 , n585269 , n57947 , n585271 , n57949 , 
     n585273 , n585274 , n57952 , n585276 , n585277 , n57955 , n57956 , n585280 , n585281 , n57959 , 
     n57960 , n585284 , n585285 , n585286 , n57964 , n585288 , n585289 , n57967 , n585291 , n585292 , 
     n57970 , n57971 , n585295 , n585296 , n57974 , n57975 , n585299 , n585300 , n57978 , n585302 , 
     n57980 , n585304 , n585305 , n57983 , n585307 , n585308 , n57986 , n57987 , n585311 , n585312 , 
     n57990 , n57991 , n585315 , n585316 , n57994 , n57995 , n57996 , n585320 , n57998 , n57999 , 
     n58000 , n585324 , n585325 , n58003 , n585327 , n58005 , n58006 , n58007 , n58008 , n58009 , 
     n58010 , n58011 , n58012 , n58013 , n58014 , n58015 , n58016 , n58017 , n58018 , n58019 , 
     n585343 , n585344 , n58022 , n585346 , n585347 , n58025 , n585349 , n585350 , n58028 , n585352 , 
     n585353 , n58031 , n58032 , n585356 , n585357 , n58035 , n585359 , n585360 , n58038 , n585362 , 
     n585363 , n58041 , n585365 , n585366 , n58044 , n585368 , n585369 , n585370 , n585371 , n58049 , 
     n585373 , n585374 , n585375 , n585376 , n58054 , n585378 , n585379 , n58057 , n585381 , n585382 , 
     n58060 , n585384 , n58062 , n585386 , n58064 , n58065 , n585389 , n585390 , n58068 , n585392 , 
     n585393 , n58071 , n585395 , n585396 , n58074 , n585398 , n585399 , n58077 , n585401 , n585402 , 
     n58080 , n585404 , n585405 , n58083 , n585407 , n585408 , n58086 , n585410 , n585411 , n58089 , 
     n58090 , n585414 , n585415 , n58093 , n585417 , n585418 , n58096 , n585420 , n585421 , n58099 , 
     n585423 , n585424 , n58102 , n585426 , n585427 , n58105 , n58106 , n58107 , n585431 , n585432 , 
     n58110 , n58111 , n585435 , n585436 , n58114 , n585438 , n585439 , n58117 , n58118 , n58119 , 
     n58120 , n58121 , n58122 , n58123 , n58124 , n58125 , n585449 , n585450 , n58128 , n585452 , 
     n58130 , n585454 , n585455 , n58133 , n585457 , n58135 , n58136 , n585460 , n585461 , n58139 , 
     n585463 , n585464 , n58142 , n585466 , n585467 , n58145 , n585469 , n58147 , n58148 , n58149 , 
     n58150 , n585474 , n58152 , n58153 , n585477 , n58155 , n585479 , n58157 , n585481 , n585482 , 
     n58160 , n585484 , n585485 , n58163 , n585487 , n58165 , n58166 , n58167 , n58168 , n58169 , 
     n58170 , n58171 , n58172 , n58173 , n585497 , n58175 , n585499 , n58177 , n58178 , n58179 , 
     n585503 , n585504 , n58182 , n585506 , n58184 , n585508 , n58186 , n585510 , n585511 , n58189 , 
     n58190 , n585514 , n585515 , n58193 , n58194 , n58195 , n58196 , n58197 , n58198 , n58199 , 
     n58200 , n58201 , n58202 , n58203 , n58204 , n58205 , n58206 , n58207 , n585531 , n58209 , 
     n585533 , n585534 , n58212 , n58213 , n58214 , n585538 , n58216 , n58217 , n58218 , n58219 , 
     n58220 , n58221 , n58222 , n585546 , n58224 , n585548 , n58226 , n58227 , n585551 , n58229 , 
     n585553 , n585554 , n585555 , n58233 , n585557 , n58235 , n58236 , n585560 , n58238 , n585562 , 
     n58240 , n58241 , n58242 , n58243 , n58244 , n58245 , n58246 , n58247 , n58248 , n58249 , 
     n58250 , n58251 , n58252 , n58253 , n58254 , n585578 , n58256 , n585580 , n58258 , n585582 , 
     n58260 , n585584 , n58262 , n585586 , n58264 , n585588 , n585589 , n58267 , n585591 , n58269 , 
     n585593 , n585594 , n58272 , n58273 , n58274 , n58275 , n585599 , n58277 , n585601 , n58279 , 
     n58280 , n58281 , n58282 , n585606 , n58284 , n58285 , n585609 , n58287 , n58288 , n585612 , 
     n58290 , n585614 , n585615 , n58293 , n585617 , n585618 , n58296 , n58297 , n585621 , n58299 , 
     n58300 , n58301 , n58302 , n585626 , n58304 , n58305 , n58306 , n58307 , n585631 , n585632 , 
     n585633 , n58311 , n585635 , n585636 , n58314 , n585638 , n58316 , n58317 , n585641 , n585642 , 
     n58320 , n585644 , n585645 , n58323 , n585647 , n585648 , n58326 , n58327 , n58328 , n58329 , 
     n585653 , n58331 , n58332 , n58333 , n58334 , n585658 , n585659 , n58337 , n585661 , n585662 , 
     n58340 , n585664 , n585665 , n585666 , n58344 , n585668 , n58346 , n58347 , n58348 , n58349 , 
     n58350 , n58351 , n58352 , n58353 , n58354 , n58355 , n58356 , n58357 , n58358 , n58359 , 
     n58360 , n58361 , n58362 , n58363 , n58364 , n58365 , n58366 , n58367 , n58368 , n58369 , 
     n58370 , n58371 , n58372 , n58373 , n58374 , n58375 , n58376 , n585700 , n58378 , n585702 , 
     n585703 , n585704 , n585705 , n58383 , n585707 , n58385 , n585709 , n58387 , n585711 , n58389 , 
     n58390 , n58391 , n58392 , n58393 , n58394 , n58395 , n58396 , n585720 , n585721 , n58399 , 
     n58400 , n58401 , n58402 , n585726 , n585727 , n58405 , n585729 , n585730 , n58408 , n585732 , 
     n585733 , n585734 , n585735 , n58413 , n585737 , n585738 , n58416 , n585740 , n585741 , n58419 , 
     n585743 , n585744 , n58422 , n585746 , n585747 , n58425 , n585749 , n585750 , n585751 , n585752 , 
     n58430 , n585754 , n585755 , n585756 , n58434 , n585758 , n58436 , n585760 , n585761 , n58439 , 
     n585763 , n58441 , n585765 , n585766 , n58444 , n585768 , n585769 , n585770 , n585771 , n58449 , 
     n585773 , n585774 , n58452 , n585776 , n585777 , n58455 , n585779 , n585780 , n58458 , n585782 , 
     n585783 , n585784 , n58462 , n585786 , n585787 , n585788 , n585789 , n58467 , n585791 , n585792 , 
     n58470 , n585794 , n585795 , n58473 , n585797 , n585798 , n58476 , n585800 , n58478 , n58479 , 
     n585803 , n58481 , n585805 , n58483 , n58484 , n58485 , n58486 , n58487 , n585811 , n58489 , 
     n58490 , n585814 , n58492 , n585816 , n585817 , n585818 , n585819 , n58497 , n585821 , n585822 , 
     n58500 , n585824 , n585825 , n58503 , n585827 , n58505 , n58506 , n585830 , n58508 , n585832 , 
     n58510 , n58511 , n585835 , n58513 , n585837 , n585838 , n58516 , n585840 , n58518 , n585842 , 
     n58520 , n58521 , n585845 , n58523 , n585847 , n585848 , n58526 , n585850 , n585851 , n585852 , 
     n585853 , n58531 , n585855 , n585856 , n58534 , n585858 , n585859 , n58537 , n585861 , n585862 , 
     n58540 , n58541 , n585865 , n585866 , n58544 , n585868 , n585869 , n58547 , n585871 , n585872 , 
     n585873 , n58551 , n585875 , n585876 , n585877 , n58555 , n585879 , n585880 , n58558 , n585882 , 
     n58560 , n58561 , n585885 , n58563 , n585887 , n58565 , n585889 , n585890 , n58568 , n585892 , 
     n585893 , n58571 , n58572 , n585896 , n58574 , n58575 , n58576 , n58577 , n585901 , n58579 , 
     n58580 , n585904 , n585905 , n585906 , n58584 , n585908 , n585909 , n585910 , n58588 , n585912 , 
     n585913 , n58591 , n585915 , n58593 , n58594 , n58595 , n58596 , n585920 , n58598 , n585922 , 
     n585923 , n58601 , n58602 , n585926 , n585927 , n58605 , n58606 , n585930 , n58608 , n58609 , 
     n58610 , n58611 , n585935 , n585936 , n585937 , n58615 , n585939 , n585940 , n585941 , n585942 , 
     n58620 , n585944 , n585945 , n58623 , n585947 , n585948 , n58626 , n585950 , n585951 , n58629 , 
     n585953 , n585954 , n58632 , n585956 , n585957 , n58635 , n585959 , n585960 , n585961 , n585962 , 
     n58640 , n585964 , n585965 , n58643 , n585967 , n585968 , n58646 , n585970 , n585971 , n58649 , 
     n585973 , n585974 , n585975 , n585976 , n58654 , n585978 , n585979 , n585980 , n585981 , n58659 , 
     n585983 , n585984 , n58662 , n585986 , n585987 , n58665 , n585989 , n585990 , n58668 , n58669 , 
     n58670 , n585994 , n585995 , n58673 , n585997 , n585998 , n58676 , n58677 , n586001 , n586002 , 
     n58680 , n58681 , n586005 , n586006 , n586007 , n586008 , n58686 , n586010 , n586011 , n58689 , 
     n586013 , n586014 , n58692 , n586016 , n586017 , n58695 , n58696 , n586020 , n586021 , n58699 , 
     n58700 , n586024 , n586025 , n58703 , n58704 , n58705 , n58706 , n58707 , n58708 , n58709 , 
     n58710 , n586034 , n58712 , n586036 , n586037 , n58715 , n58716 , n586040 , n58718 , n586042 , 
     n58720 , n586044 , n586045 , n58723 , n586047 , n58725 , n58726 , n586050 , n58728 , n586052 , 
     n586053 , n58731 , n586055 , n586056 , n58734 , n586058 , n586059 , n58737 , n58738 , n586062 , 
     n586063 , n58741 , n58742 , n586066 , n586067 , n58745 , n58746 , n586070 , n58748 , n58749 , 
     n586073 , n586074 , n58752 , n58753 , n586077 , n586078 , n58756 , n58757 , n586081 , n586082 , 
     n58760 , n586084 , n58762 , n58763 , n586087 , n586088 , n58766 , n586090 , n58768 , n586092 , 
     n58770 , n58771 , n58772 , n58773 , n58774 , n58775 , n58776 , n58777 , n58778 , n58779 , 
     n58780 , n58781 , n58782 , n58783 , n58784 , n58785 , n58786 , n58787 , n58788 , n58789 , 
     n58790 , n58791 , n58792 , n58793 , n586117 , n58795 , n586119 , n586120 , n586121 , n58799 , 
     n586123 , n586124 , n586125 , n58803 , n586127 , n586128 , n586129 , n58807 , n586131 , n586132 , 
     n58810 , n586134 , n58812 , n586136 , n586137 , n58815 , n586139 , n586140 , n58818 , n586142 , 
     n586143 , n58821 , n58822 , n58823 , n586147 , n586148 , n586149 , n58827 , n586151 , n586152 , 
     n586153 , n58831 , n586155 , n58833 , n586157 , n586158 , n58836 , n586160 , n586161 , n58839 , 
     n586163 , n586164 , n58842 , n58843 , n58844 , n586168 , n58846 , n58847 , n58848 , n58849 , 
     n58850 , n58851 , n58852 , n58853 , n58854 , n586178 , n586179 , n58857 , n586181 , n58859 , 
     n58860 , n58861 , n58862 , n58863 , n586187 , n586188 , n58866 , n586190 , n586191 , n58869 , 
     n586193 , n586194 , n58872 , n586196 , n586197 , n586198 , n586199 , n58877 , n586201 , n586202 , 
     n58880 , n586204 , n586205 , n58883 , n58884 , n586208 , n586209 , n58887 , n58888 , n586212 , 
     n586213 , n586214 , n58892 , n586216 , n586217 , n586218 , n58896 , n586220 , n586221 , n58899 , 
     n586223 , n586224 , n586225 , n586226 , n58904 , n586228 , n586229 , n58907 , n586231 , n586232 , 
     n58910 , n586234 , n586235 , n58913 , n58914 , n58915 , n586239 , n586240 , n58918 , n586242 , 
     n586243 , n58921 , n586245 , n586246 , n58924 , n586248 , n586249 , n58927 , n586251 , n586252 , 
     n586253 , n586254 , n58932 , n586256 , n586257 , n58935 , n586259 , n586260 , n58938 , n58939 , 
     n586263 , n586264 , n58942 , n58943 , n586267 , n586268 , n58946 , n58947 , n58948 , n586272 , 
     n58950 , n58951 , n58952 , n586276 , n586277 , n58955 , n586279 , n586280 , n586281 , n58959 , 
     n586283 , n58961 , n58962 , n58963 , n58964 , n58965 , n58966 , n586290 , n586291 , n58969 , 
     n586293 , n58971 , n586295 , n58973 , n58974 , n586298 , n58976 , n586300 , n586301 , n58979 , 
     n586303 , n586304 , n586305 , n586306 , n58984 , n586308 , n586309 , n58987 , n586311 , n586312 , 
     n58990 , n586314 , n586315 , n58993 , n58994 , n586318 , n586319 , n58997 , n586321 , n586322 , 
     n59000 , n586324 , n586325 , n59003 , n586327 , n586328 , n59006 , n586330 , n586331 , n59009 , 
     n586333 , n59011 , n59012 , n59013 , n59014 , n59015 , n59016 , n59017 , n59018 , n59019 , 
     n586343 , n586344 , n586345 , n59023 , n586347 , n586348 , n586349 , n586350 , n59028 , n586352 , 
     n586353 , n59031 , n586355 , n586356 , n59034 , n586358 , n586359 , n59037 , n586361 , n586362 , 
     n586363 , n586364 , n59042 , n586366 , n586367 , n59045 , n586369 , n586370 , n59048 , n586372 , 
     n586373 , n59051 , n59052 , n59053 , n586377 , n586378 , n59056 , n59057 , n586381 , n586382 , 
     n59060 , n59061 , n586385 , n586386 , n586387 , n586388 , n59066 , n586390 , n59068 , n59069 , 
     n59070 , n586394 , n586395 , n59073 , n586397 , n59075 , n586399 , n59077 , n59078 , n59079 , 
     n59080 , n59081 , n586405 , n586406 , n59084 , n586408 , n59086 , n59087 , n586411 , n59089 , 
     n586413 , n59091 , n59092 , n586416 , n586417 , n59095 , n586419 , n59097 , n586421 , n586422 , 
     n59100 , n586424 , n59102 , n59103 , n59104 , n59105 , n59106 , n59107 , n59108 , n59109 , 
     n59110 , n59111 , n59112 , n59113 , n59114 , n586438 , n59116 , n586440 , n586441 , n59119 , 
     n586443 , n586444 , n59122 , n586446 , n586447 , n586448 , n586449 , n59127 , n586451 , n586452 , 
     n59130 , n586454 , n586455 , n59133 , n586457 , n586458 , n59136 , n586460 , n586461 , n586462 , 
     n586463 , n59141 , n586465 , n586466 , n586467 , n586468 , n59146 , n586470 , n586471 , n59149 , 
     n586473 , n586474 , n59152 , n586476 , n586477 , n59155 , n586479 , n586480 , n59158 , n59159 , 
     n59160 , n586484 , n586485 , n59163 , n59164 , n59165 , n586489 , n586490 , n59168 , n586492 , 
     n586493 , n59171 , n59172 , n59173 , n59174 , n586498 , n59176 , n59177 , n59178 , n59179 , 
     n586503 , n59181 , n59182 , n59183 , n59184 , n59185 , n59186 , n59187 , n59188 , n59189 , 
     n59190 , n586514 , n59192 , n586516 , n586517 , n59195 , n586519 , n586520 , n59198 , n586522 , 
     n59200 , n59201 , n586525 , n59203 , n586527 , n59205 , n586529 , n59207 , n586531 , n586532 , 
     n59210 , n59211 , n59212 , n586536 , n586537 , n586538 , n586539 , n59217 , n586541 , n59219 , 
     n586543 , n59221 , n59222 , n586546 , n59224 , n586548 , n586549 , n59227 , n586551 , n586552 , 
     n59230 , n586554 , n586555 , n59233 , n586557 , n586558 , n59236 , n586560 , n586561 , n59239 , 
     n586563 , n586564 , n586565 , n586566 , n59244 , n586568 , n586569 , n59247 , n586571 , n586572 , 
     n59250 , n59251 , n586575 , n586576 , n59254 , n59255 , n586579 , n586580 , n59258 , n59259 , 
     n586583 , n586584 , n59262 , n59263 , n586587 , n586588 , n586589 , n59267 , n586591 , n59269 , 
     n59270 , n59271 , n59272 , n586596 , n59274 , n59275 , n586599 , n59277 , n586601 , n586602 , 
     n59280 , n59281 , n586605 , n586606 , n59284 , n59285 , n59286 , n59287 , n586611 , n586612 , 
     n59290 , n59291 , n59292 , n59293 , n59294 , n586618 , n586619 , n59297 , n586621 , n586622 , 
     n59300 , n59301 , n586625 , n59303 , n59304 , n59305 , n59306 , n586630 , n59308 , n59309 , 
     n59310 , n59311 , n59312 , n59313 , n59314 , n59315 , n59316 , n586640 , n59318 , n586642 , 
     n59320 , n586644 , n59322 , n59323 , n586647 , n59325 , n586649 , n586650 , n59328 , n586652 , 
     n586653 , n59331 , n59332 , n586656 , n586657 , n59335 , n59336 , n586660 , n59338 , n586662 , 
     n586663 , n59341 , n586665 , n586666 , n59344 , n586668 , n586669 , n59347 , n586671 , n586672 , 
     n59350 , n59351 , n586675 , n586676 , n59354 , n586678 , n586679 , n59357 , n586681 , n586682 , 
     n59360 , n586684 , n586685 , n59363 , n586687 , n586688 , n586689 , n586690 , n59368 , n586692 , 
     n586693 , n586694 , n586695 , n59373 , n586697 , n586698 , n59376 , n586700 , n586701 , n59379 , 
     n586703 , n586704 , n59382 , n59383 , n586707 , n59385 , n59386 , n59387 , n59388 , n59389 , 
     n59390 , n59391 , n59392 , n59393 , n59394 , n59395 , n59396 , n59397 , n59398 , n586722 , 
     n59400 , n586724 , n59402 , n586726 , n59404 , n59405 , n586729 , n586730 , n59408 , n59409 , 
     n59410 , n59411 , n59412 , n59413 , n586737 , n59415 , n586739 , n59417 , n59418 , n59419 , 
     n59420 , n59421 , n59422 , n59423 , n586747 , n586748 , n59426 , n586750 , n586751 , n586752 , 
     n586753 , n59431 , n586755 , n586756 , n59434 , n586758 , n59436 , n586760 , n59438 , n59439 , 
     n586763 , n586764 , n59442 , n586766 , n586767 , n59445 , n586769 , n586770 , n59448 , n586772 , 
     n586773 , n586774 , n59452 , n586776 , n586777 , n59455 , n586779 , n586780 , n59458 , n586782 , 
     n586783 , n59461 , n59462 , n586786 , n586787 , n59465 , n586789 , n586790 , n59468 , n586792 , 
     n586793 , n59471 , n586795 , n586796 , n59474 , n586798 , n59476 , n59477 , n59478 , n59479 , 
     n59480 , n59481 , n59482 , n59483 , n586807 , n59485 , n586809 , n586810 , n586811 , n59489 , 
     n586813 , n59491 , n59492 , n59493 , n59494 , n59495 , n59496 , n59497 , n586821 , n59499 , 
     n59500 , n586824 , n59502 , n59503 , n59504 , n586828 , n59506 , n59507 , n59508 , n586832 , 
     n586833 , n59511 , n586835 , n586836 , n586837 , n59515 , n586839 , n59517 , n59518 , n59519 , 
     n59520 , n59521 , n59522 , n59523 , n59524 , n59525 , n59526 , n586850 , n59528 , n59529 , 
     n586853 , n59531 , n586855 , n59533 , n586857 , n59535 , n586859 , n586860 , n59538 , n586862 , 
     n59540 , n586864 , n586865 , n59543 , n586867 , n586868 , n59546 , n59547 , n586871 , n59549 , 
     n586873 , n59551 , n586875 , n586876 , n59554 , n586878 , n586879 , n59557 , n59558 , n586882 , 
     n59560 , n59561 , n59562 , n59563 , n586887 , n586888 , n59566 , n586890 , n59568 , n586892 , 
     n59570 , n59571 , n586895 , n586896 , n59574 , n59575 , n586899 , n586900 , n59578 , n59579 , 
     n586903 , n586904 , n59582 , n59583 , n586907 , n586908 , n59586 , n59587 , n586911 , n59589 , 
     n59590 , n59591 , n59592 , n586916 , n586917 , n59595 , n586919 , n586920 , n59598 , n59599 , 
     n586923 , n59601 , n59602 , n586926 , n586927 , n586928 , n59606 , n586930 , n586931 , n586932 , 
     n59610 , n586934 , n586935 , n59613 , n586937 , n586938 , n59616 , n59617 , n59618 , n59619 , 
     n586943 , n586944 , n59622 , n586946 , n586947 , n586948 , n59626 , n586950 , n586951 , n586952 , 
     n59630 , n59631 , n586955 , n59633 , n59634 , n59635 , n59636 , n59637 , n59638 , n59639 , 
     n59640 , n59641 , n59642 , n59643 , n59644 , n59645 , n59646 , n586970 , n59648 , n586972 , 
     n59650 , n59651 , n586975 , n586976 , n59654 , n59655 , n586979 , n59657 , n59658 , n59659 , 
     n59660 , n59661 , n59662 , n586986 , n586987 , n59665 , n586989 , n586990 , n59668 , n586992 , 
     n586993 , n59671 , n586995 , n586996 , n59674 , n59675 , n586999 , n587000 , n59678 , n587002 , 
     n587003 , n59681 , n587005 , n587006 , n59684 , n587008 , n587009 , n59687 , n587011 , n587012 , 
     n587013 , n587014 , n59692 , n587016 , n587017 , n59695 , n587019 , n587020 , n59698 , n587022 , 
     n587023 , n59701 , n59702 , n587026 , n587027 , n59705 , n587029 , n587030 , n59708 , n587032 , 
     n587033 , n59711 , n587035 , n587036 , n59714 , n587038 , n587039 , n59717 , n587041 , n587042 , 
     n59720 , n587044 , n587045 , n59723 , n587047 , n587048 , n59726 , n587050 , n587051 , n59729 , 
     n59730 , n587054 , n587055 , n59733 , n587057 , n587058 , n59736 , n587060 , n587061 , n59739 , 
     n587063 , n587064 , n59742 , n587066 , n587067 , n59745 , n59746 , n59747 , n587071 , n587072 , 
     n59750 , n587074 , n587075 , n59753 , n59754 , n587078 , n587079 , n59757 , n587081 , n587082 , 
     n59760 , n587084 , n59762 , n587086 , n587087 , n59765 , n587089 , n587090 , n59768 , n59769 , 
     n587093 , n587094 , n59772 , n59773 , n587097 , n587098 , n587099 , n59777 , n587101 , n587102 , 
     n59780 , n587104 , n587105 , n59783 , n59784 , n587108 , n587109 , n59787 , n59788 , n587112 , 
     n587113 , n59791 , n587115 , n587116 , n59794 , n587118 , n587119 , n59797 , n59798 , n59799 , 
     n59800 , n59801 , n587125 , n59803 , n59804 , n587128 , n587129 , n59807 , n587131 , n587132 , 
     n59810 , n587134 , n587135 , n587136 , n59814 , n587138 , n59816 , n587140 , n587141 , n59819 , 
     n587143 , n587144 , n59822 , n587146 , n587147 , n59825 , n59826 , n59827 , n587151 , n587152 , 
     n59830 , n59831 , n59832 , n587156 , n59834 , n59835 , n59836 , n59837 , n59838 , n59839 , 
     n59840 , n59841 , n59842 , n59843 , n59844 , n59845 , n59846 , n59847 , n59848 , n59849 , 
     n59850 , n587174 , n587175 , n587176 , n59854 , n587178 , n587179 , n59857 , n587181 , n587182 , 
     n59860 , n59861 , n587185 , n587186 , n59864 , n59865 , n587189 , n587190 , n587191 , n59869 , 
     n587193 , n587194 , n59872 , n587196 , n587197 , n59875 , n59876 , n587200 , n587201 , n59879 , 
     n59880 , n587204 , n587205 , n59883 , n59884 , n59885 , n587209 , n59887 , n59888 , n59889 , 
     n587213 , n587214 , n59892 , n587216 , n587217 , n59895 , n587219 , n59897 , n587221 , n587222 , 
     n59900 , n59901 , n59902 , n587226 , n59904 , n59905 , n59906 , n59907 , n59908 , n587232 , 
     n59910 , n587234 , n59912 , n587236 , n59914 , n59915 , n587239 , n587240 , n59918 , n587242 , 
     n587243 , n59921 , n59922 , n587246 , n587247 , n59925 , n587249 , n587250 , n587251 , n587252 , 
     n59930 , n587254 , n587255 , n59933 , n587257 , n59935 , n587259 , n59937 , n59938 , n587262 , 
     n587263 , n59941 , n587265 , n587266 , n59944 , n587268 , n587269 , n59947 , n587271 , n59949 , 
     n587273 , n587274 , n59952 , n587276 , n587277 , n587278 , n59956 , n587280 , n587281 , n587282 , 
     n59960 , n587284 , n587285 , n59963 , n587287 , n587288 , n59966 , n587290 , n587291 , n59969 , 
     n59970 , n59971 , n587295 , n59973 , n59974 , n59975 , n59976 , n59977 , n59978 , n59979 , 
     n59980 , n59981 , n59982 , n59983 , n59984 , n59985 , n587309 , n59987 , n587311 , n587312 , 
     n59990 , n587314 , n587315 , n587316 , n587317 , n59995 , n587319 , n587320 , n59998 , n587322 , 
     n60000 , n587324 , n60002 , n60003 , n587327 , n587328 , n60006 , n587330 , n587331 , n60009 , 
     n587333 , n587334 , n60012 , n587336 , n587337 , n587338 , n587339 , n60017 , n587341 , n587342 , 
     n587343 , n587344 , n60022 , n587346 , n587347 , n60025 , n587349 , n60027 , n587351 , n60029 , 
     n60030 , n587354 , n587355 , n60033 , n587357 , n587358 , n60036 , n587360 , n587361 , n60039 , 
     n587363 , n587364 , n60042 , n60043 , n587367 , n60045 , n60046 , n60047 , n587371 , n587372 , 
     n60050 , n60051 , n60052 , n587376 , n587377 , n60055 , n60056 , n587380 , n587381 , n60059 , 
     n587383 , n60061 , n587385 , n587386 , n60064 , n587388 , n587389 , n60067 , n60068 , n587392 , 
     n587393 , n60071 , n60072 , n587396 , n587397 , n587398 , n60076 , n587400 , n587401 , n60079 , 
     n587403 , n587404 , n60082 , n60083 , n587407 , n587408 , n60086 , n60087 , n587411 , n587412 , 
     n60090 , n587414 , n60092 , n587416 , n587417 , n60095 , n587419 , n587420 , n60098 , n60099 , 
     n587423 , n587424 , n60102 , n60103 , n587427 , n587428 , n60106 , n60107 , n60108 , n587432 , 
     n587433 , n60111 , n60112 , n587436 , n587437 , n60115 , n60116 , n60117 , n587441 , n587442 , 
     n60120 , n60121 , n60122 , n587446 , n587447 , n60125 , n60126 , n60127 , n587451 , n587452 , 
     n60130 , n60131 , n587455 , n60133 , n60134 , n60135 , n60136 , n60137 , n60138 , n60139 , 
     n60140 , n60141 , n60142 , n587466 , n60144 , n60145 , n587469 , n60147 , n60148 , n60149 , 
     n60150 , n587474 , n587475 , n60153 , n587477 , n60155 , n60156 , n587480 , n587481 , n60159 , 
     n60160 , n587484 , n587485 , n60163 , n587487 , n60165 , n60166 , n587490 , n587491 , n60169 , 
     n60170 , n587494 , n587495 , n60173 , n587497 , n60175 , n587499 , n60177 , n60178 , n587502 , 
     n587503 , n60181 , n60182 , n587506 , n587507 , n60185 , n587509 , n60187 , n60188 , n587512 , 
     n587513 , n60191 , n60192 , n587516 , n587517 , n60195 , n60196 , n587520 , n587521 , n60199 , 
     n60200 , n60201 , n587525 , n587526 , n60204 , n587528 , n587529 , n60207 , n587531 , n587532 , 
     n60210 , n587534 , n587535 , n60213 , n587537 , n587538 , n60216 , n587540 , n587541 , n60219 , 
     n587543 , n60221 , n60222 , n60223 , n60224 , n60225 , n60226 , n60227 , n60228 , n60229 , 
     n60230 , n60231 , n60232 , n60233 , n60234 , n60235 , n587559 , n587560 , n60238 , n587562 , 
     n587563 , n60241 , n587565 , n587566 , n60244 , n587568 , n587569 , n60247 , n60248 , n587572 , 
     n587573 , n60251 , n587575 , n587576 , n60254 , n587578 , n587579 , n60257 , n587581 , n587582 , 
     n60260 , n587584 , n587585 , n60263 , n587587 , n60265 , n60266 , n587590 , n60268 , n60269 , 
     n60270 , n60271 , n60272 , n60273 , n60274 , n60275 , n60276 , n60277 , n60278 , n60279 , 
     n60280 , n60281 , n60282 , n60283 , n60284 , n587608 , n60286 , n60287 , n60288 , n587612 , 
     n587613 , n587614 , n60292 , n587616 , n587617 , n60295 , n587619 , n587620 , n60298 , n587622 , 
     n587623 , n60301 , n60302 , n587626 , n587627 , n60305 , n587629 , n587630 , n60308 , n587632 , 
     n587633 , n60311 , n587635 , n587636 , n60314 , n587638 , n587639 , n587640 , n587641 , n60319 , 
     n587643 , n587644 , n60322 , n587646 , n587647 , n60325 , n587649 , n587650 , n60328 , n60329 , 
     n587653 , n587654 , n60332 , n587656 , n587657 , n60335 , n587659 , n587660 , n60338 , n587662 , 
     n587663 , n60341 , n587665 , n587666 , n60344 , n587668 , n587669 , n60347 , n587671 , n60349 , 
     n587673 , n60351 , n60352 , n587676 , n587677 , n60355 , n60356 , n587680 , n587681 , n60359 , 
     n587683 , n60361 , n60362 , n587686 , n587687 , n60365 , n60366 , n587690 , n587691 , n60369 , 
     n60370 , n60371 , n587695 , n587696 , n60374 , n587698 , n587699 , n60377 , n60378 , n587702 , 
     n587703 , n60381 , n60382 , n60383 , n587707 , n587708 , n60386 , n60387 , n60388 , n587712 , 
     n60390 , n60391 , n60392 , n587716 , n60394 , n60395 , n60396 , n587720 , n60398 , n60399 , 
     n587723 , n587724 , n60402 , n60403 , n587727 , n587728 , n60406 , n60407 , n587731 , n60409 , 
     n60410 , n60411 , n60412 , n587736 , n60414 , n587738 , n60416 , n60417 , n587741 , n60419 , 
     n587743 , n587744 , n60422 , n60423 , n60424 , n60425 , n60426 , n60427 , n60428 , n60429 , 
     n60430 , n60431 , n60432 , n60433 , n60434 , n60435 , n587759 , n60437 , n60438 , n587762 , 
     n60440 , n587764 , n60442 , n587766 , n587767 , n60445 , n587769 , n587770 , n587771 , n60449 , 
     n587773 , n587774 , n587775 , n587776 , n60454 , n587778 , n587779 , n60457 , n587781 , n587782 , 
     n60460 , n587784 , n587785 , n60463 , n60464 , n60465 , n587789 , n587790 , n587791 , n587792 , 
     n60470 , n587794 , n587795 , n587796 , n587797 , n60475 , n587799 , n587800 , n60478 , n587802 , 
     n587803 , n60481 , n587805 , n587806 , n60484 , n60485 , n60486 , n587810 , n587811 , n60489 , 
     n60490 , n587814 , n587815 , n60493 , n587817 , n587818 , n60496 , n587820 , n60498 , n60499 , 
     n60500 , n60501 , n60502 , n60503 , n60504 , n60505 , n60506 , n60507 , n60508 , n60509 , 
     n60510 , n60511 , n60512 , n60513 , n60514 , n587838 , n587839 , n60517 , n587841 , n587842 , 
     n587843 , n60521 , n587845 , n60523 , n587847 , n587848 , n60526 , n587850 , n60528 , n60529 , 
     n60530 , n60531 , n60532 , n60533 , n60534 , n587858 , n587859 , n587860 , n60538 , n587862 , 
     n60540 , n587864 , n60542 , n60543 , n587867 , n60545 , n587869 , n587870 , n60548 , n587872 , 
     n587873 , n60551 , n60552 , n60553 , n60554 , n587878 , n587879 , n60557 , n60558 , n60559 , 
     n587883 , n60561 , n60562 , n60563 , n587887 , n587888 , n60566 , n587890 , n60568 , n60569 , 
     n60570 , n60571 , n60572 , n60573 , n60574 , n60575 , n60576 , n60577 , n60578 , n60579 , 
     n60580 , n60581 , n60582 , n60583 , n60584 , n60585 , n60586 , n60587 , n587911 , n60589 , 
     n60590 , n587914 , n60592 , n60593 , n587917 , n587918 , n60596 , n587920 , n60598 , n60599 , 
     n587923 , n587924 , n60602 , n587926 , n60604 , n587928 , n587929 , n60607 , n587931 , n60609 , 
     n60610 , n587934 , n60612 , n587936 , n60614 , n60615 , n60616 , n60617 , n60618 , n60619 , 
     n587943 , n587944 , n60622 , n587946 , n587947 , n60625 , n587949 , n60627 , n60628 , n60629 , 
     n60630 , n60631 , n60632 , n60633 , n60634 , n60635 , n60636 , n587960 , n587961 , n60639 , 
     n587963 , n587964 , n587965 , n60643 , n587967 , n60645 , n60646 , n60647 , n60648 , n60649 , 
     n60650 , n587974 , n587975 , n60653 , n587977 , n60655 , n587979 , n587980 , n60658 , n587982 , 
     n60660 , n60661 , n60662 , n60663 , n60664 , n60665 , n60666 , n60667 , n60668 , n60669 , 
     n60670 , n587994 , n60672 , n60673 , n60674 , n60675 , n60676 , n60677 , n60678 , n60679 , 
     n60680 , n60681 , n60682 , n60683 , n60684 , n60685 , n60686 , n60687 , n60688 , n60689 , 
     n60690 , n60691 , n60692 , n60693 , n60694 , n60695 , n60696 , n60697 , n60698 , n60699 , 
     n60700 , n60701 , n60702 , n60703 , n60704 , n588028 , n588029 , n60707 , n588031 , n588032 , 
     n588033 , n60711 , n588035 , n60713 , n60714 , n588038 , n588039 , n60717 , n588041 , n60719 , 
     n588043 , n588044 , n60722 , n588046 , n588047 , n60725 , n588049 , n588050 , n60728 , n588052 , 
     n588053 , n60731 , n588055 , n60733 , n588057 , n588058 , n60736 , n60737 , n60738 , n588062 , 
     n60740 , n60741 , n60742 , n588066 , n60744 , n60745 , n588069 , n60747 , n60748 , n60749 , 
     n60750 , n588074 , n588075 , n588076 , n60754 , n588078 , n588079 , n588080 , n588081 , n60759 , 
     n588083 , n588084 , n60762 , n588086 , n588087 , n60765 , n588089 , n588090 , n588091 , n588092 , 
     n60770 , n588094 , n588095 , n60773 , n588097 , n60775 , n588099 , n60777 , n60778 , n588102 , 
     n588103 , n60781 , n588105 , n588106 , n60784 , n588108 , n588109 , n60787 , n588111 , n588112 , 
     n60790 , n588114 , n588115 , n588116 , n588117 , n60795 , n588119 , n588120 , n60798 , n588122 , 
     n588123 , n60801 , n588125 , n588126 , n60804 , n60805 , n588129 , n588130 , n60808 , n60809 , 
     n588133 , n588134 , n60812 , n588136 , n588137 , n60815 , n588139 , n588140 , n60818 , n60819 , 
     n588143 , n588144 , n60822 , n60823 , n588147 , n588148 , n60826 , n588150 , n60828 , n588152 , 
     n588153 , n60831 , n588155 , n60833 , n60834 , n60835 , n60836 , n60837 , n60838 , n60839 , 
     n60840 , n60841 , n60842 , n60843 , n60844 , n60845 , n60846 , n60847 , n60848 , n60849 , 
     n60850 , n60851 , n60852 , n60853 , n60854 , n588178 , n60856 , n60857 , n60858 , n60859 , 
     n60860 , n60861 , n60862 , n588186 , n588187 , n60865 , n588189 , n588190 , n588191 , n588192 , 
     n60870 , n588194 , n588195 , n60873 , n588197 , n588198 , n60876 , n588200 , n588201 , n60879 , 
     n588203 , n588204 , n60882 , n588206 , n588207 , n60885 , n588209 , n588210 , n60888 , n588212 , 
     n60890 , n60891 , n60892 , n60893 , n60894 , n60895 , n60896 , n60897 , n60898 , n60899 , 
     n60900 , n60901 , n60902 , n60903 , n60904 , n60905 , n588229 , n588230 , n60908 , n588232 , 
     n60910 , n588234 , n60912 , n60913 , n588237 , n60915 , n588239 , n588240 , n60918 , n588242 , 
     n588243 , n588244 , n588245 , n60923 , n588247 , n60925 , n588249 , n60927 , n60928 , n588252 , 
     n60930 , n588254 , n588255 , n60933 , n588257 , n588258 , n60936 , n588260 , n588261 , n60939 , 
     n588263 , n588264 , n60942 , n588266 , n60944 , n60945 , n588269 , n588270 , n60948 , n60949 , 
     n588273 , n588274 , n60952 , n60953 , n60954 , n588278 , n60956 , n60957 , n60958 , n60959 , 
     n60960 , n60961 , n60962 , n60963 , n60964 , n60965 , n60966 , n60967 , n60968 , n60969 , 
     n60970 , n60971 , n60972 , n60973 , n588297 , n60975 , n60976 , n60977 , n60978 , n60979 , 
     n60980 , n60981 , n60982 , n60983 , n60984 , n60985 , n60986 , n588310 , n60988 , n60989 , 
     n588313 , n60991 , n588315 , n60993 , n588317 , n60995 , n60996 , n60997 , n60998 , n588322 , 
     n588323 , n61001 , n588325 , n588326 , n588327 , n588328 , n61006 , n588330 , n588331 , n588332 , 
     n588333 , n61011 , n588335 , n588336 , n61014 , n588338 , n588339 , n61017 , n588341 , n588342 , 
     n61020 , n588344 , n588345 , n61023 , n588347 , n588348 , n61026 , n588350 , n588351 , n61029 , 
     n588353 , n588354 , n61032 , n588356 , n588357 , n588358 , n588359 , n61037 , n588361 , n588362 , 
     n61040 , n588364 , n588365 , n61043 , n61044 , n588368 , n588369 , n61047 , n61048 , n588372 , 
     n588373 , n61051 , n588375 , n588376 , n588377 , n61055 , n61056 , n61057 , n588381 , n61059 , 
     n61060 , n588384 , n61062 , n588386 , n61064 , n588388 , n588389 , n61067 , n588391 , n588392 , 
     n61070 , n588394 , n588395 , n61073 , n588397 , n61075 , n588399 , n61077 , n61078 , n588402 , 
     n61080 , n588404 , n588405 , n61083 , n588407 , n588408 , n61086 , n61087 , n61088 , n61089 , 
     n61090 , n588414 , n61092 , n61093 , n61094 , n61095 , n61096 , n61097 , n588421 , n61099 , 
     n588423 , n588424 , n61102 , n588426 , n588427 , n61105 , n61106 , n588430 , n61108 , n61109 , 
     n61110 , n61111 , n588435 , n588436 , n588437 , n61115 , n588439 , n588440 , n588441 , n61119 , 
     n588443 , n61121 , n588445 , n588446 , n61124 , n588448 , n61126 , n588450 , n588451 , n61129 , 
     n588453 , n588454 , n588455 , n61133 , n588457 , n61135 , n588459 , n588460 , n61138 , n588462 , 
     n61140 , n61141 , n61142 , n588466 , n588467 , n61145 , n588469 , n588470 , n588471 , n588472 , 
     n61150 , n588474 , n588475 , n61153 , n588477 , n588478 , n61156 , n588480 , n588481 , n61159 , 
     n588483 , n61161 , n61162 , n588486 , n588487 , n588488 , n61166 , n588490 , n588491 , n588492 , 
     n588493 , n61171 , n588495 , n588496 , n61174 , n588498 , n588499 , n61177 , n588501 , n588502 , 
     n61180 , n61181 , n61182 , n588506 , n61184 , n61185 , n61186 , n588510 , n588511 , n61189 , 
     n588513 , n588514 , n588515 , n588516 , n61194 , n588518 , n588519 , n61197 , n588521 , n588522 , 
     n61200 , n588524 , n588525 , n61203 , n588527 , n61205 , n61206 , n61207 , n61208 , n61209 , 
     n588533 , n61211 , n588535 , n588536 , n61214 , n588538 , n588539 , n61217 , n588541 , n588542 , 
     n588543 , n588544 , n61222 , n588546 , n588547 , n61225 , n588549 , n61227 , n588551 , n61229 , 
     n61230 , n588554 , n61232 , n588556 , n588557 , n588558 , n61236 , n588560 , n588561 , n61239 , 
     n588563 , n588564 , n61242 , n588566 , n588567 , n588568 , n61246 , n61247 , n588571 , n61249 , 
     n588573 , n588574 , n61252 , n588576 , n61254 , n588578 , n61256 , n588580 , n588581 , n61259 , 
     n61260 , n588584 , n588585 , n61263 , n588587 , n588588 , n61266 , n588590 , n588591 , n61269 , 
     n588593 , n588594 , n61272 , n61273 , n588597 , n588598 , n61276 , n588600 , n61278 , n588602 , 
     n588603 , n61281 , n588605 , n61283 , n61284 , n61285 , n61286 , n61287 , n61288 , n61289 , 
     n61290 , n61291 , n61292 , n61293 , n61294 , n61295 , n61296 , n61297 , n61298 , n61299 , 
     n61300 , n61301 , n61302 , n61303 , n61304 , n61305 , n588629 , n61307 , n61308 , n588632 , 
     n61310 , n588634 , n61312 , n588636 , n588637 , n61315 , n588639 , n588640 , n61318 , n61319 , 
     n588643 , n588644 , n61322 , n588646 , n588647 , n61325 , n588649 , n588650 , n61328 , n61329 , 
     n61330 , n61331 , n61332 , n61333 , n61334 , n61335 , n61336 , n61337 , n61338 , n61339 , 
     n61340 , n61341 , n588665 , n61343 , n61344 , n588668 , n588669 , n61347 , n588671 , n588672 , 
     n588673 , n61351 , n588675 , n61353 , n588677 , n61355 , n61356 , n588680 , n61358 , n588682 , 
     n588683 , n61361 , n588685 , n61363 , n61364 , n61365 , n588689 , n588690 , n61368 , n588692 , 
     n588693 , n588694 , n588695 , n61373 , n588697 , n588698 , n61376 , n588700 , n588701 , n61379 , 
     n588703 , n588704 , n61382 , n588706 , n61384 , n61385 , n61386 , n61387 , n588711 , n61389 , 
     n61390 , n61391 , n61392 , n61393 , n61394 , n61395 , n61396 , n61397 , n61398 , n61399 , 
     n588723 , n588724 , n61402 , n588726 , n61404 , n61405 , n61406 , n61407 , n61408 , n61409 , 
     n61410 , n588734 , n61412 , n588736 , n61414 , n61415 , n588739 , n61417 , n588741 , n61419 , 
     n61420 , n588744 , n61422 , n61423 , n61424 , n61425 , n61426 , n61427 , n61428 , n61429 , 
     n61430 , n588754 , n588755 , n61433 , n588757 , n61435 , n588759 , n588760 , n588761 , n61439 , 
     n588763 , n61441 , n588765 , n588766 , n61444 , n588768 , n61446 , n61447 , n61448 , n61449 , 
     n588773 , n588774 , n61452 , n588776 , n588777 , n588778 , n588779 , n61457 , n588781 , n588782 , 
     n61460 , n588784 , n588785 , n61463 , n588787 , n588788 , n61466 , n588790 , n588791 , n588792 , 
     n588793 , n61471 , n588795 , n588796 , n588797 , n588798 , n61476 , n588800 , n588801 , n61479 , 
     n588803 , n588804 , n61482 , n588806 , n588807 , n61485 , n588809 , n588810 , n61488 , n588812 , 
     n61490 , n588814 , n61492 , n588816 , n61494 , n588818 , n61496 , n61497 , n588821 , n588822 , 
     n61500 , n61501 , n588825 , n588826 , n61504 , n588828 , n588829 , n61507 , n588831 , n588832 , 
     n61510 , n61511 , n588835 , n588836 , n61514 , n61515 , n588839 , n588840 , n61518 , n61519 , 
     n61520 , n61521 , n588845 , n588846 , n61524 , n588848 , n61526 , n588850 , n61528 , n61529 , 
     n588853 , n588854 , n61532 , n61533 , n588857 , n61535 , n61536 , n61537 , n61538 , n61539 , 
     n588863 , n61541 , n61542 , n61543 , n588867 , n588868 , n61546 , n588870 , n588871 , n61549 , 
     n61550 , n588874 , n61552 , n61553 , n61554 , n61555 , n588879 , n61557 , n61558 , n61559 , 
     n61560 , n588884 , n588885 , n588886 , n61564 , n588888 , n61566 , n61567 , n588891 , n588892 , 
     n61570 , n61571 , n588895 , n588896 , n61574 , n588898 , n588899 , n588900 , n588901 , n61579 , 
     n588903 , n61581 , n588905 , n588906 , n61584 , n61585 , n61586 , n61587 , n588911 , n61589 , 
     n61590 , n61591 , n61592 , n588916 , n588917 , n61595 , n61596 , n61597 , n61598 , n61599 , 
     n588923 , n588924 , n588925 , n61603 , n588927 , n588928 , n61606 , n588930 , n588931 , n61609 , 
     n61610 , n588934 , n588935 , n61613 , n61614 , n588938 , n588939 , n61617 , n61618 , n61619 , 
     n61620 , n588944 , n588945 , n61623 , n588947 , n588948 , n61626 , n588950 , n588951 , n61629 , 
     n588953 , n61631 , n61632 , n61633 , n61634 , n61635 , n588959 , n588960 , n61638 , n61639 , 
     n61640 , n61641 , n588965 , n588966 , n61644 , n588968 , n61646 , n588970 , n61648 , n588972 , 
     n588973 , n61651 , n588975 , n588976 , n61654 , n588978 , n61656 , n61657 , n61658 , n61659 , 
     n61660 , n588984 , n61662 , n588986 , n588987 , n61665 , n588989 , n588990 , n61668 , n61669 , 
     n61670 , n61671 , n588995 , n588996 , n588997 , n588998 , n61676 , n589000 , n589001 , n61679 , 
     n61680 , n61681 , n61682 , n589006 , n61684 , n61685 , n61686 , n61687 , n61688 , n589012 , 
     n589013 , n61691 , n589015 , n589016 , n589017 , n589018 , n61696 , n589020 , n589021 , n61699 , 
     n589023 , n61701 , n589025 , n61703 , n61704 , n589028 , n589029 , n61707 , n589031 , n589032 , 
     n61710 , n589034 , n589035 , n61713 , n589037 , n589038 , n589039 , n589040 , n61718 , n589042 , 
     n589043 , n589044 , n589045 , n61723 , n589047 , n589048 , n61726 , n589050 , n589051 , n61729 , 
     n589053 , n589054 , n61732 , n61733 , n61734 , n589058 , n589059 , n61737 , n589061 , n589062 , 
     n61740 , n589064 , n589065 , n589066 , n61744 , n589068 , n61746 , n589070 , n589071 , n61749 , 
     n589073 , n61751 , n61752 , n61753 , n589077 , n61755 , n61756 , n61757 , n589081 , n589082 , 
     n589083 , n61761 , n589085 , n589086 , n61764 , n589088 , n61766 , n589090 , n61768 , n589092 , 
     n589093 , n61771 , n589095 , n61773 , n61774 , n61775 , n61776 , n61777 , n61778 , n61779 , 
     n61780 , n61781 , n61782 , n61783 , n589107 , n61785 , n589109 , n61787 , n589111 , n61789 , 
     n589113 , n61791 , n589115 , n61793 , n61794 , n61795 , n589119 , n589120 , n61798 , n589122 , 
     n589123 , n61801 , n589125 , n61803 , n589127 , n61805 , n61806 , n589130 , n589131 , n61809 , 
     n589133 , n589134 , n589135 , n61813 , n589137 , n61815 , n589139 , n61817 , n61818 , n589142 , 
     n589143 , n61821 , n61822 , n589146 , n589147 , n61825 , n61826 , n589150 , n589151 , n61829 , 
     n61830 , n589154 , n589155 , n61833 , n589157 , n61835 , n589159 , n61837 , n589161 , n61839 , 
     n61840 , n589164 , n589165 , n61843 , n61844 , n589168 , n589169 , n61847 , n61848 , n589172 , 
     n589173 , n61851 , n61852 , n589176 , n589177 , n589178 , n61856 , n589180 , n589181 , n61859 , 
     n589183 , n589184 , n61862 , n61863 , n589187 , n589188 , n61866 , n61867 , n589191 , n589192 , 
     n61870 , n589194 , n589195 , n61873 , n589197 , n589198 , n589199 , n589200 , n61878 , n589202 , 
     n589203 , n61881 , n589205 , n589206 , n61884 , n61885 , n589209 , n61887 , n61888 , n589212 , 
     n589213 , n61891 , n589215 , n589216 , n61894 , n589218 , n589219 , n61897 , n61898 , n61899 , 
     n589223 , n589224 , n61902 , n61903 , n61904 , n589228 , n589229 , n61907 , n61908 , n589232 , 
     n589233 , n61911 , n61912 , n589236 , n61914 , n61915 , n61916 , n61917 , n589241 , n61919 , 
     n61920 , n61921 , n61922 , n589246 , n589247 , n589248 , n61926 , n589250 , n589251 , n589252 , 
     n589253 , n61931 , n589255 , n589256 , n61934 , n589258 , n61936 , n589260 , n61938 , n61939 , 
     n589263 , n589264 , n61942 , n589266 , n589267 , n61945 , n589269 , n589270 , n61948 , n589272 , 
     n589273 , n589274 , n589275 , n61953 , n589277 , n589278 , n589279 , n589280 , n61958 , n589282 , 
     n589283 , n61961 , n589285 , n589286 , n61964 , n589288 , n589289 , n61967 , n61968 , n61969 , 
     n589293 , n589294 , n61972 , n589296 , n61974 , n589298 , n61976 , n61977 , n589301 , n589302 , 
     n61980 , n61981 , n589305 , n589306 , n61984 , n589308 , n61986 , n61987 , n589311 , n589312 , 
     n61990 , n61991 , n589315 , n589316 , n61994 , n61995 , n61996 , n589320 , n589321 , n61999 , 
     n589323 , n589324 , n62002 , n589326 , n589327 , n62005 , n589329 , n589330 , n62008 , n589332 , 
     n589333 , n62011 , n589335 , n589336 , n62014 , n589338 , n589339 , n62017 , n589341 , n62019 , 
     n589343 , n62021 , n589345 , n589346 , n62024 , n62025 , n589349 , n62027 , n589351 , n62029 , 
     n589353 , n589354 , n62032 , n589356 , n589357 , n62035 , n62036 , n589360 , n62038 , n589362 , 
     n62040 , n589364 , n589365 , n62043 , n589367 , n589368 , n62046 , n589370 , n589371 , n62049 , 
     n62050 , n589374 , n589375 , n62053 , n589377 , n589378 , n62056 , n589380 , n589381 , n62059 , 
     n62060 , n589384 , n62062 , n62063 , n589387 , n589388 , n589389 , n62067 , n589391 , n589392 , 
     n62070 , n62071 , n589395 , n589396 , n62074 , n589398 , n589399 , n62077 , n589401 , n589402 , 
     n62080 , n589404 , n589405 , n62083 , n62084 , n589408 , n589409 , n62087 , n589411 , n589412 , 
     n62090 , n589414 , n589415 , n62093 , n62094 , n589418 , n589419 , n589420 , n589421 , n589422 , 
     n62100 , n589424 , n589425 , n62103 , n62104 , n589428 , n62106 , n589430 , n589431 , n62109 , 
     n62110 , n589434 , n589435 , n62113 , n62114 , n589438 , n62116 , n62117 , n62118 , n62119 , 
     n589443 , n589444 , n589445 , n62123 , n589447 , n589448 , n589449 , n62127 , n589451 , n62129 , 
     n589453 , n589454 , n62132 , n589456 , n62134 , n62135 , n62136 , n62137 , n62138 , n62139 , 
     n62140 , n62141 , n62142 , n62143 , n589467 , n62145 , n589469 , n589470 , n62148 , n589472 , 
     n589473 , n62151 , n62152 , n589476 , n589477 , n62155 , n62156 , n589480 , n589481 , n62159 , 
     n62160 , n589484 , n62162 , n62163 , n589487 , n589488 , n62166 , n62167 , n589491 , n62169 , 
     n62170 , n62171 , n62172 , n62173 , n62174 , n589498 , n62176 , n62177 , n62178 , n589502 , 
     n62180 , n62181 , n62182 , n62183 , n62184 , n62185 , n589509 , n62187 , n62188 , n62189 , 
     n62190 , n62191 , n589515 , n62193 , n62194 , n589518 , n589519 , n62197 , n62198 , n589522 , 
     n589523 , n62201 , n589525 , n589526 , n62204 , n589528 , n589529 , n62207 , n589531 , n589532 , 
     n589533 , n589534 , n62212 , n589536 , n589537 , n62215 , n589539 , n62217 , n589541 , n62219 , 
     n62220 , n589544 , n589545 , n62223 , n589547 , n589548 , n62226 , n589550 , n589551 , n62229 , 
     n589553 , n589554 , n589555 , n589556 , n62234 , n589558 , n589559 , n62237 , n62238 , n589562 , 
     n62240 , n62241 , n62242 , n589566 , n589567 , n62245 , n62246 , n62247 , n589571 , n589572 , 
     n589573 , n589574 , n62252 , n589576 , n62254 , n62255 , n589579 , n589580 , n62258 , n62259 , 
     n589583 , n589584 , n62262 , n62263 , n589587 , n62265 , n589589 , n589590 , n62268 , n62269 , 
     n589593 , n62271 , n589595 , n62273 , n589597 , n589598 , n62276 , n589600 , n589601 , n62279 , 
     n62280 , n589604 , n589605 , n62283 , n62284 , n589608 , n589609 , n62287 , n62288 , n62289 , 
     n589613 , n589614 , n62292 , n589616 , n62294 , n62295 , n589619 , n62297 , n589621 , n62299 , 
     n589623 , n62301 , n62302 , n62303 , n62304 , n62305 , n62306 , n62307 , n62308 , n589632 , 
     n62310 , n589634 , n62312 , n62313 , n589637 , n62315 , n62316 , n589640 , n62318 , n62319 , 
     n589643 , n62321 , n62322 , n589646 , n62324 , n62325 , n62326 , n62327 , n589651 , n62329 , 
     n62330 , n589654 , n589655 , n62333 , n589657 , n589658 , n62336 , n62337 , n589661 , n62339 , 
     n62340 , n62341 , n62342 , n62343 , n62344 , n589668 , n62346 , n62347 , n589671 , n62349 , 
     n62350 , n62351 , n62352 , n589676 , n589677 , n62355 , n589679 , n62357 , n62358 , n62359 , 
     n589683 , n589684 , n589685 , n62363 , n589687 , n589688 , n62366 , n62367 , n589691 , n589692 , 
     n589693 , n62371 , n589695 , n589696 , n589697 , n589698 , n62376 , n589700 , n589701 , n62379 , 
     n589703 , n589704 , n62382 , n589706 , n589707 , n62385 , n589709 , n589710 , n62388 , n589712 , 
     n589713 , n62391 , n589715 , n589716 , n62394 , n589718 , n589719 , n62397 , n589721 , n589722 , 
     n589723 , n589724 , n62402 , n589726 , n589727 , n62405 , n589729 , n589730 , n62408 , n62409 , 
     n589733 , n589734 , n62412 , n62413 , n589737 , n589738 , n62416 , n62417 , n589741 , n589742 , 
     n62420 , n62421 , n589745 , n589746 , n62424 , n589748 , n589749 , n62427 , n62428 , n62429 , 
     n62430 , n62431 , n589755 , n62433 , n589757 , n589758 , n62436 , n62437 , n589761 , n589762 , 
     n62440 , n589764 , n589765 , n62443 , n589767 , n62445 , n62446 , n62447 , n62448 , n62449 , 
     n62450 , n62451 , n62452 , n589776 , n589777 , n62455 , n589779 , n62457 , n62458 , n62459 , 
     n62460 , n62461 , n62462 , n62463 , n62464 , n62465 , n62466 , n62467 , n62468 , n62469 , 
     n62470 , n589794 , n62472 , n62473 , n62474 , n62475 , n589799 , n62477 , n589801 , n589802 , 
     n62480 , n589804 , n589805 , n589806 , n589807 , n62485 , n589809 , n589810 , n62488 , n589812 , 
     n589813 , n62491 , n589815 , n589816 , n62494 , n589818 , n62496 , n589820 , n62498 , n589822 , 
     n62500 , n62501 , n589825 , n589826 , n62504 , n589828 , n62506 , n589830 , n589831 , n62509 , 
     n589833 , n62511 , n62512 , n62513 , n62514 , n62515 , n62516 , n589840 , n62518 , n62519 , 
     n589843 , n62521 , n589845 , n62523 , n62524 , n589848 , n589849 , n62527 , n589851 , n62529 , 
     n62530 , n62531 , n62532 , n62533 , n62534 , n62535 , n62536 , n62537 , n62538 , n62539 , 
     n62540 , n62541 , n62542 , n62543 , n62544 , n62545 , n62546 , n62547 , n589871 , n62549 , 
     n62550 , n589874 , n589875 , n62553 , n589877 , n62555 , n589879 , n589880 , n62558 , n589882 , 
     n589883 , n589884 , n62562 , n589886 , n589887 , n62565 , n589889 , n62567 , n62568 , n589892 , 
     n589893 , n62571 , n589895 , n589896 , n62574 , n589898 , n62576 , n62577 , n62578 , n62579 , 
     n62580 , n589904 , n589905 , n62583 , n589907 , n62585 , n589909 , n62587 , n62588 , n589912 , 
     n62590 , n589914 , n589915 , n62593 , n589917 , n62595 , n62596 , n62597 , n62598 , n589922 , 
     n62600 , n62601 , n589925 , n589926 , n62604 , n589928 , n62606 , n62607 , n589931 , n62609 , 
     n589933 , n62611 , n589935 , n589936 , n62614 , n589938 , n62616 , n62617 , n589941 , n62619 , 
     n589943 , n62621 , n589945 , n589946 , n62624 , n589948 , n62626 , n62627 , n62628 , n62629 , 
     n62630 , n589954 , n62632 , n589956 , n62634 , n589958 , n62636 , n62637 , n62638 , n62639 , 
     n62640 , n62641 , n589965 , n62643 , n62644 , n589968 , n62646 , n62647 , n589971 , n62649 , 
     n62650 , n62651 , n62652 , n589976 , n62654 , n589978 , n62656 , n589980 , n589981 , n62659 , 
     n589983 , n589984 , n62662 , n62663 , n589987 , n589988 , n62666 , n62667 , n589991 , n589992 , 
     n589993 , n589994 , n589995 , n62673 , n589997 , n589998 , n62676 , n590000 , n62678 , n590002 , 
     n590003 , n62681 , n62682 , n62683 , n62684 , n62685 , n62686 , n62687 , n590011 , n62689 , 
     n590013 , n590014 , n62692 , n590016 , n590017 , n62695 , n590019 , n590020 , n590021 , n62699 , 
     n590023 , n62701 , n590025 , n590026 , n62704 , n62705 , n62706 , n62707 , n590031 , n62709 , 
     n62710 , n62711 , n62712 , n590036 , n590037 , n62715 , n62716 , n590040 , n62718 , n590042 , 
     n62720 , n62721 , n62722 , n590046 , n62724 , n590048 , n590049 , n590050 , n62728 , n590052 , 
     n590053 , n62731 , n590055 , n590056 , n62734 , n62735 , n590059 , n590060 , n62738 , n62739 , 
     n590063 , n62741 , n62742 , n62743 , n62744 , n62745 , n590069 , n62747 , n590071 , n590072 , 
     n62750 , n590074 , n590075 , n62753 , n62754 , n590078 , n590079 , n62757 , n62758 , n590082 , 
     n62760 , n62761 , n62762 , n62763 , n62764 , n62765 , n62766 , n62767 , n62768 , n62769 , 
     n590093 , n62771 , n62772 , n590096 , n62774 , n62775 , n62776 , n62777 , n590101 , n62779 , 
     n62780 , n62781 , n62782 , n62783 , n590107 , n590108 , n590109 , n62787 , n590111 , n590112 , 
     n590113 , n62791 , n590115 , n62793 , n62794 , n590118 , n590119 , n62797 , n590121 , n62799 , 
     n62800 , n62801 , n62802 , n590126 , n590127 , n590128 , n62806 , n590130 , n590131 , n590132 , 
     n590133 , n62811 , n590135 , n590136 , n62814 , n590138 , n590139 , n62817 , n590141 , n590142 , 
     n62820 , n62821 , n62822 , n590146 , n590147 , n590148 , n62826 , n590150 , n590151 , n590152 , 
     n590153 , n62831 , n590155 , n590156 , n62834 , n590158 , n590159 , n62837 , n590161 , n590162 , 
     n62840 , n62841 , n62842 , n590166 , n62844 , n62845 , n590169 , n590170 , n62848 , n590172 , 
     n62850 , n62851 , n62852 , n62853 , n62854 , n590178 , n62856 , n590180 , n590181 , n62859 , 
     n590183 , n590184 , n62862 , n62863 , n590187 , n62865 , n62866 , n590190 , n62868 , n590192 , 
     n590193 , n62871 , n62872 , n62873 , n590197 , n590198 , n590199 , n590200 , n62878 , n590202 , 
     n590203 , n62881 , n590205 , n590206 , n62884 , n590208 , n590209 , n62887 , n62888 , n590212 , 
     n590213 , n62891 , n590215 , n590216 , n62894 , n590218 , n590219 , n62897 , n590221 , n590222 , 
     n62900 , n590224 , n62902 , n62903 , n62904 , n590228 , n62906 , n590230 , n62908 , n62909 , 
     n590233 , n590234 , n62912 , n62913 , n590237 , n590238 , n62916 , n590240 , n62918 , n62919 , 
     n590243 , n590244 , n62922 , n62923 , n590247 , n62925 , n62926 , n62927 , n62928 , n62929 , 
     n62930 , n590254 , n62932 , n62933 , n62934 , n62935 , n590259 , n590260 , n62938 , n62939 , 
     n62940 , n590264 , n590265 , n62943 , n590267 , n590268 , n62946 , n62947 , n590271 , n62949 , 
     n62950 , n62951 , n62952 , n590276 , n62954 , n62955 , n590279 , n590280 , n62958 , n62959 , 
     n590283 , n590284 , n62962 , n590286 , n62964 , n62965 , n590289 , n590290 , n62968 , n62969 , 
     n590293 , n590294 , n62972 , n62973 , n590297 , n590298 , n62976 , n590300 , n590301 , n62979 , 
     n590303 , n590304 , n62982 , n590306 , n62984 , n62985 , n62986 , n590310 , n590311 , n62989 , 
     n590313 , n62991 , n590315 , n62993 , n62994 , n590318 , n62996 , n590320 , n62998 , n590322 , 
     n590323 , n63001 , n590325 , n590326 , n63004 , n63005 , n63006 , n63007 , n63008 , n590332 , 
     n63010 , n63011 , n590335 , n63013 , n63014 , n63015 , n63016 , n590340 , n63018 , n63019 , 
     n63020 , n63021 , n63022 , n590346 , n63024 , n63025 , n63026 , n63027 , n63028 , n63029 , 
     n63030 , n590354 , n63032 , n590356 , n590357 , n63035 , n590359 , n590360 , n63038 , n63039 , 
     n590363 , n590364 , n63042 , n63043 , n590367 , n63045 , n63046 , n590370 , n590371 , n63049 , 
     n590373 , n590374 , n590375 , n590376 , n63054 , n590378 , n590379 , n63057 , n590381 , n590382 , 
     n63060 , n590384 , n590385 , n63063 , n63064 , n63065 , n590389 , n63067 , n590391 , n590392 , 
     n63070 , n590394 , n590395 , n590396 , n63074 , n590398 , n63076 , n63077 , n63078 , n63079 , 
     n63080 , n63081 , n63082 , n63083 , n63084 , n63085 , n63086 , n63087 , n63088 , n63089 , 
     n63090 , n590414 , n63092 , n63093 , n590417 , n590418 , n63096 , n63097 , n590421 , n63099 , 
     n63100 , n63101 , n63102 , n590426 , n590427 , n590428 , n63106 , n590430 , n590431 , n590432 , 
     n590433 , n63111 , n590435 , n590436 , n63114 , n590438 , n590439 , n63117 , n590441 , n590442 , 
     n63120 , n63121 , n63122 , n590446 , n590447 , n63125 , n63126 , n63127 , n590451 , n63129 , 
     n590453 , n590454 , n63132 , n590456 , n590457 , n590458 , n63136 , n590460 , n63138 , n63139 , 
     n63140 , n63141 , n63142 , n63143 , n590467 , n63145 , n63146 , n63147 , n590471 , n590472 , 
     n590473 , n590474 , n63152 , n590476 , n590477 , n590478 , n590479 , n63157 , n590481 , n590482 , 
     n63160 , n590484 , n590485 , n63163 , n590487 , n590488 , n63166 , n590490 , n590491 , n63169 , 
     n63170 , n590494 , n590495 , n63173 , n590497 , n63175 , n63176 , n63177 , n63178 , n63179 , 
     n590503 , n590504 , n63182 , n590506 , n63184 , n590508 , n590509 , n63187 , n590511 , n63189 , 
     n63190 , n590514 , n590515 , n63193 , n590517 , n590518 , n63196 , n590520 , n590521 , n63199 , 
     n590523 , n63201 , n63202 , n63203 , n63204 , n590528 , n63206 , n63207 , n63208 , n63209 , 
     n63210 , n63211 , n63212 , n63213 , n63214 , n63215 , n590539 , n63217 , n63218 , n63219 , 
     n63220 , n63221 , n63222 , n590546 , n590547 , n63225 , n590549 , n63227 , n63228 , n63229 , 
     n63230 , n63231 , n63232 , n63233 , n63234 , n63235 , n63236 , n63237 , n63238 , n590562 , 
     n63240 , n63241 , n63242 , n590566 , n590567 , n590568 , n590569 , n63247 , n590571 , n590572 , 
     n590573 , n63251 , n590575 , n63253 , n590577 , n590578 , n63256 , n590580 , n63258 , n63259 , 
     n63260 , n63261 , n63262 , n63263 , n63264 , n63265 , n63266 , n63267 , n590591 , n590592 , 
     n63270 , n590594 , n63272 , n63273 , n63274 , n63275 , n63276 , n590600 , n63278 , n63279 , 
     n63280 , n63281 , n63282 , n63283 , n63284 , n63285 , n590609 , n63287 , n63288 , n590612 , 
     n63290 , n63291 , n63292 , n63293 , n590617 , n590618 , n63296 , n590620 , n63298 , n63299 , 
     n590623 , n590624 , n63302 , n590626 , n63304 , n590628 , n590629 , n63307 , n590631 , n590632 , 
     n63310 , n590634 , n590635 , n590636 , n590637 , n63315 , n590639 , n63317 , n63318 , n63319 , 
     n63320 , n63321 , n63322 , n63323 , n63324 , n63325 , n63326 , n63327 , n63328 , n590652 , 
     n63330 , n590654 , n63332 , n590656 , n590657 , n63335 , n590659 , n590660 , n63338 , n63339 , 
     n590663 , n590664 , n63342 , n63343 , n590667 , n590668 , n590669 , n63347 , n590671 , n590672 , 
     n63350 , n590674 , n590675 , n63353 , n63354 , n590678 , n590679 , n63357 , n63358 , n590682 , 
     n590683 , n63361 , n63362 , n63363 , n63364 , n63365 , n63366 , n63367 , n590691 , n63369 , 
     n63370 , n63371 , n590695 , n590696 , n63374 , n590698 , n590699 , n63377 , n63378 , n63379 , 
     n63380 , n63381 , n63382 , n63383 , n63384 , n63385 , n590709 , n63387 , n590711 , n590712 , 
     n63390 , n590714 , n590715 , n63393 , n63394 , n590718 , n590719 , n63397 , n63398 , n590722 , 
     n63400 , n63401 , n63402 , n63403 , n63404 , n63405 , n63406 , n63407 , n63408 , n63409 , 
     n63410 , n63411 , n63412 , n590736 , n63414 , n590738 , n590739 , n63417 , n63418 , n590742 , 
     n63420 , n590744 , n590745 , n590746 , n590747 , n63425 , n590749 , n63427 , n590751 , n590752 , 
     n63430 , n63431 , n63432 , n63433 , n590757 , n63435 , n63436 , n590760 , n590761 , n63439 , 
     n590763 , n63441 , n590765 , n590766 , n63444 , n590768 , n590769 , n590770 , n63448 , n590772 , 
     n63450 , n63451 , n63452 , n63453 , n63454 , n63455 , n590779 , n590780 , n590781 , n63459 , 
     n590783 , n590784 , n590785 , n590786 , n63464 , n590788 , n590789 , n63467 , n590791 , n590792 , 
     n63470 , n590794 , n590795 , n63473 , n590797 , n590798 , n63476 , n63477 , n63478 , n63479 , 
     n63480 , n63481 , n63482 , n63483 , n63484 , n63485 , n63486 , n63487 , n63488 , n63489 , 
     n63490 , n63491 , n63492 , n590816 , n63494 , n63495 , n63496 , n63497 , n63498 , n63499 , 
     n63500 , n63501 , n63502 , n63503 , n590827 , n63505 , n63506 , n63507 , n590831 , n590832 , 
     n590833 , n590834 , n63512 , n590836 , n590837 , n63515 , n63516 , n63517 , n63518 , n590842 , 
     n590843 , n63521 , n63522 , n63523 , n63524 , n63525 , n590849 , n63527 , n590851 , n590852 , 
     n63530 , n63531 , n590855 , n63533 , n63534 , n63535 , n63536 , n590860 , n63538 , n63539 , 
     n590863 , n63541 , n63542 , n590866 , n63544 , n63545 , n590869 , n63547 , n63548 , n63549 , 
     n63550 , n590874 , n63552 , n63553 , n590877 , n63555 , n63556 , n63557 , n63558 , n590882 , 
     n63560 , n63561 , n63562 , n63563 , n63564 , n63565 , n63566 , n63567 , n590891 , n63569 , 
     n63570 , n590894 , n590895 , n63573 , n590897 , n590898 , n63576 , n63577 , n590901 , n590902 , 
     n590903 , n590904 , n63582 , n590906 , n590907 , n63585 , n63586 , n63587 , n63588 , n590912 , 
     n590913 , n590914 , n63592 , n590916 , n590917 , n63595 , n63596 , n63597 , n63598 , n63599 , 
     n590923 , n590924 , n590925 , n63603 , n590927 , n590928 , n63606 , n63607 , n63608 , n63609 , 
     n590933 , n590934 , n63612 , n590936 , n63614 , n63615 , n63616 , n63617 , n63618 , n63619 , 
     n590943 , n63621 , n63622 , n63623 , n63624 , n590948 , n590949 , n590950 , n590951 , n63629 , 
     n590953 , n590954 , n590955 , n63633 , n590957 , n590958 , n590959 , n63637 , n590961 , n63639 , 
     n63640 , n63641 , n590965 , n63643 , n63644 , n590968 , n63646 , n63647 , n63648 , n63649 , 
     n590973 , n63651 , n63652 , n590976 , n63654 , n63655 , n63656 , n63657 , n590981 , n590982 , 
     n590983 , n63661 , n590985 , n590986 , n63664 , n590988 , n590989 , n63667 , n590991 , n590992 , 
     n63670 , n63671 , n590995 , n590996 , n63674 , n63675 , n590999 , n591000 , n63678 , n591002 , 
     n591003 , n63681 , n591005 , n591006 , n63684 , n63685 , n591009 , n591010 , n63688 , n63689 , 
     n591013 , n591014 , n63692 , n591016 , n591017 , n63695 , n591019 , n591020 , n63698 , n591022 , 
     n63700 , n591024 , n591025 , n63703 , n591027 , n591028 , n63706 , n591030 , n591031 , n63709 , 
     n591033 , n591034 , n591035 , n591036 , n63714 , n591038 , n591039 , n63717 , n591041 , n591042 , 
     n63720 , n591044 , n591045 , n63723 , n63724 , n63725 , n591049 , n591050 , n63728 , n63729 , 
     n591053 , n591054 , n63732 , n63733 , n591057 , n591058 , n63736 , n591060 , n591061 , n63739 , 
     n591063 , n591064 , n591065 , n591066 , n63744 , n591068 , n591069 , n63747 , n591071 , n63749 , 
     n63750 , n591074 , n63752 , n63753 , n591077 , n591078 , n63756 , n591080 , n591081 , n63759 , 
     n591083 , n591084 , n63762 , n591086 , n591087 , n63765 , n63766 , n591090 , n63768 , n591092 , 
     n591093 , n591094 , n63772 , n591096 , n591097 , n63775 , n591099 , n591100 , n63778 , n591102 , 
     n591103 , n63781 , n591105 , n591106 , n63784 , n63785 , n591109 , n591110 , n63788 , n591112 , 
     n591113 , n591114 , n591115 , n63793 , n591117 , n591118 , n63796 , n591120 , n63798 , n591122 , 
     n63800 , n63801 , n591125 , n591126 , n63804 , n591128 , n591129 , n63807 , n591131 , n591132 , 
     n63810 , n591134 , n591135 , n591136 , n591137 , n63815 , n591139 , n591140 , n63818 , n591142 , 
     n63820 , n591144 , n63822 , n63823 , n591147 , n591148 , n63826 , n63827 , n591151 , n591152 , 
     n63830 , n63831 , n63832 , n591156 , n591157 , n63835 , n591159 , n591160 , n591161 , n63839 , 
     n591163 , n63841 , n591165 , n591166 , n63844 , n591168 , n591169 , n63847 , n591171 , n591172 , 
     n63850 , n591174 , n63852 , n591176 , n591177 , n591178 , n591179 , n63857 , n591181 , n63859 , 
     n591183 , n591184 , n63862 , n63863 , n63864 , n63865 , n591189 , n63867 , n63868 , n591192 , 
     n591193 , n63871 , n591195 , n63873 , n591197 , n63875 , n63876 , n591200 , n591201 , n63879 , 
     n63880 , n591204 , n63882 , n63883 , n63884 , n63885 , n63886 , n63887 , n591211 , n63889 , 
     n591213 , n63891 , n591215 , n591216 , n63894 , n591218 , n63896 , n63897 , n63898 , n63899 , 
     n63900 , n63901 , n63902 , n63903 , n591227 , n63905 , n591229 , n591230 , n63908 , n63909 , 
     n591233 , n591234 , n591235 , n63913 , n591237 , n63915 , n591239 , n591240 , n63918 , n63919 , 
     n63920 , n63921 , n591245 , n591246 , n591247 , n63925 , n591249 , n591250 , n591251 , n63929 , 
     n591253 , n591254 , n63932 , n591256 , n63934 , n63935 , n591259 , n63937 , n63938 , n591262 , 
     n591263 , n63941 , n63942 , n63943 , n63944 , n63945 , n591269 , n63947 , n591271 , n591272 , 
     n591273 , n63951 , n591275 , n591276 , n591277 , n63955 , n591279 , n591280 , n63958 , n591282 , 
     n63960 , n63961 , n591285 , n591286 , n591287 , n63965 , n591289 , n591290 , n591291 , n591292 , 
     n63970 , n591294 , n591295 , n63973 , n63974 , n591298 , n63976 , n63977 , n63978 , n591302 , 
     n591303 , n63981 , n591305 , n63983 , n591307 , n63985 , n63986 , n591310 , n591311 , n63989 , 
     n63990 , n591314 , n591315 , n63993 , n591317 , n63995 , n63996 , n591320 , n591321 , n63999 , 
     n64000 , n591324 , n591325 , n64003 , n591327 , n591328 , n64006 , n64007 , n64008 , n64009 , 
     n64010 , n64011 , n64012 , n64013 , n64014 , n64015 , n591339 , n591340 , n64018 , n591342 , 
     n64020 , n591344 , n591345 , n64023 , n64024 , n64025 , n64026 , n591350 , n591351 , n591352 , 
     n64030 , n591354 , n591355 , n64033 , n591357 , n591358 , n64036 , n591360 , n64038 , n591362 , 
     n591363 , n591364 , n591365 , n64043 , n591367 , n64045 , n591369 , n591370 , n64048 , n64049 , 
     n64050 , n64051 , n591375 , n591376 , n591377 , n591378 , n591379 , n64057 , n64058 , n64059 , 
     n64060 , n64061 , n591385 , n591386 , n591387 , n64065 , n591389 , n64067 , n591391 , n64069 , 
     n64070 , n591394 , n64072 , n591396 , n591397 , n64075 , n591399 , n591400 , n64078 , n591402 , 
     n64080 , n591404 , n591405 , n64083 , n591407 , n591408 , n64086 , n64087 , n591411 , n591412 , 
     n64090 , n64091 , n591415 , n591416 , n64094 , n64095 , n591419 , n591420 , n64098 , n64099 , 
     n591423 , n591424 , n64102 , n591426 , n591427 , n591428 , n64106 , n591430 , n591431 , n591432 , 
     n591433 , n64111 , n591435 , n591436 , n64114 , n591438 , n591439 , n64117 , n64118 , n591442 , 
     n64120 , n64121 , n64122 , n64123 , n591447 , n64125 , n591449 , n591450 , n591451 , n64129 , 
     n591453 , n591454 , n591455 , n591456 , n64134 , n591458 , n591459 , n591460 , n591461 , n591462 , 
     n64140 , n591464 , n591465 , n591466 , n591467 , n591468 , n64146 , n591470 , n591471 , n591472 , 
     n64150 , n591474 , n591475 , n591476 , n591477 , n591478 , n64156 , n591480 , n591481 , n591482 , 
     n64160 , n591484 , n591485 , n591486 , n64164 , n591488 , n591489 , n591490 , n591491 , n591492 , 
     n64170 , n591494 , n64172 , n591496 , n64174 , n591498 , n591499 , n591500 , n64178 , n591502 , 
     n591503 , n591504 , n591505 , n591506 , n64184 , n591508 , n591509 , n591510 , n591511 , n591512 , 
     n591513 , n591514 , n591515 , n591516 , n64194 , n591518 , n591519 , n591520 , n64198 , n591522 , 
     n591523 , n591524 , n64202 , n591526 , n591527 , n591528 , n64206 , n591530 , n64208 , n591532 , 
     n64210 , n591534 , n591535 , n591536 , n64214 , n591538 , n64216 , n591540 , n64218 , n591542 , 
     n64220 , n591544 , n591545 , n591546 , n64224 , n591548 , n64226 , n591550 , n591551 , n591552 , 
     n591553 , n591554 , n591555 , n591556 , n64234 , n591558 , n591559 , n591560 , n64238 , n591562 , 
     n64240 , n591564 , n64242 , n591566 , n591567 , n591568 , n64246 , n591570 , n64248 , n591572 , 
     n591573 , n591574 , n591575 , n591576 , n591577 , n591578 , n591579 , n591580 , n64258 , n591582 , 
     n64260 , n591584 , n591585 , n591586 , n591587 , n591588 , n64266 , n591590 , n591591 , n591592 , 
     n64270 , n591594 , n64272 , n591596 , n591597 , n591598 , n64276 , n591600 , n591601 , n591602 , 
     n64280 , n591604 , n64282 , n591606 , n64284 , n591608 , n591609 , n591610 , n591611 , n591612 , 
     n591613 , n591614 , n591615 , n591616 , n591617 , n591618 , n64296 , n591620 , n591621 , n591622 , 
     n64300 , n591624 , n591625 , n591626 , n591627 , n591628 , n591629 , n591630 , n64308 , n591632 , 
     n64310 , n591634 , n591635 , n591636 , n591637 , n591638 , n591639 , n591640 , n591641 , n591642 , 
     n591643 , n591644 , n591645 , n591646 , n591647 , n591648 , n591649 , n591650 , n591651 , n591652 , 
     n591653 , n591654 , n591655 , n591656 , n591657 , n591658 , n591659 , n591660 , n591661 , n591662 , 
     n591663 , n591664 , n591665 , n591666 , n591667 , n591668 , n591669 , n591670 , n591671 , n591672 , 
     n591673 , n591674 , n591675 , n591676 , n591677 , n591678 , n591679 , n591680 , n591681 , n591682 , 
     n591683 , n591684 , n591685 , n591686 , n591687 , n591688 , n591689 , n591690 , n591691 , n591692 , 
     n591693 , n591694 , n591695 , n591696 , n591697 , n591698 , n591699 , n591700 , n591701 , n591702 , 
     n591703 , n591704 , n591705 , n591706 , n591707 , n591708 , n591709 , n591710 , n591711 , n591712 , 
     n591713 , n591714 , n591715 , n591716 , n591717 , n591718 , n591719 , n591720 , n591721 , n591722 , 
     n591723 , n591724 , n591725 , n591726 , n591727 , n591728 , n591729 , n591730 , n591731 , n591732 , 
     n591733 , n591734 , n591735 , n591736 , n591737 , n591738 , n591739 , n591740 , n591741 , n591742 , 
     n591743 , n591744 , n591745 , n591746 , n591747 , n591748 , n591749 , n591750 , n591751 , n591752 , 
     n591753 , n591754 , n591755 , n591756 , n591757 , n591758 , n591759 , n591760 , n591761 , n591762 , 
     n591763 , n591764 , n591765 , n64443 , n64444 , n64445 , n64446 , n64447 , n64448 , n64449 , 
     n64450 , n64451 , n64452 , n64453 , n64454 , n64455 , n64456 , n64457 , n64458 , n64459 , 
     n591783 , n64461 , n591785 , n591786 , n64464 , n64465 , n64466 , n64467 , n591791 , n64469 , 
     n64470 , n64471 , n64472 , n591796 , n64474 , n64475 , n64476 , n64477 , n64478 , n64479 , 
     n591803 , n64481 , n591805 , n64483 , n64484 , n64485 , n64486 , n64487 , n64488 , n64489 , 
     n64490 , n64491 , n64492 , n64493 , n64494 , n64495 , n591819 , n64497 , n64498 , n64499 , 
     n64500 , n64501 , n64502 , n591826 , n591827 , n64505 , n591829 , n591830 , n591831 , n591832 , 
     n64510 , n64511 , n64512 , n64513 , n64514 , n591838 , n64516 , n591840 , n591841 , n64519 , 
     n64520 , n64521 , n591845 , n64523 , n591847 , n64525 , n64526 , n64527 , n591851 , n64529 , 
     n591853 , n591854 , n64532 , n64533 , n64534 , n64535 , n64536 , n64537 , n64538 , n64539 , 
     n591863 , n591864 , n64542 , n64543 , n64544 , n64545 , n64546 , n64547 , n64548 , n64549 , 
     n64550 , n64551 , n64552 , n64553 , n64554 , n591878 , n64556 , n591880 , n591881 , n64559 , 
     n591883 , n591884 , n64562 , n591886 , n64564 , n64565 , n64566 , n591890 , n591891 , n64569 , 
     n591893 , n64571 , n64572 , n64573 , n64574 , n64575 , n64576 , n591900 , n64578 , n591902 , 
     n591903 , n64581 , n64582 , n64583 , n64584 , n64585 , n64586 , n64587 , n64588 , n64589 , 
     n64590 , n64591 , n64592 , n591916 , n64594 , n591918 , n591919 , n64597 , n591921 , n64599 , 
     n64600 , n64601 , n64602 , n64603 , n64604 , n64605 , n64606 , n64607 , n64608 , n64609 , 
     n64610 , n64611 , n64612 , n64613 , n64614 , n64615 , n64616 , n64617 , n64618 , n64619 , 
     n64620 , n64621 , n64622 , n64623 , n64624 , n64625 , n64626 , n64627 , n64628 , n64629 , 
     n64630 , n64631 , n64632 , n64633 , n64634 , n64635 , n64636 , n64637 , n591961 , n64639 , 
     n591963 , n591964 , n64642 , n591966 , n591967 , n64645 , n591969 , n591970 , n64648 , n64649 , 
     n64650 , n64651 , n591975 , n591976 , n64654 , n64655 , n64656 , n64657 , n591981 , n591982 , 
     n64660 , n64661 , n64662 , n64663 , n591987 , n591988 , n64666 , n591990 , n64668 , n591992 , 
     n591993 , n64671 , n591995 , n591996 , n64674 , n591998 , n591999 , n592000 , n592001 , n64679 , 
     n592003 , n592004 , n64682 , n64683 , n64684 , n64685 , n64686 , n592010 , n64688 , n592012 , 
     n592013 , n64691 , n592015 , n592016 , n64694 , n592018 , n64696 , n64697 , n64698 , n64699 , 
     n592023 , n592024 , n64702 , n592026 , n64704 , n64705 , n64706 , n64707 , n592031 , n592032 , 
     n64710 , n592034 , n64712 , n64713 , n592037 , n592038 , n64716 , n592040 , n592041 , n64719 , 
     n592043 , n64721 , n64722 , n592046 , n64724 , n592048 , n592049 , n64727 , n592051 , n64729 , 
     n592053 , n592054 , n64732 , n592056 , n64734 , n64735 , n592059 , n592060 , n64738 , n592062 , 
     n64740 , n64741 , n64742 , n64743 , n64744 , n64745 , n64746 , n64747 , n64748 , n64749 , 
     n64750 , n64751 , n64752 , n64753 , n64754 , n64755 , n592079 , n64757 , n592081 , n592082 , 
     n64760 , n64761 , n592085 , n592086 , n64764 , n592088 , n592089 , n64767 , n592091 , n592092 , 
     n64770 , n592094 , n64772 , n592096 , n592097 , n64775 , n64776 , n592100 , n64778 , n592102 , 
     n592103 , n592104 , n64782 , n592106 , n592107 , n64785 , n592109 , n592110 , n64788 , n592112 , 
     n592113 , n64791 , n592115 , n64793 , n592117 , n64795 , n592119 , n592120 , n592121 , n64799 , 
     n592123 , n592124 , n64802 , n592126 , n64804 , n592128 , n64806 , n592130 , n592131 , n592132 , 
     n64810 , n592134 , n592135 , n64813 , n592137 , n592138 , n64816 , n592140 , n592141 , n64819 , 
     n592143 , n592144 , n64822 , n592146 , n592147 , n64825 , n592149 , n64827 , n64828 , n64829 , 
     n64830 , n64831 , n592155 , n64833 , n64834 , n64835 , n64836 , n64837 , n64838 , n64839 , 
     n64840 , n64841 , n64842 , n64843 , n64844 , n64845 , n64846 , n64847 , n64848 , n64849 , 
     n64850 , n64851 , n64852 , n64853 , n64854 , n64855 , n64856 , n64857 , n64858 , n64859 , 
     n64860 , n64861 , n64862 , n592186 , n64864 , n592188 , n592189 , n64867 , n592191 , n64869 , 
     n592193 , n592194 , n64872 , n64873 , n592197 , n592198 , n64876 , n64877 , n592201 , n592202 , 
     n64880 , n592204 , n64882 , n64883 , n592207 , n592208 , n64886 , n64887 , n592211 , n64889 , 
     n592213 , n592214 , n64892 , n64893 , n64894 , n64895 , n64896 , n64897 , n64898 , n64899 , 
     n592223 , n64901 , n64902 , n64903 , n592227 , n64905 , n64906 , n64907 , n592231 , n592232 , 
     n64910 , n592234 , n64912 , n64913 , n592237 , n64915 , n592239 , n592240 , n64918 , n64919 , 
     n64920 , n64921 , n592245 , n64923 , n592247 , n592248 , n64926 , n592250 , n64928 , n64929 , 
     n592253 , n592254 , n64932 , n592256 , n592257 , n64935 , n64936 , n64937 , n64938 , n64939 , 
     n64940 , n64941 , n64942 , n64943 , n64944 , n64945 , n64946 , n64947 , n64948 , n64949 , 
     n64950 , n64951 , n592275 , n64953 , n592277 , n592278 , n64956 , n592280 , n592281 , n64959 , 
     n64960 , n64961 , n592285 , n64963 , n64964 , n64965 , n64966 , n592290 , n64968 , n592292 , 
     n592293 , n64971 , n592295 , n64973 , n64974 , n64975 , n64976 , n64977 , n64978 , n64979 , 
     n64980 , n64981 , n64982 , n64983 , n64984 , n64985 , n64986 , n64987 , n64988 , n64989 , 
     n64990 , n64991 , n64992 , n64993 , n64994 , n592318 , n592319 , n64997 , n64998 , n64999 , 
     n592323 , n65001 , n65002 , n65003 , n592327 , n592328 , n65006 , n592330 , n65008 , n65009 , 
     n65010 , n592334 , n592335 , n65013 , n592337 , n65015 , n592339 , n592340 , n65018 , n592342 , 
     n65020 , n65021 , n65022 , n65023 , n592347 , n65025 , n592349 , n65027 , n592351 , n592352 , 
     n65030 , n592354 , n65032 , n65033 , n65034 , n65035 , n65036 , n592360 , n65038 , n592362 , 
     n65040 , n65041 , n65042 , n592366 , n592367 , n65045 , n592369 , n592370 , n65048 , n592372 , 
     n65050 , n65051 , n65052 , n65053 , n65054 , n65055 , n65056 , n65057 , n65058 , n65059 , 
     n592383 , n592384 , n65062 , n592386 , n65064 , n65065 , n65066 , n65067 , n65068 , n592392 , 
     n592393 , n65071 , n592395 , n592396 , n65074 , n592398 , n592399 , n65077 , n592401 , n65079 , 
     n65080 , n592404 , n65082 , n592406 , n65084 , n592408 , n592409 , n65087 , n592411 , n65089 , 
     n65090 , n65091 , n65092 , n65093 , n592417 , n592418 , n65096 , n592420 , n592421 , n65099 , 
     n592423 , n65101 , n65102 , n65103 , n65104 , n592428 , n65106 , n592430 , n592431 , n592432 , 
     n65110 , n592434 , n592435 , n65113 , n592437 , n65115 , n65116 , n592440 , n65118 , n592442 , 
     n65120 , n65121 , n65122 , n592446 , n65124 , n592448 , n65126 , n592450 , n592451 , n592452 , 
     n65130 , n592454 , n592455 , n65133 , n592457 , n592458 , n592459 , n592460 , n592461 , n592462 , 
     n65140 , n592464 , n592465 , n65143 , n592467 , n592468 , n65146 , n592470 , n592471 , n65149 , 
     n592473 , n65151 , n592475 , n65153 , n592477 , n592478 , n65156 , n592480 , n592481 , n65159 , 
     n592483 , n592484 , n65162 , n592486 , n65164 , n65165 , n65166 , n65167 , n65168 , n65169 , 
     n65170 , n65171 , n65172 , n65173 , n65174 , n65175 , n65176 , n65177 , n65178 , n65179 , 
     n65180 , n65181 , n65182 , n65183 , n65184 , n65185 , n65186 , n65187 , n65188 , n65189 , 
     n65190 , n65191 , n65192 , n65193 , n65194 , n65195 , n65196 , n65197 , n65198 , n65199 , 
     n65200 , n65201 , n65202 , n65203 , n65204 , n65205 , n65206 , n65207 , n65208 , n65209 , 
     n65210 , n65211 , n65212 , n65213 , n65214 , n592538 , n65216 , n65217 , n65218 , n65219 , 
     n65220 , n65221 , n65222 , n65223 , n592547 , n65225 , n592549 , n65227 , n65228 , n65229 , 
     n65230 , n65231 , n65232 , n65233 , n65234 , n65235 , n65236 , n65237 , n592561 , n65239 , 
     n592563 , n592564 , n65242 , n65243 , n592567 , n65245 , n592569 , n65247 , n592571 , n592572 , 
     n65250 , n592574 , n592575 , n65253 , n65254 , n592578 , n65256 , n65257 , n592581 , n65259 , 
     n592583 , n65261 , n592585 , n65263 , n592587 , n592588 , n65266 , n592590 , n592591 , n65269 , 
     n592593 , n592594 , n65272 , n592596 , n592597 , n65275 , n65276 , n65277 , n65278 , n65279 , 
     n65280 , n65281 , n65282 , n65283 , n65284 , n592608 , n65286 , n592610 , n592611 , n65289 , 
     n592613 , n65291 , n592615 , n65293 , n592617 , n592618 , n65296 , n592620 , n65298 , n65299 , 
     n592623 , n65301 , n592625 , n592626 , n592627 , n592628 , n65306 , n592630 , n592631 , n592632 , 
     n65310 , n592634 , n592635 , n65313 , n592637 , n592638 , n592639 , n65317 , n592641 , n592642 , 
     n65320 , n592644 , n592645 , n65323 , n592647 , n592648 , n65326 , n592650 , n592651 , n65329 , 
     n592653 , n65331 , n65332 , n65333 , n65334 , n65335 , n592659 , n65337 , n592661 , n65339 , 
     n65340 , n592664 , n65342 , n65343 , n592667 , n592668 , n592669 , n65347 , n592671 , n592672 , 
     n65350 , n592674 , n592675 , n65353 , n592677 , n592678 , n65356 , n592680 , n592681 , n65359 , 
     n592683 , n592684 , n65362 , n592686 , n592687 , n65365 , n592689 , n65367 , n65368 , n65369 , 
     n65370 , n65371 , n65372 , n65373 , n65374 , n65375 , n65376 , n65377 , n65378 , n65379 , 
     n65380 , n65381 , n65382 , n65383 , n65384 , n65385 , n65386 , n65387 , n65388 , n65389 , 
     n65390 , n592714 , n65392 , n592716 , n592717 , n65395 , n65396 , n65397 , n592721 , n65399 , 
     n592723 , n65401 , n65402 , n65403 , n65404 , n592728 , n65406 , n65407 , n65408 , n65409 , 
     n592733 , n65411 , n592735 , n65413 , n65414 , n65415 , n65416 , n592740 , n65418 , n592742 , 
     n65420 , n592744 , n65422 , n592746 , n65424 , n592748 , n592749 , n592750 , n65428 , n592752 , 
     n592753 , n65431 , n65432 , n592756 , n65434 , n65435 , n592759 , n592760 , n65438 , n592762 , 
     n592763 , n65441 , n65442 , n592766 , n592767 , n65445 , n65446 , n592770 , n65448 , n65449 , 
     n592773 , n592774 , n65452 , n65453 , n592777 , n592778 , n65456 , n592780 , n65458 , n65459 , 
     n592783 , n65461 , n592785 , n65463 , n592787 , n592788 , n65466 , n592790 , n65468 , n65469 , 
     n592793 , n65471 , n65472 , n592796 , n65474 , n592798 , n592799 , n65477 , n65478 , n592802 , 
     n592803 , n65481 , n592805 , n592806 , n65484 , n592808 , n65486 , n65487 , n592811 , n592812 , 
     n65490 , n592814 , n65492 , n65493 , n65494 , n65495 , n65496 , n65497 , n65498 , n65499 , 
     n592823 , n65501 , n592825 , n65503 , n65504 , n65505 , n65506 , n65507 , n592831 , n65509 , 
     n592833 , n592834 , n592835 , n65513 , n592837 , n592838 , n65516 , n592840 , n592841 , n65519 , 
     n65520 , n65521 , n65522 , n65523 , n65524 , n65525 , n65526 , n65527 , n65528 , n65529 , 
     n65530 , n65531 , n65532 , n65533 , n592857 , n65535 , n592859 , n65537 , n592861 , n592862 , 
     n592863 , n65541 , n65542 , n65543 , n592867 , n65545 , n592869 , n65547 , n65548 , n65549 , 
     n65550 , n65551 , n65552 , n65553 , n65554 , n65555 , n65556 , n65557 , n65558 , n65559 , 
     n592883 , n65561 , n592885 , n65563 , n592887 , n65565 , n65566 , n65567 , n65568 , n65569 , 
     n65570 , n65571 , n65572 , n592896 , n592897 , n65575 , n592899 , n592900 , n65578 , n592902 , 
     n65580 , n65581 , n592905 , n592906 , n65584 , n592908 , n65586 , n592910 , n592911 , n65589 , 
     n592913 , n592914 , n65592 , n592916 , n65594 , n592918 , n592919 , n65597 , n592921 , n592922 , 
     n592923 , n65601 , n592925 , n592926 , n592927 , n65605 , n592929 , n592930 , n65608 , n592932 , 
     n592933 , n65611 , n592935 , n65613 , n65614 , n65615 , n592939 , n592940 , n65618 , n592942 , 
     n592943 , n592944 , n65622 , n592946 , n592947 , n65625 , n592949 , n592950 , n65628 , n592952 , 
     n65630 , n592954 , n592955 , n65633 , n592957 , n65635 , n65636 , n592960 , n65638 , n592962 , 
     n65640 , n65641 , n592965 , n592966 , n592967 , n65645 , n592969 , n592970 , n65648 , n65649 , 
     n65650 , n592974 , n65652 , n592976 , n65654 , n65655 , n65656 , n65657 , n65658 , n65659 , 
     n592983 , n592984 , n65662 , n592986 , n65664 , n65665 , n592989 , n65667 , n592991 , n592992 , 
     n65670 , n592994 , n592995 , n65673 , n65674 , n65675 , n65676 , n593000 , n593001 , n65679 , 
     n593003 , n593004 , n65682 , n593006 , n593007 , n65685 , n593009 , n593010 , n65688 , n593012 , 
     n65690 , n65691 , n65692 , n65693 , n65694 , n65695 , n593019 , n65697 , n593021 , n593022 , 
     n65700 , n593024 , n593025 , n65703 , n593027 , n65705 , n65706 , n593030 , n65708 , n593032 , 
     n65710 , n65711 , n65712 , n593036 , n593037 , n65715 , n593039 , n65717 , n65718 , n593042 , 
     n593043 , n65721 , n593045 , n593046 , n65724 , n593048 , n65726 , n65727 , n65728 , n65729 , 
     n593053 , n65731 , n593055 , n65733 , n65734 , n65735 , n65736 , n65737 , n65738 , n65739 , 
     n65740 , n65741 , n65742 , n65743 , n65744 , n65745 , n65746 , n65747 , n65748 , n65749 , 
     n65750 , n65751 , n65752 , n65753 , n65754 , n65755 , n65756 , n65757 , n65758 , n65759 , 
     n65760 , n65761 , n65762 , n65763 , n65764 , n65765 , n65766 , n65767 , n65768 , n65769 , 
     n65770 , n65771 , n65772 , n65773 , n65774 , n65775 , n65776 , n65777 , n65778 , n65779 , 
     n65780 , n65781 , n65782 , n593106 , n65784 , n65785 , n65786 , n65787 , n65788 , n65789 , 
     n65790 , n65791 , n65792 , n65793 , n65794 , n593118 , n65796 , n593120 , n593121 , n65799 , 
     n65800 , n65801 , n65802 , n593126 , n65804 , n593128 , n593129 , n65807 , n593131 , n593132 , 
     n65810 , n593134 , n593135 , n65813 , n593137 , n65815 , n593139 , n593140 , n65818 , n593142 , 
     n593143 , n65821 , n65822 , n65823 , n65824 , n65825 , n65826 , n65827 , n65828 , n65829 , 
     n65830 , n593154 , n65832 , n593156 , n65834 , n65835 , n593159 , n593160 , n65838 , n593162 , 
     n65840 , n65841 , n65842 , n65843 , n65844 , n65845 , n65846 , n65847 , n65848 , n593172 , 
     n593173 , n65851 , n593175 , n593176 , n593177 , n593178 , n65856 , n593180 , n593181 , n65859 , 
     n593183 , n593184 , n65862 , n593186 , n593187 , n65865 , n593189 , n65867 , n65868 , n65869 , 
     n593193 , n65871 , n593195 , n593196 , n65874 , n593198 , n65876 , n65877 , n65878 , n65879 , 
     n65880 , n65881 , n65882 , n65883 , n593207 , n65885 , n593209 , n65887 , n65888 , n593212 , 
     n65890 , n593214 , n593215 , n65893 , n593217 , n65895 , n593219 , n593220 , n65898 , n593222 , 
     n593223 , n65901 , n593225 , n593226 , n65904 , n593228 , n593229 , n65907 , n593231 , n593232 , 
     n65910 , n593234 , n593235 , n65913 , n593237 , n65915 , n65916 , n65917 , n65918 , n65919 , 
     n593243 , n593244 , n65922 , n593246 , n65924 , n65925 , n65926 , n65927 , n65928 , n65929 , 
     n65930 , n593254 , n65932 , n593256 , n65934 , n593258 , n593259 , n65937 , n593261 , n65939 , 
     n65940 , n593264 , n65942 , n593266 , n593267 , n65945 , n65946 , n593270 , n65948 , n65949 , 
     n593273 , n593274 , n65952 , n593276 , n593277 , n65955 , n593279 , n65957 , n65958 , n65959 , 
     n65960 , n593284 , n65962 , n593286 , n593287 , n593288 , n593289 , n65967 , n593291 , n593292 , 
     n65970 , n593294 , n593295 , n65973 , n593297 , n593298 , n65976 , n593300 , n65978 , n593302 , 
     n65980 , n593304 , n65982 , n65983 , n65984 , n65985 , n65986 , n65987 , n65988 , n593312 , 
     n65990 , n65991 , n593315 , n593316 , n593317 , n65995 , n593319 , n593320 , n65998 , n593322 , 
     n593323 , n66001 , n593325 , n593326 , n66004 , n593328 , n593329 , n66007 , n593331 , n66009 , 
     n66010 , n593334 , n66012 , n593336 , n593337 , n66015 , n593339 , n593340 , n66018 , n593342 , 
     n593343 , n66021 , n593345 , n66023 , n66024 , n593348 , n66026 , n593350 , n66028 , n66029 , 
     n66030 , n66031 , n66032 , n66033 , n593357 , n66035 , n593359 , n66037 , n593361 , n593362 , 
     n66040 , n593364 , n593365 , n66043 , n593367 , n593368 , n66046 , n593370 , n593371 , n66049 , 
     n593373 , n66051 , n66052 , n66053 , n66054 , n593378 , n66056 , n593380 , n66058 , n66059 , 
     n593383 , n66061 , n593385 , n66063 , n66064 , n66065 , n66066 , n66067 , n593391 , n593392 , 
     n66070 , n593394 , n593395 , n66073 , n593397 , n593398 , n593399 , n66077 , n593401 , n66079 , 
     n593403 , n66081 , n593405 , n593406 , n66084 , n593408 , n66086 , n66087 , n66088 , n593412 , 
     n66090 , n593414 , n593415 , n593416 , n593417 , n66095 , n593419 , n593420 , n66098 , n593422 , 
     n66100 , n593424 , n593425 , n593426 , n66104 , n593428 , n593429 , n66107 , n593431 , n593432 , 
     n66110 , n593434 , n66112 , n66113 , n593437 , n66115 , n593439 , n593440 , n593441 , n66119 , 
     n593443 , n66121 , n593445 , n66123 , n593447 , n66125 , n66126 , n66127 , n66128 , n593452 , 
     n593453 , n66131 , n593455 , n593456 , n66134 , n593458 , n593459 , n593460 , n66138 , n593462 , 
     n66140 , n66141 , n66142 , n66143 , n66144 , n66145 , n66146 , n66147 , n593471 , n66149 , 
     n593473 , n66151 , n593475 , n66153 , n593477 , n593478 , n593479 , n66157 , n593481 , n66159 , 
     n593483 , n66161 , n593485 , n66163 , n593487 , n66165 , n593489 , n593490 , n66168 , n593492 , 
     n66170 , n593494 , n66172 , n593496 , n593497 , n593498 , n66176 , n593500 , n66178 , n593502 , 
     n593503 , n66181 , n593505 , n66183 , n66184 , n66185 , n66186 , n66187 , n66188 , n593512 , 
     n66190 , n593514 , n593515 , n66193 , n593517 , n66195 , n593519 , n593520 , n66198 , n593522 , 
     n593523 , n593524 , n593525 , n66203 , n593527 , n593528 , n66206 , n593530 , n66208 , n593532 , 
     n593533 , n66211 , n593535 , n593536 , n66214 , n593538 , n593539 , n66217 , n593541 , n66219 , 
     n66220 , n66221 , n593545 , n593546 , n66224 , n593548 , n66226 , n593550 , n593551 , n66229 , 
     n593553 , n593554 , n66232 , n593556 , n593557 , n66235 , n593559 , n66237 , n593561 , n593562 , 
     n66240 , n593564 , n66242 , n593566 , n66244 , n593568 , n593569 , n66247 , n66248 , n66249 , 
     n66250 , n593574 , n593575 , n66253 , n593577 , n66255 , n593579 , n593580 , n66258 , n593582 , 
     n66260 , n66261 , n66262 , n66263 , n66264 , n593588 , n66266 , n593590 , n593591 , n593592 , 
     n593593 , n593594 , n66272 , n593596 , n593597 , n66275 , n66276 , n593600 , n66278 , n593602 , 
     n593603 , n66281 , n593605 , n593606 , n66284 , n593608 , n66286 , n593610 , n66288 , n593612 , 
     n593613 , n66291 , n593615 , n593616 , n66294 , n66295 , n593619 , n593620 , n66298 , n593622 , 
     n66300 , n593624 , n66302 , n593626 , n593627 , n66305 , n66306 , n593630 , n66308 , n593632 , 
     n593633 , n66311 , n593635 , n593636 , n66314 , n593638 , n593639 , n593640 , n66318 , n593642 , 
     n593643 , n593644 , n66322 , n593646 , n593647 , n66325 , n593649 , n593650 , n66328 , n593652 , 
     n593653 , n593654 , n593655 , n593656 , n66334 , n66335 , n593659 , n593660 , n66338 , n593662 , 
     n593663 , n66341 , n593665 , n66343 , n593667 , n593668 , n593669 , n593670 , n593671 , n66349 , 
     n66350 , n66351 , n66352 , n66353 , n593677 , n593678 , n593679 , n593680 , n66358 , n593682 , 
     n593683 , n66361 , n593685 , n593686 , n593687 , n66365 , n593689 , n593690 , n66368 , n593692 , 
     n593693 , n593694 , n593695 , n66373 , n593697 , n593698 , n593699 , n66377 , n593701 , n593702 , 
     n593703 , n66381 , n593705 , n66383 , n66384 , n593708 , n593709 , n593710 , n66388 , n593712 , 
     n66390 , n593714 , n593715 , n593716 , n66394 , n593718 , n66396 , n593720 , n66398 , n593722 , 
     n593723 , n593724 , n66402 , n593726 , n66404 , n66405 , n66406 , n66407 , n66408 , n593732 , 
     n66410 , n593734 , n593735 , n593736 , n66414 , n593738 , n593739 , n593740 , n593741 , n66419 , 
     n593743 , n593744 , n593745 , n593746 , n66424 , n593748 , n593749 , n593750 , n593751 , n66429 , 
     n593753 , n593754 , n593755 , n66433 , n593757 , n66435 , n593759 , n66437 , n593761 , n593762 , 
     n593763 , n593764 , n66442 , n593766 , n593767 , n593768 , n66446 , n593770 , n66448 , n66449 , 
     n593773 , n66451 , n593775 , n593776 , n66454 , n593778 , n593779 , n66457 , n593781 , n593782 , 
     n593783 , n66461 , n593785 , n593786 , n593787 , n66465 , n593789 , n593790 , n66468 , n593792 , 
     n593793 , n66471 , n593795 , n66473 , n593797 , n593798 , n66476 , n593800 , n593801 , n66479 , 
     n593803 , n66481 , n593805 , n593806 , n593807 , n66485 , n593809 , n593810 , n66488 , n66489 , 
     n593813 , n593814 , n593815 , n66493 , n593817 , n66495 , n593819 , n593820 , n593821 , n66499 , 
     n593823 , n593824 , n66502 , n66503 , n593827 , n593828 , n593829 , n66507 , n593831 , n593832 , 
     n66510 , n593834 , n593835 , n66513 , n66514 , n66515 , n66516 , n66517 , n66518 , n593842 , 
     n593843 , n66521 , n593845 , n593846 , n593847 , n66525 , n593849 , n593850 , n66528 , n66529 , 
     n66530 , n66531 , n593855 , n593856 , n66534 , n593858 , n66536 , n593860 , n593861 , n593862 , 
     n66540 , n593864 , n593865 , n66543 , n593867 , n593868 , n66546 , n593870 , n593871 , n593872 , 
     n66550 , n593874 , n66552 , n593876 , n66554 , n593878 , n593879 , n593880 , n66558 , n593882 , 
     n66560 , n593884 , n593885 , n66563 , n593887 , n66565 , n593889 , n66567 , n66568 , n66569 , 
     n66570 , n593894 , n593895 , n66573 , n593897 , n66575 , n593899 , n593900 , n593901 , n66579 , 
     n593903 , n593904 , n593905 , n66583 , n593907 , n66585 , n593909 , n593910 , n593911 , n593912 , 
     n593913 , n66591 , n593915 , n593916 , n66594 , n593918 , n593919 , n593920 , n66598 , n593922 , 
     n593923 , n593924 , n593925 , n66603 , n593927 , n593928 , n66606 , n66607 , n66608 , n66609 , 
     n593933 , n593934 , n593935 , n593936 , n66614 , n66615 , n593939 , n593940 , n593941 , n66619 , 
     n593943 , n593944 , n593945 , n66623 , n593947 , n593948 , n66626 , n593950 , n593951 , n593952 , 
     n66630 , n593954 , n593955 , n66633 , n593957 , n593958 , n593959 , n66637 , n593961 , n593962 , 
     n66640 , n593964 , n66642 , n66643 , n593967 , n66645 , n593969 , n593970 , n66648 , n593972 , 
     n66650 , n593974 , n593975 , n66653 , n593977 , n593978 , n66656 , n66657 , n66658 , n66659 , 
     n66660 , n593984 , n66662 , n593986 , n593987 , n593988 , n593989 , n66667 , n593991 , n66669 , 
     n66670 , n593994 , n66672 , n593996 , n593997 , n66675 , n593999 , n594000 , n594001 , n66679 , 
     n594003 , n594004 , n594005 , n66683 , n594007 , n594008 , n594009 , n66687 , n594011 , n594012 , 
     n594013 , n66691 , n594015 , n66693 , n594017 , n594018 , n66696 , n594020 , n66698 , n66699 , 
     n594023 , n594024 , n66702 , n594026 , n594027 , n594028 , n66706 , n594030 , n594031 , n594032 , 
     n66710 , n594034 , n594035 , n594036 , n66714 , n594038 , n594039 , n66717 , n66718 , n594042 , 
     n66720 , n594044 , n594045 , n594046 , n66724 , n594048 , n594049 , n66727 , n594051 , n594052 , 
     n66730 , n66731 , n594055 , n66733 , n66734 , n66735 , n66736 , n66737 , n66738 , n66739 , 
     n66740 , n66741 , n66742 , n66743 , n594067 , n66745 , n66746 , n66747 , n66748 , n66749 , 
     n66750 , n66751 , n66752 , n66753 , n66754 , n66755 , n66756 , n66757 , n66758 , n66759 , 
     n66760 , n66761 , n66762 , n66763 , n66764 , n66765 , n66766 , n66767 , n66768 , n66769 , 
     n66770 , n66771 , n66772 , n66773 , n66774 , n66775 , n66776 , n594100 , n66778 , n594102 , 
     n594103 , n66781 , n594105 , n594106 , n66784 , n66785 , n66786 , n66787 , n594111 , n66789 , 
     n594113 , n594114 , n594115 , n66793 , n594117 , n594118 , n66796 , n594120 , n594121 , n66799 , 
     n594123 , n594124 , n66802 , n66803 , n594127 , n594128 , n66806 , n594130 , n66808 , n66809 , 
     n594133 , n594134 , n66812 , n594136 , n66814 , n594138 , n66816 , n66817 , n594141 , n594142 , 
     n66820 , n594144 , n594145 , n66823 , n594147 , n594148 , n594149 , n66827 , n594151 , n594152 , 
     n66830 , n594154 , n594155 , n66833 , n594157 , n594158 , n66836 , n594160 , n66838 , n594162 , 
     n594163 , n66841 , n594165 , n66843 , n66844 , n66845 , n66846 , n66847 , n66848 , n66849 , 
     n594173 , n66851 , n594175 , n66853 , n594177 , n594178 , n594179 , n66857 , n594181 , n594182 , 
     n66860 , n66861 , n594185 , n66863 , n594187 , n66865 , n66866 , n594190 , n66868 , n66869 , 
     n66870 , n66871 , n594195 , n594196 , n594197 , n66875 , n66876 , n66877 , n594201 , n594202 , 
     n66880 , n594204 , n594205 , n66883 , n66884 , n66885 , n66886 , n594210 , n594211 , n66889 , 
     n594213 , n594214 , n66892 , n594216 , n594217 , n66895 , n594219 , n594220 , n66898 , n594222 , 
     n594223 , n594224 , n66902 , n594226 , n66904 , n66905 , n66906 , n66907 , n66908 , n66909 , 
     n594233 , n66911 , n594235 , n66913 , n66914 , n594238 , n594239 , n66917 , n594241 , n594242 , 
     n66920 , n594244 , n594245 , n66923 , n594247 , n594248 , n66926 , n594250 , n594251 , n66929 , 
     n66930 , n594254 , n594255 , n66933 , n594257 , n594258 , n594259 , n594260 , n66938 , n594262 , 
     n66940 , n66941 , n594265 , n66943 , n594267 , n594268 , n66946 , n66947 , n594271 , n594272 , 
     n594273 , n66951 , n594275 , n594276 , n66954 , n594278 , n594279 , n594280 , n66958 , n594282 , 
     n594283 , n594284 , n66962 , n594286 , n66964 , n594288 , n594289 , n66967 , n594291 , n594292 , 
     n66970 , n594294 , n594295 , n66973 , n594297 , n594298 , n66976 , n594300 , n594301 , n594302 , 
     n66980 , n594304 , n594305 , n594306 , n66984 , n594308 , n594309 , n66987 , n66988 , n594312 , 
     n594313 , n66991 , n594315 , n594316 , n594317 , n594318 , n66996 , n66997 , n594321 , n594322 , 
     n594323 , n594324 , n67002 , n594326 , n594327 , n67005 , n67006 , n594330 , n67008 , n67009 , 
     n594333 , n67011 , n594335 , n594336 , n594337 , n67015 , n594339 , n594340 , n67018 , n67019 , 
     n67020 , n67021 , n67022 , n594346 , n67024 , n594348 , n594349 , n67027 , n594351 , n594352 , 
     n594353 , n67031 , n594355 , n594356 , n594357 , n67035 , n594359 , n594360 , n67038 , n594362 , 
     n67040 , n67041 , n67042 , n594366 , n67044 , n594368 , n594369 , n67047 , n594371 , n594372 , 
     n67050 , n594374 , n594375 , n67053 , n594377 , n67055 , n594379 , n594380 , n67058 , n594382 , 
     n594383 , n67061 , n594385 , n594386 , n594387 , n67065 , n594389 , n594390 , n594391 , n67069 , 
     n594393 , n594394 , n594395 , n67073 , n594397 , n594398 , n67076 , n594400 , n594401 , n594402 , 
     n67080 , n594404 , n594405 , n67083 , n594407 , n594408 , n594409 , n67087 , n594411 , n594412 , 
     n594413 , n67091 , n594415 , n594416 , n594417 , n67095 , n594419 , n594420 , n67098 , n594422 , 
     n594423 , n67101 , n594425 , n594426 , n67104 , n594428 , n594429 , n67107 , n594431 , n594432 , 
     n67110 , n594434 , n594435 , n67113 , n594437 , n594438 , n67116 , n594440 , n594441 , n67119 , 
     n594443 , n594444 , n67122 , n594446 , n594447 , n67125 , n67126 , n67127 , n67128 , n594452 , 
     n594453 , n594454 , n594455 , n67133 , n67134 , n594458 , n594459 , n594460 , n67138 , n67139 , 
     n594463 , n594464 , n594465 , n67143 , n67144 , n594468 , n594469 , n594470 , n67148 , n67149 , 
     n594473 , n594474 , n594475 , n67153 , n67154 , n594478 , n594479 , n594480 , n67158 , n67159 , 
     n594483 , n594484 , n594485 , n67163 , n67164 , n594488 , n594489 , n594490 , n67168 , n67169 , 
     n594493 , n594494 , n594495 , n67173 , n67174 , n594498 , n594499 , n594500 , n67178 , n67179 , 
     n594503 , n67181 , n67182 , n67183 , n67184 , n594508 , n67186 , n594510 , n594511 , n67189 , 
     n594513 , n594514 , n67192 , n594516 , n67194 , n67195 , n67196 , n67197 , n67198 , n67199 , 
     n67200 , n67201 , n67202 , n594526 , n67204 , n594528 , n594529 , n67207 , n67208 , n594532 , 
     n67210 , n594534 , n594535 , n67213 , n594537 , n67215 , n594539 , n594540 , n67218 , n594542 , 
     n594543 , n67221 , n67222 , n594546 , n67224 , n67225 , n67226 , n67227 , n67228 , n67229 , 
     n67230 , n67231 , n67232 , n67233 , n67234 , n594558 , n67236 , n594560 , n594561 , n67239 , 
     n67240 , n67241 , n67242 , n67243 , n67244 , n67245 , n594569 , n67247 , n594571 , n594572 , 
     n67250 , n594574 , n594575 , n67253 , n594577 , n594578 , n67256 , n67257 , n67258 , n594582 , 
     n67260 , n594584 , n594585 , n67263 , n594587 , n67265 , n67266 , n67267 , n67268 , n67269 , 
     n67270 , n67271 , n67272 , n67273 , n67274 , n67275 , n67276 , n67277 , n594601 , n67279 , 
     n594603 , n594604 , n67282 , n594606 , n594607 , n67285 , n594609 , n594610 , n67288 , n594612 , 
     n594613 , n67291 , n67292 , n594616 , n67294 , n594618 , n594619 , n67297 , n594621 , n594622 , 
     n594623 , n67301 , n594625 , n594626 , n67304 , n594628 , n594629 , n67307 , n67308 , n594632 , 
     n67310 , n67311 , n67312 , n67313 , n67314 , n67315 , n67316 , n67317 , n67318 , n67319 , 
     n67320 , n67321 , n594645 , n67323 , n594647 , n594648 , n67326 , n67327 , n594651 , n594652 , 
     n67330 , n594654 , n594655 , n67333 , n594657 , n594658 , n594659 , n594660 , n67338 , n594662 , 
     n594663 , n594664 , n67342 , n594666 , n594667 , n67345 , n594669 , n594670 , n67348 , n594672 , 
     n594673 , n67351 , n594675 , n594676 , n67354 , n594678 , n594679 , n67357 , n67358 , n67359 , 
     n67360 , n67361 , n67362 , n67363 , n67364 , n67365 , n67366 , n594690 , n67368 , n594692 , 
     n67370 , n594694 , n67372 , n67373 , n67374 , n67375 , n67376 , n67377 , n67378 , n67379 , 
     n67380 , n67381 , n67382 , n67383 , n67384 , n67385 , n67386 , n594710 , n67388 , n67389 , 
     n67390 , n67391 , n594715 , n67393 , n594717 , n67395 , n594719 , n594720 , n67398 , n594722 , 
     n67400 , n67401 , n594725 , n67403 , n67404 , n67405 , n67406 , n67407 , n67408 , n67409 , 
     n67410 , n67411 , n67412 , n67413 , n594737 , n67415 , n594739 , n594740 , n67418 , n594742 , 
     n594743 , n67421 , n67422 , n594746 , n67424 , n594748 , n594749 , n594750 , n67428 , n594752 , 
     n594753 , n67431 , n594755 , n67433 , n594757 , n67435 , n594759 , n67437 , n67438 , n594762 , 
     n67440 , n594764 , n594765 , n67443 , n67444 , n67445 , n67446 , n67447 , n67448 , n67449 , 
     n594773 , n67451 , n594775 , n594776 , n67454 , n594778 , n67456 , n67457 , n67458 , n67459 , 
     n67460 , n67461 , n67462 , n67463 , n67464 , n67465 , n67466 , n67467 , n67468 , n67469 , 
     n67470 , n594794 , n67472 , n67473 , n67474 , n594798 , n594799 , n67477 , n594801 , n594802 , 
     n67480 , n594804 , n594805 , n67483 , n594807 , n594808 , n67486 , n67487 , n67488 , n67489 , 
     n594813 , n67491 , n594815 , n594816 , n67494 , n594818 , n594819 , n67497 , n594821 , n594822 , 
     n67500 , n594824 , n67502 , n67503 , n67504 , n67505 , n67506 , n67507 , n67508 , n67509 , 
     n67510 , n67511 , n67512 , n594836 , n67514 , n67515 , n67516 , n594840 , n594841 , n67519 , 
     n594843 , n594844 , n67522 , n594846 , n594847 , n67525 , n594849 , n594850 , n67528 , n594852 , 
     n594853 , n67531 , n594855 , n594856 , n67534 , n594858 , n594859 , n67537 , n594861 , n594862 , 
     n67540 , n594864 , n594865 , n67543 , n594867 , n594868 , n67546 , n67547 , n594871 , n594872 , 
     n67550 , n594874 , n594875 , n67553 , n594877 , n594878 , n67556 , n67557 , n67558 , n594882 , 
     n67560 , n67561 , n67562 , n67563 , n67564 , n67565 , n67566 , n67567 , n67568 , n67569 , 
     n594893 , n67571 , n67572 , n67573 , n594897 , n67575 , n594899 , n594900 , n67578 , n67579 , 
     n594903 , n594904 , n67582 , n67583 , n594907 , n67585 , n67586 , n67587 , n67588 , n67589 , 
     n67590 , n594914 , n67592 , n594916 , n67594 , n67595 , n594919 , n67597 , n594921 , n67599 , 
     n67600 , n67601 , n67602 , n67603 , n67604 , n67605 , n594929 , n67607 , n594931 , n594932 , 
     n67610 , n594934 , n594935 , n67613 , n67614 , n594938 , n67616 , n594940 , n594941 , n594942 , 
     n67620 , n594944 , n594945 , n67623 , n594947 , n594948 , n594949 , n67627 , n594951 , n594952 , 
     n67630 , n594954 , n594955 , n67633 , n594957 , n594958 , n67636 , n594960 , n594961 , n67639 , 
     n67640 , n594964 , n594965 , n67643 , n67644 , n67645 , n594969 , n594970 , n67648 , n67649 , 
     n594973 , n67651 , n67652 , n594976 , n67654 , n67655 , n594979 , n67657 , n594981 , n594982 , 
     n67660 , n594984 , n67662 , n594986 , n67664 , n594988 , n67666 , n67667 , n594991 , n67669 , 
     n594993 , n594994 , n67672 , n67673 , n67674 , n594998 , n67676 , n67677 , n595001 , n67679 , 
     n595003 , n595004 , n67682 , n595006 , n595007 , n67685 , n595009 , n595010 , n67688 , n67689 , 
     n595013 , n67691 , n595015 , n595016 , n67694 , n67695 , n595019 , n67697 , n595021 , n595022 , 
     n67700 , n595024 , n595025 , n67703 , n67704 , n67705 , n595029 , n67707 , n595031 , n595032 , 
     n595033 , n67711 , n595035 , n595036 , n67714 , n595038 , n595039 , n67717 , n595041 , n595042 , 
     n67720 , n595044 , n595045 , n67723 , n595047 , n67725 , n595049 , n67727 , n67728 , n595052 , 
     n67730 , n595054 , n67732 , n67733 , n595057 , n67735 , n595059 , n67737 , n595061 , n595062 , 
     n67740 , n595064 , n595065 , n595066 , n67744 , n595068 , n595069 , n67747 , n595071 , n595072 , 
     n67750 , n595074 , n595075 , n67753 , n67754 , n595078 , n67756 , n67757 , n595081 , n595082 , 
     n67760 , n595084 , n595085 , n67763 , n595087 , n595088 , n67766 , n595090 , n67768 , n595092 , 
     n67770 , n595094 , n595095 , n67773 , n595097 , n595098 , n67776 , n67777 , n595101 , n67779 , 
     n595103 , n595104 , n67782 , n595106 , n67784 , n595108 , n595109 , n67787 , n595111 , n595112 , 
     n67790 , n67791 , n595115 , n67793 , n595117 , n67795 , n67796 , n595120 , n595121 , n67799 , 
     n595123 , n595124 , n67802 , n595126 , n595127 , n595128 , n595129 , n67807 , n595131 , n595132 , 
     n595133 , n67811 , n595135 , n595136 , n67814 , n595138 , n595139 , n67817 , n595141 , n595142 , 
     n67820 , n595144 , n595145 , n67823 , n595147 , n595148 , n67826 , n595150 , n595151 , n67829 , 
     n67830 , n67831 , n595155 , n595156 , n67834 , n595158 , n595159 , n67837 , n67838 , n595162 , 
     n67840 , n67841 , n595165 , n595166 , n595167 , n595168 , n67846 , n595170 , n595171 , n67849 , 
     n595173 , n595174 , n67852 , n595176 , n595177 , n67855 , n595179 , n67857 , n595181 , n67859 , 
     n595183 , n595184 , n595185 , n595186 , n67864 , n595188 , n595189 , n67867 , n595191 , n595192 , 
     n67870 , n595194 , n595195 , n67873 , n595197 , n67875 , n595199 , n67877 , n67878 , n67879 , 
     n67880 , n67881 , n67882 , n67883 , n67884 , n67885 , n67886 , n67887 , n67888 , n595212 , 
     n67890 , n595214 , n595215 , n67893 , n67894 , n67895 , n67896 , n67897 , n595221 , n67899 , 
     n595223 , n67901 , n595225 , n595226 , n67904 , n595228 , n595229 , n67907 , n67908 , n595232 , 
     n67910 , n595234 , n595235 , n595236 , n67914 , n595238 , n595239 , n67917 , n67918 , n595242 , 
     n595243 , n67921 , n67922 , n67923 , n595247 , n67925 , n595249 , n67927 , n595251 , n595252 , 
     n67930 , n67931 , n67932 , n595256 , n595257 , n595258 , n595259 , n67937 , n595261 , n595262 , 
     n67940 , n67941 , n595265 , n67943 , n67944 , n595268 , n595269 , n595270 , n595271 , n67949 , 
     n595273 , n595274 , n67952 , n595276 , n595277 , n67955 , n595279 , n67957 , n67958 , n595282 , 
     n67960 , n595284 , n595285 , n67963 , n595287 , n67965 , n67966 , n595290 , n67968 , n595292 , 
     n67970 , n595294 , n67972 , n67973 , n67974 , n67975 , n595299 , n67977 , n595301 , n595302 , 
     n595303 , n67981 , n595305 , n67983 , n595307 , n595308 , n67986 , n595310 , n67988 , n595312 , 
     n67990 , n67991 , n595315 , n67993 , n595317 , n595318 , n67996 , n595320 , n595321 , n595322 , 
     n68000 , n595324 , n595325 , n68003 , n595327 , n595328 , n68006 , n68007 , n595331 , n68009 , 
     n595333 , n68011 , n595335 , n595336 , n68014 , n595338 , n595339 , n68017 , n68018 , n595342 , 
     n595343 , n68021 , n595345 , n595346 , n68024 , n595348 , n595349 , n595350 , n68028 , n595352 , 
     n595353 , n68031 , n595355 , n595356 , n68034 , n595358 , n68036 , n595360 , n68038 , n68039 , 
     n595363 , n595364 , n68042 , n595366 , n595367 , n68045 , n595369 , n595370 , n595371 , n68049 , 
     n595373 , n68051 , n595375 , n68053 , n595377 , n595378 , n68056 , n595380 , n595381 , n68059 , 
     n595383 , n595384 , n68062 , n595386 , n595387 , n595388 , n68066 , n595390 , n68068 , n68069 , 
     n595393 , n595394 , n68072 , n595396 , n595397 , n68075 , n595399 , n595400 , n595401 , n68079 , 
     n595403 , n68081 , n68082 , n68083 , n68084 , n68085 , n68086 , n68087 , n68088 , n68089 , 
     n68090 , n68091 , n68092 , n68093 , n68094 , n68095 , n68096 , n68097 , n68098 , n68099 , 
     n68100 , n68101 , n595425 , n68103 , n595427 , n595428 , n68106 , n595430 , n595431 , n68109 , 
     n595433 , n595434 , n68112 , n68113 , n595437 , n68115 , n595439 , n595440 , n68118 , n595442 , 
     n595443 , n595444 , n68122 , n595446 , n595447 , n68125 , n595449 , n595450 , n68128 , n68129 , 
     n595453 , n595454 , n68132 , n595456 , n595457 , n68135 , n595459 , n595460 , n68138 , n68139 , 
     n68140 , n68141 , n68142 , n68143 , n595467 , n68145 , n595469 , n595470 , n68148 , n595472 , 
     n68150 , n595474 , n68152 , n595476 , n68154 , n68155 , n68156 , n68157 , n68158 , n68159 , 
     n68160 , n68161 , n68162 , n595486 , n595487 , n595488 , n68166 , n595490 , n595491 , n68169 , 
     n595493 , n595494 , n68172 , n68173 , n595497 , n68175 , n68176 , n595500 , n595501 , n68179 , 
     n595503 , n595504 , n68182 , n68183 , n68184 , n68185 , n68186 , n68187 , n68188 , n68189 , 
     n68190 , n595514 , n68192 , n595516 , n595517 , n68195 , n595519 , n595520 , n595521 , n68199 , 
     n595523 , n595524 , n68202 , n595526 , n595527 , n68205 , n68206 , n68207 , n68208 , n68209 , 
     n68210 , n595534 , n68212 , n595536 , n595537 , n68215 , n595539 , n595540 , n595541 , n68219 , 
     n68220 , n68221 , n68222 , n68223 , n68224 , n68225 , n68226 , n68227 , n68228 , n595552 , 
     n68230 , n595554 , n595555 , n68233 , n595557 , n595558 , n68236 , n595560 , n595561 , n68239 , 
     n68240 , n595564 , n595565 , n68243 , n595567 , n595568 , n68246 , n595570 , n595571 , n68249 , 
     n595573 , n595574 , n68252 , n595576 , n595577 , n68255 , n68256 , n68257 , n595581 , n595582 , 
     n68260 , n68261 , n595585 , n595586 , n68264 , n595588 , n595589 , n68267 , n595591 , n68269 , 
     n595593 , n68271 , n595595 , n68273 , n68274 , n595598 , n68276 , n68277 , n595601 , n595602 , 
     n68280 , n595604 , n595605 , n68283 , n595607 , n595608 , n68286 , n68287 , n595611 , n68289 , 
     n595613 , n595614 , n595615 , n68293 , n595617 , n595618 , n68296 , n595620 , n595621 , n595622 , 
     n68300 , n595624 , n595625 , n68303 , n595627 , n68305 , n68306 , n68307 , n595631 , n68309 , 
     n595633 , n595634 , n68312 , n68313 , n595637 , n68315 , n68316 , n595640 , n68318 , n595642 , 
     n68320 , n595644 , n68322 , n68323 , n68324 , n68325 , n68326 , n68327 , n68328 , n68329 , 
     n68330 , n68331 , n68332 , n68333 , n68334 , n68335 , n68336 , n68337 , n68338 , n68339 , 
     n68340 , n68341 , n68342 , n68343 , n68344 , n68345 , n68346 , n68347 , n68348 , n68349 , 
     n595673 , n68351 , n595675 , n595676 , n68354 , n595678 , n68356 , n68357 , n68358 , n68359 , 
     n68360 , n68361 , n68362 , n68363 , n68364 , n595688 , n68366 , n595690 , n595691 , n68369 , 
     n595693 , n68371 , n68372 , n68373 , n68374 , n68375 , n68376 , n68377 , n68378 , n68379 , 
     n68380 , n68381 , n68382 , n68383 , n68384 , n68385 , n68386 , n68387 , n595711 , n68389 , 
     n595713 , n68391 , n68392 , n68393 , n68394 , n68395 , n595719 , n68397 , n595721 , n68399 , 
     n595723 , n595724 , n68402 , n595726 , n68404 , n595728 , n68406 , n595730 , n595731 , n68409 , 
     n595733 , n595734 , n68412 , n595736 , n595737 , n595738 , n595739 , n68417 , n68418 , n595742 , 
     n68420 , n68421 , n595745 , n595746 , n68424 , n595748 , n595749 , n68427 , n595751 , n595752 , 
     n68430 , n68431 , n68432 , n68433 , n68434 , n68435 , n595759 , n68437 , n595761 , n68439 , 
     n595763 , n595764 , n68442 , n595766 , n595767 , n68445 , n68446 , n595770 , n68448 , n595772 , 
     n595773 , n68451 , n595775 , n595776 , n68454 , n595778 , n68456 , n595780 , n595781 , n68459 , 
     n595783 , n595784 , n68462 , n68463 , n595787 , n68465 , n68466 , n68467 , n68468 , n68469 , 
     n595793 , n595794 , n68472 , n595796 , n595797 , n595798 , n68476 , n595800 , n68478 , n68479 , 
     n68480 , n68481 , n68482 , n68483 , n68484 , n68485 , n68486 , n595810 , n68488 , n595812 , 
     n595813 , n68491 , n68492 , n595816 , n68494 , n595818 , n595819 , n595820 , n68498 , n595822 , 
     n595823 , n68501 , n595825 , n595826 , n595827 , n68505 , n595829 , n595830 , n68508 , n595832 , 
     n595833 , n68511 , n595835 , n595836 , n68514 , n595838 , n595839 , n68517 , n68518 , n68519 , 
     n595843 , n595844 , n68522 , n595846 , n595847 , n68525 , n595849 , n68527 , n595851 , n68529 , 
     n595853 , n68531 , n595855 , n595856 , n68534 , n68535 , n595859 , n595860 , n68538 , n595862 , 
     n595863 , n68541 , n595865 , n595866 , n68544 , n68545 , n595869 , n595870 , n68548 , n595872 , 
     n595873 , n68551 , n595875 , n68553 , n68554 , n595878 , n68556 , n68557 , n68558 , n68559 , 
     n68560 , n595884 , n68562 , n68563 , n595887 , n595888 , n68566 , n595890 , n595891 , n68569 , 
     n595893 , n68571 , n68572 , n68573 , n68574 , n68575 , n68576 , n68577 , n68578 , n68579 , 
     n68580 , n68581 , n68582 , n68583 , n68584 , n68585 , n68586 , n595910 , n68588 , n595912 , 
     n68590 , n68591 , n68592 , n68593 , n68594 , n595918 , n68596 , n595920 , n68598 , n595922 , 
     n595923 , n68601 , n595925 , n68603 , n68604 , n68605 , n68606 , n68607 , n68608 , n595932 , 
     n68610 , n68611 , n595935 , n595936 , n68614 , n595938 , n595939 , n68617 , n595941 , n68619 , 
     n595943 , n595944 , n68622 , n595946 , n595947 , n68625 , n595949 , n68627 , n595951 , n595952 , 
     n68630 , n595954 , n595955 , n68633 , n68634 , n595958 , n595959 , n68637 , n595961 , n595962 , 
     n68640 , n595964 , n595965 , n68643 , n595967 , n595968 , n68646 , n595970 , n68648 , n595972 , 
     n595973 , n68651 , n595975 , n68653 , n595977 , n595978 , n68656 , n68657 , n595981 , n595982 , 
     n68660 , n68661 , n595985 , n68663 , n595987 , n68665 , n595989 , n595990 , n68668 , n595992 , 
     n595993 , n68671 , n595995 , n595996 , n68674 , n68675 , n595999 , n68677 , n68678 , n596002 , 
     n596003 , n68681 , n596005 , n596006 , n68684 , n68685 , n596009 , n596010 , n68688 , n596012 , 
     n596013 , n68691 , n596015 , n68693 , n596017 , n68695 , n68696 , n68697 , n596021 , n596022 , 
     n68700 , n596024 , n596025 , n596026 , n68704 , n596028 , n68706 , n68707 , n596031 , n68709 , 
     n596033 , n596034 , n68712 , n596036 , n596037 , n596038 , n68716 , n596040 , n596041 , n68719 , 
     n596043 , n596044 , n68722 , n596046 , n596047 , n68725 , n596049 , n68727 , n68728 , n596052 , 
     n68730 , n596054 , n68732 , n596056 , n596057 , n68735 , n68736 , n596060 , n68738 , n596062 , 
     n68740 , n596064 , n596065 , n68743 , n596067 , n596068 , n596069 , n68747 , n68748 , n596072 , 
     n68750 , n596074 , n68752 , n68753 , n596077 , n68755 , n68756 , n596080 , n68758 , n68759 , 
     n68760 , n596084 , n68762 , n68763 , n596087 , n596088 , n68766 , n596090 , n596091 , n68769 , 
     n596093 , n68771 , n596095 , n68773 , n596097 , n596098 , n68776 , n596100 , n68778 , n596102 , 
     n68780 , n68781 , n68782 , n596106 , n68784 , n596108 , n68786 , n68787 , n596111 , n68789 , 
     n68790 , n596114 , n596115 , n68793 , n596117 , n596118 , n68796 , n596120 , n596121 , n68799 , 
     n68800 , n596124 , n68802 , n68803 , n596127 , n68805 , n596129 , n596130 , n68808 , n68809 , 
     n596133 , n596134 , n68812 , n596136 , n596137 , n68815 , n596139 , n596140 , n596141 , n68819 , 
     n596143 , n596144 , n68822 , n596146 , n596147 , n68825 , n68826 , n68827 , n596151 , n68829 , 
     n596153 , n68831 , n68832 , n596156 , n68834 , n596158 , n68836 , n68837 , n68838 , n68839 , 
     n68840 , n68841 , n68842 , n68843 , n68844 , n68845 , n596169 , n68847 , n596171 , n596172 , 
     n596173 , n68851 , n596175 , n596176 , n68854 , n596178 , n596179 , n68857 , n596181 , n68859 , 
     n596183 , n68861 , n596185 , n68863 , n596187 , n596188 , n68866 , n596190 , n596191 , n68869 , 
     n596193 , n596194 , n68872 , n68873 , n596197 , n596198 , n68876 , n596200 , n596201 , n68879 , 
     n596203 , n596204 , n68882 , n68883 , n596207 , n596208 , n68886 , n596210 , n68888 , n596212 , 
     n596213 , n68891 , n68892 , n596216 , n596217 , n68895 , n596219 , n596220 , n68898 , n596222 , 
     n596223 , n68901 , n596225 , n596226 , n68904 , n596228 , n596229 , n68907 , n596231 , n596232 , 
     n68910 , n596234 , n596235 , n68913 , n68914 , n596238 , n68916 , n596240 , n68918 , n596242 , 
     n596243 , n68921 , n596245 , n68923 , n596247 , n596248 , n68926 , n68927 , n596251 , n68929 , 
     n596253 , n596254 , n68932 , n596256 , n596257 , n596258 , n68936 , n596260 , n68938 , n596262 , 
     n68940 , n596264 , n596265 , n68943 , n596267 , n596268 , n68946 , n68947 , n596271 , n596272 , 
     n68950 , n596274 , n596275 , n68953 , n596277 , n596278 , n68956 , n68957 , n596281 , n68959 , 
     n596283 , n68961 , n68962 , n596286 , n596287 , n68965 , n596289 , n596290 , n68968 , n596292 , 
     n596293 , n596294 , n68972 , n596296 , n596297 , n68975 , n596299 , n596300 , n68978 , n596302 , 
     n68980 , n596304 , n68982 , n596306 , n68984 , n596308 , n596309 , n68987 , n596311 , n596312 , 
     n68990 , n68991 , n596315 , n596316 , n68994 , n596318 , n596319 , n68997 , n596321 , n596322 , 
     n69000 , n69001 , n596325 , n69003 , n596327 , n69005 , n69006 , n596330 , n596331 , n69009 , 
     n596333 , n596334 , n69012 , n596336 , n596337 , n596338 , n69016 , n596340 , n596341 , n69019 , 
     n596343 , n596344 , n69022 , n69023 , n596347 , n69025 , n596349 , n596350 , n69028 , n596352 , 
     n69030 , n596354 , n596355 , n69033 , n69034 , n69035 , n69036 , n69037 , n69038 , n69039 , 
     n69040 , n69041 , n69042 , n69043 , n69044 , n596368 , n69046 , n596370 , n596371 , n69049 , 
     n596373 , n596374 , n69052 , n596376 , n596377 , n69055 , n596379 , n596380 , n596381 , n69059 , 
     n596383 , n596384 , n596385 , n69063 , n596387 , n69065 , n69066 , n69067 , n596391 , n596392 , 
     n596393 , n69071 , n596395 , n596396 , n69074 , n596398 , n596399 , n69077 , n596401 , n69079 , 
     n596403 , n69081 , n596405 , n69083 , n596407 , n596408 , n69086 , n69087 , n596411 , n596412 , 
     n69090 , n596414 , n596415 , n69093 , n596417 , n596418 , n69096 , n69097 , n596421 , n596422 , 
     n69100 , n596424 , n596425 , n69103 , n596427 , n596428 , n69106 , n596430 , n596431 , n69109 , 
     n596433 , n596434 , n69112 , n596436 , n596437 , n69115 , n69116 , n69117 , n596441 , n69119 , 
     n596443 , n69121 , n596445 , n596446 , n69124 , n69125 , n596449 , n596450 , n69128 , n596452 , 
     n596453 , n69131 , n596455 , n69133 , n69134 , n596458 , n69136 , n596460 , n69138 , n69139 , 
     n596463 , n596464 , n69142 , n596466 , n596467 , n69145 , n596469 , n596470 , n596471 , n69149 , 
     n596473 , n69151 , n69152 , n596476 , n69154 , n69155 , n596479 , n69157 , n69158 , n596482 , 
     n596483 , n69161 , n596485 , n596486 , n69164 , n596488 , n69166 , n69167 , n596491 , n69169 , 
     n596493 , n69171 , n69172 , n69173 , n69174 , n596498 , n596499 , n69177 , n596501 , n69179 , 
     n69180 , n69181 , n596505 , n69183 , n596507 , n69185 , n69186 , n596510 , n596511 , n69189 , 
     n596513 , n596514 , n69192 , n596516 , n69194 , n69195 , n596519 , n69197 , n596521 , n69199 , 
     n596523 , n596524 , n69202 , n69203 , n596527 , n596528 , n69206 , n596530 , n596531 , n69209 , 
     n596533 , n596534 , n596535 , n69213 , n596537 , n69215 , n69216 , n596540 , n69218 , n596542 , 
     n69220 , n596544 , n596545 , n69223 , n69224 , n69225 , n596549 , n69227 , n69228 , n69229 , 
     n69230 , n69231 , n596555 , n596556 , n596557 , n69235 , n596559 , n69237 , n596561 , n69239 , 
     n69240 , n596564 , n69242 , n596566 , n596567 , n69245 , n596569 , n596570 , n596571 , n69249 , 
     n596573 , n596574 , n69252 , n596576 , n596577 , n69255 , n69256 , n596580 , n596581 , n69259 , 
     n596583 , n596584 , n69262 , n596586 , n596587 , n596588 , n69266 , n596590 , n69268 , n69269 , 
     n596593 , n596594 , n69272 , n596596 , n596597 , n69275 , n596599 , n596600 , n69278 , n596602 , 
     n69280 , n596604 , n69282 , n69283 , n596607 , n596608 , n69286 , n596610 , n596611 , n69289 , 
     n596613 , n596614 , n69292 , n596616 , n596617 , n69295 , n596619 , n69297 , n596621 , n596622 , 
     n596623 , n596624 , n69302 , n69303 , n596627 , n69305 , n69306 , n596630 , n69308 , n596632 , 
     n596633 , n69311 , n596635 , n596636 , n69314 , n596638 , n596639 , n69317 , n69318 , n596642 , 
     n69320 , n596644 , n69322 , n69323 , n69324 , n69325 , n69326 , n69327 , n69328 , n69329 , 
     n69330 , n69331 , n69332 , n596656 , n69334 , n596658 , n69336 , n69337 , n596661 , n69339 , 
     n596663 , n69341 , n596665 , n69343 , n69344 , n596668 , n69346 , n596670 , n69348 , n596672 , 
     n596673 , n69351 , n596675 , n596676 , n69354 , n596678 , n596679 , n69357 , n69358 , n596682 , 
     n596683 , n69361 , n596685 , n596686 , n69364 , n596688 , n596689 , n596690 , n69368 , n596692 , 
     n596693 , n69371 , n596695 , n596696 , n69374 , n69375 , n69376 , n69377 , n596701 , n69379 , 
     n596703 , n596704 , n69382 , n596706 , n69384 , n596708 , n69386 , n596710 , n69388 , n69389 , 
     n69390 , n69391 , n596715 , n69393 , n596717 , n69395 , n596719 , n596720 , n69398 , n596722 , 
     n596723 , n69401 , n69402 , n69403 , n69404 , n69405 , n596729 , n69407 , n596731 , n69409 , 
     n69410 , n596734 , n596735 , n69413 , n596737 , n596738 , n69416 , n596740 , n596741 , n69419 , 
     n69420 , n69421 , n596745 , n596746 , n69424 , n69425 , n69426 , n596750 , n596751 , n69429 , 
     n69430 , n69431 , n69432 , n69433 , n69434 , n69435 , n596759 , n69437 , n596761 , n69439 , 
     n596763 , n69441 , n596765 , n69443 , n596767 , n596768 , n69446 , n596770 , n596771 , n69449 , 
     n69450 , n596774 , n69452 , n596776 , n596777 , n596778 , n69456 , n596780 , n596781 , n69459 , 
     n596783 , n596784 , n69462 , n69463 , n69464 , n596788 , n69466 , n596790 , n69468 , n69469 , 
     n596793 , n69471 , n596795 , n69473 , n69474 , n596798 , n69476 , n596800 , n69478 , n596802 , 
     n69480 , n596804 , n69482 , n596806 , n69484 , n596808 , n69486 , n596810 , n69488 , n596812 , 
     n69490 , n69491 , n596815 , n596816 , n69494 , n596818 , n69496 , n69497 , n69498 , n69499 , 
     n69500 , n69501 , n596825 , n69503 , n69504 , n69505 , n69506 , n69507 , n596831 , n69509 , 
     n596833 , n596834 , n69512 , n596836 , n69514 , n69515 , n596839 , n596840 , n69518 , n69519 , 
     n596843 , n596844 , n69522 , n596846 , n596847 , n69525 , n596849 , n69527 , n596851 , n69529 , 
     n69530 , n596854 , n596855 , n69533 , n596857 , n596858 , n69536 , n596860 , n596861 , n69539 , 
     n69540 , n596864 , n69542 , n596866 , n69544 , n596868 , n596869 , n69547 , n69548 , n596872 , 
     n69550 , n596874 , n69552 , n69553 , n596877 , n596878 , n69556 , n596880 , n596881 , n69559 , 
     n596883 , n69561 , n596885 , n69563 , n596887 , n596888 , n69566 , n596890 , n596891 , n69569 , 
     n596893 , n69571 , n69572 , n596896 , n596897 , n69575 , n596899 , n69577 , n596901 , n69579 , 
     n69580 , n69581 , n69582 , n69583 , n69584 , n69585 , n69586 , n596910 , n596911 , n596912 , 
     n69590 , n596914 , n69592 , n69593 , n596917 , n596918 , n69596 , n596920 , n596921 , n69599 , 
     n596923 , n596924 , n69602 , n596926 , n69604 , n596928 , n69606 , n69607 , n596931 , n596932 , 
     n69610 , n596934 , n596935 , n69613 , n596937 , n596938 , n69616 , n69617 , n69618 , n596942 , 
     n69620 , n69621 , n69622 , n69623 , n69624 , n69625 , n69626 , n596950 , n69628 , n596952 , 
     n596953 , n69631 , n69632 , n69633 , n596957 , n69635 , n596959 , n69637 , n596961 , n69639 , 
     n69640 , n596964 , n596965 , n69643 , n596967 , n596968 , n69646 , n596970 , n69648 , n596972 , 
     n69650 , n596974 , n596975 , n69653 , n596977 , n69655 , n596979 , n596980 , n69658 , n69659 , 
     n596983 , n69661 , n596985 , n69663 , n69664 , n596988 , n596989 , n69667 , n596991 , n596992 , 
     n69670 , n596994 , n596995 , n596996 , n69674 , n69675 , n596999 , n69677 , n69678 , n597002 , 
     n69680 , n597004 , n69682 , n69683 , n597007 , n597008 , n69686 , n597010 , n597011 , n69689 , 
     n597013 , n69691 , n69692 , n597016 , n69694 , n597018 , n597019 , n597020 , n69698 , n597022 , 
     n69700 , n69701 , n69702 , n69703 , n69704 , n69705 , n69706 , n69707 , n69708 , n69709 , 
     n69710 , n69711 , n69712 , n69713 , n69714 , n597038 , n69716 , n597040 , n69718 , n69719 , 
     n597043 , n69721 , n597045 , n69723 , n69724 , n597048 , n69726 , n597050 , n69728 , n597052 , 
     n69730 , n69731 , n597055 , n597056 , n69734 , n597058 , n69736 , n597060 , n597061 , n69739 , 
     n597063 , n597064 , n69742 , n597066 , n597067 , n69745 , n597069 , n69747 , n597071 , n597072 , 
     n69750 , n597074 , n597075 , n69753 , n69754 , n597078 , n69756 , n597080 , n69758 , n69759 , 
     n69760 , n69761 , n597085 , n597086 , n69764 , n597088 , n597089 , n69767 , n597091 , n597092 , 
     n69770 , n597094 , n597095 , n597096 , n69774 , n597098 , n69776 , n597100 , n597101 , n69779 , 
     n597103 , n597104 , n69782 , n597106 , n597107 , n69785 , n69786 , n597110 , n69788 , n597112 , 
     n69790 , n597114 , n597115 , n69793 , n597117 , n597118 , n69796 , n69797 , n597121 , n69799 , 
     n597123 , n69801 , n597125 , n69803 , n69804 , n597128 , n69806 , n597130 , n69808 , n597132 , 
     n69810 , n597134 , n597135 , n69813 , n597137 , n69815 , n69816 , n597140 , n69818 , n597142 , 
     n69820 , n69821 , n597145 , n597146 , n69824 , n597148 , n597149 , n69827 , n597151 , n597152 , 
     n597153 , n69831 , n597155 , n597156 , n69834 , n597158 , n597159 , n69837 , n597161 , n597162 , 
     n69840 , n69841 , n69842 , n69843 , n69844 , n597168 , n597169 , n69847 , n597171 , n597172 , 
     n69850 , n597174 , n597175 , n69853 , n597177 , n597178 , n69856 , n69857 , n597181 , n69859 , 
     n69860 , n597184 , n597185 , n69863 , n69864 , n597188 , n69866 , n597190 , n69868 , n597192 , 
     n597193 , n69871 , n597195 , n597196 , n69874 , n597198 , n69876 , n69877 , n69878 , n69879 , 
     n597203 , n69881 , n69882 , n597206 , n597207 , n69885 , n69886 , n597210 , n597211 , n69889 , 
     n69890 , n597214 , n69892 , n597216 , n69894 , n69895 , n597219 , n597220 , n69898 , n597222 , 
     n69900 , n69901 , n69902 , n69903 , n69904 , n69905 , n597229 , n69907 , n597231 , n597232 , 
     n69910 , n597234 , n597235 , n69913 , n597237 , n597238 , n69916 , n69917 , n597241 , n69919 , 
     n69920 , n597244 , n597245 , n69923 , n69924 , n597248 , n597249 , n69927 , n597251 , n597252 , 
     n69930 , n597254 , n69932 , n597256 , n69934 , n597258 , n69936 , n597260 , n597261 , n69939 , 
     n69940 , n597264 , n597265 , n69943 , n597267 , n597268 , n69946 , n597270 , n597271 , n597272 , 
     n69950 , n597274 , n597275 , n69953 , n597277 , n597278 , n69956 , n597280 , n597281 , n69959 , 
     n597283 , n69961 , n69962 , n597286 , n69964 , n69965 , n69966 , n69967 , n69968 , n597292 , 
     n597293 , n597294 , n597295 , n69973 , n597297 , n597298 , n597299 , n69977 , n597301 , n69979 , 
     n597303 , n69981 , n597305 , n597306 , n69984 , n69985 , n597309 , n597310 , n69988 , n597312 , 
     n597313 , n69991 , n597315 , n597316 , n69994 , n69995 , n597319 , n597320 , n69998 , n597322 , 
     n597323 , n70001 , n597325 , n597326 , n70004 , n597328 , n70006 , n597330 , n70008 , n597332 , 
     n70010 , n70011 , n597335 , n597336 , n70014 , n597338 , n597339 , n70017 , n597341 , n597342 , 
     n70020 , n70021 , n597345 , n597346 , n70024 , n597348 , n597349 , n70027 , n597351 , n597352 , 
     n70030 , n597354 , n597355 , n70033 , n597357 , n70035 , n597359 , n597360 , n597361 , n70039 , 
     n597363 , n70041 , n597365 , n597366 , n597367 , n597368 , n70046 , n597370 , n597371 , n70049 , 
     n597373 , n597374 , n70052 , n597376 , n597377 , n70055 , n597379 , n597380 , n70058 , n70059 , 
     n70060 , n597384 , n597385 , n70063 , n70064 , n597388 , n70066 , n597390 , n70068 , n70069 , 
     n70070 , n597394 , n70072 , n597396 , n70074 , n597398 , n70076 , n70077 , n70078 , n597402 , 
     n597403 , n70081 , n70082 , n70083 , n597407 , n597408 , n70086 , n597410 , n597411 , n70089 , 
     n597413 , n597414 , n70092 , n597416 , n597417 , n70095 , n70096 , n597420 , n597421 , n597422 , 
     n70100 , n597424 , n70102 , n597426 , n70104 , n70105 , n597429 , n597430 , n70108 , n597432 , 
     n597433 , n70111 , n597435 , n597436 , n70114 , n70115 , n597439 , n597440 , n70118 , n597442 , 
     n597443 , n70121 , n597445 , n597446 , n70124 , n70125 , n70126 , n597450 , n70128 , n597452 , 
     n70130 , n70131 , n70132 , n597456 , n70134 , n597458 , n597459 , n597460 , n70138 , n597462 , 
     n597463 , n70141 , n597465 , n597466 , n597467 , n70145 , n597469 , n70147 , n70148 , n70149 , 
     n70150 , n70151 , n70152 , n70153 , n70154 , n70155 , n597479 , n597480 , n70158 , n597482 , 
     n70160 , n70161 , n597485 , n70163 , n597487 , n70165 , n597489 , n70167 , n597491 , n597492 , 
     n70170 , n70171 , n597495 , n597496 , n70174 , n597498 , n597499 , n70177 , n597501 , n597502 , 
     n70180 , n70181 , n597505 , n597506 , n70184 , n597508 , n597509 , n70187 , n597511 , n597512 , 
     n70190 , n597514 , n70192 , n597516 , n597517 , n70195 , n70196 , n597520 , n70198 , n70199 , 
     n597523 , n597524 , n70202 , n597526 , n597527 , n70205 , n70206 , n70207 , n597531 , n597532 , 
     n70210 , n597534 , n597535 , n70213 , n597537 , n597538 , n70216 , n70217 , n597541 , n597542 , 
     n70220 , n597544 , n597545 , n70223 , n597547 , n70225 , n597549 , n70227 , n597551 , n70229 , 
     n597553 , n70231 , n70232 , n597556 , n597557 , n70235 , n597559 , n597560 , n70238 , n597562 , 
     n597563 , n70241 , n70242 , n597566 , n597567 , n70245 , n597569 , n597570 , n70248 , n597572 , 
     n70250 , n70251 , n70252 , n70253 , n70254 , n70255 , n597579 , n70257 , n70258 , n70259 , 
     n70260 , n70261 , n70262 , n70263 , n597587 , n597588 , n70266 , n597590 , n70268 , n70269 , 
     n597593 , n70271 , n597595 , n70273 , n597597 , n597598 , n70276 , n70277 , n597601 , n597602 , 
     n70280 , n597604 , n597605 , n70283 , n597607 , n597608 , n597609 , n70287 , n597611 , n597612 , 
     n70290 , n597614 , n597615 , n70293 , n597617 , n70295 , n597619 , n70297 , n70298 , n597622 , 
     n70300 , n597624 , n70302 , n70303 , n597627 , n70305 , n597629 , n70307 , n597631 , n597632 , 
     n70310 , n597634 , n597635 , n597636 , n70314 , n597638 , n597639 , n70317 , n597641 , n597642 , 
     n70320 , n70321 , n70322 , n597646 , n597647 , n70325 , n70326 , n70327 , n597651 , n597652 , 
     n70330 , n70331 , n597655 , n597656 , n70334 , n70335 , n70336 , n597660 , n70338 , n597662 , 
     n70340 , n597664 , n70342 , n70343 , n70344 , n597668 , n70346 , n597670 , n70348 , n70349 , 
     n597673 , n70351 , n597675 , n597676 , n70354 , n597678 , n70356 , n597680 , n597681 , n70359 , 
     n597683 , n70361 , n70362 , n70363 , n70364 , n70365 , n597689 , n597690 , n70368 , n70369 , 
     n597693 , n70371 , n70372 , n597696 , n70374 , n70375 , n597699 , n597700 , n70378 , n597702 , 
     n70380 , n70381 , n70382 , n70383 , n597707 , n597708 , n70386 , n597710 , n597711 , n70389 , 
     n597713 , n597714 , n70392 , n70393 , n597717 , n597718 , n597719 , n597720 , n70398 , n597722 , 
     n597723 , n70401 , n597725 , n597726 , n597727 , n70405 , n597729 , n597730 , n70408 , n597732 , 
     n70410 , n597734 , n597735 , n597736 , n597737 , n597738 , n70416 , n597740 , n70418 , n70419 , 
     n70420 , n70421 , n70422 , n70423 , n70424 , n597748 , n70426 , n597750 , n597751 , n70429 , 
     n597753 , n597754 , n70432 , n597756 , n597757 , n597758 , n70436 , n597760 , n597761 , n70439 , 
     n597763 , n597764 , n70442 , n597766 , n70444 , n70445 , n70446 , n70447 , n70448 , n70449 , 
     n70450 , n70451 , n70452 , n70453 , n597777 , n70455 , n597779 , n597780 , n70458 , n597782 , 
     n597783 , n70461 , n597785 , n597786 , n70464 , n70465 , n70466 , n597790 , n70468 , n597792 , 
     n70470 , n597794 , n70472 , n70473 , n597797 , n70475 , n597799 , n70477 , n597801 , n597802 , 
     n70480 , n70481 , n597805 , n597806 , n70484 , n597808 , n597809 , n70487 , n597811 , n597812 , 
     n597813 , n70491 , n597815 , n597816 , n70494 , n597818 , n70496 , n70497 , n70498 , n70499 , 
     n70500 , n70501 , n597825 , n70503 , n597827 , n70505 , n597829 , n70507 , n70508 , n597832 , 
     n70510 , n597834 , n70512 , n597836 , n597837 , n70515 , n597839 , n597840 , n70518 , n70519 , 
     n597843 , n597844 , n70522 , n597846 , n597847 , n70525 , n597849 , n597850 , n70528 , n70529 , 
     n597853 , n70531 , n597855 , n70533 , n597857 , n70535 , n70536 , n597860 , n70538 , n597862 , 
     n70540 , n597864 , n597865 , n70543 , n70544 , n597868 , n70546 , n597870 , n70548 , n597872 , 
     n597873 , n70551 , n597875 , n597876 , n597877 , n70555 , n597879 , n597880 , n70558 , n597882 , 
     n597883 , n70561 , n70562 , n70563 , n597887 , n70565 , n70566 , n70567 , n597891 , n70569 , 
     n70570 , n70571 , n597895 , n597896 , n597897 , n70575 , n597899 , n597900 , n70578 , n70579 , 
     n70580 , n70581 , n70582 , n70583 , n597907 , n70585 , n70586 , n597910 , n597911 , n70589 , 
     n70590 , n597914 , n597915 , n70593 , n70594 , n70595 , n597919 , n70597 , n70598 , n70599 , 
     n70600 , n597924 , n70602 , n597926 , n70604 , n70605 , n597929 , n597930 , n70608 , n597932 , 
     n597933 , n70611 , n597935 , n70613 , n70614 , n70615 , n70616 , n70617 , n70618 , n70619 , 
     n70620 , n597944 , n70622 , n597946 , n70624 , n70625 , n597949 , n597950 , n70628 , n70629 , 
     n597953 , n70631 , n597955 , n70633 , n597957 , n70635 , n70636 , n70637 , n70638 , n70639 , 
     n70640 , n597964 , n70642 , n597966 , n70644 , n70645 , n70646 , n70647 , n70648 , n70649 , 
     n597973 , n70651 , n70652 , n70653 , n597977 , n597978 , n70656 , n597980 , n70658 , n597982 , 
     n70660 , n597984 , n70662 , n70663 , n597987 , n597988 , n70666 , n70667 , n597991 , n597992 , 
     n70670 , n70671 , n597995 , n597996 , n70674 , n70675 , n597999 , n598000 , n70678 , n70679 , 
     n70680 , n598004 , n598005 , n70683 , n598007 , n598008 , n70686 , n598010 , n70688 , n70689 , 
     n70690 , n598014 , n598015 , n70693 , n598017 , n598018 , n598019 , n70697 , n598021 , n70699 , 
     n598023 , n70701 , n70702 , n598026 , n598027 , n70705 , n70706 , n598030 , n598031 , n70709 , 
     n70710 , n598034 , n598035 , n70713 , n70714 , n598038 , n598039 , n598040 , n70718 , n598042 , 
     n70720 , n70721 , n598045 , n70723 , n598047 , n70725 , n70726 , n598050 , n70728 , n598052 , 
     n598053 , n70731 , n598055 , n70733 , n598057 , n598058 , n70736 , n598060 , n598061 , n598062 , 
     n70740 , n598064 , n598065 , n70743 , n598067 , n598068 , n70746 , n598070 , n70748 , n598072 , 
     n70750 , n70751 , n598075 , n70753 , n598077 , n70755 , n70756 , n598080 , n598081 , n70759 , 
     n598083 , n598084 , n70762 , n598086 , n598087 , n598088 , n70766 , n598090 , n598091 , n70769 , 
     n598093 , n598094 , n70772 , n70773 , n598097 , n598098 , n70776 , n598100 , n70778 , n598102 , 
     n70780 , n70781 , n70782 , n70783 , n70784 , n70785 , n70786 , n70787 , n70788 , n598112 , 
     n598113 , n70791 , n598115 , n70793 , n70794 , n70795 , n598119 , n70797 , n598121 , n598122 , 
     n598123 , n70801 , n598125 , n70803 , n70804 , n598128 , n70806 , n598130 , n70808 , n598132 , 
     n598133 , n70811 , n70812 , n598136 , n598137 , n70815 , n598139 , n598140 , n70818 , n598142 , 
     n598143 , n598144 , n70822 , n598146 , n598147 , n70825 , n598149 , n598150 , n70828 , n70829 , 
     n70830 , n70831 , n70832 , n70833 , n70834 , n70835 , n70836 , n70837 , n598161 , n70839 , 
     n70840 , n70841 , n598165 , n598166 , n70844 , n598168 , n598169 , n70847 , n598171 , n598172 , 
     n598173 , n70851 , n598175 , n70853 , n598177 , n70855 , n70856 , n598180 , n598181 , n70859 , 
     n598183 , n598184 , n70862 , n598186 , n598187 , n70865 , n70866 , n598190 , n598191 , n70869 , 
     n598193 , n598194 , n70872 , n598196 , n598197 , n70875 , n598199 , n70877 , n598201 , n70879 , 
     n598203 , n70881 , n70882 , n598206 , n70884 , n598208 , n70886 , n598210 , n598211 , n70889 , 
     n598213 , n598214 , n70892 , n70893 , n598217 , n598218 , n70896 , n598220 , n598221 , n70899 , 
     n598223 , n598224 , n70902 , n70903 , n70904 , n70905 , n70906 , n70907 , n70908 , n70909 , 
     n70910 , n70911 , n598235 , n598236 , n70914 , n598238 , n70916 , n598240 , n70918 , n70919 , 
     n598243 , n598244 , n70922 , n70923 , n70924 , n598248 , n70926 , n598250 , n598251 , n70929 , 
     n598253 , n598254 , n70932 , n70933 , n70934 , n598258 , n598259 , n70937 , n70938 , n598262 , 
     n598263 , n70941 , n70942 , n70943 , n598267 , n70945 , n598269 , n598270 , n70948 , n70949 , 
     n70950 , n598274 , n598275 , n70953 , n598277 , n598278 , n70956 , n70957 , n70958 , n70959 , 
     n598283 , n598284 , n70962 , n598286 , n598287 , n598288 , n70966 , n70967 , n598291 , n70969 , 
     n598293 , n598294 , n70972 , n598296 , n598297 , n70975 , n70976 , n70977 , n598301 , n598302 , 
     n70980 , n70981 , n598305 , n598306 , n70984 , n70985 , n70986 , n598310 , n70988 , n598312 , 
     n70990 , n598314 , n70992 , n598316 , n598317 , n70995 , n70996 , n598320 , n70998 , n70999 , 
     n598323 , n71001 , n598325 , n598326 , n71004 , n598328 , n71006 , n71007 , n598331 , n598332 , 
     n71010 , n598334 , n71012 , n71013 , n598337 , n71015 , n598339 , n598340 , n71018 , n71019 , 
     n71020 , n598344 , n71022 , n71023 , n598347 , n598348 , n71026 , n71027 , n598351 , n598352 , 
     n71030 , n598354 , n598355 , n71033 , n598357 , n71035 , n71036 , n71037 , n71038 , n598362 , 
     n71040 , n598364 , n71042 , n71043 , n598367 , n598368 , n71046 , n598370 , n598371 , n71049 , 
     n598373 , n71051 , n71052 , n71053 , n71054 , n71055 , n71056 , n598380 , n598381 , n71059 , 
     n598383 , n71061 , n598385 , n71063 , n598387 , n598388 , n71066 , n71067 , n71068 , n71069 , 
     n71070 , n71071 , n71072 , n71073 , n71074 , n598398 , n71076 , n598400 , n71078 , n71079 , 
     n71080 , n71081 , n598405 , n71083 , n71084 , n71085 , n71086 , n71087 , n71088 , n598412 , 
     n598413 , n598414 , n71092 , n598416 , n71094 , n71095 , n598419 , n71097 , n598421 , n71099 , 
     n71100 , n71101 , n598425 , n598426 , n71104 , n598428 , n598429 , n71107 , n598431 , n598432 , 
     n598433 , n71111 , n598435 , n598436 , n71114 , n598438 , n598439 , n71117 , n598441 , n71119 , 
     n598443 , n71121 , n71122 , n598446 , n71124 , n598448 , n71126 , n71127 , n598451 , n598452 , 
     n71130 , n598454 , n598455 , n71133 , n598457 , n598458 , n598459 , n71137 , n598461 , n598462 , 
     n71140 , n598464 , n598465 , n71143 , n71144 , n71145 , n598469 , n71147 , n598471 , n71149 , 
     n598473 , n71151 , n71152 , n71153 , n71154 , n71155 , n71156 , n598480 , n598481 , n71159 , 
     n598483 , n598484 , n71162 , n598486 , n71164 , n71165 , n71166 , n598490 , n71168 , n598492 , 
     n598493 , n71171 , n71172 , n598496 , n71174 , n598498 , n598499 , n71177 , n71178 , n71179 , 
     n71180 , n71181 , n71182 , n71183 , n71184 , n71185 , n71186 , n71187 , n71188 , n71189 , 
     n71190 , n71191 , n71192 , n71193 , n71194 , n598518 , n71196 , n71197 , n71198 , n598522 , 
     n598523 , n71201 , n71202 , n71203 , n598527 , n598528 , n71206 , n71207 , n71208 , n598532 , 
     n598533 , n71211 , n71212 , n71213 , n598537 , n598538 , n71216 , n598540 , n598541 , n71219 , 
     n598543 , n71221 , n71222 , n598546 , n598547 , n71225 , n598549 , n71227 , n71228 , n71229 , 
     n598553 , n598554 , n71232 , n598556 , n71234 , n71235 , n71236 , n598560 , n598561 , n71239 , 
     n598563 , n71241 , n71242 , n71243 , n598567 , n71245 , n598569 , n71247 , n71248 , n598572 , 
     n598573 , n71251 , n598575 , n71253 , n598577 , n71255 , n71256 , n598580 , n71258 , n598582 , 
     n71260 , n71261 , n598585 , n598586 , n71264 , n598588 , n598589 , n71267 , n598591 , n598592 , 
     n598593 , n71271 , n598595 , n598596 , n71274 , n598598 , n598599 , n598600 , n598601 , n71279 , 
     n598603 , n71281 , n598605 , n71283 , n71284 , n71285 , n71286 , n71287 , n71288 , n71289 , 
     n71290 , n71291 , n71292 , n71293 , n71294 , n598618 , n71296 , n598620 , n598621 , n71299 , 
     n598623 , n598624 , n71302 , n598626 , n598627 , n598628 , n71306 , n598630 , n598631 , n71309 , 
     n598633 , n71311 , n598635 , n71313 , n71314 , n598638 , n71316 , n598640 , n598641 , n598642 , 
     n598643 , n71321 , n598645 , n598646 , n71324 , n598648 , n598649 , n71327 , n71328 , n598652 , 
     n71330 , n71331 , n598655 , n598656 , n71334 , n598658 , n598659 , n71337 , n598661 , n598662 , 
     n71340 , n598664 , n598665 , n598666 , n71344 , n598668 , n598669 , n71347 , n71348 , n71349 , 
     n71350 , n71351 , n71352 , n71353 , n71354 , n598678 , n598679 , n71357 , n598681 , n598682 , 
     n71360 , n598684 , n598685 , n71363 , n598687 , n71365 , n598689 , n598690 , n71368 , n598692 , 
     n598693 , n598694 , n71372 , n598696 , n71374 , n598698 , n598699 , n71377 , n598701 , n598702 , 
     n71380 , n598704 , n598705 , n71383 , n598707 , n71385 , n598709 , n71387 , n71388 , n71389 , 
     n598713 , n598714 , n598715 , n71393 , n598717 , n598718 , n71396 , n598720 , n598721 , n71399 , 
     n71400 , n71401 , n598725 , n71403 , n71404 , n71405 , n71406 , n71407 , n71408 , n71409 , 
     n71410 , n598734 , n71412 , n598736 , n71414 , n71415 , n71416 , n71417 , n71418 , n71419 , 
     n71420 , n71421 , n71422 , n71423 , n598747 , n71425 , n71426 , n71427 , n71428 , n71429 , 
     n71430 , n598754 , n71432 , n71433 , n71434 , n71435 , n71436 , n71437 , n598761 , n71439 , 
     n598763 , n598764 , n71442 , n598766 , n598767 , n71445 , n598769 , n71447 , n71448 , n71449 , 
     n71450 , n598774 , n71452 , n598776 , n71454 , n71455 , n71456 , n71457 , n71458 , n71459 , 
     n598783 , n598784 , n71462 , n598786 , n71464 , n71465 , n71466 , n71467 , n71468 , n71469 , 
     n71470 , n71471 , n71472 , n71473 , n598797 , n598798 , n71476 , n598800 , n71478 , n71479 , 
     n71480 , n71481 , n71482 , n71483 , n598807 , n71485 , n598809 , n71487 , n598811 , n71489 , 
     n71490 , n71491 , n71492 , n71493 , n71494 , n598818 , n598819 , n71497 , n598821 , n598822 , 
     n71500 , n598824 , n598825 , n598826 , n71504 , n598828 , n71506 , n71507 , n598831 , n71509 , 
     n598833 , n71511 , n71512 , n71513 , n71514 , n598838 , n598839 , n71517 , n598841 , n598842 , 
     n71520 , n598844 , n598845 , n71523 , n598847 , n598848 , n598849 , n598850 , n71528 , n71529 , 
     n71530 , n598854 , n598855 , n71533 , n598857 , n598858 , n71536 , n598860 , n598861 , n71539 , 
     n71540 , n71541 , n598865 , n598866 , n71544 , n598868 , n598869 , n71547 , n71548 , n71549 , 
     n598873 , n598874 , n71552 , n598876 , n598877 , n71555 , n71556 , n598880 , n71558 , n598882 , 
     n71560 , n71561 , n598885 , n71563 , n71564 , n71565 , n598889 , n71567 , n598891 , n598892 , 
     n71570 , n71571 , n598895 , n71573 , n598897 , n71575 , n598899 , n598900 , n71578 , n71579 , 
     n598903 , n71581 , n598905 , n71583 , n598907 , n71585 , n71586 , n598910 , n598911 , n71589 , 
     n598913 , n598914 , n71592 , n598916 , n598917 , n71595 , n71596 , n598920 , n598921 , n71599 , 
     n598923 , n598924 , n71602 , n598926 , n598927 , n71605 , n71606 , n598930 , n598931 , n71609 , 
     n598933 , n71611 , n598935 , n71613 , n598937 , n71615 , n598939 , n598940 , n71618 , n598942 , 
     n598943 , n71621 , n71622 , n598946 , n71624 , n598948 , n71626 , n598950 , n598951 , n71629 , 
     n598953 , n598954 , n71632 , n71633 , n598957 , n598958 , n71636 , n598960 , n598961 , n71639 , 
     n598963 , n598964 , n71642 , n71643 , n71644 , n598968 , n598969 , n71647 , n598971 , n598972 , 
     n71650 , n598974 , n598975 , n71653 , n598977 , n598978 , n598979 , n71657 , n598981 , n71659 , 
     n598983 , n598984 , n71662 , n598986 , n598987 , n71665 , n71666 , n598990 , n598991 , n71669 , 
     n71670 , n598994 , n71672 , n598996 , n71674 , n71675 , n71676 , n599000 , n599001 , n71679 , 
     n599003 , n71681 , n71682 , n599006 , n599007 , n599008 , n71686 , n599010 , n71688 , n599012 , 
     n599013 , n71691 , n599015 , n599016 , n71694 , n599018 , n71696 , n599020 , n71698 , n71699 , 
     n599023 , n71701 , n599025 , n71703 , n71704 , n599028 , n599029 , n71707 , n599031 , n599032 , 
     n71710 , n599034 , n599035 , n599036 , n71714 , n599038 , n599039 , n71717 , n599041 , n599042 , 
     n599043 , n71721 , n599045 , n71723 , n599047 , n71725 , n71726 , n599050 , n71728 , n599052 , 
     n71730 , n599054 , n599055 , n71733 , n599057 , n599058 , n71736 , n71737 , n599061 , n599062 , 
     n71740 , n599064 , n599065 , n71743 , n599067 , n599068 , n71746 , n599070 , n599071 , n71749 , 
     n599073 , n71751 , n599075 , n71753 , n71754 , n599078 , n71756 , n599080 , n71758 , n71759 , 
     n599083 , n599084 , n71762 , n599086 , n599087 , n71765 , n599089 , n599090 , n599091 , n71769 , 
     n599093 , n599094 , n71772 , n599096 , n599097 , n71775 , n71776 , n71777 , n599101 , n71779 , 
     n71780 , n71781 , n71782 , n71783 , n71784 , n599108 , n71786 , n599110 , n599111 , n71789 , 
     n599113 , n71791 , n71792 , n71793 , n71794 , n599118 , n71796 , n599120 , n71798 , n599122 , 
     n71800 , n599124 , n599125 , n599126 , n599127 , n71805 , n599129 , n599130 , n71808 , n599132 , 
     n599133 , n71811 , n71812 , n71813 , n599137 , n599138 , n71816 , n599140 , n71818 , n71819 , 
     n71820 , n599144 , n71822 , n71823 , n71824 , n71825 , n71826 , n71827 , n71828 , n599152 , 
     n599153 , n71831 , n71832 , n71833 , n71834 , n599158 , n599159 , n71837 , n71838 , n71839 , 
     n71840 , n71841 , n599165 , n599166 , n599167 , n71845 , n599169 , n71847 , n71848 , n599172 , 
     n71850 , n599174 , n71852 , n71853 , n599177 , n71855 , n599179 , n599180 , n599181 , n71859 , 
     n599183 , n599184 , n71862 , n599186 , n599187 , n599188 , n71866 , n599190 , n599191 , n71869 , 
     n599193 , n599194 , n71872 , n599196 , n71874 , n599198 , n71876 , n71877 , n599201 , n599202 , 
     n71880 , n599204 , n599205 , n71883 , n599207 , n599208 , n71886 , n71887 , n599211 , n599212 , 
     n71890 , n599214 , n599215 , n71893 , n599217 , n71895 , n599219 , n71897 , n599221 , n71899 , 
     n71900 , n599224 , n71902 , n599226 , n71904 , n599228 , n599229 , n71907 , n71908 , n599232 , 
     n599233 , n71911 , n599235 , n599236 , n71914 , n599238 , n599239 , n599240 , n71918 , n599242 , 
     n599243 , n71921 , n599245 , n71923 , n599247 , n71925 , n599249 , n599250 , n71928 , n71929 , 
     n71930 , n71931 , n599255 , n599256 , n71934 , n599258 , n71936 , n71937 , n599261 , n599262 , 
     n71940 , n599264 , n599265 , n71943 , n599267 , n599268 , n71946 , n599270 , n71948 , n599272 , 
     n599273 , n599274 , n71952 , n599276 , n71954 , n599278 , n599279 , n71957 , n599281 , n599282 , 
     n71960 , n599284 , n71962 , n599286 , n71964 , n599288 , n71966 , n71967 , n599291 , n599292 , 
     n71970 , n599294 , n599295 , n71973 , n599297 , n599298 , n71976 , n71977 , n599301 , n599302 , 
     n71980 , n599304 , n599305 , n71983 , n599307 , n599308 , n71986 , n599310 , n599311 , n71989 , 
     n599313 , n71991 , n599315 , n71993 , n599317 , n71995 , n71996 , n599320 , n599321 , n71999 , 
     n599323 , n599324 , n72002 , n599326 , n599327 , n72005 , n72006 , n599330 , n599331 , n72009 , 
     n599333 , n599334 , n72012 , n599336 , n599337 , n72015 , n599339 , n599340 , n72018 , n72019 , 
     n599343 , n72021 , n599345 , n599346 , n599347 , n72025 , n599349 , n599350 , n72028 , n599352 , 
     n599353 , n72031 , n72032 , n72033 , n72034 , n599358 , n599359 , n72037 , n599361 , n599362 , 
     n72040 , n599364 , n72042 , n599366 , n72044 , n72045 , n599369 , n72047 , n599371 , n72049 , 
     n72050 , n599374 , n599375 , n72053 , n599377 , n599378 , n72056 , n599380 , n599381 , n599382 , 
     n72060 , n599384 , n599385 , n72063 , n599387 , n599388 , n72066 , n72067 , n72068 , n72069 , 
     n599393 , n599394 , n72072 , n599396 , n72074 , n599398 , n599399 , n599400 , n72078 , n599402 , 
     n72080 , n72081 , n599405 , n72083 , n599407 , n72085 , n72086 , n599410 , n72088 , n599412 , 
     n599413 , n599414 , n72092 , n599416 , n599417 , n72095 , n599419 , n599420 , n599421 , n72099 , 
     n599423 , n599424 , n72102 , n599426 , n599427 , n72105 , n599429 , n72107 , n599431 , n72109 , 
     n72110 , n599434 , n72112 , n72113 , n599437 , n72115 , n72116 , n72117 , n599441 , n72119 , 
     n72120 , n599444 , n599445 , n599446 , n72124 , n599448 , n599449 , n72127 , n599451 , n599452 , 
     n72130 , n599454 , n599455 , n72133 , n599457 , n599458 , n599459 , n72137 , n599461 , n72139 , 
     n72140 , n599464 , n599465 , n72143 , n599467 , n72145 , n599469 , n599470 , n72148 , n599472 , 
     n599473 , n72151 , n72152 , n72153 , n72154 , n599478 , n599479 , n72157 , n599481 , n72159 , 
     n72160 , n599484 , n72162 , n599486 , n599487 , n72165 , n72166 , n72167 , n72168 , n72169 , 
     n72170 , n72171 , n599495 , n72173 , n72174 , n72175 , n72176 , n599500 , n599501 , n72179 , 
     n599503 , n72181 , n599505 , n599506 , n72184 , n599508 , n72186 , n599510 , n72188 , n599512 , 
     n599513 , n72191 , n599515 , n599516 , n72194 , n599518 , n599519 , n72197 , n599521 , n599522 , 
     n72200 , n599524 , n72202 , n72203 , n72204 , n72205 , n599529 , n72207 , n72208 , n72209 , 
     n72210 , n72211 , n72212 , n72213 , n72214 , n72215 , n72216 , n599540 , n599541 , n72219 , 
     n599543 , n599544 , n72222 , n72223 , n72224 , n72225 , n72226 , n599550 , n599551 , n72229 , 
     n72230 , n72231 , n72232 , n72233 , n599557 , n72235 , n599559 , n599560 , n599561 , n72239 , 
     n599563 , n72241 , n72242 , n599566 , n72244 , n599568 , n599569 , n72247 , n599571 , n599572 , 
     n72250 , n72251 , n599575 , n599576 , n72254 , n599578 , n599579 , n72257 , n599581 , n599582 , 
     n599583 , n72261 , n599585 , n72263 , n599587 , n72265 , n599589 , n599590 , n72268 , n72269 , 
     n599593 , n599594 , n72272 , n599596 , n599597 , n72275 , n599599 , n599600 , n72278 , n72279 , 
     n599603 , n599604 , n72282 , n599606 , n599607 , n72285 , n599609 , n599610 , n72288 , n599612 , 
     n599613 , n72291 , n599615 , n72293 , n599617 , n599618 , n599619 , n72297 , n599621 , n599622 , 
     n72300 , n599624 , n599625 , n72303 , n599627 , n599628 , n72306 , n599630 , n72308 , n599632 , 
     n599633 , n72311 , n599635 , n599636 , n599637 , n72315 , n599639 , n72317 , n72318 , n599642 , 
     n72320 , n599644 , n72322 , n72323 , n72324 , n72325 , n599649 , n72327 , n599651 , n599652 , 
     n599653 , n72331 , n599655 , n599656 , n72334 , n599658 , n599659 , n72337 , n599661 , n72339 , 
     n599663 , n72341 , n72342 , n599666 , n599667 , n72345 , n72346 , n599670 , n72348 , n72349 , 
     n599673 , n599674 , n599675 , n72353 , n599677 , n599678 , n72356 , n599680 , n599681 , n72359 , 
     n599683 , n599684 , n72362 , n599686 , n72364 , n599688 , n72366 , n599690 , n599691 , n72369 , 
     n599693 , n599694 , n599695 , n72373 , n599697 , n72375 , n72376 , n72377 , n72378 , n72379 , 
     n72380 , n72381 , n599705 , n599706 , n599707 , n72385 , n72386 , n72387 , n72388 , n72389 , 
     n599713 , n72391 , n72392 , n599716 , n599717 , n72395 , n599719 , n599720 , n72398 , n599722 , 
     n599723 , n72401 , n72402 , n72403 , n72404 , n72405 , n599729 , n599730 , n72408 , n72409 , 
     n72410 , n599734 , n599735 , n599736 , n72414 , n599738 , n72416 , n72417 , n599741 , n72419 , 
     n599743 , n72421 , n72422 , n599746 , n72424 , n599748 , n599749 , n72427 , n599751 , n599752 , 
     n72430 , n599754 , n72432 , n599756 , n599757 , n72435 , n599759 , n72437 , n599761 , n599762 , 
     n72440 , n72441 , n599765 , n72443 , n599767 , n599768 , n599769 , n72447 , n599771 , n72449 , 
     n599773 , n599774 , n72452 , n599776 , n599777 , n599778 , n72456 , n599780 , n72458 , n599782 , 
     n599783 , n72461 , n72462 , n599786 , n72464 , n599788 , n599789 , n599790 , n72468 , n599792 , 
     n72470 , n599794 , n599795 , n72473 , n599797 , n599798 , n72476 , n599800 , n72478 , n599802 , 
     n72480 , n72481 , n599805 , n72483 , n599807 , n72485 , n72486 , n599810 , n72488 , n599812 , 
     n72490 , n599814 , n599815 , n72493 , n599817 , n599818 , n599819 , n72497 , n599821 , n599822 , 
     n72500 , n599824 , n72502 , n72503 , n72504 , n72505 , n72506 , n599830 , n72508 , n599832 , 
     n72510 , n72511 , n599835 , n599836 , n72514 , n72515 , n599839 , n72517 , n72518 , n72519 , 
     n599843 , n72521 , n599845 , n599846 , n72524 , n599848 , n72526 , n72527 , n599851 , n72529 , 
     n599853 , n72531 , n72532 , n599856 , n599857 , n72535 , n599859 , n72537 , n599861 , n599862 , 
     n72540 , n599864 , n599865 , n599866 , n72544 , n599868 , n72546 , n72547 , n599871 , n72549 , 
     n599873 , n72551 , n72552 , n599876 , n72554 , n599878 , n599879 , n599880 , n72558 , n599882 , 
     n599883 , n72561 , n599885 , n599886 , n599887 , n72565 , n599889 , n599890 , n72568 , n599892 , 
     n599893 , n599894 , n72572 , n599896 , n72574 , n599898 , n72576 , n72577 , n599901 , n72579 , 
     n599903 , n599904 , n599905 , n72583 , n599907 , n599908 , n72586 , n599910 , n599911 , n72589 , 
     n72590 , n599914 , n599915 , n72593 , n599917 , n599918 , n72596 , n599920 , n599921 , n72599 , 
     n599923 , n72601 , n599925 , n72603 , n72604 , n599928 , n72606 , n599930 , n72608 , n599932 , 
     n599933 , n72611 , n72612 , n599936 , n599937 , n72615 , n599939 , n599940 , n72618 , n599942 , 
     n599943 , n599944 , n72622 , n599946 , n599947 , n72625 , n599949 , n599950 , n72628 , n599952 , 
     n599953 , n72631 , n72632 , n72633 , n599957 , n599958 , n72636 , n72637 , n72638 , n599962 , 
     n599963 , n72641 , n72642 , n72643 , n72644 , n599968 , n599969 , n599970 , n72648 , n599972 , 
     n72650 , n72651 , n599975 , n599976 , n72654 , n72655 , n599979 , n72657 , n72658 , n599982 , 
     n599983 , n599984 , n72662 , n599986 , n599987 , n72665 , n599989 , n599990 , n599991 , n72669 , 
     n599993 , n72671 , n72672 , n599996 , n72674 , n599998 , n72676 , n72677 , n600001 , n600002 , 
     n72680 , n600004 , n600005 , n72683 , n600007 , n600008 , n600009 , n72687 , n600011 , n600012 , 
     n72690 , n600014 , n600015 , n72693 , n600017 , n72695 , n600019 , n72697 , n600021 , n72699 , 
     n72700 , n600024 , n600025 , n72703 , n600027 , n600028 , n72706 , n600030 , n600031 , n72709 , 
     n72710 , n600034 , n600035 , n72713 , n600037 , n600038 , n72716 , n600040 , n600041 , n72719 , 
     n600043 , n600044 , n72722 , n72723 , n72724 , n72725 , n600049 , n600050 , n72728 , n600052 , 
     n72730 , n72731 , n600055 , n600056 , n72734 , n600058 , n72736 , n600060 , n600061 , n72739 , 
     n600063 , n600064 , n72742 , n600066 , n72744 , n600068 , n600069 , n72747 , n72748 , n600072 , 
     n600073 , n72751 , n72752 , n600076 , n600077 , n72755 , n600079 , n600080 , n600081 , n72759 , 
     n600083 , n72761 , n72762 , n600086 , n72764 , n600088 , n72766 , n72767 , n600091 , n600092 , 
     n72770 , n600094 , n600095 , n72773 , n600097 , n600098 , n600099 , n72777 , n600101 , n600102 , 
     n72780 , n600104 , n600105 , n72783 , n600107 , n72785 , n600109 , n72787 , n72788 , n600112 , 
     n72790 , n600114 , n72792 , n72793 , n600117 , n72795 , n600119 , n600120 , n600121 , n72799 , 
     n600123 , n600124 , n72802 , n600126 , n600127 , n600128 , n72806 , n600130 , n600131 , n72809 , 
     n600133 , n600134 , n72812 , n600136 , n600137 , n72815 , n600139 , n600140 , n72818 , n600142 , 
     n72820 , n72821 , n72822 , n600146 , n600147 , n72825 , n600149 , n72827 , n72828 , n72829 , 
     n72830 , n72831 , n72832 , n600156 , n72834 , n72835 , n72836 , n72837 , n600161 , n72839 , 
     n600163 , n72841 , n72842 , n600166 , n72844 , n600168 , n72846 , n72847 , n72848 , n72849 , 
     n72850 , n72851 , n72852 , n72853 , n72854 , n600178 , n600179 , n72857 , n600181 , n72859 , 
     n72860 , n72861 , n72862 , n72863 , n72864 , n72865 , n72866 , n72867 , n72868 , n72869 , 
     n72870 , n600194 , n600195 , n72873 , n600197 , n72875 , n72876 , n72877 , n72878 , n600202 , 
     n72880 , n600204 , n600205 , n72883 , n600207 , n72885 , n600209 , n600210 , n72888 , n600212 , 
     n72890 , n72891 , n600215 , n72893 , n600217 , n72895 , n600219 , n600220 , n72898 , n600222 , 
     n72900 , n72901 , n72902 , n72903 , n72904 , n72905 , n72906 , n600230 , n72908 , n600232 , 
     n72910 , n72911 , n600235 , n600236 , n72914 , n600238 , n600239 , n72917 , n600241 , n600242 , 
     n600243 , n72921 , n600245 , n72923 , n600247 , n72925 , n72926 , n72927 , n600251 , n72929 , 
     n600253 , n72931 , n72932 , n600256 , n72934 , n72935 , n600259 , n600260 , n72938 , n600262 , 
     n600263 , n72941 , n600265 , n600266 , n72944 , n600268 , n72946 , n600270 , n72948 , n72949 , 
     n600273 , n72951 , n600275 , n72953 , n72954 , n600278 , n600279 , n72957 , n600281 , n600282 , 
     n72960 , n600284 , n600285 , n600286 , n72964 , n600288 , n600289 , n72967 , n600291 , n600292 , 
     n72970 , n600294 , n72972 , n600296 , n72974 , n600298 , n600299 , n72977 , n72978 , n600302 , 
     n72980 , n72981 , n600305 , n72983 , n72984 , n72985 , n72986 , n600310 , n600311 , n72989 , 
     n72990 , n600314 , n600315 , n72993 , n600317 , n600318 , n600319 , n72997 , n600321 , n72999 , 
     n600323 , n73001 , n73002 , n600326 , n600327 , n73005 , n600329 , n600330 , n73008 , n600332 , 
     n600333 , n73011 , n73012 , n600336 , n600337 , n73015 , n600339 , n600340 , n73018 , n600342 , 
     n600343 , n73021 , n73022 , n73023 , n73024 , n600348 , n73026 , n600350 , n73028 , n73029 , 
     n600353 , n600354 , n73032 , n600356 , n600357 , n73035 , n600359 , n73037 , n73038 , n600362 , 
     n73040 , n600364 , n600365 , n73043 , n73044 , n73045 , n73046 , n600370 , n600371 , n73049 , 
     n600373 , n73051 , n600375 , n73053 , n73054 , n600378 , n73056 , n600380 , n73058 , n73059 , 
     n600383 , n73061 , n600385 , n73063 , n600387 , n600388 , n73066 , n600390 , n600391 , n600392 , 
     n73070 , n600394 , n600395 , n73073 , n600397 , n600398 , n73076 , n600400 , n73078 , n600402 , 
     n73080 , n600404 , n73082 , n73083 , n600407 , n73085 , n600409 , n73087 , n73088 , n600412 , 
     n73090 , n600414 , n600415 , n73093 , n600417 , n600418 , n600419 , n73097 , n600421 , n600422 , 
     n73100 , n600424 , n600425 , n600426 , n73104 , n600428 , n600429 , n73107 , n600431 , n73109 , 
     n73110 , n600434 , n73112 , n600436 , n73114 , n73115 , n73116 , n600440 , n73118 , n600442 , 
     n73120 , n73121 , n600445 , n73123 , n600447 , n73125 , n600449 , n600450 , n73128 , n600452 , 
     n73130 , n73131 , n600455 , n73133 , n600457 , n73135 , n600459 , n73137 , n73138 , n73139 , 
     n73140 , n73141 , n73142 , n600466 , n73144 , n600468 , n600469 , n73147 , n600471 , n600472 , 
     n73150 , n73151 , n600475 , n600476 , n73154 , n600478 , n600479 , n73157 , n600481 , n600482 , 
     n73160 , n600484 , n600485 , n600486 , n73164 , n600488 , n73166 , n600490 , n600491 , n73169 , 
     n73170 , n600494 , n600495 , n73173 , n600497 , n73175 , n600499 , n600500 , n73178 , n600502 , 
     n600503 , n73181 , n600505 , n73183 , n600507 , n600508 , n600509 , n73187 , n600511 , n600512 , 
     n73190 , n73191 , n600515 , n600516 , n73194 , n600518 , n73196 , n73197 , n600521 , n73199 , 
     n600523 , n73201 , n73202 , n600526 , n600527 , n73205 , n600529 , n73207 , n600531 , n600532 , 
     n73210 , n600534 , n600535 , n600536 , n73214 , n600538 , n73216 , n73217 , n600541 , n73219 , 
     n600543 , n73221 , n73222 , n600546 , n600547 , n73225 , n600549 , n600550 , n73228 , n600552 , 
     n600553 , n600554 , n73232 , n600556 , n600557 , n73235 , n600559 , n600560 , n73238 , n600562 , 
     n73240 , n600564 , n73242 , n73243 , n600567 , n73245 , n600569 , n73247 , n73248 , n600572 , 
     n600573 , n73251 , n600575 , n600576 , n73254 , n600578 , n600579 , n600580 , n73258 , n600582 , 
     n600583 , n73261 , n600585 , n600586 , n73264 , n600588 , n73266 , n600590 , n73268 , n600592 , 
     n73270 , n73271 , n600595 , n73273 , n600597 , n73275 , n73276 , n600600 , n600601 , n73279 , 
     n600603 , n600604 , n73282 , n600606 , n600607 , n600608 , n73286 , n600610 , n600611 , n73289 , 
     n600613 , n73291 , n73292 , n73293 , n73294 , n600618 , n73296 , n600620 , n600621 , n73299 , 
     n600623 , n73301 , n600625 , n600626 , n73304 , n600628 , n600629 , n73307 , n600631 , n73309 , 
     n600633 , n600634 , n73312 , n600636 , n600637 , n73315 , n73316 , n600640 , n600641 , n73319 , 
     n600643 , n600644 , n73322 , n600646 , n600647 , n73325 , n600649 , n73327 , n73328 , n73329 , 
     n73330 , n73331 , n73332 , n600656 , n600657 , n600658 , n600659 , n73337 , n600661 , n73339 , 
     n73340 , n73341 , n73342 , n73343 , n73344 , n73345 , n600669 , n73347 , n73348 , n600672 , 
     n73350 , n600674 , n73352 , n73353 , n600677 , n600678 , n73356 , n600680 , n73358 , n600682 , 
     n73360 , n73361 , n600685 , n600686 , n73364 , n600688 , n600689 , n73367 , n600691 , n600692 , 
     n73370 , n73371 , n600695 , n600696 , n73374 , n600698 , n600699 , n73377 , n600701 , n600702 , 
     n73380 , n73381 , n73382 , n73383 , n73384 , n600708 , n73386 , n73387 , n600711 , n600712 , 
     n73390 , n600714 , n600715 , n73393 , n600717 , n73395 , n600719 , n73397 , n600721 , n73399 , 
     n73400 , n73401 , n73402 , n73403 , n600727 , n600728 , n73406 , n600730 , n73408 , n600732 , 
     n600733 , n73411 , n600735 , n600736 , n73414 , n600738 , n600739 , n73417 , n600741 , n73419 , 
     n600743 , n73421 , n600745 , n600746 , n73424 , n73425 , n600749 , n73427 , n73428 , n600752 , 
     n600753 , n73431 , n73432 , n73433 , n73434 , n73435 , n73436 , n73437 , n73438 , n73439 , 
     n600763 , n73441 , n600765 , n73443 , n73444 , n600768 , n600769 , n73447 , n600771 , n73449 , 
     n73450 , n600774 , n600775 , n73453 , n600777 , n73455 , n73456 , n73457 , n73458 , n73459 , 
     n73460 , n73461 , n600785 , n600786 , n73464 , n600788 , n73466 , n73467 , n600791 , n73469 , 
     n600793 , n600794 , n73472 , n600796 , n73474 , n600798 , n73476 , n600800 , n600801 , n73479 , 
     n600803 , n73481 , n600805 , n73483 , n73484 , n73485 , n73486 , n73487 , n73488 , n73489 , 
     n73490 , n73491 , n73492 , n73493 , n73494 , n73495 , n73496 , n73497 , n73498 , n73499 , 
     n73500 , n73501 , n73502 , n73503 , n73504 , n73505 , n600829 , n73507 , n73508 , n73509 , 
     n73510 , n73511 , n73512 , n73513 , n73514 , n73515 , n73516 , n73517 , n73518 , n73519 , 
     n73520 , n73521 , n73522 , n73523 , n73524 , n73525 , n600849 , n73527 , n600851 , n600852 , 
     n600853 , n73531 , n600855 , n600856 , n73534 , n600858 , n600859 , n600860 , n73538 , n600862 , 
     n600863 , n73541 , n600865 , n600866 , n73544 , n600868 , n73546 , n73547 , n73548 , n73549 , 
     n73550 , n73551 , n600875 , n73553 , n600877 , n73555 , n600879 , n600880 , n73558 , n600882 , 
     n600883 , n73561 , n600885 , n600886 , n73564 , n600888 , n600889 , n73567 , n600891 , n73569 , 
     n73570 , n73571 , n73572 , n73573 , n73574 , n73575 , n73576 , n73577 , n73578 , n73579 , 
     n73580 , n73581 , n600905 , n73583 , n600907 , n600908 , n73586 , n73587 , n73588 , n73589 , 
     n600913 , n73591 , n600915 , n73593 , n600917 , n600918 , n73596 , n73597 , n600921 , n73599 , 
     n73600 , n600924 , n73602 , n600926 , n600927 , n73605 , n600929 , n600930 , n73608 , n73609 , 
     n600933 , n600934 , n73612 , n600936 , n600937 , n73615 , n600939 , n73617 , n73618 , n73619 , 
     n73620 , n73621 , n73622 , n73623 , n73624 , n73625 , n73626 , n600950 , n73628 , n600952 , 
     n73630 , n600954 , n600955 , n73633 , n600957 , n600958 , n73636 , n73637 , n600961 , n73639 , 
     n600963 , n73641 , n600965 , n600966 , n73644 , n600968 , n73646 , n73647 , n73648 , n600972 , 
     n73650 , n600974 , n73652 , n600976 , n73654 , n73655 , n600979 , n600980 , n73658 , n600982 , 
     n600983 , n73661 , n600985 , n600986 , n600987 , n73665 , n73666 , n600990 , n73668 , n600992 , 
     n73670 , n73671 , n600995 , n600996 , n73674 , n600998 , n600999 , n73677 , n601001 , n73679 , 
     n601003 , n73681 , n601005 , n601006 , n73684 , n601008 , n601009 , n73687 , n73688 , n601012 , 
     n73690 , n601014 , n73692 , n73693 , n601017 , n73695 , n601019 , n73697 , n601021 , n73699 , 
     n73700 , n601024 , n73702 , n601026 , n73704 , n601028 , n601029 , n73707 , n601031 , n601032 , 
     n73710 , n73711 , n73712 , n73713 , n73714 , n73715 , n73716 , n601040 , n601041 , n73719 , 
     n601043 , n601044 , n73722 , n601046 , n601047 , n73725 , n601049 , n601050 , n73728 , n601052 , 
     n73730 , n601054 , n73732 , n601056 , n73734 , n601058 , n73736 , n73737 , n601061 , n601062 , 
     n73740 , n601064 , n601065 , n73743 , n601067 , n73745 , n73746 , n601070 , n73748 , n601072 , 
     n73750 , n73751 , n601075 , n601076 , n73754 , n601078 , n601079 , n73757 , n601081 , n73759 , 
     n73760 , n601084 , n73762 , n73763 , n73764 , n601088 , n73766 , n73767 , n601091 , n601092 , 
     n601093 , n73771 , n601095 , n601096 , n73774 , n73775 , n73776 , n73777 , n601101 , n73779 , 
     n601103 , n73781 , n601105 , n601106 , n73784 , n73785 , n601109 , n601110 , n73788 , n601112 , 
     n601113 , n73791 , n601115 , n601116 , n73794 , n73795 , n601119 , n73797 , n601121 , n73799 , 
     n73800 , n601124 , n73802 , n601126 , n73804 , n601128 , n601129 , n73807 , n601131 , n601132 , 
     n601133 , n73811 , n601135 , n601136 , n73814 , n601138 , n601139 , n73817 , n601141 , n601142 , 
     n73820 , n601144 , n73822 , n601146 , n601147 , n73825 , n601149 , n73827 , n601151 , n73829 , 
     n73830 , n601154 , n73832 , n601156 , n73834 , n601158 , n601159 , n73837 , n601161 , n601162 , 
     n73840 , n73841 , n73842 , n73843 , n73844 , n601168 , n73846 , n601170 , n73848 , n601172 , 
     n73850 , n601174 , n601175 , n73853 , n601177 , n601178 , n73856 , n601180 , n601181 , n73859 , 
     n601183 , n601184 , n73862 , n73863 , n601187 , n601188 , n73866 , n601190 , n73868 , n601192 , 
     n73870 , n601194 , n73872 , n73873 , n601197 , n601198 , n73876 , n601200 , n601201 , n73879 , 
     n601203 , n601204 , n73882 , n73883 , n601207 , n73885 , n601209 , n73887 , n73888 , n601212 , 
     n601213 , n73891 , n601215 , n601216 , n73894 , n601218 , n601219 , n601220 , n73898 , n601222 , 
     n601223 , n73901 , n601225 , n601226 , n73904 , n601228 , n601229 , n73907 , n601231 , n601232 , 
     n73910 , n601234 , n73912 , n601236 , n73914 , n601238 , n73916 , n73917 , n601241 , n601242 , 
     n73920 , n601244 , n601245 , n73923 , n601247 , n601248 , n73926 , n73927 , n601251 , n73929 , 
     n601253 , n73931 , n73932 , n601256 , n601257 , n73935 , n601259 , n601260 , n73938 , n601262 , 
     n601263 , n601264 , n73942 , n601266 , n601267 , n73945 , n601269 , n601270 , n73948 , n601272 , 
     n73950 , n73951 , n601275 , n601276 , n73954 , n601278 , n601279 , n73957 , n601281 , n601282 , 
     n73960 , n601284 , n601285 , n73963 , n601287 , n73965 , n73966 , n601290 , n73968 , n601292 , 
     n73970 , n73971 , n73972 , n601296 , n601297 , n73975 , n601299 , n601300 , n73978 , n601302 , 
     n601303 , n601304 , n73982 , n73983 , n601307 , n73985 , n601309 , n73987 , n601311 , n73989 , 
     n73990 , n601314 , n73992 , n601316 , n601317 , n601318 , n73996 , n601320 , n73998 , n601322 , 
     n601323 , n74001 , n601325 , n601326 , n74004 , n74005 , n601329 , n74007 , n74008 , n601332 , 
     n601333 , n74011 , n601335 , n601336 , n601337 , n74015 , n601339 , n601340 , n74018 , n74019 , 
     n74020 , n74021 , n74022 , n74023 , n74024 , n74025 , n74026 , n74027 , n74028 , n74029 , 
     n74030 , n74031 , n74032 , n74033 , n74034 , n74035 , n74036 , n74037 , n74038 , n74039 , 
     n74040 , n74041 , n74042 , n74043 , n74044 , n74045 , n74046 , n74047 , n74048 , n74049 , 
     n74050 , n74051 , n74052 , n74053 , n74054 , n74055 , n74056 , n601380 , n74058 , n601382 , 
     n74060 , n74061 , n74062 , n74063 , n74064 , n74065 , n74066 , n74067 , n74068 , n74069 , 
     n74070 , n74071 , n74072 , n74073 , n74074 , n74075 , n74076 , n74077 , n74078 , n74079 , 
     n601403 , n74081 , n601405 , n601406 , n74084 , n601408 , n601409 , n601410 , n74088 , n601412 , 
     n74090 , n74091 , n74092 , n601416 , n74094 , n601418 , n74096 , n601420 , n74098 , n601422 , 
     n74100 , n601424 , n601425 , n74103 , n74104 , n74105 , n601429 , n74107 , n601431 , n601432 , 
     n74110 , n74111 , n601435 , n74113 , n601437 , n601438 , n74116 , n74117 , n601441 , n74119 , 
     n74120 , n601444 , n601445 , n74123 , n601447 , n601448 , n74126 , n601450 , n601451 , n74129 , 
     n74130 , n601454 , n74132 , n601456 , n601457 , n74135 , n601459 , n601460 , n601461 , n74139 , 
     n601463 , n601464 , n74142 , n601466 , n601467 , n601468 , n74146 , n601470 , n601471 , n74149 , 
     n601473 , n601474 , n74152 , n601476 , n601477 , n601478 , n74156 , n601480 , n74158 , n601482 , 
     n74160 , n74161 , n601485 , n601486 , n74164 , n601488 , n601489 , n74167 , n601491 , n601492 , 
     n74170 , n74171 , n601495 , n74173 , n601497 , n74175 , n74176 , n601500 , n601501 , n74179 , 
     n601503 , n601504 , n74182 , n601506 , n601507 , n601508 , n74186 , n601510 , n601511 , n74189 , 
     n601513 , n601514 , n74192 , n601516 , n74194 , n74195 , n74196 , n74197 , n74198 , n601522 , 
     n74200 , n74201 , n601525 , n601526 , n74204 , n601528 , n601529 , n74207 , n601531 , n601532 , 
     n74210 , n601534 , n74212 , n601536 , n74214 , n601538 , n601539 , n601540 , n74218 , n601542 , 
     n74220 , n601544 , n74222 , n74223 , n601547 , n74225 , n601549 , n74227 , n601551 , n601552 , 
     n74230 , n601554 , n601555 , n74233 , n74234 , n601558 , n601559 , n74237 , n601561 , n601562 , 
     n74240 , n601564 , n601565 , n74243 , n601567 , n74245 , n601569 , n74247 , n601571 , n601572 , 
     n74250 , n74251 , n601575 , n74253 , n74254 , n601578 , n601579 , n74257 , n74258 , n601582 , 
     n74260 , n601584 , n74262 , n601586 , n74264 , n601588 , n74266 , n601590 , n74268 , n601592 , 
     n601593 , n601594 , n74272 , n601596 , n74274 , n601598 , n74276 , n74277 , n601601 , n74279 , 
     n601603 , n74281 , n601605 , n601606 , n74284 , n74285 , n601609 , n601610 , n74288 , n601612 , 
     n601613 , n74291 , n601615 , n601616 , n601617 , n74295 , n601619 , n601620 , n74298 , n601622 , 
     n601623 , n74301 , n601625 , n74303 , n601627 , n74305 , n601629 , n74307 , n601631 , n74309 , 
     n74310 , n601634 , n74312 , n601636 , n601637 , n601638 , n74316 , n601640 , n74318 , n601642 , 
     n74320 , n601644 , n74322 , n74323 , n601647 , n74325 , n601649 , n601650 , n74328 , n601652 , 
     n74330 , n74331 , n601655 , n74333 , n601657 , n74335 , n74336 , n601660 , n601661 , n74339 , 
     n601663 , n74341 , n74342 , n601666 , n601667 , n74345 , n601669 , n601670 , n74348 , n601672 , 
     n601673 , n74351 , n601675 , n601676 , n74354 , n601678 , n601679 , n74357 , n601681 , n74359 , 
     n601683 , n601684 , n74362 , n601686 , n601687 , n74365 , n74366 , n601690 , n601691 , n74369 , 
     n74370 , n601694 , n74372 , n74373 , n74374 , n74375 , n74376 , n74377 , n74378 , n74379 , 
     n601703 , n74381 , n601705 , n601706 , n601707 , n74385 , n601709 , n74387 , n74388 , n74389 , 
     n74390 , n601714 , n74392 , n601716 , n601717 , n74395 , n601719 , n74397 , n601721 , n601722 , 
     n74400 , n74401 , n601725 , n601726 , n74404 , n74405 , n601729 , n74407 , n601731 , n601732 , 
     n74410 , n74411 , n601735 , n601736 , n601737 , n74415 , n74416 , n601740 , n601741 , n74419 , 
     n601743 , n601744 , n74422 , n74423 , n601747 , n74425 , n601749 , n74427 , n74428 , n601752 , 
     n601753 , n74431 , n74432 , n601756 , n601757 , n74435 , n74436 , n601760 , n601761 , n601762 , 
     n601763 , n74441 , n601765 , n74443 , n74444 , n601768 , n74446 , n74447 , n601771 , n601772 , 
     n74450 , n601774 , n601775 , n74453 , n601777 , n601778 , n74456 , n601780 , n74458 , n601782 , 
     n601783 , n74461 , n601785 , n74463 , n74464 , n74465 , n74466 , n74467 , n74468 , n74469 , 
     n74470 , n74471 , n74472 , n74473 , n74474 , n74475 , n74476 , n74477 , n74478 , n74479 , 
     n74480 , n74481 , n74482 , n601806 , n601807 , n74485 , n601809 , n74487 , n74488 , n74489 , 
     n74490 , n74491 , n74492 , n74493 , n74494 , n74495 , n74496 , n74497 , n74498 , n74499 , 
     n74500 , n74501 , n74502 , n74503 , n74504 , n74505 , n74506 , n74507 , n74508 , n74509 , 
     n74510 , n74511 , n74512 , n74513 , n74514 , n74515 , n74516 , n74517 , n74518 , n74519 , 
     n74520 , n74521 , n74522 , n74523 , n74524 , n74525 , n601849 , n74527 , n601851 , n74529 , 
     n74530 , n601854 , n74532 , n74533 , n601857 , n74535 , n74536 , n601860 , n601861 , n74539 , 
     n601863 , n601864 , n74542 , n601866 , n601867 , n601868 , n74546 , n601870 , n601871 , n74549 , 
     n601873 , n74551 , n74552 , n74553 , n601877 , n74555 , n601879 , n74557 , n601881 , n74559 , 
     n74560 , n601884 , n601885 , n74563 , n601887 , n601888 , n74566 , n601890 , n74568 , n601892 , 
     n74570 , n601894 , n601895 , n74573 , n74574 , n601898 , n74576 , n601900 , n601901 , n74579 , 
     n74580 , n601904 , n601905 , n601906 , n74584 , n74585 , n74586 , n74587 , n74588 , n74589 , 
     n601913 , n74591 , n74592 , n601916 , n74594 , n601918 , n74596 , n74597 , n601921 , n601922 , 
     n74600 , n601924 , n601925 , n74603 , n601927 , n601928 , n601929 , n74607 , n601931 , n601932 , 
     n74610 , n601934 , n601935 , n74613 , n74614 , n74615 , n74616 , n74617 , n74618 , n74619 , 
     n74620 , n601944 , n74622 , n601946 , n74624 , n74625 , n601949 , n601950 , n74628 , n601952 , 
     n601953 , n74631 , n601955 , n601956 , n601957 , n74635 , n601959 , n74637 , n74638 , n74639 , 
     n74640 , n74641 , n74642 , n74643 , n74644 , n74645 , n74646 , n74647 , n601971 , n601972 , 
     n601973 , n74651 , n74652 , n601976 , n74654 , n74655 , n601979 , n601980 , n74658 , n601982 , 
     n601983 , n74661 , n601985 , n74663 , n74664 , n601988 , n74666 , n601990 , n74668 , n74669 , 
     n74670 , n74671 , n601995 , n601996 , n74674 , n74675 , n601999 , n602000 , n74678 , n74679 , 
     n74680 , n74681 , n74682 , n74683 , n74684 , n74685 , n74686 , n602010 , n74688 , n602012 , 
     n74690 , n602014 , n74692 , n602016 , n602017 , n74695 , n74696 , n602020 , n602021 , n74699 , 
     n602023 , n602024 , n74702 , n602026 , n602027 , n74705 , n74706 , n602030 , n74708 , n602032 , 
     n74710 , n74711 , n602035 , n74713 , n74714 , n74715 , n74716 , n74717 , n74718 , n74719 , 
     n74720 , n74721 , n74722 , n74723 , n74724 , n74725 , n74726 , n74727 , n74728 , n74729 , 
     n602053 , n74731 , n74732 , n602056 , n602057 , n74735 , n602059 , n602060 , n74738 , n602062 , 
     n602063 , n602064 , n74742 , n602066 , n602067 , n74745 , n602069 , n602070 , n74748 , n74749 , 
     n74750 , n74751 , n74752 , n74753 , n74754 , n74755 , n74756 , n74757 , n74758 , n74759 , 
     n74760 , n74761 , n74762 , n74763 , n74764 , n74765 , n74766 , n74767 , n74768 , n74769 , 
     n74770 , n74771 , n74772 , n74773 , n74774 , n74775 , n602099 , n74777 , n602101 , n74779 , 
     n74780 , n602104 , n74782 , n602106 , n74784 , n74785 , n74786 , n74787 , n74788 , n74789 , 
     n74790 , n74791 , n74792 , n74793 , n74794 , n74795 , n74796 , n602120 , n74798 , n74799 , 
     n74800 , n74801 , n74802 , n74803 , n74804 , n74805 , n74806 , n74807 , n74808 , n74809 , 
     n602133 , n74811 , n602135 , n74813 , n74814 , n74815 , n602139 , n74817 , n74818 , n74819 , 
     n602143 , n602144 , n74822 , n602146 , n602147 , n74825 , n602149 , n602150 , n602151 , n74829 , 
     n602153 , n602154 , n74832 , n602156 , n74834 , n74835 , n74836 , n74837 , n602161 , n74839 , 
     n74840 , n74841 , n602165 , n74843 , n602167 , n74845 , n74846 , n74847 , n74848 , n74849 , 
     n74850 , n602174 , n74852 , n74853 , n602177 , n602178 , n74856 , n602180 , n602181 , n74859 , 
     n602183 , n74861 , n602185 , n74863 , n602187 , n602188 , n74866 , n602190 , n602191 , n74869 , 
     n602193 , n602194 , n74872 , n74873 , n74874 , n74875 , n602199 , n602200 , n74878 , n602202 , 
     n74880 , n602204 , n74882 , n74883 , n602207 , n602208 , n74886 , n602210 , n602211 , n74889 , 
     n602213 , n602214 , n74892 , n74893 , n602217 , n602218 , n74896 , n602220 , n602221 , n74899 , 
     n602223 , n602224 , n602225 , n74903 , n74904 , n74905 , n74906 , n74907 , n602231 , n74909 , 
     n74910 , n602234 , n74912 , n602236 , n74914 , n74915 , n602239 , n74917 , n602241 , n74919 , 
     n602243 , n602244 , n74922 , n602246 , n602247 , n602248 , n74926 , n602250 , n602251 , n74929 , 
     n602253 , n602254 , n74932 , n602256 , n74934 , n602258 , n74936 , n602260 , n74938 , n74939 , 
     n602263 , n602264 , n74942 , n602266 , n602267 , n74945 , n602269 , n602270 , n74948 , n74949 , 
     n602273 , n602274 , n74952 , n602276 , n602277 , n74955 , n602279 , n602280 , n74958 , n602282 , 
     n602283 , n74961 , n602285 , n74963 , n602287 , n74965 , n74966 , n602290 , n74968 , n602292 , 
     n74970 , n602294 , n602295 , n74973 , n602297 , n602298 , n74976 , n74977 , n74978 , n602302 , 
     n74980 , n602304 , n602305 , n602306 , n74984 , n602308 , n602309 , n74987 , n602311 , n602312 , 
     n602313 , n74991 , n602315 , n74993 , n602317 , n74995 , n602319 , n602320 , n74998 , n74999 , 
     n602323 , n602324 , n75002 , n602326 , n602327 , n75005 , n602329 , n602330 , n75008 , n75009 , 
     n602333 , n602334 , n75012 , n602336 , n602337 , n75015 , n602339 , n602340 , n75018 , n75019 , 
     n75020 , n75021 , n75022 , n75023 , n75024 , n75025 , n75026 , n75027 , n75028 , n75029 , 
     n75030 , n75031 , n75032 , n75033 , n75034 , n75035 , n602359 , n75037 , n602361 , n75039 , 
     n602363 , n75041 , n602365 , n75043 , n602367 , n602368 , n75046 , n75047 , n602371 , n75049 , 
     n602373 , n602374 , n602375 , n75053 , n602377 , n602378 , n75056 , n602380 , n602381 , n75059 , 
     n75060 , n602384 , n602385 , n75063 , n602387 , n602388 , n75066 , n602390 , n602391 , n75069 , 
     n75070 , n75071 , n75072 , n75073 , n75074 , n75075 , n75076 , n602400 , n75078 , n602402 , 
     n602403 , n75081 , n75082 , n75083 , n602407 , n602408 , n602409 , n75087 , n602411 , n75089 , 
     n602413 , n75091 , n75092 , n602416 , n602417 , n75095 , n602419 , n602420 , n75098 , n602422 , 
     n602423 , n75101 , n75102 , n602426 , n602427 , n75105 , n602429 , n602430 , n75108 , n602432 , 
     n602433 , n75111 , n602435 , n75113 , n602437 , n75115 , n602439 , n75117 , n75118 , n602442 , 
     n602443 , n75121 , n602445 , n602446 , n75124 , n602448 , n602449 , n75127 , n75128 , n602452 , 
     n602453 , n75131 , n602455 , n602456 , n75134 , n602458 , n602459 , n75137 , n602461 , n602462 , 
     n602463 , n75141 , n602465 , n75143 , n602467 , n75145 , n75146 , n602470 , n602471 , n75149 , 
     n602473 , n602474 , n75152 , n602476 , n602477 , n75155 , n75156 , n602480 , n602481 , n75159 , 
     n602483 , n602484 , n75162 , n602486 , n602487 , n75165 , n75166 , n75167 , n602491 , n75169 , 
     n602493 , n75171 , n602495 , n75173 , n602497 , n75175 , n75176 , n602500 , n75178 , n602502 , 
     n602503 , n602504 , n75182 , n602506 , n602507 , n75185 , n602509 , n602510 , n75188 , n75189 , 
     n602513 , n602514 , n75192 , n602516 , n602517 , n75195 , n602519 , n75197 , n75198 , n75199 , 
     n75200 , n75201 , n75202 , n75203 , n75204 , n75205 , n602529 , n75207 , n75208 , n75209 , 
     n75210 , n75211 , n602535 , n602536 , n75214 , n602538 , n602539 , n75217 , n602541 , n602542 , 
     n75220 , n602544 , n602545 , n75223 , n75224 , n602548 , n75226 , n602550 , n75228 , n602552 , 
     n602553 , n75231 , n75232 , n602556 , n602557 , n75235 , n602559 , n602560 , n602561 , n602562 , 
     n602563 , n602564 , n602565 , n75243 , n602567 , n602568 , n602569 , n602570 , n602571 , n602572 , 
     n602573 , n75251 , n602575 , n75253 , n602577 , n75255 , n602579 , n75257 , n602581 , n75259 , 
     n602583 , n75261 , n602585 , n75263 , n602587 , n602588 , n602589 , n75267 , n602591 , n75269 , 
     n602593 , n75271 , n602595 , n75273 , n602597 , n75275 , n602599 , n602600 , n602601 , n75279 , 
     n602603 , n602604 , n602605 , n602606 , n602607 , n75285 , n602609 , n75287 , n602611 , n602612 , 
     n602613 , n602614 , n602615 , n75293 , n602617 , n75295 , n602619 , n75297 , n602621 , n75299 , 
     n602623 , n75301 , n602625 , n75303 , n602627 , n602628 , n602629 , n602630 , n602631 , n75309 , 
     n602633 , n602634 , n602635 , n602636 , n602637 , n75315 , n602639 , n602640 , n602641 , n75319 , 
     n602643 , n75321 , n602645 , n75323 , n602647 , n75325 , n602649 , n75327 , n602651 , n75329 , 
     n602653 , n602654 , n602655 , n602656 , n602657 , n75335 , n602659 , n602660 , n602661 , n75339 , 
     n602663 , n602664 , n602665 , n75343 , n602667 , n602668 , n602669 , n75347 , n602671 , n75349 , 
     n602673 , n602674 , n602675 , n75353 , n602677 , n75355 , n602679 , n75357 , n602681 , n602682 , 
     n602683 , n75361 , n602685 , n602686 , n602687 , n602688 , n602689 , n602690 , n602691 , n602692 , 
     n602693 , n75371 , n602695 , n75373 , n602697 , n75375 , n602699 , n75377 , n602701 , n75379 , 
     n602703 , n75381 , n602705 , n602706 , n602707 , n602708 , n602709 , n75387 , n602711 , n602712 , 
     n602713 , n602714 , n602715 , n75393 , n602717 , n602718 , n602719 , n75397 , n602721 , n602722 , 
     n602723 , n602724 , n602725 , n75403 , n602727 , n602728 , n602729 , n602730 , n602731 , n602732 , 
     n602733 , n602734 , n602735 , n75413 , n602737 , n602738 , n602739 , n602740 , n602741 , n75419 , 
     n602743 , n602744 , n602745 , n75423 , n602747 , n602748 , n602749 , n75427 , n602751 , n602752 , 
     n602753 , n602754 , n602755 , n602756 , n602757 , n75435 , n75436 , n602760 , n75438 , n602762 , 
     n602763 , n75441 , n75442 , n602766 , n75444 , n75445 , n75446 , n602770 , n75448 , n602772 , 
     n75450 , n75451 , n75452 , n602776 , n75454 , n602778 , n75456 , n75457 , n602781 , n75459 , 
     n602783 , n602784 , n75462 , n75463 , n75464 , n75465 , n75466 , n75467 , n75468 , n75469 , 
     n75470 , n75471 , n75472 , n602796 , n75474 , n602798 , n75476 , n75477 , n75478 , n602802 , 
     n602803 , n75481 , n602805 , n75483 , n602807 , n75485 , n602809 , n602810 , n602811 , n602812 , 
     n75490 , n602814 , n602815 , n75493 , n602817 , n602818 , n602819 , n75497 , n602821 , n75499 , 
     n75500 , n75501 , n75502 , n75503 ;
buf ( n1090  , n0 );
buf ( n1091  , n1 );
buf ( n1092  , n2 );
buf ( n1093  , n3 );
buf ( n1094  , n4 );
buf ( n1095  , n5 );
buf ( n1096  , n6 );
buf ( n1097  , n7 );
buf ( n1098  , n8 );
buf ( n1099  , n9 );
buf ( n1100  , n10 );
buf ( n1101  , n11 );
buf ( n1102  , n12 );
buf ( n1103  , n13 );
buf ( n1104  , n14 );
buf ( n1105  , n15 );
buf ( n1106  , n16 );
buf ( n1107  , n17 );
buf ( n1108  , n18 );
buf ( n1109  , n19 );
buf ( n1110  , n20 );
buf ( n1111  , n21 );
buf ( n1112  , n22 );
buf ( n1113  , n23 );
buf ( n1114  , n24 );
buf ( n1115  , n25 );
buf ( n1116  , n26 );
buf ( n1117  , n27 );
buf ( n1118  , n28 );
buf ( n1119  , n29 );
buf ( n1120  , n30 );
buf ( n1121  , n31 );
buf ( n1122  , n32 );
buf ( n1123  , n33 );
buf ( n1124  , n34 );
buf ( n1125  , n35 );
buf ( n1126  , n36 );
buf ( n1127  , n37 );
buf ( n1128  , n38 );
buf ( n1129  , n39 );
buf ( n1130  , n40 );
buf ( n1131  , n41 );
buf ( n1132  , n42 );
buf ( n1133  , n43 );
buf ( n1134  , n44 );
buf ( n1135  , n45 );
buf ( n1136  , n46 );
buf ( n1137  , n47 );
buf ( n1138  , n48 );
buf ( n1139  , n49 );
buf ( n1140  , n50 );
buf ( n1141  , n51 );
buf ( n1142  , n52 );
buf ( n1143  , n53 );
buf ( n1144  , n54 );
buf ( n1145  , n55 );
buf ( n1146  , n56 );
buf ( n1147  , n57 );
buf ( n1148  , n58 );
buf ( n1149  , n59 );
buf ( n1150  , n60 );
buf ( n1151  , n61 );
buf ( n1152  , n62 );
buf ( n1153  , n63 );
buf ( n1154  , n64 );
buf ( n1155  , n65 );
buf ( n1156  , n66 );
buf ( n1157  , n67 );
buf ( n1158  , n68 );
buf ( n1159  , n69 );
buf ( n1160  , n70 );
buf ( n1161  , n71 );
buf ( n1162  , n72 );
buf ( n1163  , n73 );
buf ( n1164  , n74 );
buf ( n1165  , n75 );
buf ( n1166  , n76 );
buf ( n1167  , n77 );
buf ( n1168  , n78 );
buf ( n1169  , n79 );
buf ( n1170  , n80 );
buf ( n1171  , n81 );
buf ( n1172  , n82 );
buf ( n1173  , n83 );
buf ( n1174  , n84 );
buf ( n1175  , n85 );
buf ( n1176  , n86 );
buf ( n1177  , n87 );
buf ( n1178  , n88 );
buf ( n1179  , n89 );
buf ( n1180  , n90 );
buf ( n1181  , n91 );
buf ( n1182  , n92 );
buf ( n1183  , n93 );
buf ( n1184  , n94 );
buf ( n1185  , n95 );
buf ( n1186  , n96 );
buf ( n1187  , n97 );
buf ( n1188  , n98 );
buf ( n1189  , n99 );
buf ( n1190  , n100 );
buf ( n1191  , n101 );
buf ( n1192  , n102 );
buf ( n1193  , n103 );
buf ( n1194  , n104 );
buf ( n1195  , n105 );
buf ( n1196  , n106 );
buf ( n1197  , n107 );
buf ( n1198  , n108 );
buf ( n1199  , n109 );
buf ( n1200  , n110 );
buf ( n1201  , n111 );
buf ( n1202  , n112 );
buf ( n1203  , n113 );
buf ( n1204  , n114 );
buf ( n1205  , n115 );
buf ( n1206  , n116 );
buf ( n1207  , n117 );
buf ( n1208  , n118 );
buf ( n1209  , n119 );
buf ( n1210  , n120 );
buf ( n1211  , n121 );
buf ( n1212  , n122 );
buf ( n1213  , n123 );
buf ( n1214  , n124 );
buf ( n1215  , n125 );
buf ( n1216  , n126 );
buf ( n1217  , n127 );
buf ( n1218  , n128 );
buf ( n1219  , n129 );
buf ( n1220  , n130 );
buf ( n1221  , n131 );
buf ( n1222  , n132 );
buf ( n1223  , n133 );
buf ( n1224  , n134 );
buf ( n1225  , n135 );
buf ( n1226  , n136 );
buf ( n1227  , n137 );
buf ( n1228  , n138 );
buf ( n1229  , n139 );
buf ( n1230  , n140 );
buf ( n1231  , n141 );
buf ( n1232  , n142 );
buf ( n1233  , n143 );
buf ( n1234  , n144 );
buf ( n1235  , n145 );
buf ( n1236  , n146 );
buf ( n1237  , n147 );
buf ( n1238  , n148 );
buf ( n1239  , n149 );
buf ( n1240  , n150 );
buf ( n1241  , n151 );
buf ( n1242  , n152 );
buf ( n1243  , n153 );
buf ( n1244  , n154 );
buf ( n1245  , n155 );
buf ( n1246  , n156 );
buf ( n1247  , n157 );
buf ( n1248  , n158 );
buf ( n1249  , n159 );
buf ( n160 , n1250 );
buf ( n161 , n1251 );
buf ( n162 , n1252 );
buf ( n163 , n1253 );
buf ( n164 , n1254 );
buf ( n165 , n1255 );
buf ( n166 , n1256 );
buf ( n167 , n1257 );
buf ( n168 , n1258 );
buf ( n169 , n1259 );
buf ( n170 , n1260 );
buf ( n171 , n1261 );
buf ( n172 , n1262 );
buf ( n173 , n1263 );
buf ( n174 , n1264 );
buf ( n175 , n1265 );
buf ( n176 , n1266 );
buf ( n177 , n1267 );
buf ( n178 , n1268 );
buf ( n179 , n1269 );
buf ( n180 , n1270 );
buf ( n181 , n1271 );
buf ( n182 , n1272 );
buf ( n183 , n1273 );
buf ( n184 , n1274 );
buf ( n185 , n1275 );
buf ( n186 , n1276 );
buf ( n187 , n1277 );
buf ( n188 , n1278 );
buf ( n189 , n1279 );
buf ( n190 , n1280 );
buf ( n191 , n1281 );
buf ( n192 , n1282 );
buf ( n193 , n1283 );
buf ( n194 , n1284 );
buf ( n195 , n1285 );
buf ( n196 , n1286 );
buf ( n197 , n1287 );
buf ( n198 , n1288 );
buf ( n199 , n1289 );
buf ( n200 , n1290 );
buf ( n201 , n1291 );
buf ( n202 , n1292 );
buf ( n203 , n1293 );
buf ( n204 , n1294 );
buf ( n205 , n1295 );
buf ( n206 , n1296 );
buf ( n207 , n1297 );
buf ( n208 , n1298 );
buf ( n209 , n1299 );
buf ( n210 , n1300 );
buf ( n211 , n1301 );
buf ( n212 , n1302 );
buf ( n213 , n1303 );
buf ( n214 , n1304 );
buf ( n215 , n1305 );
buf ( n216 , n1306 );
buf ( n217 , n1307 );
buf ( n218 , n1308 );
buf ( n219 , n1309 );
buf ( n220 , n1310 );
buf ( n221 , n1311 );
buf ( n222 , n1312 );
buf ( n223 , n1313 );
buf ( n224 , n1314 );
buf ( n225 , n1315 );
buf ( n226 , n1316 );
buf ( n227 , n1317 );
buf ( n228 , n1318 );
buf ( n229 , n1319 );
buf ( n230 , n1320 );
buf ( n231 , n1321 );
buf ( n232 , n1322 );
buf ( n233 , n1323 );
buf ( n234 , n1324 );
buf ( n235 , n1325 );
buf ( n236 , n1326 );
buf ( n237 , n1327 );
buf ( n238 , n1328 );
buf ( n239 , n1329 );
buf ( n240 , n1330 );
buf ( n241 , n1331 );
buf ( n242 , n1332 );
buf ( n243 , n1333 );
buf ( n244 , n1334 );
buf ( n245 , n1335 );
buf ( n246 , n1336 );
buf ( n247 , n1337 );
buf ( n248 , n1338 );
buf ( n249 , n1339 );
buf ( n250 , n1340 );
buf ( n251 , n1341 );
buf ( n252 , n1342 );
buf ( n253 , n1343 );
buf ( n254 , n1344 );
buf ( n255 , n1345 );
buf ( n256 , n1346 );
buf ( n257 , n1347 );
buf ( n258 , n1348 );
buf ( n259 , n1349 );
buf ( n260 , n1350 );
buf ( n261 , n1351 );
buf ( n262 , n1352 );
buf ( n263 , n1353 );
buf ( n264 , n1354 );
buf ( n265 , n1355 );
buf ( n266 , n1356 );
buf ( n267 , n1357 );
buf ( n268 , n1358 );
buf ( n269 , n1359 );
buf ( n270 , n1360 );
buf ( n271 , n1361 );
buf ( n272 , n1362 );
buf ( n273 , n1363 );
buf ( n274 , n1364 );
buf ( n275 , n1365 );
buf ( n276 , n1366 );
buf ( n277 , n1367 );
buf ( n278 , n1368 );
buf ( n279 , n1369 );
buf ( n280 , n1370 );
buf ( n281 , n1371 );
buf ( n282 , n1372 );
buf ( n283 , n1373 );
buf ( n284 , n1374 );
buf ( n285 , n1375 );
buf ( n286 , n1376 );
buf ( n287 , n1377 );
buf ( n288 , n1378 );
buf ( n289 , n1379 );
buf ( n290 , n1380 );
buf ( n291 , n1381 );
buf ( n292 , n1382 );
buf ( n293 , n1383 );
buf ( n294 , n1384 );
buf ( n295 , n1385 );
buf ( n296 , n1386 );
buf ( n297 , n1387 );
buf ( n298 , n1388 );
buf ( n299 , n1389 );
buf ( n300 , n1390 );
buf ( n301 , n1391 );
buf ( n302 , n1392 );
buf ( n303 , n1393 );
buf ( n304 , n1394 );
buf ( n305 , n1395 );
buf ( n306 , n1396 );
buf ( n307 , n1397 );
buf ( n308 , n1398 );
buf ( n309 , n1399 );
buf ( n310 , n1400 );
buf ( n311 , n1401 );
buf ( n312 , n1402 );
buf ( n313 , n1403 );
buf ( n314 , n1404 );
buf ( n315 , n1405 );
buf ( n316 , n1406 );
buf ( n317 , n1407 );
buf ( n318 , n1408 );
buf ( n319 , n1409 );
buf ( n320 , n1410 );
buf ( n321 , n1411 );
buf ( n322 , n1412 );
buf ( n323 , n1413 );
buf ( n324 , n1414 );
buf ( n325 , n1415 );
buf ( n326 , n1416 );
buf ( n327 , n1417 );
buf ( n328 , n1418 );
buf ( n329 , n1419 );
buf ( n330 , n1420 );
buf ( n331 , n1421 );
buf ( n332 , n1422 );
buf ( n333 , n1423 );
buf ( n334 , n1424 );
buf ( n335 , n1425 );
buf ( n336 , n1426 );
buf ( n337 , n1427 );
buf ( n338 , n1428 );
buf ( n339 , n1429 );
buf ( n340 , n1430 );
buf ( n341 , n1431 );
buf ( n342 , n1432 );
buf ( n343 , n1433 );
buf ( n344 , n1434 );
buf ( n345 , n1435 );
buf ( n346 , n1436 );
buf ( n347 , n1437 );
buf ( n348 , n1438 );
buf ( n349 , n1439 );
buf ( n350 , n1440 );
buf ( n351 , n1441 );
buf ( n352 , n1442 );
buf ( n353 , n1443 );
buf ( n354 , n1444 );
buf ( n355 , n1445 );
buf ( n356 , n1446 );
buf ( n357 , n1447 );
buf ( n358 , n1448 );
buf ( n359 , n1449 );
buf ( n360 , n1450 );
buf ( n361 , n1451 );
buf ( n362 , n1452 );
buf ( n363 , n1453 );
buf ( n364 , n1454 );
buf ( n365 , n1455 );
buf ( n366 , n1456 );
buf ( n367 , n1457 );
buf ( n368 , n1458 );
buf ( n369 , n1459 );
buf ( n370 , n1460 );
buf ( n371 , n1461 );
buf ( n372 , n1462 );
buf ( n373 , n1463 );
buf ( n374 , n1464 );
buf ( n375 , n1465 );
buf ( n376 , n1466 );
buf ( n377 , n1467 );
buf ( n378 , n1468 );
buf ( n379 , n1469 );
buf ( n380 , n1470 );
buf ( n381 , n1471 );
buf ( n382 , n1472 );
buf ( n383 , n1473 );
buf ( n384 , n1474 );
buf ( n385 , n1475 );
buf ( n386 , n1476 );
buf ( n387 , n1477 );
buf ( n388 , n1478 );
buf ( n389 , n1479 );
buf ( n390 , n1480 );
buf ( n391 , n1481 );
buf ( n392 , n1482 );
buf ( n393 , n1483 );
buf ( n394 , n1484 );
buf ( n395 , n1485 );
buf ( n396 , n1486 );
buf ( n397 , n1487 );
buf ( n398 , n1488 );
buf ( n399 , n1489 );
buf ( n400 , n1490 );
buf ( n401 , n1491 );
buf ( n402 , n1492 );
buf ( n403 , n1493 );
buf ( n404 , n1494 );
buf ( n405 , n1495 );
buf ( n406 , n1496 );
buf ( n407 , n1497 );
buf ( n408 , n1498 );
buf ( n409 , n1499 );
buf ( n410 , n1500 );
buf ( n411 , n1501 );
buf ( n412 , n1502 );
buf ( n413 , n1503 );
buf ( n414 , n1504 );
buf ( n415 , n1505 );
buf ( n416 , n1506 );
buf ( n417 , n1507 );
buf ( n418 , n1508 );
buf ( n419 , n1509 );
buf ( n420 , n1510 );
buf ( n421 , n1511 );
buf ( n422 , n1512 );
buf ( n423 , n1513 );
buf ( n424 , n1514 );
buf ( n425 , n1515 );
buf ( n426 , n1516 );
buf ( n427 , n1517 );
buf ( n428 , n1518 );
buf ( n429 , n1519 );
buf ( n430 , n1520 );
buf ( n431 , n1521 );
buf ( n432 , n1522 );
buf ( n433 , n1523 );
buf ( n434 , n1524 );
buf ( n435 , n1525 );
buf ( n436 , n1526 );
buf ( n437 , n1527 );
buf ( n438 , n1528 );
buf ( n439 , n1529 );
buf ( n440 , n1530 );
buf ( n441 , n1531 );
buf ( n442 , n1532 );
buf ( n443 , n1533 );
buf ( n444 , n1534 );
buf ( n445 , n1535 );
buf ( n446 , n1536 );
buf ( n447 , n1537 );
buf ( n448 , n1538 );
buf ( n449 , n1539 );
buf ( n450 , n1540 );
buf ( n451 , n1541 );
buf ( n452 , n1542 );
buf ( n453 , n1543 );
buf ( n454 , n1544 );
buf ( n455 , n1545 );
buf ( n456 , n1546 );
buf ( n457 , n1547 );
buf ( n458 , n1548 );
buf ( n459 , n1549 );
buf ( n460 , n1550 );
buf ( n461 , n1551 );
buf ( n462 , n1552 );
buf ( n463 , n1553 );
buf ( n464 , n1554 );
buf ( n465 , n1555 );
buf ( n466 , n1556 );
buf ( n467 , n1557 );
buf ( n468 , n1558 );
buf ( n469 , n1559 );
buf ( n470 , n1560 );
buf ( n471 , n1561 );
buf ( n472 , n1562 );
buf ( n473 , n1563 );
buf ( n474 , n1564 );
buf ( n475 , n1565 );
buf ( n476 , n1566 );
buf ( n477 , n1567 );
buf ( n478 , n1568 );
buf ( n479 , n1569 );
buf ( n480 , n1570 );
buf ( n481 , n1571 );
buf ( n482 , n1572 );
buf ( n483 , n1573 );
buf ( n484 , n1574 );
buf ( n485 , n1575 );
buf ( n486 , n1576 );
buf ( n487 , n1577 );
buf ( n488 , n1578 );
buf ( n489 , n1579 );
buf ( n490 , n1580 );
buf ( n491 , n1581 );
buf ( n492 , n1582 );
buf ( n493 , n1583 );
buf ( n494 , n1584 );
buf ( n495 , n1585 );
buf ( n496 , n1586 );
buf ( n497 , n1587 );
buf ( n498 , n1588 );
buf ( n499 , n1589 );
buf ( n500 , n1590 );
buf ( n501 , n1591 );
buf ( n502 , n1592 );
buf ( n503 , n1593 );
buf ( n504 , n1594 );
buf ( n505 , n1595 );
buf ( n506 , n1596 );
buf ( n507 , n1597 );
buf ( n508 , n1598 );
buf ( n509 , n1599 );
buf ( n510 , n1600 );
buf ( n511 , n1601 );
buf ( n512 , n1602 );
buf ( n513 , n1603 );
buf ( n514 , n1604 );
buf ( n515 , n1605 );
buf ( n516 , n1606 );
buf ( n517 , n1607 );
buf ( n518 , n1608 );
buf ( n519 , n1609 );
buf ( n520 , n1610 );
buf ( n521 , n1611 );
buf ( n522 , n1612 );
buf ( n523 , n1613 );
buf ( n524 , n1614 );
buf ( n525 , n1615 );
buf ( n526 , n1616 );
buf ( n527 , n1617 );
buf ( n528 , n1618 );
buf ( n529 , n1619 );
buf ( n530 , n1620 );
buf ( n531 , n1621 );
buf ( n532 , n1622 );
buf ( n533 , n1623 );
buf ( n534 , n1624 );
buf ( n535 , n1625 );
buf ( n536 , n1626 );
buf ( n537 , n1627 );
buf ( n538 , n1628 );
buf ( n539 , n1629 );
buf ( n540 , n1630 );
buf ( n541 , n1631 );
buf ( n542 , n1632 );
buf ( n543 , n1633 );
buf ( n544 , n1634 );
buf ( n1250 , 1'b0 );
buf ( n1251 , 1'b0 );
buf ( n1252 , 1'b0 );
buf ( n1253 , 1'b0 );
buf ( n1254 , 1'b0 );
buf ( n1255 , 1'b0 );
buf ( n1256 , 1'b0 );
buf ( n1257 , 1'b0 );
buf ( n1258 , 1'b0 );
buf ( n1259 , 1'b0 );
buf ( n1260 , 1'b0 );
buf ( n1261 , 1'b0 );
buf ( n1262 , 1'b0 );
buf ( n1263 , 1'b0 );
buf ( n1264 , 1'b0 );
buf ( n1265 , 1'b0 );
buf ( n1266 , 1'b0 );
buf ( n1267 , 1'b0 );
buf ( n1268 , 1'b0 );
buf ( n1269 , 1'b0 );
buf ( n1270 , 1'b0 );
buf ( n1271 , 1'b0 );
buf ( n1272 , 1'b0 );
buf ( n1273 , 1'b0 );
buf ( n1274 , 1'b0 );
buf ( n1275 , 1'b0 );
buf ( n1276 , 1'b0 );
buf ( n1277 , 1'b0 );
buf ( n1278 , 1'b0 );
buf ( n1279 , 1'b0 );
buf ( n1280 , 1'b0 );
buf ( n1281 , n602561 );
buf ( n1282 , n602563 );
buf ( n1283 , n602565 );
buf ( n1284 , n602567 );
buf ( n1285 , n602569 );
buf ( n1286 , n602571 );
buf ( n1287 , n602573 );
buf ( n1288 , n602575 );
buf ( n1289 , n602577 );
buf ( n1290 , n602579 );
buf ( n1291 , n602581 );
buf ( n1292 , n602583 );
buf ( n1293 , n602585 );
buf ( n1294 , n602587 );
buf ( n1295 , n602589 );
buf ( n1296 , n602591 );
buf ( n1297 , n602593 );
buf ( n1298 , n602595 );
buf ( n1299 , n602597 );
buf ( n1300 , n602599 );
buf ( n1301 , n602601 );
buf ( n1302 , n602603 );
buf ( n1303 , n602605 );
buf ( n1304 , n602607 );
buf ( n1305 , n602609 );
buf ( n1306 , n602611 );
buf ( n1307 , n602613 );
buf ( n1308 , n602615 );
buf ( n1309 , n602617 );
buf ( n1310 , n602619 );
buf ( n1311 , n602621 );
buf ( n1312 , n602623 );
buf ( n1313 , n602625 );
buf ( n1314 , n602627 );
buf ( n1315 , n602629 );
buf ( n1316 , n602631 );
buf ( n1317 , n602633 );
buf ( n1318 , n602635 );
buf ( n1319 , n602637 );
buf ( n1320 , n602639 );
buf ( n1321 , n602641 );
buf ( n1322 , n602643 );
buf ( n1323 , n602645 );
buf ( n1324 , n602647 );
buf ( n1325 , n602649 );
buf ( n1326 , n602651 );
buf ( n1327 , n602653 );
buf ( n1328 , n602655 );
buf ( n1329 , n602657 );
buf ( n1330 , n602659 );
buf ( n1331 , n602661 );
buf ( n1332 , n602663 );
buf ( n1333 , n602665 );
buf ( n1334 , n602667 );
buf ( n1335 , n602669 );
buf ( n1336 , n602671 );
buf ( n1337 , n602673 );
buf ( n1338 , n602675 );
buf ( n1339 , n602677 );
buf ( n1340 , n602679 );
buf ( n1341 , n602681 );
buf ( n1342 , n602683 );
buf ( n1343 , n602685 );
buf ( n1344 , n602687 );
buf ( n1345 , n602689 );
buf ( n1346 , n602691 );
buf ( n1347 , n602693 );
buf ( n1348 , n602695 );
buf ( n1349 , n602697 );
buf ( n1350 , n602699 );
buf ( n1351 , n602701 );
buf ( n1352 , n602703 );
buf ( n1353 , n602705 );
buf ( n1354 , n602707 );
buf ( n1355 , n602709 );
buf ( n1356 , n602711 );
buf ( n1357 , n602713 );
buf ( n1358 , n602715 );
buf ( n1359 , n602717 );
buf ( n1360 , n602719 );
buf ( n1361 , n602721 );
buf ( n1362 , n602723 );
buf ( n1363 , n602725 );
buf ( n1364 , n602727 );
buf ( n1365 , n602729 );
buf ( n1366 , n602731 );
buf ( n1367 , n602733 );
buf ( n1368 , n602735 );
buf ( n1369 , n602737 );
buf ( n1370 , n602739 );
buf ( n1371 , n602741 );
buf ( n1372 , n602743 );
buf ( n1373 , n602745 );
buf ( n1374 , n602747 );
buf ( n1375 , n602749 );
buf ( n1376 , n602751 );
buf ( n1377 , n602753 );
buf ( n1378 , 1'b0 );
buf ( n1379 , 1'b0 );
buf ( n1380 , 1'b0 );
buf ( n1381 , 1'b0 );
buf ( n1382 , 1'b0 );
buf ( n1383 , 1'b0 );
buf ( n1384 , 1'b0 );
buf ( n1385 , 1'b0 );
buf ( n1386 , 1'b0 );
buf ( n1387 , 1'b0 );
buf ( n1388 , 1'b0 );
buf ( n1389 , 1'b0 );
buf ( n1390 , 1'b0 );
buf ( n1391 , 1'b0 );
buf ( n1392 , 1'b0 );
buf ( n1393 , 1'b0 );
buf ( n1394 , 1'b0 );
buf ( n1395 , 1'b0 );
buf ( n1396 , 1'b0 );
buf ( n1397 , 1'b0 );
buf ( n1398 , 1'b0 );
buf ( n1399 , 1'b0 );
buf ( n1400 , n591458 );
buf ( n1401 , n591460 );
buf ( n1402 , n591462 );
buf ( n1403 , n591464 );
buf ( n1404 , n591466 );
buf ( n1405 , n591468 );
buf ( n1406 , n591470 );
buf ( n1407 , n591472 );
buf ( n1408 , n591474 );
buf ( n1409 , n591476 );
buf ( n1410 , n591478 );
buf ( n1411 , n591480 );
buf ( n1412 , n591482 );
buf ( n1413 , n591484 );
buf ( n1414 , n591486 );
buf ( n1415 , n591488 );
buf ( n1416 , n591490 );
buf ( n1417 , n591492 );
buf ( n1418 , n591494 );
buf ( n1419 , n591496 );
buf ( n1420 , n591498 );
buf ( n1421 , n591500 );
buf ( n1422 , n591502 );
buf ( n1423 , n591504 );
buf ( n1424 , n591506 );
buf ( n1425 , n591508 );
buf ( n1426 , n591510 );
buf ( n1427 , n591512 );
buf ( n1428 , n591514 );
buf ( n1429 , n591516 );
buf ( n1430 , n591518 );
buf ( n1431 , n591520 );
buf ( n1432 , n591522 );
buf ( n1433 , n591524 );
buf ( n1434 , n591526 );
buf ( n1435 , n591528 );
buf ( n1436 , n591530 );
buf ( n1437 , n591532 );
buf ( n1438 , n591534 );
buf ( n1439 , n591536 );
buf ( n1440 , n591538 );
buf ( n1441 , n591540 );
buf ( n1442 , n591542 );
buf ( n1443 , n591544 );
buf ( n1444 , n591546 );
buf ( n1445 , n591548 );
buf ( n1446 , n591550 );
buf ( n1447 , n591552 );
buf ( n1448 , n591554 );
buf ( n1449 , n591556 );
buf ( n1450 , n591558 );
buf ( n1451 , n591560 );
buf ( n1452 , n591562 );
buf ( n1453 , n591564 );
buf ( n1454 , n591566 );
buf ( n1455 , n591568 );
buf ( n1456 , n591570 );
buf ( n1457 , n591572 );
buf ( n1458 , n591574 );
buf ( n1459 , n591576 );
buf ( n1460 , n591578 );
buf ( n1461 , n591580 );
buf ( n1462 , n591582 );
buf ( n1463 , n591584 );
buf ( n1464 , n591586 );
buf ( n1465 , n591588 );
buf ( n1466 , n591590 );
buf ( n1467 , n591592 );
buf ( n1468 , n591594 );
buf ( n1469 , n591596 );
buf ( n1470 , n591598 );
buf ( n1471 , n591600 );
buf ( n1472 , n591602 );
buf ( n1473 , n591604 );
buf ( n1474 , n591606 );
buf ( n1475 , n591608 );
buf ( n1476 , n591610 );
buf ( n1477 , n591612 );
buf ( n1478 , n591614 );
buf ( n1479 , n591616 );
buf ( n1480 , n591618 );
buf ( n1481 , n591620 );
buf ( n1482 , n591622 );
buf ( n1483 , n591624 );
buf ( n1484 , n591626 );
buf ( n1485 , n591628 );
buf ( n1486 , n591630 );
buf ( n1487 , n591632 );
buf ( n1488 , n591634 );
buf ( n1489 , n591636 );
buf ( n1490 , n591638 );
buf ( n1491 , n591640 );
buf ( n1492 , n591642 );
buf ( n1493 , n591644 );
buf ( n1494 , n591646 );
buf ( n1495 , n591648 );
buf ( n1496 , n591650 );
buf ( n1497 , n591652 );
buf ( n1498 , n591654 );
buf ( n1499 , n591656 );
buf ( n1500 , n591658 );
buf ( n1501 , n591660 );
buf ( n1502 , n591662 );
buf ( n1503 , n591664 );
buf ( n1504 , n591666 );
buf ( n1505 , n591668 );
buf ( n1506 , n578582 );
buf ( n1507 , n578584 );
buf ( n1508 , n578586 );
buf ( n1509 , n578588 );
buf ( n1510 , n578590 );
buf ( n1511 , n578592 );
buf ( n1512 , n578594 );
buf ( n1513 , n578596 );
buf ( n1514 , n578598 );
buf ( n1515 , n578600 );
buf ( n1516 , n578602 );
buf ( n1517 , n578604 );
buf ( n1518 , n578606 );
buf ( n1519 , n578608 );
buf ( n1520 , n578610 );
buf ( n1521 , n578612 );
buf ( n1522 , n578614 );
buf ( n1523 , n578616 );
buf ( n1524 , n578618 );
buf ( n1525 , n578620 );
buf ( n1526 , n578622 );
buf ( n1527 , n578624 );
buf ( n1528 , n578626 );
buf ( n1529 , n578628 );
buf ( n1530 , n578630 );
buf ( n1531 , n578632 );
buf ( n1532 , n578634 );
buf ( n1533 , n578636 );
buf ( n1534 , n578638 );
buf ( n1535 , n578639 );
buf ( n1536 , n578641 );
buf ( n1537 , n578643 );
buf ( n1538 , n578645 );
buf ( n1539 , n578647 );
buf ( n1540 , n578649 );
buf ( n1541 , n578651 );
buf ( n1542 , n578653 );
buf ( n1543 , n578655 );
buf ( n1544 , n578657 );
buf ( n1545 , n578659 );
buf ( n1546 , n578661 );
buf ( n1547 , n578663 );
buf ( n1548 , n578665 );
buf ( n1549 , n578667 );
buf ( n1550 , n578669 );
buf ( n1551 , n578671 );
buf ( n1552 , n578673 );
buf ( n1553 , n578675 );
buf ( n1554 , n578677 );
buf ( n1555 , n578679 );
buf ( n1556 , n578681 );
buf ( n1557 , n578683 );
buf ( n1558 , n578685 );
buf ( n1559 , n578687 );
buf ( n1560 , n578689 );
buf ( n1561 , n578691 );
buf ( n1562 , n578693 );
buf ( n1563 , n578695 );
buf ( n1564 , n578697 );
buf ( n1565 , n578699 );
buf ( n1566 , n578701 );
buf ( n1567 , n578703 );
buf ( n1568 , n578705 );
buf ( n1569 , n578707 );
buf ( n1570 , n578709 );
buf ( n1571 , n578711 );
buf ( n1572 , n578713 );
buf ( n1573 , n578715 );
buf ( n1574 , n578717 );
buf ( n1575 , n578719 );
buf ( n1576 , n578721 );
buf ( n1577 , n578723 );
buf ( n1578 , n578725 );
buf ( n1579 , n578727 );
buf ( n1580 , n578729 );
buf ( n1581 , n578731 );
buf ( n1582 , n578733 );
buf ( n1583 , n578735 );
buf ( n1584 , n578737 );
buf ( n1585 , n578739 );
buf ( n1586 , n578741 );
buf ( n1587 , n578743 );
buf ( n1588 , n578745 );
buf ( n1589 , n578747 );
buf ( n1590 , n578749 );
buf ( n1591 , n578751 );
buf ( n1592 , n578753 );
buf ( n1593 , n578755 );
buf ( n1594 , n578757 );
buf ( n1595 , n578759 );
buf ( n1596 , n578761 );
buf ( n1597 , n578763 );
buf ( n1598 , n578765 );
buf ( n1599 , n578767 );
buf ( n1600 , n578769 );
buf ( n1601 , n578771 );
buf ( n1602 , n578773 );
buf ( n1603 , n578775 );
buf ( n1604 , n578777 );
buf ( n1605 , n578779 );
buf ( n1606 , n578781 );
buf ( n1607 , n578783 );
buf ( n1608 , n578785 );
buf ( n1609 , n578787 );
buf ( n1610 , n578789 );
buf ( n1611 , n578791 );
buf ( n1612 , n578793 );
buf ( n1613 , n578795 );
buf ( n1614 , n578797 );
buf ( n1615 , n578800 );
buf ( n1616 , n578803 );
buf ( n1617 , n578806 );
buf ( n1618 , n578809 );
buf ( n1619 , n578812 );
buf ( n1620 , n578815 );
buf ( n1621 , n578818 );
buf ( n1622 , n578821 );
buf ( n1623 , n578824 );
buf ( n1624 , n578827 );
buf ( n1625 , n578830 );
buf ( n1626 , n578833 );
buf ( n1627 , n578836 );
buf ( n1628 , n578839 );
buf ( n1629 , n578842 );
buf ( n1630 , n578845 );
buf ( n1631 , n578848 );
buf ( n1632 , n578851 );
buf ( n1633 , n578854 );
buf ( n1634 , n578856 );
buf ( n529140 , n1131 );
buf ( n1883 , n529140 );
buf ( n529142 , n1164 );
buf ( n1885 , n529142 );
buf ( n529144 , n1165 );
buf ( n1887 , n529144 );
xor ( n1888 , n1885 , n1887 );
buf ( n529147 , n1166 );
buf ( n1890 , n529147 );
xor ( n1891 , n1887 , n1890 );
not ( n1892 , n1891 );
and ( n1893 , n1888 , n1892 );
and ( n1894 , n1883 , n1893 );
buf ( n529153 , n1130 );
buf ( n1896 , n529153 );
and ( n1897 , n1896 , n1891 );
nor ( n1898 , n1894 , n1897 );
and ( n1899 , n1887 , n1890 );
not ( n1900 , n1899 );
and ( n1901 , n1885 , n1900 );
xnor ( n1902 , n1898 , n1901 );
buf ( n529161 , n1133 );
buf ( n1904 , n529161 );
buf ( n529163 , n1162 );
buf ( n1906 , n529163 );
buf ( n529165 , n1163 );
buf ( n1908 , n529165 );
xor ( n1909 , n1906 , n1908 );
xor ( n1910 , n1908 , n1885 );
not ( n1911 , n1910 );
and ( n1912 , n1909 , n1911 );
and ( n1913 , n1904 , n1912 );
buf ( n529172 , n1132 );
buf ( n1915 , n529172 );
and ( n1916 , n1915 , n1910 );
nor ( n1917 , n1913 , n1916 );
and ( n1918 , n1908 , n1885 );
not ( n1919 , n1918 );
and ( n1920 , n1906 , n1919 );
xnor ( n1921 , n1917 , n1920 );
and ( n1922 , n1902 , n1921 );
buf ( n529181 , n1142 );
buf ( n1924 , n529181 );
buf ( n529183 , n1154 );
buf ( n1926 , n529183 );
and ( n1927 , n1924 , n1926 );
and ( n1928 , n1921 , n1927 );
and ( n1929 , n1902 , n1927 );
or ( n1930 , n1922 , n1928 , n1929 );
buf ( n529189 , n1174 );
buf ( n1932 , n529189 );
buf ( n529191 , n1175 );
buf ( n1934 , n529191 );
buf ( n529193 , n1176 );
buf ( n1936 , n529193 );
and ( n1937 , n1934 , n1936 );
not ( n1938 , n1937 );
and ( n1939 , n1932 , n1938 );
not ( n1940 , n1939 );
buf ( n529199 , n1123 );
buf ( n1942 , n529199 );
buf ( n529201 , n1172 );
buf ( n1944 , n529201 );
buf ( n529203 , n1173 );
buf ( n1946 , n529203 );
xor ( n1947 , n1944 , n1946 );
xor ( n1948 , n1946 , n1932 );
not ( n1949 , n1948 );
and ( n1950 , n1947 , n1949 );
and ( n1951 , n1942 , n1950 );
buf ( n529210 , n1122 );
buf ( n1953 , n529210 );
and ( n1954 , n1953 , n1948 );
nor ( n1955 , n1951 , n1954 );
and ( n1956 , n1946 , n1932 );
not ( n1957 , n1956 );
and ( n1958 , n1944 , n1957 );
xnor ( n1959 , n1955 , n1958 );
and ( n1960 , n1940 , n1959 );
buf ( n529219 , n1127 );
buf ( n1962 , n529219 );
buf ( n529221 , n1168 );
buf ( n1964 , n529221 );
buf ( n529223 , n1169 );
buf ( n1966 , n529223 );
xor ( n1967 , n1964 , n1966 );
buf ( n529226 , n1170 );
buf ( n1969 , n529226 );
xor ( n1970 , n1966 , n1969 );
not ( n1971 , n1970 );
and ( n1972 , n1967 , n1971 );
and ( n1973 , n1962 , n1972 );
buf ( n529232 , n1126 );
buf ( n1975 , n529232 );
and ( n1976 , n1975 , n1970 );
nor ( n1977 , n1973 , n1976 );
and ( n1978 , n1966 , n1969 );
not ( n1979 , n1978 );
and ( n1980 , n1964 , n1979 );
xnor ( n1981 , n1977 , n1980 );
and ( n1982 , n1959 , n1981 );
and ( n1983 , n1940 , n1981 );
or ( n1984 , n1960 , n1982 , n1983 );
and ( n1985 , n1930 , n1984 );
buf ( n529244 , n1129 );
buf ( n1987 , n529244 );
buf ( n529246 , n1167 );
buf ( n1989 , n529246 );
xor ( n1990 , n1890 , n1989 );
xor ( n1991 , n1989 , n1964 );
not ( n1992 , n1991 );
and ( n1993 , n1990 , n1992 );
and ( n1994 , n1987 , n1993 );
buf ( n529253 , n1128 );
buf ( n1996 , n529253 );
and ( n1997 , n1996 , n1991 );
nor ( n1998 , n1994 , n1997 );
and ( n1999 , n1989 , n1964 );
not ( n2000 , n1999 );
and ( n2001 , n1890 , n2000 );
xnor ( n2002 , n1998 , n2001 );
buf ( n529261 , n1135 );
buf ( n2004 , n529261 );
buf ( n529263 , n1160 );
buf ( n2006 , n529263 );
buf ( n529265 , n1161 );
buf ( n2008 , n529265 );
xor ( n2009 , n2006 , n2008 );
xor ( n2010 , n2008 , n1906 );
not ( n2011 , n2010 );
and ( n2012 , n2009 , n2011 );
and ( n2013 , n2004 , n2012 );
buf ( n529272 , n1134 );
buf ( n2015 , n529272 );
and ( n2016 , n2015 , n2010 );
nor ( n2017 , n2013 , n2016 );
and ( n2018 , n2008 , n1906 );
not ( n2019 , n2018 );
and ( n2020 , n2006 , n2019 );
xnor ( n2021 , n2017 , n2020 );
and ( n2022 , n2002 , n2021 );
buf ( n529281 , n1137 );
buf ( n2024 , n529281 );
buf ( n529283 , n1158 );
buf ( n2026 , n529283 );
buf ( n529285 , n1159 );
buf ( n2028 , n529285 );
xor ( n2029 , n2026 , n2028 );
xor ( n2030 , n2028 , n2006 );
not ( n2031 , n2030 );
and ( n2032 , n2029 , n2031 );
and ( n2033 , n2024 , n2032 );
buf ( n529292 , n1136 );
buf ( n2035 , n529292 );
and ( n2036 , n2035 , n2030 );
nor ( n2037 , n2033 , n2036 );
and ( n2038 , n2028 , n2006 );
not ( n2039 , n2038 );
and ( n2040 , n2026 , n2039 );
xnor ( n2041 , n2037 , n2040 );
and ( n2042 , n2021 , n2041 );
and ( n2043 , n2002 , n2041 );
or ( n2044 , n2022 , n2042 , n2043 );
and ( n2045 , n1984 , n2044 );
and ( n2046 , n1930 , n2044 );
or ( n2047 , n1985 , n2045 , n2046 );
buf ( n529306 , n1125 );
buf ( n2049 , n529306 );
buf ( n529308 , n1171 );
buf ( n2050 , n529308 );
xor ( n2051 , n1969 , n2050 );
xor ( n2052 , n2050 , n1944 );
not ( n2053 , n2052 );
and ( n2054 , n2051 , n2053 );
and ( n2055 , n2049 , n2054 );
buf ( n529315 , n1124 );
buf ( n2057 , n529315 );
and ( n2058 , n2057 , n2052 );
nor ( n2059 , n2055 , n2058 );
and ( n2060 , n2050 , n1944 );
not ( n2061 , n2060 );
and ( n2062 , n1969 , n2061 );
xnor ( n2063 , n2059 , n2062 );
buf ( n529323 , n1139 );
buf ( n2065 , n529323 );
buf ( n529325 , n1156 );
buf ( n2067 , n529325 );
buf ( n529327 , n1157 );
buf ( n2069 , n529327 );
xor ( n2070 , n2067 , n2069 );
xor ( n2071 , n2069 , n2026 );
not ( n2072 , n2071 );
and ( n2073 , n2070 , n2072 );
and ( n2074 , n2065 , n2073 );
buf ( n529334 , n1138 );
buf ( n2076 , n529334 );
and ( n2077 , n2076 , n2071 );
nor ( n2078 , n2074 , n2077 );
and ( n2079 , n2069 , n2026 );
not ( n2080 , n2079 );
and ( n2081 , n2067 , n2080 );
xnor ( n2082 , n2078 , n2081 );
and ( n2083 , n2063 , n2082 );
buf ( n529343 , n1141 );
buf ( n2085 , n529343 );
buf ( n529345 , n1155 );
buf ( n2087 , n529345 );
xor ( n2088 , n1926 , n2087 );
xor ( n2089 , n2087 , n2067 );
not ( n2090 , n2089 );
and ( n2091 , n2088 , n2090 );
and ( n2092 , n2085 , n2091 );
buf ( n529352 , n1140 );
buf ( n2094 , n529352 );
and ( n2095 , n2094 , n2089 );
nor ( n2096 , n2092 , n2095 );
and ( n2097 , n2087 , n2067 );
not ( n2098 , n2097 );
and ( n2099 , n1926 , n2098 );
xnor ( n2100 , n2096 , n2099 );
and ( n2101 , n2082 , n2100 );
and ( n2102 , n2063 , n2100 );
or ( n2103 , n2083 , n2101 , n2102 );
and ( n2104 , n2057 , n2054 );
and ( n2105 , n1942 , n2052 );
nor ( n2106 , n2104 , n2105 );
xnor ( n2107 , n2106 , n2062 );
not ( n2108 , n2107 );
and ( n2109 , n2103 , n2108 );
and ( n2110 , n2015 , n2012 );
and ( n2111 , n1904 , n2010 );
nor ( n2112 , n2110 , n2111 );
xnor ( n2113 , n2112 , n2020 );
and ( n2114 , n2108 , n2113 );
and ( n2115 , n2103 , n2113 );
or ( n2116 , n2109 , n2114 , n2115 );
and ( n2117 , n2047 , n2116 );
buf ( n2118 , n2107 );
and ( n2119 , n1883 , n1912 );
and ( n2120 , n1896 , n1910 );
nor ( n2121 , n2119 , n2120 );
xnor ( n2122 , n2121 , n1920 );
xor ( n2123 , n2118 , n2122 );
and ( n2124 , n1904 , n2012 );
and ( n2125 , n1915 , n2010 );
nor ( n2126 , n2124 , n2125 );
xnor ( n2127 , n2126 , n2020 );
xor ( n2128 , n2123 , n2127 );
and ( n2129 , n2116 , n2128 );
and ( n2130 , n2047 , n2128 );
or ( n2131 , n2117 , n2129 , n2130 );
and ( n2132 , n1953 , n1950 );
not ( n2133 , n2132 );
xnor ( n2134 , n2133 , n1958 );
and ( n2135 , n1975 , n1972 );
and ( n2136 , n2049 , n1970 );
nor ( n2137 , n2135 , n2136 );
xnor ( n2138 , n2137 , n1980 );
xor ( n2139 , n2134 , n2138 );
and ( n2140 , n1915 , n1912 );
and ( n2141 , n1883 , n1910 );
nor ( n2142 , n2140 , n2141 );
xnor ( n2143 , n2142 , n1920 );
xor ( n2144 , n2139 , n2143 );
and ( n2145 , n1896 , n1893 );
and ( n2146 , n1987 , n1891 );
nor ( n2147 , n2145 , n2146 );
xnor ( n2148 , n2147 , n1901 );
and ( n2149 , n2094 , n2091 );
and ( n2150 , n2065 , n2089 );
nor ( n2151 , n2149 , n2150 );
xnor ( n2152 , n2151 , n2099 );
xor ( n2153 , n2148 , n2152 );
and ( n2154 , n2085 , n1926 );
xor ( n2155 , n2153 , n2154 );
and ( n2156 , n2144 , n2155 );
and ( n2157 , n1996 , n1993 );
and ( n2158 , n1962 , n1991 );
nor ( n2159 , n2157 , n2158 );
xnor ( n2160 , n2159 , n2001 );
and ( n2161 , n2035 , n2032 );
and ( n2162 , n2004 , n2030 );
nor ( n2163 , n2161 , n2162 );
xnor ( n2164 , n2163 , n2040 );
xor ( n2165 , n2160 , n2164 );
and ( n2166 , n2076 , n2073 );
and ( n2167 , n2024 , n2071 );
nor ( n2168 , n2166 , n2167 );
xnor ( n2169 , n2168 , n2081 );
xor ( n2170 , n2165 , n2169 );
and ( n2171 , n2155 , n2170 );
and ( n2172 , n2144 , n2170 );
or ( n2173 , n2156 , n2171 , n2172 );
and ( n2174 , n2134 , n2138 );
and ( n2175 , n2138 , n2143 );
and ( n2176 , n2134 , n2143 );
or ( n2177 , n2174 , n2175 , n2176 );
and ( n2178 , n2148 , n2152 );
and ( n2179 , n2152 , n2154 );
and ( n2180 , n2148 , n2154 );
or ( n2181 , n2178 , n2179 , n2180 );
xor ( n2182 , n2177 , n2181 );
and ( n2183 , n2160 , n2164 );
and ( n2184 , n2164 , n2169 );
and ( n2185 , n2160 , n2169 );
or ( n2186 , n2183 , n2184 , n2185 );
xor ( n2187 , n2182 , n2186 );
and ( n2188 , n2173 , n2187 );
and ( n2189 , n1987 , n1893 );
and ( n2190 , n1996 , n1891 );
nor ( n2191 , n2189 , n2190 );
xnor ( n2192 , n2191 , n1901 );
and ( n2193 , n2004 , n2032 );
and ( n2194 , n2015 , n2030 );
nor ( n2195 , n2193 , n2194 );
xnor ( n2196 , n2195 , n2040 );
xor ( n2197 , n2192 , n2196 );
and ( n2198 , n2024 , n2073 );
and ( n2199 , n2035 , n2071 );
nor ( n2200 , n2198 , n2199 );
xnor ( n2201 , n2200 , n2081 );
xor ( n2202 , n2197 , n2201 );
and ( n2203 , n2049 , n1972 );
and ( n2204 , n2057 , n1970 );
nor ( n2205 , n2203 , n2204 );
xnor ( n2206 , n2205 , n1980 );
and ( n2207 , n2065 , n2091 );
and ( n2208 , n2076 , n2089 );
nor ( n2209 , n2207 , n2208 );
xnor ( n2210 , n2209 , n2099 );
xor ( n2211 , n2206 , n2210 );
and ( n2212 , n2094 , n1926 );
xor ( n2213 , n2211 , n2212 );
xor ( n2214 , n2202 , n2213 );
not ( n2215 , n1958 );
and ( n2216 , n1942 , n2054 );
and ( n2217 , n1953 , n2052 );
nor ( n2218 , n2216 , n2217 );
xnor ( n2219 , n2218 , n2062 );
xor ( n2220 , n2215 , n2219 );
and ( n2221 , n1962 , n1993 );
and ( n2222 , n1975 , n1991 );
nor ( n2223 , n2221 , n2222 );
xnor ( n2224 , n2223 , n2001 );
xor ( n2225 , n2220 , n2224 );
xor ( n2226 , n2214 , n2225 );
and ( n2227 , n2187 , n2226 );
and ( n2228 , n2173 , n2226 );
or ( n2229 , n2188 , n2227 , n2228 );
and ( n2230 , n2131 , n2229 );
and ( n2231 , n2177 , n2181 );
and ( n2232 , n2181 , n2186 );
and ( n2233 , n2177 , n2186 );
or ( n2234 , n2231 , n2232 , n2233 );
and ( n2235 , n2118 , n2122 );
and ( n2236 , n2122 , n2127 );
and ( n2237 , n2118 , n2127 );
or ( n2238 , n2235 , n2236 , n2237 );
xor ( n2239 , n2234 , n2238 );
and ( n2240 , n1975 , n1993 );
and ( n2241 , n2049 , n1991 );
nor ( n2242 , n2240 , n2241 );
xnor ( n2243 , n2242 , n2001 );
and ( n2244 , n1915 , n2012 );
and ( n2245 , n1883 , n2010 );
nor ( n2246 , n2244 , n2245 );
xnor ( n2247 , n2246 , n2020 );
xor ( n2248 , n2243 , n2247 );
and ( n2249 , n2015 , n2032 );
and ( n2250 , n1904 , n2030 );
nor ( n2251 , n2249 , n2250 );
xnor ( n2252 , n2251 , n2040 );
xor ( n2253 , n2248 , n2252 );
xor ( n2254 , n2239 , n2253 );
and ( n2255 , n2229 , n2254 );
and ( n2256 , n2131 , n2254 );
or ( n2257 , n2230 , n2255 , n2256 );
and ( n2258 , n2192 , n2196 );
and ( n2259 , n2196 , n2201 );
and ( n2260 , n2192 , n2201 );
or ( n2261 , n2258 , n2259 , n2260 );
and ( n2262 , n2215 , n2219 );
and ( n2263 , n2219 , n2224 );
and ( n2264 , n2215 , n2224 );
or ( n2265 , n2262 , n2263 , n2264 );
and ( n2266 , n2261 , n2265 );
and ( n2267 , n1953 , n2054 );
not ( n2268 , n2267 );
xnor ( n2269 , n2268 , n2062 );
not ( n2270 , n2269 );
and ( n2271 , n2265 , n2270 );
and ( n2272 , n2261 , n2270 );
or ( n2273 , n2266 , n2271 , n2272 );
and ( n2274 , n2206 , n2210 );
and ( n2275 , n2210 , n2212 );
and ( n2276 , n2206 , n2212 );
or ( n2277 , n2274 , n2275 , n2276 );
and ( n2278 , n1996 , n1893 );
and ( n2279 , n1962 , n1891 );
nor ( n2280 , n2278 , n2279 );
xnor ( n2281 , n2280 , n1901 );
and ( n2282 , n2035 , n2073 );
and ( n2283 , n2004 , n2071 );
nor ( n2284 , n2282 , n2283 );
xnor ( n2285 , n2284 , n2081 );
xor ( n2286 , n2281 , n2285 );
and ( n2287 , n2076 , n2091 );
and ( n2288 , n2024 , n2089 );
nor ( n2289 , n2287 , n2288 );
xnor ( n2290 , n2289 , n2099 );
xor ( n2291 , n2286 , n2290 );
and ( n2292 , n2277 , n2291 );
and ( n2293 , n2057 , n1972 );
and ( n2294 , n1942 , n1970 );
nor ( n2295 , n2293 , n2294 );
xnor ( n2296 , n2295 , n1980 );
and ( n2297 , n1896 , n1912 );
and ( n2298 , n1987 , n1910 );
nor ( n2299 , n2297 , n2298 );
xnor ( n2300 , n2299 , n1920 );
xor ( n2301 , n2296 , n2300 );
and ( n2302 , n2065 , n1926 );
xor ( n2303 , n2301 , n2302 );
and ( n2304 , n2291 , n2303 );
and ( n2305 , n2277 , n2303 );
or ( n2306 , n2292 , n2304 , n2305 );
xor ( n2307 , n2273 , n2306 );
and ( n2308 , n2296 , n2300 );
and ( n2309 , n2300 , n2302 );
and ( n2310 , n2296 , n2302 );
or ( n2311 , n2308 , n2309 , n2310 );
and ( n2312 , n2243 , n2247 );
and ( n2313 , n2247 , n2252 );
and ( n2314 , n2243 , n2252 );
or ( n2315 , n2312 , n2313 , n2314 );
xor ( n2316 , n2311 , n2315 );
and ( n2317 , n2049 , n1993 );
and ( n2318 , n2057 , n1991 );
nor ( n2319 , n2317 , n2318 );
xnor ( n2320 , n2319 , n2001 );
and ( n2321 , n1883 , n2012 );
and ( n2322 , n1896 , n2010 );
nor ( n2323 , n2321 , n2322 );
xnor ( n2324 , n2323 , n2020 );
xor ( n2325 , n2320 , n2324 );
and ( n2326 , n2076 , n1926 );
xor ( n2327 , n2325 , n2326 );
xor ( n2328 , n2316 , n2327 );
xor ( n2329 , n2307 , n2328 );
xor ( n2330 , n2257 , n2329 );
and ( n2331 , n2234 , n2238 );
and ( n2332 , n2238 , n2253 );
and ( n2333 , n2234 , n2253 );
or ( n2334 , n2331 , n2332 , n2333 );
and ( n2335 , n2202 , n2213 );
and ( n2336 , n2213 , n2225 );
and ( n2337 , n2202 , n2225 );
or ( n2338 , n2335 , n2336 , n2337 );
xor ( n2339 , n2261 , n2265 );
xor ( n2340 , n2339 , n2270 );
and ( n2341 , n2338 , n2340 );
xor ( n2342 , n2277 , n2291 );
xor ( n2343 , n2342 , n2303 );
and ( n2344 , n2340 , n2343 );
and ( n2345 , n2338 , n2343 );
or ( n2346 , n2341 , n2344 , n2345 );
xor ( n2347 , n2334 , n2346 );
not ( n2348 , n2062 );
and ( n2349 , n1942 , n1972 );
and ( n2350 , n1953 , n1970 );
nor ( n2351 , n2349 , n2350 );
xnor ( n2352 , n2351 , n1980 );
xor ( n2353 , n2348 , n2352 );
and ( n2354 , n1962 , n1893 );
and ( n2355 , n1975 , n1891 );
nor ( n2356 , n2354 , n2355 );
xnor ( n2357 , n2356 , n1901 );
xor ( n2358 , n2353 , n2357 );
and ( n2359 , n1987 , n1912 );
and ( n2360 , n1996 , n1910 );
nor ( n2361 , n2359 , n2360 );
xnor ( n2362 , n2361 , n1920 );
and ( n2363 , n2004 , n2073 );
and ( n2364 , n2015 , n2071 );
nor ( n2365 , n2363 , n2364 );
xnor ( n2366 , n2365 , n2081 );
xor ( n2367 , n2362 , n2366 );
and ( n2368 , n2024 , n2091 );
and ( n2369 , n2035 , n2089 );
nor ( n2370 , n2368 , n2369 );
xnor ( n2371 , n2370 , n2099 );
xor ( n2372 , n2367 , n2371 );
xor ( n2373 , n2358 , n2372 );
and ( n2374 , n2281 , n2285 );
and ( n2375 , n2285 , n2290 );
and ( n2376 , n2281 , n2290 );
or ( n2377 , n2374 , n2375 , n2376 );
buf ( n2378 , n2269 );
xor ( n2379 , n2377 , n2378 );
and ( n2380 , n1904 , n2032 );
and ( n2381 , n1915 , n2030 );
nor ( n2382 , n2380 , n2381 );
xnor ( n2383 , n2382 , n2040 );
xor ( n2384 , n2379 , n2383 );
xor ( n2385 , n2373 , n2384 );
xor ( n2386 , n2347 , n2385 );
xor ( n2387 , n2330 , n2386 );
xor ( n2388 , n1932 , n1934 );
xor ( n2389 , n1934 , n1936 );
not ( n2390 , n2389 );
and ( n2391 , n2388 , n2390 );
and ( n2392 , n1953 , n2391 );
not ( n2393 , n2392 );
xnor ( n2394 , n2393 , n1939 );
and ( n2395 , n1975 , n2054 );
and ( n2396 , n2049 , n2052 );
nor ( n2397 , n2395 , n2396 );
xnor ( n2398 , n2397 , n2062 );
and ( n2399 , n2394 , n2398 );
buf ( n529659 , n1143 );
buf ( n2401 , n529659 );
and ( n2402 , n2401 , n1926 );
and ( n2403 , n2398 , n2402 );
and ( n2404 , n2394 , n2402 );
or ( n2405 , n2399 , n2403 , n2404 );
and ( n2406 , n1996 , n1972 );
and ( n2407 , n1962 , n1970 );
nor ( n2408 , n2406 , n2407 );
xnor ( n2409 , n2408 , n1980 );
and ( n2410 , n2035 , n2012 );
and ( n2411 , n2004 , n2010 );
nor ( n2412 , n2410 , n2411 );
xnor ( n2413 , n2412 , n2020 );
and ( n2414 , n2409 , n2413 );
and ( n2415 , n2076 , n2032 );
and ( n2416 , n2024 , n2030 );
nor ( n2417 , n2415 , n2416 );
xnor ( n2418 , n2417 , n2040 );
and ( n2419 , n2413 , n2418 );
and ( n2420 , n2409 , n2418 );
or ( n2421 , n2414 , n2419 , n2420 );
and ( n2422 , n2405 , n2421 );
and ( n2423 , n2057 , n1950 );
and ( n2424 , n1942 , n1948 );
nor ( n2425 , n2423 , n2424 );
xnor ( n2426 , n2425 , n1958 );
buf ( n2427 , n2426 );
and ( n2428 , n2421 , n2427 );
and ( n2429 , n2405 , n2427 );
or ( n2430 , n2422 , n2428 , n2429 );
xor ( n2431 , n1930 , n1984 );
xor ( n2432 , n2431 , n2044 );
and ( n2433 , n2430 , n2432 );
xor ( n2434 , n2103 , n2108 );
xor ( n2435 , n2434 , n2113 );
and ( n2436 , n2432 , n2435 );
and ( n2437 , n2430 , n2435 );
or ( n2438 , n2433 , n2436 , n2437 );
xor ( n2439 , n2047 , n2116 );
xor ( n2440 , n2439 , n2128 );
and ( n2441 , n2438 , n2440 );
xor ( n2442 , n2173 , n2187 );
xor ( n2443 , n2442 , n2226 );
and ( n2444 , n2440 , n2443 );
and ( n2445 , n2438 , n2443 );
or ( n2446 , n2441 , n2444 , n2445 );
xor ( n2447 , n2338 , n2340 );
xor ( n2448 , n2447 , n2343 );
and ( n2449 , n2446 , n2448 );
xor ( n2450 , n2131 , n2229 );
xor ( n2451 , n2450 , n2254 );
and ( n2452 , n2448 , n2451 );
and ( n2453 , n2446 , n2451 );
or ( n2454 , n2449 , n2452 , n2453 );
xor ( n2455 , n2387 , n2454 );
xor ( n2456 , n2446 , n2448 );
xor ( n2457 , n2456 , n2451 );
and ( n2458 , n1896 , n1993 );
and ( n2459 , n1987 , n1991 );
nor ( n2460 , n2458 , n2459 );
xnor ( n2461 , n2460 , n2001 );
and ( n2462 , n2094 , n2073 );
and ( n2463 , n2065 , n2071 );
nor ( n2464 , n2462 , n2463 );
xnor ( n2465 , n2464 , n2081 );
and ( n2466 , n2461 , n2465 );
and ( n2467 , n1924 , n2091 );
and ( n2468 , n2085 , n2089 );
nor ( n2469 , n2467 , n2468 );
xnor ( n2470 , n2469 , n2099 );
and ( n2471 , n2465 , n2470 );
and ( n2472 , n2461 , n2470 );
or ( n2473 , n2466 , n2471 , n2472 );
xor ( n2474 , n2063 , n2082 );
xor ( n2475 , n2474 , n2100 );
and ( n2476 , n2473 , n2475 );
xor ( n2477 , n1902 , n1921 );
xor ( n2478 , n2477 , n1927 );
and ( n2479 , n2475 , n2478 );
and ( n2480 , n2473 , n2478 );
or ( n2481 , n2476 , n2479 , n2480 );
not ( n2482 , n2426 );
and ( n2483 , n1915 , n1893 );
and ( n2484 , n1883 , n1891 );
nor ( n2485 , n2483 , n2484 );
xnor ( n2486 , n2485 , n1901 );
and ( n2487 , n2482 , n2486 );
and ( n2488 , n2015 , n1912 );
and ( n2489 , n1904 , n1910 );
nor ( n2490 , n2488 , n2489 );
xnor ( n2491 , n2490 , n1920 );
and ( n2492 , n2486 , n2491 );
and ( n2493 , n2482 , n2491 );
or ( n2494 , n2487 , n2492 , n2493 );
xor ( n2495 , n1940 , n1959 );
xor ( n2496 , n2495 , n1981 );
and ( n2497 , n2494 , n2496 );
xor ( n2498 , n2002 , n2021 );
xor ( n2499 , n2498 , n2041 );
and ( n2500 , n2496 , n2499 );
and ( n2501 , n2494 , n2499 );
or ( n2502 , n2497 , n2500 , n2501 );
and ( n2503 , n2481 , n2502 );
xor ( n2504 , n2144 , n2155 );
xor ( n2505 , n2504 , n2170 );
and ( n2506 , n2502 , n2505 );
and ( n2507 , n2481 , n2505 );
or ( n2508 , n2503 , n2506 , n2507 );
buf ( n529768 , n1177 );
buf ( n2510 , n529768 );
buf ( n529770 , n1178 );
buf ( n2512 , n529770 );
and ( n2513 , n2510 , n2512 );
not ( n2514 , n2513 );
and ( n2515 , n1936 , n2514 );
not ( n2516 , n2515 );
and ( n2517 , n1942 , n2391 );
and ( n2518 , n1953 , n2389 );
nor ( n2519 , n2517 , n2518 );
xnor ( n2520 , n2519 , n1939 );
and ( n2521 , n2516 , n2520 );
and ( n2522 , n1962 , n2054 );
and ( n2523 , n1975 , n2052 );
nor ( n2524 , n2522 , n2523 );
xnor ( n2525 , n2524 , n2062 );
and ( n2526 , n2520 , n2525 );
and ( n2527 , n2516 , n2525 );
or ( n2528 , n2521 , n2526 , n2527 );
and ( n2529 , n2049 , n1950 );
and ( n2530 , n2057 , n1948 );
nor ( n2531 , n2529 , n2530 );
xnor ( n2532 , n2531 , n1958 );
and ( n2533 , n2065 , n2032 );
and ( n2534 , n2076 , n2030 );
nor ( n2535 , n2533 , n2534 );
xnor ( n2536 , n2535 , n2040 );
and ( n2537 , n2532 , n2536 );
and ( n2538 , n2085 , n2073 );
and ( n2539 , n2094 , n2071 );
nor ( n2540 , n2538 , n2539 );
xnor ( n2541 , n2540 , n2081 );
and ( n2542 , n2536 , n2541 );
and ( n2543 , n2532 , n2541 );
or ( n2544 , n2537 , n2542 , n2543 );
and ( n2545 , n2528 , n2544 );
and ( n2546 , n1883 , n1993 );
and ( n2547 , n1896 , n1991 );
nor ( n2548 , n2546 , n2547 );
xnor ( n2549 , n2548 , n2001 );
and ( n2550 , n2401 , n2091 );
and ( n2551 , n1924 , n2089 );
nor ( n2552 , n2550 , n2551 );
xnor ( n2553 , n2552 , n2099 );
and ( n2554 , n2549 , n2553 );
buf ( n529814 , n1144 );
buf ( n2556 , n529814 );
and ( n2557 , n2556 , n1926 );
and ( n2558 , n2553 , n2557 );
and ( n2559 , n2549 , n2557 );
or ( n2560 , n2554 , n2558 , n2559 );
and ( n2561 , n2544 , n2560 );
and ( n2562 , n2528 , n2560 );
or ( n2563 , n2545 , n2561 , n2562 );
and ( n2564 , n1987 , n1972 );
and ( n2565 , n1996 , n1970 );
nor ( n2566 , n2564 , n2565 );
xnor ( n2567 , n2566 , n1980 );
and ( n2568 , n2004 , n1912 );
and ( n2569 , n2015 , n1910 );
nor ( n2570 , n2568 , n2569 );
xnor ( n2571 , n2570 , n1920 );
and ( n2572 , n2567 , n2571 );
and ( n2573 , n2024 , n2012 );
and ( n2574 , n2035 , n2010 );
nor ( n2575 , n2573 , n2574 );
xnor ( n2576 , n2575 , n2020 );
and ( n2577 , n2571 , n2576 );
and ( n2578 , n2567 , n2576 );
or ( n2579 , n2572 , n2577 , n2578 );
xor ( n2580 , n2394 , n2398 );
xor ( n2581 , n2580 , n2402 );
and ( n2582 , n2579 , n2581 );
xor ( n2583 , n2409 , n2413 );
xor ( n2584 , n2583 , n2418 );
and ( n2585 , n2581 , n2584 );
and ( n2586 , n2579 , n2584 );
or ( n2587 , n2582 , n2585 , n2586 );
and ( n2588 , n2563 , n2587 );
xor ( n2589 , n2405 , n2421 );
xor ( n2590 , n2589 , n2427 );
and ( n2591 , n2587 , n2590 );
and ( n2592 , n2563 , n2590 );
or ( n2593 , n2588 , n2591 , n2592 );
and ( n2594 , n1996 , n2054 );
and ( n2595 , n1962 , n2052 );
nor ( n2596 , n2594 , n2595 );
xnor ( n2597 , n2596 , n2062 );
and ( n2598 , n2035 , n1912 );
and ( n2599 , n2004 , n1910 );
nor ( n2600 , n2598 , n2599 );
xnor ( n2601 , n2600 , n1920 );
and ( n2602 , n2597 , n2601 );
and ( n2603 , n2076 , n2012 );
and ( n529863 , n2024 , n2010 );
nor ( n2604 , n2603 , n529863 );
xnor ( n2605 , n2604 , n2020 );
and ( n2606 , n2601 , n2605 );
and ( n2607 , n2597 , n2605 );
or ( n2608 , n2602 , n2606 , n2607 );
xor ( n2609 , n1936 , n2510 );
xor ( n2610 , n2510 , n2512 );
not ( n2611 , n2610 );
and ( n2612 , n2609 , n2611 );
and ( n2613 , n1953 , n2612 );
not ( n2614 , n2613 );
xnor ( n2615 , n2614 , n2515 );
and ( n2616 , n1915 , n1993 );
and ( n2617 , n1883 , n1991 );
nor ( n2618 , n2616 , n2617 );
xnor ( n2619 , n2618 , n2001 );
and ( n2620 , n2615 , n2619 );
and ( n2621 , n2556 , n2091 );
and ( n2622 , n2401 , n2089 );
nor ( n2623 , n2621 , n2622 );
xnor ( n2624 , n2623 , n2099 );
and ( n2625 , n2619 , n2624 );
and ( n2626 , n2615 , n2624 );
or ( n2627 , n2620 , n2625 , n2626 );
and ( n2628 , n2608 , n2627 );
and ( n2629 , n1975 , n1950 );
and ( n2630 , n2049 , n1948 );
nor ( n2631 , n2629 , n2630 );
xnor ( n2632 , n2631 , n1958 );
and ( n2633 , n2015 , n1893 );
and ( n2634 , n1904 , n1891 );
nor ( n2635 , n2633 , n2634 );
xnor ( n2636 , n2635 , n1901 );
and ( n2637 , n2632 , n2636 );
buf ( n529898 , n1145 );
buf ( n2639 , n529898 );
and ( n2640 , n2639 , n1926 );
and ( n2641 , n2636 , n2640 );
and ( n2642 , n2632 , n2640 );
or ( n2643 , n2637 , n2641 , n2642 );
and ( n2644 , n2627 , n2643 );
and ( n2645 , n2608 , n2643 );
or ( n2646 , n2628 , n2644 , n2645 );
xor ( n2647 , n2461 , n2465 );
xor ( n2648 , n2647 , n2470 );
and ( n2649 , n2646 , n2648 );
xor ( n2650 , n2482 , n2486 );
xor ( n2651 , n2650 , n2491 );
and ( n2652 , n2648 , n2651 );
and ( n2653 , n2646 , n2651 );
or ( n2654 , n2649 , n2652 , n2653 );
xor ( n2655 , n2473 , n2475 );
xor ( n2656 , n2655 , n2478 );
and ( n2657 , n2654 , n2656 );
xor ( n2658 , n2494 , n2496 );
xor ( n2659 , n2658 , n2499 );
and ( n2660 , n2656 , n2659 );
and ( n2661 , n2654 , n2659 );
or ( n2662 , n2657 , n2660 , n2661 );
and ( n2663 , n2593 , n2662 );
xor ( n2664 , n2430 , n2432 );
xor ( n2665 , n2664 , n2435 );
and ( n2666 , n2662 , n2665 );
and ( n2667 , n2593 , n2665 );
or ( n2668 , n2663 , n2666 , n2667 );
and ( n2669 , n2508 , n2668 );
xor ( n2670 , n2438 , n2440 );
xor ( n2671 , n2670 , n2443 );
and ( n2672 , n2668 , n2671 );
and ( n2673 , n2508 , n2671 );
or ( n2674 , n2669 , n2672 , n2673 );
and ( n2675 , n2457 , n2674 );
xor ( n2676 , n2457 , n2674 );
xor ( n2677 , n2508 , n2668 );
xor ( n2678 , n2677 , n2671 );
and ( n2679 , n1896 , n1972 );
and ( n2680 , n1987 , n1970 );
nor ( n2681 , n2679 , n2680 );
xnor ( n2682 , n2681 , n1980 );
and ( n2683 , n2094 , n2032 );
and ( n2684 , n2065 , n2030 );
nor ( n2685 , n2683 , n2684 );
xnor ( n2686 , n2685 , n2040 );
and ( n2687 , n2682 , n2686 );
and ( n2688 , n1924 , n2073 );
and ( n2689 , n2085 , n2071 );
nor ( n2690 , n2688 , n2689 );
xnor ( n2691 , n2690 , n2081 );
and ( n2692 , n2686 , n2691 );
and ( n2693 , n2682 , n2691 );
or ( n2694 , n2687 , n2692 , n2693 );
and ( n2695 , n2057 , n2391 );
and ( n2696 , n1942 , n2389 );
nor ( n2697 , n2695 , n2696 );
xnor ( n2698 , n2697 , n1939 );
buf ( n2699 , n2698 );
and ( n2700 , n2694 , n2699 );
and ( n2701 , n1904 , n1893 );
and ( n2702 , n1915 , n1891 );
nor ( n2703 , n2701 , n2702 );
xnor ( n2704 , n2703 , n1901 );
and ( n2705 , n2699 , n2704 );
and ( n2706 , n2694 , n2704 );
or ( n2707 , n2700 , n2705 , n2706 );
xor ( n2708 , n2516 , n2520 );
xor ( n2709 , n2708 , n2525 );
xor ( n2710 , n2532 , n2536 );
xor ( n2711 , n2710 , n2541 );
and ( n2712 , n2709 , n2711 );
xor ( n2713 , n2567 , n2571 );
xor ( n2714 , n2713 , n2576 );
and ( n2715 , n2711 , n2714 );
and ( n2716 , n2709 , n2714 );
or ( n2717 , n2712 , n2715 , n2716 );
and ( n2718 , n2707 , n2717 );
xor ( n2719 , n2528 , n2544 );
xor ( n529980 , n2719 , n2560 );
and ( n2721 , n2717 , n529980 );
and ( n529982 , n2707 , n529980 );
or ( n2723 , n2718 , n2721 , n529982 );
and ( n2724 , n1987 , n2054 );
and ( n2725 , n1996 , n2052 );
nor ( n2726 , n2724 , n2725 );
xnor ( n2727 , n2726 , n2062 );
and ( n2728 , n2004 , n1893 );
and ( n2729 , n2015 , n1891 );
nor ( n2730 , n2728 , n2729 );
xnor ( n2731 , n2730 , n1901 );
and ( n2732 , n2727 , n2731 );
and ( n2733 , n2024 , n1912 );
and ( n2734 , n2035 , n1910 );
nor ( n2735 , n2733 , n2734 );
xnor ( n2736 , n2735 , n1920 );
and ( n2737 , n2731 , n2736 );
and ( n2738 , n2727 , n2736 );
or ( n2739 , n2732 , n2737 , n2738 );
and ( n2740 , n2049 , n2391 );
and ( n2741 , n2057 , n2389 );
nor ( n2742 , n2740 , n2741 );
xnor ( n2743 , n2742 , n1939 );
and ( n2744 , n2065 , n2012 );
and ( n2745 , n2076 , n2010 );
nor ( n2746 , n2744 , n2745 );
xnor ( n2747 , n2746 , n2020 );
and ( n2748 , n2743 , n2747 );
and ( n2749 , n2085 , n2032 );
and ( n2750 , n2094 , n2030 );
nor ( n2751 , n2749 , n2750 );
xnor ( n2752 , n2751 , n2040 );
and ( n2753 , n2747 , n2752 );
and ( n2754 , n2743 , n2752 );
or ( n2755 , n2748 , n2753 , n2754 );
and ( n2756 , n2739 , n2755 );
not ( n2757 , n2698 );
and ( n2758 , n2755 , n2757 );
and ( n2759 , n2739 , n2757 );
or ( n2760 , n2756 , n2758 , n2759 );
xor ( n2761 , n2549 , n2553 );
xor ( n2762 , n2761 , n2557 );
and ( n2763 , n2760 , n2762 );
xor ( n2764 , n2694 , n2699 );
xor ( n2765 , n2764 , n2704 );
and ( n2766 , n2762 , n2765 );
and ( n2767 , n2760 , n2765 );
or ( n2768 , n2763 , n2766 , n2767 );
xor ( n2769 , n2579 , n2581 );
xor ( n2770 , n2769 , n2584 );
and ( n2771 , n2768 , n2770 );
xor ( n2772 , n2646 , n2648 );
xor ( n2773 , n2772 , n2651 );
and ( n2774 , n2770 , n2773 );
and ( n2775 , n2768 , n2773 );
or ( n2776 , n2771 , n2774 , n2775 );
and ( n2777 , n2723 , n2776 );
xor ( n2778 , n2563 , n2587 );
xor ( n2779 , n2778 , n2590 );
and ( n2780 , n2776 , n2779 );
and ( n2781 , n2723 , n2779 );
or ( n2782 , n2777 , n2780 , n2781 );
xor ( n2783 , n2481 , n2502 );
xor ( n2784 , n2783 , n2505 );
and ( n2785 , n2782 , n2784 );
xor ( n2786 , n2593 , n2662 );
xor ( n2787 , n2786 , n2665 );
and ( n2788 , n2784 , n2787 );
and ( n2789 , n2782 , n2787 );
or ( n2790 , n2785 , n2788 , n2789 );
and ( n2791 , n2678 , n2790 );
xor ( n2792 , n2678 , n2790 );
xor ( n2793 , n2782 , n2784 );
xor ( n2794 , n2793 , n2787 );
xor ( n2795 , n2597 , n2601 );
xor ( n2796 , n2795 , n2605 );
xor ( n2797 , n2615 , n2619 );
xor ( n2798 , n2797 , n2624 );
and ( n2799 , n2796 , n2798 );
xor ( n2800 , n2682 , n2686 );
xor ( n2801 , n2800 , n2691 );
and ( n2802 , n2798 , n2801 );
and ( n2803 , n2796 , n2801 );
or ( n2804 , n2799 , n2802 , n2803 );
buf ( n530065 , n1179 );
buf ( n2806 , n530065 );
buf ( n530067 , n1180 );
buf ( n2808 , n530067 );
and ( n2809 , n2806 , n2808 );
not ( n2810 , n2809 );
and ( n2811 , n2512 , n2810 );
not ( n2812 , n2811 );
and ( n2813 , n1942 , n2612 );
and ( n2814 , n1953 , n2610 );
nor ( n2815 , n2813 , n2814 );
xnor ( n2816 , n2815 , n2515 );
and ( n2817 , n2812 , n2816 );
and ( n2818 , n1962 , n1950 );
and ( n2819 , n1975 , n1948 );
nor ( n2820 , n2818 , n2819 );
xnor ( n2821 , n2820 , n1958 );
and ( n2822 , n2816 , n2821 );
and ( n2823 , n2812 , n2821 );
or ( n2824 , n2817 , n2822 , n2823 );
and ( n2825 , n1883 , n1972 );
and ( n2826 , n1896 , n1970 );
nor ( n2827 , n2825 , n2826 );
xnor ( n2828 , n2827 , n1980 );
and ( n2829 , n2401 , n2073 );
and ( n2830 , n1924 , n2071 );
nor ( n2831 , n2829 , n2830 );
xnor ( n2832 , n2831 , n2081 );
and ( n2833 , n2828 , n2832 );
and ( n2834 , n2639 , n2091 );
and ( n2835 , n2556 , n2089 );
nor ( n2836 , n2834 , n2835 );
xnor ( n2837 , n2836 , n2099 );
and ( n2838 , n2832 , n2837 );
and ( n2839 , n2828 , n2837 );
or ( n2840 , n2833 , n2838 , n2839 );
and ( n2841 , n2824 , n2840 );
xor ( n2842 , n2632 , n2636 );
xor ( n2843 , n2842 , n2640 );
and ( n2844 , n2840 , n2843 );
and ( n2845 , n2824 , n2843 );
or ( n2846 , n2841 , n2844 , n2845 );
and ( n2847 , n2804 , n2846 );
xor ( n2848 , n2608 , n2627 );
xor ( n2849 , n2848 , n2643 );
and ( n2850 , n2846 , n2849 );
and ( n2851 , n2804 , n2849 );
or ( n2852 , n2847 , n2850 , n2851 );
and ( n2853 , n1996 , n1950 );
and ( n2854 , n1962 , n1948 );
nor ( n2855 , n2853 , n2854 );
xnor ( n2856 , n2855 , n1958 );
and ( n530117 , n2035 , n1893 );
and ( n2858 , n2004 , n1891 );
nor ( n530119 , n530117 , n2858 );
xnor ( n2860 , n530119 , n1901 );
and ( n2861 , n2856 , n2860 );
and ( n2862 , n2076 , n1912 );
and ( n2863 , n2024 , n1910 );
nor ( n2864 , n2862 , n2863 );
xnor ( n2865 , n2864 , n1920 );
and ( n2866 , n2860 , n2865 );
and ( n2867 , n2856 , n2865 );
or ( n2868 , n2861 , n2866 , n2867 );
xor ( n2869 , n2512 , n2806 );
xor ( n2870 , n2806 , n2808 );
not ( n2871 , n2870 );
and ( n2872 , n2869 , n2871 );
and ( n2873 , n1953 , n2872 );
not ( n2874 , n2873 );
xnor ( n2875 , n2874 , n2811 );
and ( n2876 , n1915 , n1972 );
and ( n2877 , n1883 , n1970 );
nor ( n2878 , n2876 , n2877 );
xnor ( n2879 , n2878 , n1980 );
and ( n2880 , n2875 , n2879 );
and ( n2881 , n2556 , n2073 );
and ( n2882 , n2401 , n2071 );
nor ( n2883 , n2881 , n2882 );
xnor ( n2884 , n2883 , n2081 );
and ( n530145 , n2879 , n2884 );
and ( n2886 , n2875 , n2884 );
or ( n2887 , n2880 , n530145 , n2886 );
and ( n2888 , n2868 , n2887 );
and ( n2889 , n1896 , n2054 );
and ( n2890 , n1987 , n2052 );
nor ( n2891 , n2889 , n2890 );
xnor ( n2892 , n2891 , n2062 );
and ( n2893 , n2094 , n2012 );
and ( n2894 , n2065 , n2010 );
nor ( n2895 , n2893 , n2894 );
xnor ( n2896 , n2895 , n2020 );
and ( n2897 , n2892 , n2896 );
and ( n2898 , n1924 , n2032 );
and ( n2899 , n2085 , n2030 );
nor ( n2900 , n2898 , n2899 );
xnor ( n2901 , n2900 , n2040 );
and ( n2902 , n2896 , n2901 );
and ( n2903 , n2892 , n2901 );
or ( n2904 , n2897 , n2902 , n2903 );
and ( n2905 , n2887 , n2904 );
and ( n2906 , n2868 , n2904 );
or ( n2907 , n2888 , n2905 , n2906 );
and ( n2908 , n2057 , n2612 );
and ( n2909 , n1942 , n2610 );
nor ( n2910 , n2908 , n2909 );
xnor ( n2911 , n2910 , n2515 );
buf ( n2912 , n2911 );
and ( n2913 , n1904 , n1993 );
and ( n2914 , n1915 , n1991 );
nor ( n2915 , n2913 , n2914 );
xnor ( n2916 , n2915 , n2001 );
and ( n2917 , n2912 , n2916 );
buf ( n530178 , n1146 );
buf ( n2919 , n530178 );
and ( n2920 , n2919 , n1926 );
and ( n2921 , n2916 , n2920 );
and ( n2922 , n2912 , n2920 );
or ( n2923 , n2917 , n2921 , n2922 );
and ( n2924 , n2907 , n2923 );
xor ( n2925 , n2739 , n2755 );
xor ( n2926 , n2925 , n2757 );
and ( n2927 , n2923 , n2926 );
and ( n2928 , n2907 , n2926 );
or ( n2929 , n2924 , n2927 , n2928 );
xor ( n2930 , n2709 , n2711 );
xor ( n2931 , n2930 , n2714 );
and ( n2932 , n2929 , n2931 );
xor ( n2933 , n2760 , n2762 );
xor ( n2934 , n2933 , n2765 );
and ( n2935 , n2931 , n2934 );
and ( n2936 , n2929 , n2934 );
or ( n2937 , n2932 , n2935 , n2936 );
and ( n2938 , n2852 , n2937 );
xor ( n2939 , n2707 , n2717 );
xor ( n2940 , n2939 , n529980 );
and ( n2941 , n2937 , n2940 );
and ( n2942 , n2852 , n2940 );
or ( n2943 , n2938 , n2941 , n2942 );
xor ( n2944 , n2654 , n2656 );
xor ( n2945 , n2944 , n2659 );
and ( n2946 , n2943 , n2945 );
xor ( n2947 , n2723 , n2776 );
xor ( n2948 , n2947 , n2779 );
and ( n2949 , n2945 , n2948 );
and ( n2950 , n2943 , n2948 );
or ( n2951 , n2946 , n2949 , n2950 );
and ( n2952 , n2794 , n2951 );
xor ( n2953 , n2794 , n2951 );
xor ( n2954 , n2943 , n2945 );
xor ( n2955 , n2954 , n2948 );
and ( n2956 , n1987 , n1950 );
and ( n2957 , n1996 , n1948 );
nor ( n2958 , n2956 , n2957 );
xnor ( n2959 , n2958 , n1958 );
and ( n2960 , n2004 , n1993 );
and ( n2961 , n2015 , n1991 );
nor ( n2962 , n2960 , n2961 );
xnor ( n2963 , n2962 , n2001 );
and ( n2964 , n2959 , n2963 );
and ( n2965 , n2024 , n1893 );
and ( n2966 , n2035 , n1891 );
nor ( n2967 , n2965 , n2966 );
xnor ( n2968 , n2967 , n1901 );
and ( n2969 , n2963 , n2968 );
and ( n2970 , n2959 , n2968 );
or ( n2971 , n2964 , n2969 , n2970 );
buf ( n530232 , n1181 );
buf ( n2973 , n530232 );
buf ( n530234 , n1182 );
buf ( n2975 , n530234 );
and ( n2976 , n2973 , n2975 );
not ( n2977 , n2976 );
and ( n2978 , n2808 , n2977 );
not ( n2979 , n2978 );
and ( n2980 , n1942 , n2872 );
and ( n2981 , n1953 , n2870 );
nor ( n2982 , n2980 , n2981 );
xnor ( n2983 , n2982 , n2811 );
and ( n2984 , n2979 , n2983 );
and ( n2985 , n1962 , n2391 );
and ( n2986 , n1975 , n2389 );
nor ( n2987 , n2985 , n2986 );
xnor ( n2988 , n2987 , n1939 );
and ( n2989 , n2983 , n2988 );
and ( n2990 , n2979 , n2988 );
or ( n2991 , n2984 , n2989 , n2990 );
and ( n2992 , n2971 , n2991 );
and ( n2993 , n2049 , n2612 );
and ( n2994 , n2057 , n2610 );
nor ( n2995 , n2993 , n2994 );
xnor ( n2996 , n2995 , n2515 );
and ( n2997 , n2065 , n1912 );
and ( n2998 , n2076 , n1910 );
nor ( n2999 , n2997 , n2998 );
xnor ( n3000 , n2999 , n1920 );
and ( n3001 , n2996 , n3000 );
and ( n3002 , n2085 , n2012 );
and ( n3003 , n2094 , n2010 );
nor ( n3004 , n3002 , n3003 );
xnor ( n3005 , n3004 , n2020 );
and ( n3006 , n3000 , n3005 );
and ( n3007 , n2996 , n3005 );
or ( n3008 , n3001 , n3006 , n3007 );
and ( n3009 , n2991 , n3008 );
and ( n3010 , n2971 , n3008 );
or ( n3011 , n2992 , n3009 , n3010 );
and ( n3012 , n1883 , n2054 );
and ( n3013 , n1896 , n2052 );
nor ( n3014 , n3012 , n3013 );
xnor ( n3015 , n3014 , n2062 );
and ( n3016 , n2401 , n2032 );
and ( n3017 , n1924 , n2030 );
nor ( n3018 , n3016 , n3017 );
xnor ( n3019 , n3018 , n2040 );
and ( n3020 , n3015 , n3019 );
and ( n3021 , n2639 , n2073 );
and ( n3022 , n2556 , n2071 );
nor ( n3023 , n3021 , n3022 );
xnor ( n3024 , n3023 , n2081 );
and ( n3025 , n3019 , n3024 );
and ( n3026 , n3015 , n3024 );
or ( n3027 , n3020 , n3025 , n3026 );
not ( n3028 , n2911 );
and ( n3029 , n3027 , n3028 );
and ( n3030 , n2015 , n1993 );
and ( n3031 , n1904 , n1991 );
nor ( n3032 , n3030 , n3031 );
xnor ( n3033 , n3032 , n2001 );
and ( n3034 , n3028 , n3033 );
and ( n3035 , n3027 , n3033 );
or ( n3036 , n3029 , n3034 , n3035 );
and ( n3037 , n3011 , n3036 );
xor ( n3038 , n2868 , n2887 );
xor ( n3039 , n3038 , n2904 );
and ( n3040 , n3036 , n3039 );
and ( n3041 , n3011 , n3039 );
or ( n3042 , n3037 , n3040 , n3041 );
xor ( n3043 , n2796 , n2798 );
xor ( n3044 , n3043 , n2801 );
and ( n3045 , n3042 , n3044 );
xor ( n3046 , n2907 , n2923 );
xor ( n3047 , n3046 , n2926 );
and ( n3048 , n3044 , n3047 );
and ( n3049 , n3042 , n3047 );
or ( n3050 , n3045 , n3048 , n3049 );
and ( n3051 , n1975 , n2391 );
and ( n3052 , n2049 , n2389 );
nor ( n3053 , n3051 , n3052 );
xnor ( n3054 , n3053 , n1939 );
and ( n3055 , n2919 , n2091 );
and ( n3056 , n2639 , n2089 );
nor ( n3057 , n3055 , n3056 );
xnor ( n3058 , n3057 , n2099 );
and ( n3059 , n3054 , n3058 );
buf ( n530320 , n1147 );
buf ( n3061 , n530320 );
and ( n3062 , n3061 , n1926 );
and ( n3063 , n3058 , n3062 );
and ( n3064 , n3054 , n3062 );
or ( n3065 , n3059 , n3063 , n3064 );
xor ( n3066 , n2727 , n2731 );
xor ( n3067 , n3066 , n2736 );
and ( n3068 , n3065 , n3067 );
xor ( n3069 , n2812 , n2816 );
xor ( n3070 , n3069 , n2821 );
and ( n3071 , n3067 , n3070 );
and ( n3072 , n3065 , n3070 );
or ( n3073 , n3068 , n3071 , n3072 );
xor ( n3074 , n2828 , n2832 );
xor ( n3075 , n3074 , n2837 );
xor ( n3076 , n2743 , n2747 );
xor ( n3077 , n3076 , n2752 );
and ( n3078 , n3075 , n3077 );
xor ( n3079 , n2912 , n2916 );
xor ( n3080 , n3079 , n2920 );
and ( n3081 , n3077 , n3080 );
and ( n3082 , n3075 , n3080 );
or ( n3083 , n3078 , n3081 , n3082 );
and ( n3084 , n3073 , n3083 );
xor ( n3085 , n2824 , n2840 );
xor ( n3086 , n3085 , n2843 );
and ( n3087 , n3083 , n3086 );
and ( n3088 , n3073 , n3086 );
or ( n3089 , n3084 , n3087 , n3088 );
and ( n3090 , n3050 , n3089 );
xor ( n3091 , n2804 , n2846 );
xor ( n3092 , n3091 , n2849 );
and ( n3093 , n3089 , n3092 );
and ( n3094 , n3050 , n3092 );
or ( n3095 , n3090 , n3093 , n3094 );
xor ( n3096 , n2768 , n2770 );
xor ( n3097 , n3096 , n2773 );
and ( n3098 , n3095 , n3097 );
xor ( n3099 , n2852 , n2937 );
xor ( n3100 , n3099 , n2940 );
and ( n3101 , n3097 , n3100 );
and ( n3102 , n3095 , n3100 );
or ( n3103 , n3098 , n3101 , n3102 );
and ( n3104 , n2955 , n3103 );
xor ( n3105 , n2955 , n3103 );
xor ( n3106 , n3095 , n3097 );
xor ( n3107 , n3106 , n3100 );
xor ( n3108 , n2875 , n2879 );
xor ( n3109 , n3108 , n2884 );
xor ( n3110 , n2892 , n2896 );
xor ( n3111 , n3110 , n2901 );
and ( n3112 , n3109 , n3111 );
xor ( n3113 , n3027 , n3028 );
xor ( n3114 , n3113 , n3033 );
and ( n3115 , n3111 , n3114 );
and ( n3116 , n3109 , n3114 );
or ( n3117 , n3112 , n3115 , n3116 );
and ( n3118 , n2057 , n2872 );
and ( n3119 , n1942 , n2870 );
nor ( n3120 , n3118 , n3119 );
xnor ( n3121 , n3120 , n2811 );
and ( n3122 , n1996 , n2391 );
and ( n3123 , n1962 , n2389 );
nor ( n3124 , n3122 , n3123 );
xnor ( n3125 , n3124 , n1939 );
and ( n3126 , n3121 , n3125 );
and ( n3127 , n2035 , n1993 );
and ( n3128 , n2004 , n1991 );
nor ( n3129 , n3127 , n3128 );
xnor ( n3130 , n3129 , n2001 );
and ( n3131 , n3125 , n3130 );
and ( n3132 , n3121 , n3130 );
or ( n3133 , n3126 , n3131 , n3132 );
and ( n3134 , n1896 , n1950 );
and ( n3135 , n1987 , n1948 );
nor ( n3136 , n3134 , n3135 );
xnor ( n3137 , n3136 , n1958 );
and ( n3138 , n2076 , n1893 );
and ( n3139 , n2024 , n1891 );
nor ( n3140 , n3138 , n3139 );
xnor ( n3141 , n3140 , n1901 );
and ( n3142 , n3137 , n3141 );
and ( n3143 , n2094 , n1912 );
and ( n3144 , n2065 , n1910 );
nor ( n3145 , n3143 , n3144 );
xnor ( n3146 , n3145 , n1920 );
and ( n3147 , n3141 , n3146 );
and ( n3148 , n3137 , n3146 );
or ( n3149 , n3142 , n3147 , n3148 );
and ( n3150 , n3133 , n3149 );
xor ( n3151 , n2808 , n2973 );
xor ( n3152 , n2973 , n2975 );
not ( n3153 , n3152 );
and ( n3154 , n3151 , n3153 );
and ( n3155 , n1953 , n3154 );
not ( n3156 , n3155 );
xnor ( n3157 , n3156 , n2978 );
buf ( n3158 , n3157 );
and ( n3159 , n3149 , n3158 );
and ( n3160 , n3133 , n3158 );
or ( n3161 , n3150 , n3159 , n3160 );
and ( n3162 , n2015 , n1972 );
and ( n3163 , n1904 , n1970 );
nor ( n3164 , n3162 , n3163 );
xnor ( n3165 , n3164 , n1980 );
and ( n3166 , n2556 , n2032 );
and ( n3167 , n2401 , n2030 );
nor ( n3168 , n3166 , n3167 );
xnor ( n3169 , n3168 , n2040 );
and ( n3170 , n3165 , n3169 );
and ( n3171 , n2919 , n2073 );
and ( n3172 , n2639 , n2071 );
nor ( n3173 , n3171 , n3172 );
xnor ( n3174 , n3173 , n2081 );
and ( n3175 , n3169 , n3174 );
and ( n3176 , n3165 , n3174 );
or ( n3177 , n3170 , n3175 , n3176 );
and ( n3178 , n1975 , n2612 );
and ( n3179 , n2049 , n2610 );
nor ( n3180 , n3178 , n3179 );
xnor ( n3181 , n3180 , n2515 );
and ( n3182 , n1915 , n2054 );
and ( n3183 , n1883 , n2052 );
nor ( n3184 , n3182 , n3183 );
xnor ( n3185 , n3184 , n2062 );
and ( n3186 , n3181 , n3185 );
and ( n3187 , n1924 , n2012 );
and ( n3188 , n2085 , n2010 );
nor ( n3189 , n3187 , n3188 );
xnor ( n3190 , n3189 , n2020 );
and ( n3191 , n3185 , n3190 );
and ( n3192 , n3181 , n3190 );
or ( n3193 , n3186 , n3191 , n3192 );
and ( n3194 , n3177 , n3193 );
xor ( n3195 , n2959 , n2963 );
xor ( n3196 , n3195 , n2968 );
and ( n3197 , n3193 , n3196 );
and ( n3198 , n3177 , n3196 );
or ( n3199 , n3194 , n3197 , n3198 );
and ( n3200 , n3161 , n3199 );
xor ( n3201 , n2971 , n2991 );
xor ( n3202 , n3201 , n3008 );
and ( n3203 , n3199 , n3202 );
and ( n3204 , n3161 , n3202 );
or ( n3205 , n3200 , n3203 , n3204 );
and ( n3206 , n3117 , n3205 );
xor ( n3207 , n3011 , n3036 );
xor ( n3208 , n3207 , n3039 );
and ( n3209 , n3205 , n3208 );
and ( n3210 , n3117 , n3208 );
or ( n3211 , n3206 , n3209 , n3210 );
and ( n3212 , n1904 , n1972 );
and ( n3213 , n1915 , n1970 );
nor ( n3214 , n3212 , n3213 );
xnor ( n3215 , n3214 , n1980 );
and ( n3216 , n3061 , n2091 );
and ( n3217 , n2919 , n2089 );
nor ( n3218 , n3216 , n3217 );
xnor ( n3219 , n3218 , n2099 );
and ( n3220 , n3215 , n3219 );
buf ( n530481 , n1148 );
buf ( n3222 , n530481 );
and ( n3223 , n3222 , n1926 );
and ( n3224 , n3219 , n3223 );
and ( n3225 , n3215 , n3223 );
or ( n3226 , n3220 , n3224 , n3225 );
xor ( n3227 , n3054 , n3058 );
xor ( n3228 , n3227 , n3062 );
and ( n3229 , n3226 , n3228 );
xor ( n3230 , n2856 , n2860 );
xor ( n3231 , n3230 , n2865 );
and ( n3232 , n3228 , n3231 );
and ( n3233 , n3226 , n3231 );
or ( n3234 , n3229 , n3232 , n3233 );
xor ( n3235 , n3065 , n3067 );
xor ( n3236 , n3235 , n3070 );
and ( n3237 , n3234 , n3236 );
xor ( n3238 , n3075 , n3077 );
xor ( n3239 , n3238 , n3080 );
and ( n3240 , n3236 , n3239 );
and ( n3241 , n3234 , n3239 );
or ( n3242 , n3237 , n3240 , n3241 );
and ( n3243 , n3211 , n3242 );
xor ( n3244 , n3073 , n3083 );
xor ( n3245 , n3244 , n3086 );
and ( n3246 , n3242 , n3245 );
and ( n3247 , n3211 , n3245 );
or ( n3248 , n3243 , n3246 , n3247 );
xor ( n3249 , n2929 , n2931 );
xor ( n3250 , n3249 , n2934 );
and ( n3251 , n3248 , n3250 );
xor ( n3252 , n3050 , n3089 );
xor ( n3253 , n3252 , n3092 );
and ( n3254 , n3250 , n3253 );
and ( n3255 , n3248 , n3253 );
or ( n3256 , n3251 , n3254 , n3255 );
and ( n3257 , n3107 , n3256 );
xor ( n3258 , n3107 , n3256 );
xor ( n3259 , n3248 , n3250 );
xor ( n3260 , n3259 , n3253 );
xor ( n3261 , n3215 , n3219 );
xor ( n3262 , n3261 , n3223 );
xor ( n3263 , n2979 , n2983 );
xor ( n3264 , n3263 , n2988 );
and ( n3265 , n3262 , n3264 );
xor ( n3266 , n3015 , n3019 );
xor ( n3267 , n3266 , n3024 );
and ( n3268 , n3264 , n3267 );
and ( n3269 , n3262 , n3267 );
or ( n3270 , n3265 , n3268 , n3269 );
and ( n3271 , n2004 , n1972 );
and ( n3272 , n2015 , n1970 );
nor ( n3273 , n3271 , n3272 );
xnor ( n3274 , n3273 , n1980 );
and ( n3275 , n2024 , n1993 );
and ( n3276 , n2035 , n1991 );
nor ( n3277 , n3275 , n3276 );
xnor ( n3278 , n3277 , n2001 );
and ( n3279 , n3274 , n3278 );
buf ( n530540 , n1150 );
buf ( n3281 , n530540 );
and ( n3282 , n3281 , n1926 );
and ( n3283 , n3278 , n3282 );
and ( n3284 , n3274 , n3282 );
or ( n3285 , n3279 , n3283 , n3284 );
buf ( n530546 , n1183 );
buf ( n3287 , n530546 );
buf ( n530548 , n1184 );
buf ( n3289 , n530548 );
and ( n3290 , n3287 , n3289 );
not ( n3291 , n3290 );
and ( n3292 , n2975 , n3291 );
not ( n3293 , n3292 );
and ( n3294 , n1942 , n3154 );
and ( n3295 , n1953 , n3152 );
nor ( n3296 , n3294 , n3295 );
xnor ( n3297 , n3296 , n2978 );
and ( n3298 , n3293 , n3297 );
and ( n3299 , n1962 , n2612 );
and ( n3300 , n1975 , n2610 );
nor ( n3301 , n3299 , n3300 );
xnor ( n3302 , n3301 , n2515 );
and ( n3303 , n3297 , n3302 );
and ( n3304 , n3293 , n3302 );
or ( n3305 , n3298 , n3303 , n3304 );
and ( n3306 , n3285 , n3305 );
and ( n3307 , n1987 , n2391 );
and ( n3308 , n1996 , n2389 );
nor ( n3309 , n3307 , n3308 );
xnor ( n3310 , n3309 , n1939 );
and ( n3311 , n2065 , n1893 );
and ( n3312 , n2076 , n1891 );
nor ( n3313 , n3311 , n3312 );
xnor ( n3314 , n3313 , n1901 );
and ( n3315 , n3310 , n3314 );
and ( n3316 , n2085 , n1912 );
and ( n3317 , n2094 , n1910 );
nor ( n3318 , n3316 , n3317 );
xnor ( n3319 , n3318 , n1920 );
and ( n3320 , n3314 , n3319 );
and ( n3321 , n3310 , n3319 );
or ( n3322 , n3315 , n3320 , n3321 );
and ( n3323 , n3305 , n3322 );
and ( n3324 , n3285 , n3322 );
or ( n3325 , n3306 , n3323 , n3324 );
not ( n3326 , n3157 );
and ( n3327 , n3222 , n2091 );
and ( n3328 , n3061 , n2089 );
nor ( n3329 , n3327 , n3328 );
xnor ( n3330 , n3329 , n2099 );
and ( n3331 , n3326 , n3330 );
buf ( n530592 , n1149 );
buf ( n3333 , n530592 );
and ( n3334 , n3333 , n1926 );
and ( n3335 , n3330 , n3334 );
and ( n3336 , n3326 , n3334 );
or ( n3337 , n3331 , n3335 , n3336 );
and ( n3338 , n3325 , n3337 );
xor ( n3339 , n2996 , n3000 );
xor ( n3340 , n3339 , n3005 );
and ( n3341 , n3337 , n3340 );
and ( n3342 , n3325 , n3340 );
or ( n3343 , n3338 , n3341 , n3342 );
and ( n3344 , n3270 , n3343 );
xor ( n3345 , n3226 , n3228 );
xor ( n3346 , n3345 , n3231 );
and ( n3347 , n3343 , n3346 );
and ( n3348 , n3270 , n3346 );
or ( n3349 , n3344 , n3347 , n3348 );
xor ( n3350 , n3117 , n3205 );
xor ( n3351 , n3350 , n3208 );
and ( n3352 , n3349 , n3351 );
xor ( n3353 , n3234 , n3236 );
xor ( n3354 , n3353 , n3239 );
and ( n3355 , n3351 , n3354 );
and ( n3356 , n3349 , n3354 );
or ( n3357 , n3352 , n3355 , n3356 );
xor ( n3358 , n3042 , n3044 );
xor ( n3359 , n3358 , n3047 );
and ( n3360 , n3357 , n3359 );
xor ( n3361 , n3211 , n3242 );
xor ( n3362 , n3361 , n3245 );
and ( n3363 , n3359 , n3362 );
and ( n3364 , n3357 , n3362 );
or ( n3365 , n3360 , n3363 , n3364 );
and ( n3366 , n3260 , n3365 );
xor ( n3367 , n3260 , n3365 );
xor ( n3368 , n3357 , n3359 );
xor ( n3369 , n3368 , n3362 );
and ( n3370 , n1904 , n2054 );
and ( n3371 , n1915 , n2052 );
nor ( n3372 , n3370 , n3371 );
xnor ( n3373 , n3372 , n2062 );
and ( n3374 , n2639 , n2032 );
and ( n3375 , n2556 , n2030 );
nor ( n3376 , n3374 , n3375 );
xnor ( n3377 , n3376 , n2040 );
and ( n3378 , n3373 , n3377 );
and ( n3379 , n3061 , n2073 );
and ( n3380 , n2919 , n2071 );
nor ( n3381 , n3379 , n3380 );
xnor ( n3382 , n3381 , n2081 );
and ( n3383 , n3377 , n3382 );
and ( n3384 , n3373 , n3382 );
or ( n3385 , n3378 , n3383 , n3384 );
and ( n3386 , n2049 , n2872 );
and ( n3387 , n2057 , n2870 );
nor ( n3388 , n3386 , n3387 );
xnor ( n3389 , n3388 , n2811 );
and ( n3390 , n1883 , n1950 );
and ( n3391 , n1896 , n1948 );
nor ( n3392 , n3390 , n3391 );
xnor ( n3393 , n3392 , n1958 );
and ( n3394 , n3389 , n3393 );
and ( n3395 , n2401 , n2012 );
and ( n3396 , n1924 , n2010 );
nor ( n3397 , n3395 , n3396 );
xnor ( n3398 , n3397 , n2020 );
and ( n3399 , n3393 , n3398 );
and ( n3400 , n3389 , n3398 );
or ( n3401 , n3394 , n3399 , n3400 );
and ( n3402 , n3385 , n3401 );
xor ( n3403 , n3121 , n3125 );
xor ( n3404 , n3403 , n3130 );
and ( n3405 , n3401 , n3404 );
and ( n3406 , n3385 , n3404 );
or ( n3407 , n3402 , n3405 , n3406 );
xor ( n3408 , n3133 , n3149 );
xor ( n3409 , n3408 , n3158 );
and ( n3410 , n3407 , n3409 );
xor ( n3411 , n3177 , n3193 );
xor ( n3412 , n3411 , n3196 );
and ( n3413 , n3409 , n3412 );
and ( n3414 , n3407 , n3412 );
or ( n3415 , n3410 , n3413 , n3414 );
xor ( n3416 , n3109 , n3111 );
xor ( n3417 , n3416 , n3114 );
and ( n3418 , n3415 , n3417 );
xor ( n3419 , n3161 , n3199 );
xor ( n3420 , n3419 , n3202 );
and ( n3421 , n3417 , n3420 );
and ( n3422 , n3415 , n3420 );
or ( n3423 , n3418 , n3421 , n3422 );
xor ( n3424 , n3165 , n3169 );
xor ( n3425 , n3424 , n3174 );
xor ( n3426 , n3137 , n3141 );
xor ( n3427 , n3426 , n3146 );
and ( n3428 , n3425 , n3427 );
xor ( n3429 , n3181 , n3185 );
xor ( n3430 , n3429 , n3190 );
and ( n3431 , n3427 , n3430 );
and ( n3432 , n3425 , n3430 );
or ( n3433 , n3428 , n3431 , n3432 );
xor ( n3434 , n3262 , n3264 );
xor ( n3435 , n3434 , n3267 );
and ( n3436 , n3433 , n3435 );
xor ( n3437 , n3325 , n3337 );
xor ( n3438 , n3437 , n3340 );
and ( n3439 , n3435 , n3438 );
and ( n3440 , n3433 , n3438 );
or ( n3441 , n3436 , n3439 , n3440 );
xor ( n3442 , n3270 , n3343 );
xor ( n3443 , n3442 , n3346 );
and ( n3444 , n3441 , n3443 );
xor ( n3445 , n3415 , n3417 );
xor ( n3446 , n3445 , n3420 );
and ( n3447 , n3443 , n3446 );
and ( n3448 , n3441 , n3446 );
or ( n3449 , n3444 , n3447 , n3448 );
and ( n3450 , n3423 , n3449 );
xor ( n3451 , n3349 , n3351 );
xor ( n3452 , n3451 , n3354 );
and ( n3453 , n3449 , n3452 );
and ( n3454 , n3423 , n3452 );
or ( n3455 , n3450 , n3453 , n3454 );
and ( n3456 , n3369 , n3455 );
xor ( n3457 , n3369 , n3455 );
xor ( n3458 , n3423 , n3449 );
xor ( n3459 , n3458 , n3452 );
and ( n3460 , n1896 , n2391 );
and ( n3461 , n1987 , n2389 );
nor ( n3462 , n3460 , n3461 );
xnor ( n3463 , n3462 , n1939 );
and ( n3464 , n2035 , n1972 );
and ( n3465 , n2004 , n1970 );
nor ( n3466 , n3464 , n3465 );
xnor ( n3467 , n3466 , n1980 );
and ( n3468 , n3463 , n3467 );
and ( n3469 , n2076 , n1993 );
and ( n3470 , n2024 , n1991 );
nor ( n3471 , n3469 , n3470 );
xnor ( n3472 , n3471 , n2001 );
and ( n3473 , n3467 , n3472 );
and ( n3474 , n3463 , n3472 );
or ( n3475 , n3468 , n3473 , n3474 );
and ( n3476 , n1975 , n2872 );
and ( n3477 , n2049 , n2870 );
nor ( n3478 , n3476 , n3477 );
xnor ( n3479 , n3478 , n2811 );
and ( n3480 , n2094 , n1893 );
and ( n3481 , n2065 , n1891 );
nor ( n3482 , n3480 , n3481 );
xnor ( n3483 , n3482 , n1901 );
and ( n3484 , n3479 , n3483 );
and ( n3485 , n1924 , n1912 );
and ( n3486 , n2085 , n1910 );
nor ( n3487 , n3485 , n3486 );
xnor ( n3488 , n3487 , n1920 );
and ( n3489 , n3483 , n3488 );
and ( n3490 , n3479 , n3488 );
or ( n3491 , n3484 , n3489 , n3490 );
and ( n3492 , n3475 , n3491 );
and ( n3493 , n1915 , n1950 );
and ( n3494 , n1883 , n1948 );
nor ( n3495 , n3493 , n3494 );
xnor ( n3496 , n3495 , n1958 );
and ( n3497 , n2556 , n2012 );
and ( n3498 , n2401 , n2010 );
nor ( n3499 , n3497 , n3498 );
xnor ( n3500 , n3499 , n2020 );
and ( n3501 , n3496 , n3500 );
and ( n3502 , n2919 , n2032 );
and ( n3503 , n2639 , n2030 );
nor ( n3504 , n3502 , n3503 );
xnor ( n3505 , n3504 , n2040 );
and ( n3506 , n3500 , n3505 );
and ( n3507 , n3496 , n3505 );
or ( n3508 , n3501 , n3506 , n3507 );
and ( n3509 , n3491 , n3508 );
and ( n3510 , n3475 , n3508 );
or ( n3511 , n3492 , n3509 , n3510 );
and ( n3512 , n2057 , n3154 );
and ( n3513 , n1942 , n3152 );
nor ( n3514 , n3512 , n3513 );
xnor ( n3515 , n3514 , n2978 );
and ( n3516 , n1996 , n2612 );
and ( n3517 , n1962 , n2610 );
nor ( n3518 , n3516 , n3517 );
xnor ( n3519 , n3518 , n2515 );
and ( n3520 , n3515 , n3519 );
buf ( n530781 , n1151 );
buf ( n3522 , n530781 );
and ( n3523 , n3522 , n1926 );
and ( n3524 , n3519 , n3523 );
and ( n3525 , n3515 , n3523 );
or ( n3526 , n3520 , n3524 , n3525 );
xor ( n3527 , n2975 , n3287 );
xor ( n3528 , n3287 , n3289 );
not ( n3529 , n3528 );
and ( n3530 , n3527 , n3529 );
and ( n3531 , n1953 , n3530 );
not ( n3532 , n3531 );
xnor ( n3533 , n3532 , n3292 );
buf ( n3534 , n3533 );
and ( n3535 , n3526 , n3534 );
and ( n3536 , n3333 , n2091 );
and ( n3537 , n3222 , n2089 );
nor ( n3538 , n3536 , n3537 );
xnor ( n3539 , n3538 , n2099 );
and ( n3540 , n3534 , n3539 );
and ( n3541 , n3526 , n3539 );
or ( n3542 , n3535 , n3540 , n3541 );
and ( n3543 , n3511 , n3542 );
xor ( n3544 , n3326 , n3330 );
xor ( n3545 , n3544 , n3334 );
and ( n3546 , n3542 , n3545 );
and ( n3547 , n3511 , n3545 );
or ( n3548 , n3543 , n3546 , n3547 );
and ( n3549 , n2015 , n2054 );
and ( n3550 , n1904 , n2052 );
nor ( n3551 , n3549 , n3550 );
xnor ( n3552 , n3551 , n2062 );
and ( n3553 , n3222 , n2073 );
and ( n3554 , n3061 , n2071 );
nor ( n3555 , n3553 , n3554 );
xnor ( n3556 , n3555 , n2081 );
and ( n3557 , n3552 , n3556 );
and ( n3558 , n3281 , n2091 );
and ( n3559 , n3333 , n2089 );
nor ( n3560 , n3558 , n3559 );
xnor ( n3561 , n3560 , n2099 );
and ( n3562 , n3556 , n3561 );
and ( n3563 , n3552 , n3561 );
or ( n3564 , n3557 , n3562 , n3563 );
xor ( n3565 , n3274 , n3278 );
xor ( n3566 , n3565 , n3282 );
and ( n3567 , n3564 , n3566 );
xor ( n3568 , n3293 , n3297 );
xor ( n3569 , n3568 , n3302 );
and ( n3570 , n3566 , n3569 );
and ( n3571 , n3564 , n3569 );
or ( n3572 , n3567 , n3570 , n3571 );
xor ( n3573 , n3285 , n3305 );
xor ( n3574 , n3573 , n3322 );
and ( n3575 , n3572 , n3574 );
xor ( n3576 , n3385 , n3401 );
xor ( n3577 , n3576 , n3404 );
and ( n3578 , n3574 , n3577 );
and ( n3579 , n3572 , n3577 );
or ( n3580 , n3575 , n3578 , n3579 );
and ( n3581 , n3548 , n3580 );
xor ( n3582 , n3407 , n3409 );
xor ( n3583 , n3582 , n3412 );
and ( n3584 , n3580 , n3583 );
and ( n3585 , n3548 , n3583 );
or ( n3586 , n3581 , n3584 , n3585 );
xor ( n3587 , n3373 , n3377 );
xor ( n3588 , n3587 , n3382 );
xor ( n3589 , n3310 , n3314 );
xor ( n3590 , n3589 , n3319 );
and ( n3591 , n3588 , n3590 );
xor ( n3592 , n3389 , n3393 );
xor ( n3593 , n3592 , n3398 );
and ( n3594 , n3590 , n3593 );
and ( n3595 , n3588 , n3593 );
or ( n3596 , n3591 , n3594 , n3595 );
and ( n3597 , n1942 , n3530 );
and ( n3598 , n1953 , n3528 );
nor ( n3599 , n3597 , n3598 );
xnor ( n3600 , n3599 , n3292 );
and ( n3601 , n1962 , n2872 );
and ( n3602 , n1975 , n2870 );
nor ( n3603 , n3601 , n3602 );
xnor ( n3604 , n3603 , n2811 );
and ( n3605 , n3600 , n3604 );
and ( n3606 , n2024 , n1972 );
and ( n3607 , n2035 , n1970 );
nor ( n3608 , n3606 , n3607 );
xnor ( n3609 , n3608 , n1980 );
and ( n3610 , n3604 , n3609 );
and ( n3611 , n3600 , n3609 );
or ( n3612 , n3605 , n3610 , n3611 );
and ( n3613 , n2049 , n3154 );
and ( n3614 , n2057 , n3152 );
nor ( n3615 , n3613 , n3614 );
xnor ( n3616 , n3615 , n2978 );
and ( n3617 , n1883 , n2391 );
and ( n3618 , n1896 , n2389 );
nor ( n3619 , n3617 , n3618 );
xnor ( n3620 , n3619 , n1939 );
and ( n3621 , n3616 , n3620 );
and ( n3622 , n2401 , n1912 );
and ( n3623 , n1924 , n1910 );
nor ( n3624 , n3622 , n3623 );
xnor ( n3625 , n3624 , n1920 );
and ( n3626 , n3620 , n3625 );
and ( n3627 , n3616 , n3625 );
or ( n3628 , n3621 , n3626 , n3627 );
and ( n3629 , n3612 , n3628 );
and ( n3630 , n1987 , n2612 );
and ( n3631 , n1996 , n2610 );
nor ( n3632 , n3630 , n3631 );
xnor ( n3633 , n3632 , n2515 );
and ( n3634 , n2065 , n1993 );
and ( n3635 , n2076 , n1991 );
nor ( n3636 , n3634 , n3635 );
xnor ( n3637 , n3636 , n2001 );
and ( n3638 , n3633 , n3637 );
and ( n3639 , n2085 , n1893 );
and ( n3640 , n2094 , n1891 );
nor ( n3641 , n3639 , n3640 );
xnor ( n3642 , n3641 , n1901 );
and ( n3643 , n3637 , n3642 );
and ( n3644 , n3633 , n3642 );
or ( n3645 , n3638 , n3643 , n3644 );
and ( n3646 , n3628 , n3645 );
and ( n3647 , n3612 , n3645 );
or ( n3648 , n3629 , n3646 , n3647 );
and ( n3649 , n2004 , n2054 );
and ( n3650 , n2015 , n2052 );
nor ( n3651 , n3649 , n3650 );
xnor ( n3652 , n3651 , n2062 );
and ( n3653 , n3522 , n2091 );
and ( n3654 , n3281 , n2089 );
nor ( n3655 , n3653 , n3654 );
xnor ( n3656 , n3655 , n2099 );
and ( n3657 , n3652 , n3656 );
buf ( n530918 , n1152 );
buf ( n3659 , n530918 );
and ( n3660 , n3659 , n1926 );
and ( n3661 , n3656 , n3660 );
and ( n3662 , n3652 , n3660 );
or ( n3663 , n3657 , n3661 , n3662 );
not ( n3664 , n3289 );
buf ( n3665 , n3664 );
and ( n3666 , n3663 , n3665 );
not ( n3667 , n3533 );
and ( n3668 , n3665 , n3667 );
and ( n3669 , n3663 , n3667 );
or ( n3670 , n3666 , n3668 , n3669 );
and ( n3671 , n3648 , n3670 );
xor ( n3672 , n3526 , n3534 );
xor ( n3673 , n3672 , n3539 );
and ( n3674 , n3670 , n3673 );
and ( n3675 , n3648 , n3673 );
or ( n3676 , n3671 , n3674 , n3675 );
and ( n3677 , n3596 , n3676 );
xor ( n3678 , n3425 , n3427 );
xor ( n3679 , n3678 , n3430 );
and ( n3680 , n3676 , n3679 );
and ( n3681 , n3596 , n3679 );
or ( n3682 , n3677 , n3680 , n3681 );
and ( n3683 , n1904 , n1950 );
and ( n3684 , n1915 , n1948 );
nor ( n3685 , n3683 , n3684 );
xnor ( n3686 , n3685 , n1958 );
and ( n3687 , n2639 , n2012 );
and ( n3688 , n2556 , n2010 );
nor ( n3689 , n3687 , n3688 );
xnor ( n3690 , n3689 , n2020 );
and ( n3691 , n3686 , n3690 );
and ( n3692 , n3061 , n2032 );
and ( n3693 , n2919 , n2030 );
nor ( n3694 , n3692 , n3693 );
xnor ( n3695 , n3694 , n2040 );
and ( n3696 , n3690 , n3695 );
and ( n3697 , n3686 , n3695 );
or ( n3698 , n3691 , n3696 , n3697 );
xor ( n3699 , n3552 , n3556 );
xor ( n3700 , n3699 , n3561 );
and ( n3701 , n3698 , n3700 );
xor ( n3702 , n3463 , n3467 );
xor ( n3703 , n3702 , n3472 );
and ( n3704 , n3700 , n3703 );
and ( n3705 , n3698 , n3703 );
or ( n3706 , n3701 , n3704 , n3705 );
xor ( n3707 , n3515 , n3519 );
xor ( n3708 , n3707 , n3523 );
xor ( n3709 , n3479 , n3483 );
xor ( n3710 , n3709 , n3488 );
and ( n3711 , n3708 , n3710 );
xor ( n3712 , n3496 , n3500 );
xor ( n3713 , n3712 , n3505 );
and ( n3714 , n3710 , n3713 );
and ( n3715 , n3708 , n3713 );
or ( n3716 , n3711 , n3714 , n3715 );
and ( n3717 , n3706 , n3716 );
xor ( n3718 , n3475 , n3491 );
xor ( n3719 , n3718 , n3508 );
and ( n3720 , n3716 , n3719 );
and ( n3721 , n3706 , n3719 );
or ( n3722 , n3717 , n3720 , n3721 );
xor ( n3723 , n3511 , n3542 );
xor ( n3724 , n3723 , n3545 );
and ( n3725 , n3722 , n3724 );
xor ( n3726 , n3572 , n3574 );
xor ( n3727 , n3726 , n3577 );
and ( n3728 , n3724 , n3727 );
and ( n3729 , n3722 , n3727 );
or ( n3730 , n3725 , n3728 , n3729 );
and ( n3731 , n3682 , n3730 );
xor ( n3732 , n3433 , n3435 );
xor ( n3733 , n3732 , n3438 );
and ( n3734 , n3730 , n3733 );
and ( n3735 , n3682 , n3733 );
or ( n3736 , n3731 , n3734 , n3735 );
and ( n3737 , n3586 , n3736 );
xor ( n3738 , n3441 , n3443 );
xor ( n3739 , n3738 , n3446 );
and ( n3740 , n3736 , n3739 );
and ( n3741 , n3586 , n3739 );
or ( n3742 , n3737 , n3740 , n3741 );
and ( n3743 , n3459 , n3742 );
xor ( n3744 , n3459 , n3742 );
xor ( n3745 , n3586 , n3736 );
xor ( n3746 , n3745 , n3739 );
and ( n3747 , n1996 , n2872 );
and ( n3748 , n1962 , n2870 );
nor ( n3749 , n3747 , n3748 );
xnor ( n3750 , n3749 , n2811 );
and ( n3751 , n2035 , n2054 );
and ( n3752 , n2004 , n2052 );
nor ( n3753 , n3751 , n3752 );
xnor ( n3754 , n3753 , n2062 );
and ( n3755 , n3750 , n3754 );
and ( n3756 , n3659 , n2091 );
and ( n3757 , n3522 , n2089 );
nor ( n3758 , n3756 , n3757 );
xnor ( n3759 , n3758 , n2099 );
and ( n3760 , n3754 , n3759 );
and ( n3761 , n3750 , n3759 );
or ( n3762 , n3755 , n3760 , n3761 );
and ( n3763 , n1896 , n2612 );
and ( n3764 , n1987 , n2610 );
nor ( n3765 , n3763 , n3764 );
xnor ( n3766 , n3765 , n2515 );
and ( n3767 , n2076 , n1972 );
and ( n3768 , n2024 , n1970 );
nor ( n3769 , n3767 , n3768 );
xnor ( n3770 , n3769 , n1980 );
and ( n3771 , n3766 , n3770 );
and ( n3772 , n2094 , n1993 );
and ( n3773 , n2065 , n1991 );
nor ( n3774 , n3772 , n3773 );
xnor ( n3775 , n3774 , n2001 );
and ( n3776 , n3770 , n3775 );
and ( n3777 , n3766 , n3775 );
or ( n3778 , n3771 , n3776 , n3777 );
and ( n3779 , n3762 , n3778 );
and ( n3780 , n2015 , n1950 );
and ( n3781 , n1904 , n1948 );
nor ( n3782 , n3780 , n3781 );
xnor ( n3783 , n3782 , n1958 );
and ( n3784 , n2556 , n1912 );
and ( n3785 , n2401 , n1910 );
nor ( n3786 , n3784 , n3785 );
xnor ( n3787 , n3786 , n1920 );
and ( n3788 , n3783 , n3787 );
and ( n3789 , n2919 , n2012 );
and ( n3790 , n2639 , n2010 );
nor ( n3791 , n3789 , n3790 );
xnor ( n3792 , n3791 , n2020 );
and ( n3793 , n3787 , n3792 );
and ( n3794 , n3783 , n3792 );
or ( n3795 , n3788 , n3793 , n3794 );
and ( n3796 , n3778 , n3795 );
and ( n3797 , n3762 , n3795 );
or ( n3798 , n3779 , n3796 , n3797 );
buf ( n531059 , n1185 );
buf ( n3800 , n531059 );
xor ( n3801 , n3289 , n3800 );
not ( n3802 , n3800 );
and ( n3803 , n3801 , n3802 );
and ( n3804 , n1953 , n3803 );
not ( n3805 , n3804 );
xnor ( n3806 , n3805 , n3289 );
and ( n3807 , n2057 , n3530 );
and ( n3808 , n1942 , n3528 );
nor ( n3809 , n3807 , n3808 );
xnor ( n3810 , n3809 , n3292 );
and ( n3811 , n3806 , n3810 );
buf ( n531072 , n1153 );
buf ( n3813 , n531072 );
and ( n3814 , n3813 , n1926 );
and ( n3815 , n3810 , n3814 );
and ( n3816 , n3806 , n3814 );
or ( n3817 , n3811 , n3815 , n3816 );
and ( n3818 , n3817 , n3289 );
and ( n3819 , n3333 , n2073 );
and ( n3820 , n3222 , n2071 );
nor ( n3821 , n3819 , n3820 );
xnor ( n3822 , n3821 , n2081 );
and ( n3823 , n3289 , n3822 );
and ( n3824 , n3817 , n3822 );
or ( n3825 , n3818 , n3823 , n3824 );
and ( n3826 , n3798 , n3825 );
xor ( n3827 , n3612 , n3628 );
xor ( n3828 , n3827 , n3645 );
and ( n3829 , n3825 , n3828 );
and ( n3830 , n3798 , n3828 );
or ( n3831 , n3826 , n3829 , n3830 );
and ( n3832 , n1975 , n3154 );
and ( n3833 , n2049 , n3152 );
nor ( n3834 , n3832 , n3833 );
xnor ( n3835 , n3834 , n2978 );
and ( n3836 , n1915 , n2391 );
and ( n3837 , n1883 , n2389 );
nor ( n3838 , n3836 , n3837 );
xnor ( n3839 , n3838 , n1939 );
and ( n3840 , n3835 , n3839 );
and ( n3841 , n1924 , n1893 );
and ( n3842 , n2085 , n1891 );
nor ( n3843 , n3841 , n3842 );
xnor ( n3844 , n3843 , n1901 );
and ( n3845 , n3839 , n3844 );
and ( n3846 , n3835 , n3844 );
or ( n3847 , n3840 , n3845 , n3846 );
xor ( n3848 , n3652 , n3656 );
xor ( n3849 , n3848 , n3660 );
and ( n3850 , n3847 , n3849 );
xor ( n3851 , n3686 , n3690 );
xor ( n3852 , n3851 , n3695 );
and ( n3853 , n3849 , n3852 );
and ( n3854 , n3847 , n3852 );
or ( n3855 , n3850 , n3853 , n3854 );
xor ( n3856 , n3600 , n3604 );
xor ( n3857 , n3856 , n3609 );
xor ( n3858 , n3616 , n3620 );
xor ( n3859 , n3858 , n3625 );
and ( n3860 , n3857 , n3859 );
xor ( n3861 , n3633 , n3637 );
xor ( n3862 , n3861 , n3642 );
and ( n3863 , n3859 , n3862 );
and ( n3864 , n3857 , n3862 );
or ( n3865 , n3860 , n3863 , n3864 );
and ( n3866 , n3855 , n3865 );
xor ( n3867 , n3663 , n3665 );
xor ( n3868 , n3867 , n3667 );
and ( n3869 , n3865 , n3868 );
and ( n3870 , n3855 , n3868 );
or ( n3871 , n3866 , n3869 , n3870 );
and ( n3872 , n3831 , n3871 );
xor ( n3873 , n3706 , n3716 );
xor ( n3874 , n3873 , n3719 );
and ( n3875 , n3871 , n3874 );
and ( n3876 , n3831 , n3874 );
or ( n3877 , n3872 , n3875 , n3876 );
xor ( n3878 , n3564 , n3566 );
xor ( n3879 , n3878 , n3569 );
xor ( n3880 , n3588 , n3590 );
xor ( n3881 , n3880 , n3593 );
and ( n3882 , n3879 , n3881 );
xor ( n3883 , n3648 , n3670 );
xor ( n3884 , n3883 , n3673 );
and ( n3885 , n3881 , n3884 );
and ( n3886 , n3879 , n3884 );
or ( n3887 , n3882 , n3885 , n3886 );
and ( n3888 , n3877 , n3887 );
xor ( n3889 , n3596 , n3676 );
xor ( n3890 , n3889 , n3679 );
and ( n3891 , n3887 , n3890 );
and ( n3892 , n3877 , n3890 );
or ( n3893 , n3888 , n3891 , n3892 );
xor ( n3894 , n3548 , n3580 );
xor ( n3895 , n3894 , n3583 );
and ( n3896 , n3893 , n3895 );
xor ( n3897 , n3682 , n3730 );
xor ( n3898 , n3897 , n3733 );
and ( n3899 , n3895 , n3898 );
and ( n3900 , n3893 , n3898 );
or ( n3901 , n3896 , n3899 , n3900 );
and ( n3902 , n3746 , n3901 );
xor ( n3903 , n3746 , n3901 );
xor ( n3904 , n3893 , n3895 );
xor ( n3905 , n3904 , n3898 );
xor ( n3906 , n3766 , n3770 );
xor ( n3907 , n3906 , n3775 );
xor ( n3908 , n3835 , n3839 );
xor ( n3909 , n3908 , n3844 );
and ( n3910 , n3907 , n3909 );
xor ( n3911 , n3783 , n3787 );
xor ( n3912 , n3911 , n3792 );
and ( n3913 , n3909 , n3912 );
and ( n3914 , n3907 , n3912 );
or ( n3915 , n3910 , n3913 , n3914 );
xor ( n3916 , n3762 , n3778 );
xor ( n3917 , n3916 , n3795 );
and ( n3918 , n3915 , n3917 );
xor ( n3919 , n3817 , n3289 );
xor ( n3920 , n3919 , n3822 );
and ( n3921 , n3917 , n3920 );
and ( n3922 , n3915 , n3920 );
or ( n3923 , n3918 , n3921 , n3922 );
xor ( n3924 , n3698 , n3700 );
xor ( n3925 , n3924 , n3703 );
and ( n3926 , n3923 , n3925 );
xor ( n3927 , n3708 , n3710 );
xor ( n3928 , n3927 , n3713 );
and ( n3929 , n3925 , n3928 );
and ( n3930 , n3923 , n3928 );
or ( n3931 , n3926 , n3929 , n3930 );
and ( n3932 , n1942 , n3803 );
and ( n3933 , n1953 , n3800 );
nor ( n3934 , n3932 , n3933 );
xnor ( n3935 , n3934 , n3289 );
and ( n3936 , n3813 , n2089 );
not ( n3937 , n3936 );
and ( n3938 , n3937 , n2099 );
and ( n3939 , n3935 , n3938 );
and ( n3940 , n3222 , n2032 );
and ( n3941 , n3061 , n2030 );
nor ( n3942 , n3940 , n3941 );
xnor ( n3943 , n3942 , n2040 );
and ( n3944 , n3939 , n3943 );
and ( n3945 , n3281 , n2073 );
and ( n3946 , n3333 , n2071 );
nor ( n3947 , n3945 , n3946 );
xnor ( n3948 , n3947 , n2081 );
and ( n3949 , n3943 , n3948 );
and ( n3950 , n3939 , n3948 );
or ( n3951 , n3944 , n3949 , n3950 );
and ( n3952 , n2049 , n3530 );
and ( n3953 , n2057 , n3528 );
nor ( n3954 , n3952 , n3953 );
xnor ( n3955 , n3954 , n3292 );
and ( n3956 , n1987 , n2872 );
and ( n3957 , n1996 , n2870 );
nor ( n3958 , n3956 , n3957 );
xnor ( n3959 , n3958 , n2811 );
and ( n3960 , n3955 , n3959 );
and ( n3961 , n3813 , n2091 );
and ( n3962 , n3659 , n2089 );
nor ( n3963 , n3961 , n3962 );
xnor ( n3964 , n3963 , n2099 );
and ( n3965 , n3959 , n3964 );
and ( n3966 , n3955 , n3964 );
or ( n3967 , n3960 , n3965 , n3966 );
and ( n3968 , n1883 , n2612 );
and ( n3969 , n1896 , n2610 );
nor ( n3970 , n3968 , n3969 );
xnor ( n3971 , n3970 , n2515 );
and ( n3972 , n2024 , n2054 );
and ( n3973 , n2035 , n2052 );
nor ( n3974 , n3972 , n3973 );
xnor ( n3975 , n3974 , n2062 );
and ( n3976 , n3971 , n3975 );
and ( n3977 , n2065 , n1972 );
and ( n3978 , n2076 , n1970 );
nor ( n3979 , n3977 , n3978 );
xnor ( n3980 , n3979 , n1980 );
and ( n3981 , n3975 , n3980 );
and ( n3982 , n3971 , n3980 );
or ( n3983 , n3976 , n3981 , n3982 );
and ( n3984 , n3967 , n3983 );
and ( n3985 , n1962 , n3154 );
and ( n3986 , n1975 , n3152 );
nor ( n3987 , n3985 , n3986 );
xnor ( n3988 , n3987 , n2978 );
and ( n3989 , n2085 , n1993 );
and ( n3990 , n2094 , n1991 );
nor ( n3991 , n3989 , n3990 );
xnor ( n3992 , n3991 , n2001 );
and ( n3993 , n3988 , n3992 );
and ( n3994 , n2401 , n1893 );
and ( n3995 , n1924 , n1891 );
nor ( n3996 , n3994 , n3995 );
xnor ( n3997 , n3996 , n1901 );
and ( n3998 , n3992 , n3997 );
and ( n3999 , n3988 , n3997 );
or ( n4000 , n3993 , n3998 , n3999 );
and ( n4001 , n3983 , n4000 );
and ( n4002 , n3967 , n4000 );
or ( n4003 , n3984 , n4001 , n4002 );
and ( n4004 , n3951 , n4003 );
and ( n4005 , n2004 , n1950 );
and ( n4006 , n2015 , n1948 );
nor ( n4007 , n4005 , n4006 );
xnor ( n4008 , n4007 , n1958 );
and ( n4009 , n3333 , n2032 );
and ( n4010 , n3222 , n2030 );
nor ( n4011 , n4009 , n4010 );
xnor ( n4012 , n4011 , n2040 );
and ( n4013 , n4008 , n4012 );
and ( n4014 , n3522 , n2073 );
and ( n4015 , n3281 , n2071 );
nor ( n4016 , n4014 , n4015 );
xnor ( n4017 , n4016 , n2081 );
and ( n4018 , n4012 , n4017 );
and ( n4019 , n4008 , n4017 );
or ( n4020 , n4013 , n4018 , n4019 );
and ( n4021 , n1904 , n2391 );
and ( n4022 , n1915 , n2389 );
nor ( n4023 , n4021 , n4022 );
xnor ( n4024 , n4023 , n1939 );
and ( n4025 , n2639 , n1912 );
and ( n4026 , n2556 , n1910 );
nor ( n4027 , n4025 , n4026 );
xnor ( n4028 , n4027 , n1920 );
and ( n4029 , n4024 , n4028 );
and ( n4030 , n3061 , n2012 );
and ( n4031 , n2919 , n2010 );
nor ( n4032 , n4030 , n4031 );
xnor ( n4033 , n4032 , n2020 );
and ( n4034 , n4028 , n4033 );
and ( n4035 , n4024 , n4033 );
or ( n4036 , n4029 , n4034 , n4035 );
and ( n4037 , n4020 , n4036 );
xor ( n4038 , n3806 , n3810 );
xor ( n4039 , n4038 , n3814 );
and ( n4040 , n4036 , n4039 );
and ( n4041 , n4020 , n4039 );
or ( n4042 , n4037 , n4040 , n4041 );
and ( n4043 , n4003 , n4042 );
and ( n4044 , n3951 , n4042 );
or ( n4045 , n4004 , n4043 , n4044 );
xor ( n4046 , n3798 , n3825 );
xor ( n4047 , n4046 , n3828 );
and ( n4048 , n4045 , n4047 );
xor ( n4049 , n3855 , n3865 );
xor ( n4050 , n4049 , n3868 );
and ( n4051 , n4047 , n4050 );
and ( n4052 , n4045 , n4050 );
or ( n4053 , n4048 , n4051 , n4052 );
and ( n4054 , n3931 , n4053 );
xor ( n4055 , n3879 , n3881 );
xor ( n4056 , n4055 , n3884 );
and ( n4057 , n4053 , n4056 );
and ( n4058 , n3931 , n4056 );
or ( n4059 , n4054 , n4057 , n4058 );
xor ( n4060 , n3722 , n3724 );
xor ( n4061 , n4060 , n3727 );
and ( n4062 , n4059 , n4061 );
xor ( n4063 , n3877 , n3887 );
xor ( n4064 , n4063 , n3890 );
and ( n4065 , n4061 , n4064 );
and ( n4066 , n4059 , n4064 );
or ( n4067 , n4062 , n4065 , n4066 );
and ( n4068 , n3905 , n4067 );
xor ( n4069 , n3905 , n4067 );
xor ( n4070 , n4059 , n4061 );
xor ( n4071 , n4070 , n4064 );
and ( n4072 , n2035 , n1950 );
and ( n4073 , n2004 , n1948 );
nor ( n4074 , n4072 , n4073 );
xnor ( n4075 , n4074 , n1958 );
and ( n4076 , n3222 , n2012 );
and ( n4077 , n3061 , n2010 );
nor ( n4078 , n4076 , n4077 );
xnor ( n4079 , n4078 , n2020 );
and ( n4080 , n4075 , n4079 );
and ( n4081 , n3281 , n2032 );
and ( n4082 , n3333 , n2030 );
nor ( n4083 , n4081 , n4082 );
xnor ( n4084 , n4083 , n2040 );
and ( n4085 , n4079 , n4084 );
and ( n4086 , n4075 , n4084 );
or ( n4087 , n4080 , n4085 , n4086 );
and ( n4088 , n1996 , n3154 );
and ( n4089 , n1962 , n3152 );
nor ( n4090 , n4088 , n4089 );
xnor ( n4091 , n4090 , n2978 );
and ( n4092 , n2015 , n2391 );
and ( n4093 , n1904 , n2389 );
nor ( n4094 , n4092 , n4093 );
xnor ( n4095 , n4094 , n1939 );
and ( n4096 , n4091 , n4095 );
and ( n4097 , n2919 , n1912 );
and ( n4098 , n2639 , n1910 );
nor ( n4099 , n4097 , n4098 );
xnor ( n4100 , n4099 , n1920 );
and ( n4101 , n4095 , n4100 );
and ( n4102 , n4091 , n4100 );
or ( n4103 , n4096 , n4101 , n4102 );
and ( n4104 , n4087 , n4103 );
and ( n4105 , n1915 , n2612 );
and ( n4106 , n1883 , n2610 );
nor ( n4107 , n4105 , n4106 );
xnor ( n4108 , n4107 , n2515 );
and ( n4109 , n1924 , n1993 );
and ( n4110 , n2085 , n1991 );
nor ( n4111 , n4109 , n4110 );
xnor ( n4112 , n4111 , n2001 );
and ( n4113 , n4108 , n4112 );
and ( n4114 , n2556 , n1893 );
and ( n4115 , n2401 , n1891 );
nor ( n4116 , n4114 , n4115 );
xnor ( n4117 , n4116 , n1901 );
and ( n4118 , n4112 , n4117 );
and ( n4119 , n4108 , n4117 );
or ( n4120 , n4113 , n4118 , n4119 );
and ( n4121 , n4103 , n4120 );
and ( n4122 , n4087 , n4120 );
or ( n4123 , n4104 , n4121 , n4122 );
xor ( n4124 , n3750 , n3754 );
xor ( n4125 , n4124 , n3759 );
and ( n4126 , n4123 , n4125 );
xor ( n4127 , n3939 , n3943 );
xor ( n4128 , n4127 , n3948 );
and ( n4129 , n4125 , n4128 );
and ( n4130 , n4123 , n4128 );
or ( n4131 , n4126 , n4129 , n4130 );
xor ( n4132 , n3847 , n3849 );
xor ( n4133 , n4132 , n3852 );
and ( n4134 , n4131 , n4133 );
xor ( n4135 , n3857 , n3859 );
xor ( n4136 , n4135 , n3862 );
and ( n4137 , n4133 , n4136 );
and ( n4138 , n4131 , n4136 );
or ( n4139 , n4134 , n4137 , n4138 );
xor ( n4140 , n3935 , n3938 );
and ( n4141 , n2057 , n3803 );
and ( n4142 , n1942 , n3800 );
nor ( n4143 , n4141 , n4142 );
xnor ( n4144 , n4143 , n3289 );
and ( n4145 , n1975 , n3530 );
and ( n4146 , n2049 , n3528 );
nor ( n4147 , n4145 , n4146 );
xnor ( n4148 , n4147 , n3292 );
and ( n4149 , n4144 , n4148 );
and ( n4150 , n4148 , n3936 );
and ( n4151 , n4144 , n3936 );
or ( n4152 , n4149 , n4150 , n4151 );
and ( n4153 , n4140 , n4152 );
and ( n4154 , n1896 , n2872 );
and ( n4155 , n1987 , n2870 );
nor ( n4156 , n4154 , n4155 );
xnor ( n4157 , n4156 , n2811 );
and ( n4158 , n2076 , n2054 );
and ( n4159 , n2024 , n2052 );
nor ( n4160 , n4158 , n4159 );
xnor ( n4161 , n4160 , n2062 );
and ( n4162 , n4157 , n4161 );
and ( n4163 , n2094 , n1972 );
and ( n4164 , n2065 , n1970 );
nor ( n4165 , n4163 , n4164 );
xnor ( n4166 , n4165 , n1980 );
and ( n4167 , n4161 , n4166 );
and ( n4168 , n4157 , n4166 );
or ( n4169 , n4162 , n4167 , n4168 );
and ( n4170 , n4152 , n4169 );
and ( n4171 , n4140 , n4169 );
or ( n4172 , n4153 , n4170 , n4171 );
xor ( n4173 , n4008 , n4012 );
xor ( n4174 , n4173 , n4017 );
xor ( n4175 , n3955 , n3959 );
xor ( n4176 , n4175 , n3964 );
and ( n4177 , n4174 , n4176 );
xor ( n4178 , n3971 , n3975 );
xor ( n4179 , n4178 , n3980 );
and ( n4180 , n4176 , n4179 );
and ( n4181 , n4174 , n4179 );
or ( n4182 , n4177 , n4180 , n4181 );
and ( n4183 , n4172 , n4182 );
xor ( n4184 , n4020 , n4036 );
xor ( n4185 , n4184 , n4039 );
and ( n4186 , n4182 , n4185 );
and ( n4187 , n4172 , n4185 );
or ( n4188 , n4183 , n4186 , n4187 );
xor ( n4189 , n3951 , n4003 );
xor ( n4190 , n4189 , n4042 );
and ( n4191 , n4188 , n4190 );
xor ( n4192 , n3915 , n3917 );
xor ( n4193 , n4192 , n3920 );
and ( n4194 , n4190 , n4193 );
and ( n4195 , n4188 , n4193 );
or ( n4196 , n4191 , n4194 , n4195 );
and ( n4197 , n4139 , n4196 );
xor ( n4198 , n3923 , n3925 );
xor ( n4199 , n4198 , n3928 );
and ( n4200 , n4196 , n4199 );
and ( n4201 , n4139 , n4199 );
or ( n4202 , n4197 , n4200 , n4201 );
xor ( n4203 , n3831 , n3871 );
xor ( n4204 , n4203 , n3874 );
and ( n4205 , n4202 , n4204 );
xor ( n4206 , n3931 , n4053 );
xor ( n4207 , n4206 , n4056 );
and ( n4208 , n4204 , n4207 );
and ( n4209 , n4202 , n4207 );
or ( n4210 , n4205 , n4208 , n4209 );
and ( n4211 , n4071 , n4210 );
xor ( n4212 , n4071 , n4210 );
and ( n4213 , n2024 , n1950 );
and ( n4214 , n2035 , n1948 );
nor ( n4215 , n4213 , n4214 );
xnor ( n4216 , n4215 , n1958 );
and ( n4217 , n3061 , n1912 );
and ( n4218 , n2919 , n1910 );
nor ( n4219 , n4217 , n4218 );
xnor ( n4220 , n4219 , n1920 );
and ( n4221 , n4216 , n4220 );
and ( n4222 , n3333 , n2012 );
and ( n4223 , n3222 , n2010 );
nor ( n4224 , n4222 , n4223 );
xnor ( n4225 , n4224 , n2020 );
and ( n4226 , n4220 , n4225 );
and ( n4227 , n4216 , n4225 );
or ( n4228 , n4221 , n4226 , n4227 );
and ( n4229 , n1904 , n2612 );
and ( n4230 , n1915 , n2610 );
nor ( n4231 , n4229 , n4230 );
xnor ( n4232 , n4231 , n2515 );
and ( n4233 , n2085 , n1972 );
and ( n4234 , n2094 , n1970 );
nor ( n4235 , n4233 , n4234 );
xnor ( n4236 , n4235 , n1980 );
and ( n4237 , n4232 , n4236 );
and ( n4238 , n2401 , n1993 );
and ( n4239 , n1924 , n1991 );
nor ( n4240 , n4238 , n4239 );
xnor ( n4241 , n4240 , n2001 );
and ( n4242 , n4236 , n4241 );
and ( n4243 , n4232 , n4241 );
or ( n4244 , n4237 , n4242 , n4243 );
and ( n4245 , n4228 , n4244 );
and ( n4246 , n1987 , n3154 );
and ( n4247 , n1996 , n3152 );
nor ( n4248 , n4246 , n4247 );
xnor ( n4249 , n4248 , n2978 );
and ( n4250 , n2004 , n2391 );
and ( n4251 , n2015 , n2389 );
nor ( n4252 , n4250 , n4251 );
xnor ( n4253 , n4252 , n1939 );
and ( n4254 , n4249 , n4253 );
and ( n4255 , n2639 , n1893 );
and ( n4256 , n2556 , n1891 );
nor ( n4257 , n4255 , n4256 );
xnor ( n4258 , n4257 , n1901 );
and ( n4259 , n4253 , n4258 );
and ( n4260 , n4249 , n4258 );
or ( n4261 , n4254 , n4259 , n4260 );
and ( n4262 , n4244 , n4261 );
and ( n4263 , n4228 , n4261 );
or ( n4264 , n4245 , n4262 , n4263 );
xor ( n4265 , n3988 , n3992 );
xor ( n4266 , n4265 , n3997 );
and ( n4267 , n4264 , n4266 );
xor ( n4268 , n4024 , n4028 );
xor ( n4269 , n4268 , n4033 );
and ( n4270 , n4266 , n4269 );
and ( n4271 , n4264 , n4269 );
or ( n4272 , n4267 , n4270 , n4271 );
xor ( n4273 , n3967 , n3983 );
xor ( n4274 , n4273 , n4000 );
and ( n4275 , n4272 , n4274 );
xor ( n4276 , n3907 , n3909 );
xor ( n4277 , n4276 , n3912 );
and ( n4278 , n4274 , n4277 );
and ( n4279 , n4272 , n4277 );
or ( n4280 , n4275 , n4278 , n4279 );
and ( n4281 , n1962 , n3530 );
and ( n4282 , n1975 , n3528 );
nor ( n4283 , n4281 , n4282 );
xnor ( n4284 , n4283 , n3292 );
and ( n4285 , n1883 , n2872 );
and ( n4286 , n1896 , n2870 );
nor ( n4287 , n4285 , n4286 );
xnor ( n4288 , n4287 , n2811 );
and ( n4289 , n4284 , n4288 );
and ( n4290 , n2065 , n2054 );
and ( n4291 , n2076 , n2052 );
nor ( n4292 , n4290 , n4291 );
xnor ( n4293 , n4292 , n2062 );
and ( n4294 , n4288 , n4293 );
and ( n4295 , n4284 , n4293 );
or ( n4296 , n4289 , n4294 , n4295 );
and ( n4297 , n2049 , n3803 );
and ( n4298 , n2057 , n3800 );
nor ( n4299 , n4297 , n4298 );
xnor ( n4300 , n4299 , n3289 );
and ( n4301 , n3813 , n2071 );
not ( n4302 , n4301 );
and ( n4303 , n4302 , n2081 );
and ( n4304 , n4300 , n4303 );
and ( n4305 , n4296 , n4304 );
and ( n4306 , n3659 , n2073 );
and ( n4307 , n3522 , n2071 );
nor ( n4308 , n4306 , n4307 );
xnor ( n4309 , n4308 , n2081 );
and ( n4310 , n4304 , n4309 );
and ( n4311 , n4296 , n4309 );
or ( n4312 , n4305 , n4310 , n4311 );
xor ( n4313 , n4087 , n4103 );
xor ( n4314 , n4313 , n4120 );
and ( n4315 , n4312 , n4314 );
xor ( n4316 , n4140 , n4152 );
xor ( n4317 , n4316 , n4169 );
and ( n4318 , n4314 , n4317 );
and ( n4319 , n4312 , n4317 );
or ( n4320 , n4315 , n4318 , n4319 );
xor ( n4321 , n4144 , n4148 );
xor ( n4322 , n4321 , n3936 );
xor ( n4323 , n4075 , n4079 );
xor ( n4324 , n4323 , n4084 );
and ( n4325 , n4322 , n4324 );
xor ( n4326 , n4091 , n4095 );
xor ( n4327 , n4326 , n4100 );
and ( n4328 , n4324 , n4327 );
and ( n4329 , n4322 , n4327 );
or ( n4330 , n4325 , n4328 , n4329 );
xor ( n4331 , n4300 , n4303 );
and ( n4332 , n3522 , n2032 );
and ( n4333 , n3281 , n2030 );
nor ( n4334 , n4332 , n4333 );
xnor ( n4335 , n4334 , n2040 );
and ( n4336 , n4331 , n4335 );
and ( n4337 , n3813 , n2073 );
and ( n4338 , n3659 , n2071 );
nor ( n4339 , n4337 , n4338 );
xnor ( n4340 , n4339 , n2081 );
and ( n4341 , n4335 , n4340 );
and ( n4342 , n4331 , n4340 );
or ( n4343 , n4336 , n4341 , n4342 );
xor ( n4344 , n4108 , n4112 );
xor ( n4345 , n4344 , n4117 );
and ( n4346 , n4343 , n4345 );
xor ( n4347 , n4157 , n4161 );
xor ( n4348 , n4347 , n4166 );
and ( n4349 , n4345 , n4348 );
and ( n4350 , n4343 , n4348 );
or ( n4351 , n4346 , n4349 , n4350 );
and ( n4352 , n4330 , n4351 );
xor ( n4353 , n4174 , n4176 );
xor ( n4354 , n4353 , n4179 );
and ( n4355 , n4351 , n4354 );
and ( n4356 , n4330 , n4354 );
or ( n4357 , n4352 , n4355 , n4356 );
and ( n4358 , n4320 , n4357 );
xor ( n4359 , n4123 , n4125 );
xor ( n4360 , n4359 , n4128 );
and ( n4361 , n4357 , n4360 );
and ( n4362 , n4320 , n4360 );
or ( n4363 , n4358 , n4361 , n4362 );
and ( n4364 , n4280 , n4363 );
xor ( n4365 , n4131 , n4133 );
xor ( n4366 , n4365 , n4136 );
and ( n4367 , n4363 , n4366 );
and ( n4368 , n4280 , n4366 );
or ( n4369 , n4364 , n4367 , n4368 );
xor ( n4370 , n4045 , n4047 );
xor ( n4371 , n4370 , n4050 );
and ( n4372 , n4369 , n4371 );
xor ( n4373 , n4139 , n4196 );
xor ( n4374 , n4373 , n4199 );
and ( n4375 , n4371 , n4374 );
and ( n4376 , n4369 , n4374 );
or ( n4377 , n4372 , n4375 , n4376 );
xor ( n4378 , n4202 , n4204 );
xor ( n4379 , n4378 , n4207 );
and ( n4380 , n4377 , n4379 );
xor ( n4381 , n4377 , n4379 );
xor ( n4382 , n4369 , n4371 );
xor ( n4383 , n4382 , n4374 );
xor ( n4384 , n4172 , n4182 );
xor ( n4385 , n4384 , n4185 );
xor ( n4386 , n4272 , n4274 );
xor ( n4387 , n4386 , n4277 );
and ( n4388 , n4385 , n4387 );
xor ( n4389 , n4320 , n4357 );
xor ( n4390 , n4389 , n4360 );
and ( n4391 , n4387 , n4390 );
and ( n4392 , n4385 , n4390 );
or ( n4393 , n4388 , n4391 , n4392 );
xor ( n4394 , n4188 , n4190 );
xor ( n4395 , n4394 , n4193 );
and ( n4396 , n4393 , n4395 );
xor ( n4397 , n4280 , n4363 );
xor ( n4398 , n4397 , n4366 );
and ( n4399 , n4395 , n4398 );
and ( n4400 , n4393 , n4398 );
or ( n4401 , n4396 , n4399 , n4400 );
and ( n4402 , n4383 , n4401 );
xor ( n4403 , n4383 , n4401 );
xor ( n4404 , n4393 , n4395 );
xor ( n4405 , n4404 , n4398 );
and ( n4406 , n1996 , n3530 );
and ( n4407 , n1962 , n3528 );
nor ( n4408 , n4406 , n4407 );
xnor ( n4409 , n4408 , n3292 );
and ( n4410 , n1915 , n2872 );
and ( n4411 , n1883 , n2870 );
nor ( n4412 , n4410 , n4411 );
xnor ( n4413 , n4412 , n2811 );
and ( n4414 , n4409 , n4413 );
and ( n4415 , n4413 , n4301 );
and ( n4416 , n4409 , n4301 );
or ( n4417 , n4414 , n4415 , n4416 );
and ( n4418 , n1975 , n3803 );
and ( n4419 , n2049 , n3800 );
nor ( n4420 , n4418 , n4419 );
xnor ( n4421 , n4420 , n3289 );
and ( n4422 , n2556 , n1993 );
and ( n4423 , n2401 , n1991 );
nor ( n4424 , n4422 , n4423 );
xnor ( n4425 , n4424 , n2001 );
and ( n4426 , n4421 , n4425 );
and ( n4427 , n2919 , n1893 );
and ( n4428 , n2639 , n1891 );
nor ( n4429 , n4427 , n4428 );
xnor ( n4430 , n4429 , n1901 );
and ( n4431 , n4425 , n4430 );
and ( n4432 , n4421 , n4430 );
or ( n4433 , n4426 , n4431 , n4432 );
and ( n4434 , n4417 , n4433 );
and ( n4435 , n2015 , n2612 );
and ( n4436 , n1904 , n2610 );
nor ( n4437 , n4435 , n4436 );
xnor ( n4438 , n4437 , n2515 );
and ( n4439 , n2094 , n2054 );
and ( n4440 , n2065 , n2052 );
nor ( n4441 , n4439 , n4440 );
xnor ( n4442 , n4441 , n2062 );
and ( n4443 , n4438 , n4442 );
and ( n4444 , n1924 , n1972 );
and ( n4445 , n2085 , n1970 );
nor ( n4446 , n4444 , n4445 );
xnor ( n4447 , n4446 , n1980 );
and ( n4448 , n4442 , n4447 );
and ( n4449 , n4438 , n4447 );
or ( n4450 , n4443 , n4448 , n4449 );
and ( n4451 , n4433 , n4450 );
and ( n4452 , n4417 , n4450 );
or ( n4453 , n4434 , n4451 , n4452 );
xor ( n4454 , n4216 , n4220 );
xor ( n4455 , n4454 , n4225 );
xor ( n4456 , n4232 , n4236 );
xor ( n4457 , n4456 , n4241 );
and ( n4458 , n4455 , n4457 );
xor ( n4459 , n4249 , n4253 );
xor ( n4460 , n4459 , n4258 );
and ( n4461 , n4457 , n4460 );
and ( n4462 , n4455 , n4460 );
or ( n4463 , n4458 , n4461 , n4462 );
and ( n4464 , n4453 , n4463 );
xor ( n4465 , n4296 , n4304 );
xor ( n4466 , n4465 , n4309 );
and ( n4467 , n4463 , n4466 );
and ( n4468 , n4453 , n4466 );
or ( n4469 , n4464 , n4467 , n4468 );
and ( n4470 , n1896 , n3154 );
and ( n4471 , n1987 , n3152 );
nor ( n4472 , n4470 , n4471 );
xnor ( n4473 , n4472 , n2978 );
and ( n4474 , n2076 , n1950 );
and ( n4475 , n2024 , n1948 );
nor ( n4476 , n4474 , n4475 );
xnor ( n4477 , n4476 , n1958 );
and ( n4478 , n4473 , n4477 );
and ( n4479 , n3659 , n2032 );
and ( n4480 , n3522 , n2030 );
nor ( n4481 , n4479 , n4480 );
xnor ( n4482 , n4481 , n2040 );
and ( n4483 , n4477 , n4482 );
and ( n4484 , n4473 , n4482 );
or ( n4485 , n4478 , n4483 , n4484 );
and ( n4486 , n2035 , n2391 );
and ( n4487 , n2004 , n2389 );
nor ( n4488 , n4486 , n4487 );
xnor ( n4489 , n4488 , n1939 );
and ( n4490 , n3222 , n1912 );
and ( n4491 , n3061 , n1910 );
nor ( n4492 , n4490 , n4491 );
xnor ( n4493 , n4492 , n1920 );
and ( n4494 , n4489 , n4493 );
and ( n4495 , n3281 , n2012 );
and ( n4496 , n3333 , n2010 );
nor ( n4497 , n4495 , n4496 );
xnor ( n4498 , n4497 , n2020 );
and ( n4499 , n4493 , n4498 );
and ( n4500 , n4489 , n4498 );
or ( n4501 , n4494 , n4499 , n4500 );
and ( n4502 , n4485 , n4501 );
xor ( n4503 , n4284 , n4288 );
xor ( n4504 , n4503 , n4293 );
and ( n4505 , n4501 , n4504 );
and ( n4506 , n4485 , n4504 );
or ( n4507 , n4502 , n4505 , n4506 );
xor ( n4508 , n4228 , n4244 );
xor ( n4509 , n4508 , n4261 );
and ( n4510 , n4507 , n4509 );
xor ( n4511 , n4343 , n4345 );
xor ( n4512 , n4511 , n4348 );
and ( n4513 , n4509 , n4512 );
and ( n4514 , n4507 , n4512 );
or ( n4515 , n4510 , n4513 , n4514 );
and ( n4516 , n4469 , n4515 );
xor ( n4517 , n4264 , n4266 );
xor ( n4518 , n4517 , n4269 );
and ( n4519 , n4515 , n4518 );
and ( n4520 , n4469 , n4518 );
or ( n4521 , n4516 , n4519 , n4520 );
and ( n4522 , n1904 , n2872 );
and ( n4523 , n1915 , n2870 );
nor ( n4524 , n4522 , n4523 );
xnor ( n4525 , n4524 , n2811 );
and ( n4526 , n2085 , n2054 );
and ( n4527 , n2094 , n2052 );
nor ( n4528 , n4526 , n4527 );
xnor ( n4529 , n4528 , n2062 );
and ( n4530 , n4525 , n4529 );
and ( n4531 , n2401 , n1972 );
and ( n4532 , n1924 , n1970 );
nor ( n4533 , n4531 , n4532 );
xnor ( n4534 , n4533 , n1980 );
and ( n4535 , n4529 , n4534 );
and ( n4536 , n4525 , n4534 );
or ( n4537 , n4530 , n4535 , n4536 );
and ( n4538 , n2004 , n2612 );
and ( n4539 , n2015 , n2610 );
nor ( n4540 , n4538 , n4539 );
xnor ( n4541 , n4540 , n2515 );
and ( n4542 , n2639 , n1993 );
and ( n4543 , n2556 , n1991 );
nor ( n4544 , n4542 , n4543 );
xnor ( n4545 , n4544 , n2001 );
and ( n4546 , n4541 , n4545 );
and ( n4547 , n3061 , n1893 );
and ( n4548 , n2919 , n1891 );
nor ( n4549 , n4547 , n4548 );
xnor ( n4550 , n4549 , n1901 );
and ( n4551 , n4545 , n4550 );
and ( n4552 , n4541 , n4550 );
or ( n4553 , n4546 , n4551 , n4552 );
and ( n4554 , n4537 , n4553 );
and ( n4555 , n1987 , n3530 );
and ( n4556 , n1996 , n3528 );
nor ( n4557 , n4555 , n4556 );
xnor ( n4558 , n4557 , n3292 );
and ( n4559 , n3813 , n2030 );
not ( n4560 , n4559 );
and ( n4561 , n4560 , n2040 );
and ( n4562 , n4558 , n4561 );
and ( n4563 , n4553 , n4562 );
and ( n4564 , n4537 , n4562 );
or ( n4565 , n4554 , n4563 , n4564 );
xor ( n4566 , n4473 , n4477 );
xor ( n4567 , n4566 , n4482 );
xor ( n4568 , n4409 , n4413 );
xor ( n4569 , n4568 , n4301 );
and ( n4570 , n4567 , n4569 );
xor ( n4571 , n4421 , n4425 );
xor ( n4572 , n4571 , n4430 );
and ( n4573 , n4569 , n4572 );
and ( n4574 , n4567 , n4572 );
or ( n4575 , n4570 , n4573 , n4574 );
and ( n4576 , n4565 , n4575 );
xor ( n4577 , n4331 , n4335 );
xor ( n4578 , n4577 , n4340 );
and ( n4579 , n4575 , n4578 );
and ( n4580 , n4565 , n4578 );
or ( n4581 , n4576 , n4579 , n4580 );
and ( n4582 , n1883 , n3154 );
and ( n4583 , n1896 , n3152 );
nor ( n4584 , n4582 , n4583 );
xnor ( n4585 , n4584 , n2978 );
and ( n4586 , n3522 , n2012 );
and ( n4587 , n3281 , n2010 );
nor ( n4588 , n4586 , n4587 );
xnor ( n4589 , n4588 , n2020 );
and ( n4590 , n4585 , n4589 );
and ( n4591 , n3813 , n2032 );
and ( n4592 , n3659 , n2030 );
nor ( n4593 , n4591 , n4592 );
xnor ( n4594 , n4593 , n2040 );
and ( n4595 , n4589 , n4594 );
and ( n4596 , n4585 , n4594 );
or ( n4597 , n4590 , n4595 , n4596 );
and ( n4598 , n1962 , n3803 );
and ( n4599 , n1975 , n3800 );
nor ( n4600 , n4598 , n4599 );
xnor ( n4601 , n4600 , n3289 );
and ( n4602 , n2024 , n2391 );
and ( n4603 , n2035 , n2389 );
nor ( n4604 , n4602 , n4603 );
xnor ( n4605 , n4604 , n1939 );
and ( n4606 , n4601 , n4605 );
and ( n4607 , n3333 , n1912 );
and ( n4608 , n3222 , n1910 );
nor ( n4609 , n4607 , n4608 );
xnor ( n4610 , n4609 , n1920 );
and ( n4611 , n4605 , n4610 );
and ( n4612 , n4601 , n4610 );
or ( n4613 , n4606 , n4611 , n4612 );
and ( n4614 , n4597 , n4613 );
xor ( n4615 , n4438 , n4442 );
xor ( n4616 , n4615 , n4447 );
and ( n4617 , n4613 , n4616 );
and ( n4618 , n4597 , n4616 );
or ( n4619 , n4614 , n4617 , n4618 );
xor ( n4620 , n4417 , n4433 );
xor ( n4621 , n4620 , n4450 );
and ( n4622 , n4619 , n4621 );
xor ( n4623 , n4485 , n4501 );
xor ( n4624 , n4623 , n4504 );
and ( n4625 , n4621 , n4624 );
and ( n4626 , n4619 , n4624 );
or ( n4627 , n4622 , n4625 , n4626 );
and ( n4628 , n4581 , n4627 );
xor ( n4629 , n4322 , n4324 );
xor ( n4630 , n4629 , n4327 );
and ( n4631 , n4627 , n4630 );
and ( n4632 , n4581 , n4630 );
or ( n4633 , n4628 , n4631 , n4632 );
xor ( n4634 , n4312 , n4314 );
xor ( n4635 , n4634 , n4317 );
and ( n4636 , n4633 , n4635 );
xor ( n4637 , n4330 , n4351 );
xor ( n4638 , n4637 , n4354 );
and ( n4639 , n4635 , n4638 );
and ( n4640 , n4633 , n4638 );
or ( n4641 , n4636 , n4639 , n4640 );
and ( n4642 , n4521 , n4641 );
xor ( n4643 , n4385 , n4387 );
xor ( n4644 , n4643 , n4390 );
and ( n4645 , n4641 , n4644 );
and ( n4646 , n4521 , n4644 );
or ( n4647 , n4642 , n4645 , n4646 );
and ( n4648 , n4405 , n4647 );
xor ( n4649 , n4405 , n4647 );
and ( n4650 , n2035 , n2612 );
and ( n4651 , n2004 , n2610 );
nor ( n4652 , n4650 , n4651 );
xnor ( n4653 , n4652 , n2515 );
and ( n4654 , n1924 , n2054 );
and ( n4655 , n2085 , n2052 );
nor ( n4656 , n4654 , n4655 );
xnor ( n4657 , n4656 , n2062 );
and ( n4658 , n4653 , n4657 );
and ( n4659 , n2556 , n1972 );
and ( n4660 , n2401 , n1970 );
nor ( n4661 , n4659 , n4660 );
xnor ( n4662 , n4661 , n1980 );
and ( n4663 , n4657 , n4662 );
and ( n4664 , n4653 , n4662 );
or ( n4665 , n4658 , n4663 , n4664 );
and ( n4666 , n2076 , n2391 );
and ( n4667 , n2024 , n2389 );
nor ( n4668 , n4666 , n4667 );
xnor ( n4669 , n4668 , n1939 );
and ( n4670 , n3281 , n1912 );
and ( n4671 , n3333 , n1910 );
nor ( n4672 , n4670 , n4671 );
xnor ( n4673 , n4672 , n1920 );
and ( n4674 , n4669 , n4673 );
and ( n4675 , n3659 , n2012 );
and ( n4676 , n3522 , n2010 );
nor ( n4677 , n4675 , n4676 );
xnor ( n4678 , n4677 , n2020 );
and ( n4679 , n4673 , n4678 );
and ( n4680 , n4669 , n4678 );
or ( n4681 , n4674 , n4679 , n4680 );
and ( n4682 , n4665 , n4681 );
and ( n4683 , n1996 , n3803 );
and ( n4684 , n1962 , n3800 );
nor ( n4685 , n4683 , n4684 );
xnor ( n4686 , n4685 , n3289 );
and ( n4687 , n2919 , n1993 );
and ( n4688 , n2639 , n1991 );
nor ( n4689 , n4687 , n4688 );
xnor ( n4690 , n4689 , n2001 );
and ( n4691 , n4686 , n4690 );
and ( n4692 , n3222 , n1893 );
and ( n4693 , n3061 , n1891 );
nor ( n4694 , n4692 , n4693 );
xnor ( n4695 , n4694 , n1901 );
and ( n4696 , n4690 , n4695 );
and ( n4697 , n4686 , n4695 );
or ( n4698 , n4691 , n4696 , n4697 );
and ( n4699 , n4681 , n4698 );
and ( n4700 , n4665 , n4698 );
or ( n4701 , n4682 , n4699 , n4700 );
xor ( n4702 , n4558 , n4561 );
and ( n4703 , n1896 , n3530 );
and ( n4704 , n1987 , n3528 );
nor ( n4705 , n4703 , n4704 );
xnor ( n4706 , n4705 , n3292 );
and ( n4707 , n2015 , n2872 );
and ( n4708 , n1904 , n2870 );
nor ( n4709 , n4707 , n4708 );
xnor ( n4710 , n4709 , n2811 );
and ( n4711 , n4706 , n4710 );
and ( n4712 , n4710 , n4559 );
and ( n4713 , n4706 , n4559 );
or ( n4714 , n4711 , n4712 , n4713 );
and ( n4715 , n4702 , n4714 );
and ( n4716 , n2065 , n1950 );
and ( n4717 , n2076 , n1948 );
nor ( n4718 , n4716 , n4717 );
xnor ( n4719 , n4718 , n1958 );
and ( n4720 , n4714 , n4719 );
and ( n4721 , n4702 , n4719 );
or ( n4722 , n4715 , n4720 , n4721 );
and ( n4723 , n4701 , n4722 );
xor ( n4724 , n4489 , n4493 );
xor ( n4725 , n4724 , n4498 );
and ( n4726 , n4722 , n4725 );
and ( n4727 , n4701 , n4725 );
or ( n4728 , n4723 , n4726 , n4727 );
xor ( n4729 , n4585 , n4589 );
xor ( n4730 , n4729 , n4594 );
xor ( n4731 , n4525 , n4529 );
xor ( n4732 , n4731 , n4534 );
and ( n4733 , n4730 , n4732 );
xor ( n4734 , n4601 , n4605 );
xor ( n4735 , n4734 , n4610 );
and ( n4736 , n4732 , n4735 );
and ( n4737 , n4730 , n4735 );
or ( n4738 , n4733 , n4736 , n4737 );
xor ( n4739 , n4537 , n4553 );
xor ( n4740 , n4739 , n4562 );
and ( n4741 , n4738 , n4740 );
xor ( n4742 , n4597 , n4613 );
xor ( n4743 , n4742 , n4616 );
and ( n4744 , n4740 , n4743 );
and ( n4745 , n4738 , n4743 );
or ( n4746 , n4741 , n4744 , n4745 );
and ( n4747 , n4728 , n4746 );
xor ( n4748 , n4455 , n4457 );
xor ( n4749 , n4748 , n4460 );
and ( n4750 , n4746 , n4749 );
and ( n4751 , n4728 , n4749 );
or ( n4752 , n4747 , n4750 , n4751 );
xor ( n4753 , n4453 , n4463 );
xor ( n4754 , n4753 , n4466 );
and ( n4755 , n4752 , n4754 );
xor ( n4756 , n4507 , n4509 );
xor ( n4757 , n4756 , n4512 );
and ( n4758 , n4754 , n4757 );
and ( n4759 , n4752 , n4757 );
or ( n4760 , n4755 , n4758 , n4759 );
xor ( n4761 , n4469 , n4515 );
xor ( n4762 , n4761 , n4518 );
and ( n4763 , n4760 , n4762 );
xor ( n4764 , n4633 , n4635 );
xor ( n4765 , n4764 , n4638 );
and ( n4766 , n4762 , n4765 );
and ( n4767 , n4760 , n4765 );
or ( n4768 , n4763 , n4766 , n4767 );
xor ( n4769 , n4521 , n4641 );
xor ( n4770 , n4769 , n4644 );
and ( n4771 , n4768 , n4770 );
xor ( n4772 , n4768 , n4770 );
xor ( n4773 , n4760 , n4762 );
xor ( n4774 , n4773 , n4765 );
xor ( n4775 , n4565 , n4575 );
xor ( n4776 , n4775 , n4578 );
xor ( n4777 , n4619 , n4621 );
xor ( n4778 , n4777 , n4624 );
and ( n4779 , n4776 , n4778 );
xor ( n4780 , n4728 , n4746 );
xor ( n4781 , n4780 , n4749 );
and ( n4782 , n4778 , n4781 );
and ( n4783 , n4776 , n4781 );
or ( n4784 , n4779 , n4782 , n4783 );
xor ( n4785 , n4581 , n4627 );
xor ( n4786 , n4785 , n4630 );
and ( n4787 , n4784 , n4786 );
xor ( n4788 , n4752 , n4754 );
xor ( n4789 , n4788 , n4757 );
and ( n4790 , n4786 , n4789 );
and ( n4791 , n4784 , n4789 );
or ( n4792 , n4787 , n4790 , n4791 );
and ( n4793 , n4774 , n4792 );
xor ( n4794 , n4774 , n4792 );
xor ( n4795 , n4784 , n4786 );
xor ( n4796 , n4795 , n4789 );
and ( n4797 , n1883 , n3530 );
and ( n4798 , n1896 , n3528 );
nor ( n4799 , n4797 , n4798 );
xnor ( n4800 , n4799 , n3292 );
and ( n4801 , n3813 , n2010 );
not ( n4802 , n4801 );
and ( n4803 , n4802 , n2020 );
and ( n4804 , n4800 , n4803 );
and ( n4805 , n1915 , n3154 );
and ( n4806 , n1883 , n3152 );
nor ( n4807 , n4805 , n4806 );
xnor ( n4808 , n4807 , n2978 );
and ( n4809 , n4804 , n4808 );
and ( n4810 , n2094 , n1950 );
and ( n4811 , n2065 , n1948 );
nor ( n4812 , n4810 , n4811 );
xnor ( n4813 , n4812 , n1958 );
and ( n4814 , n4808 , n4813 );
and ( n4815 , n4804 , n4813 );
or ( n4816 , n4809 , n4814 , n4815 );
xor ( n4817 , n4541 , n4545 );
xor ( n4818 , n4817 , n4550 );
and ( n4819 , n4816 , n4818 );
xor ( n4820 , n4702 , n4714 );
xor ( n4821 , n4820 , n4719 );
and ( n4822 , n4818 , n4821 );
and ( n4823 , n4816 , n4821 );
or ( n4824 , n4819 , n4822 , n4823 );
and ( n4825 , n2004 , n2872 );
and ( n4826 , n2015 , n2870 );
nor ( n4827 , n4825 , n4826 );
xnor ( n4828 , n4827 , n2811 );
and ( n4829 , n2401 , n2054 );
and ( n4830 , n1924 , n2052 );
nor ( n4831 , n4829 , n4830 );
xnor ( n4832 , n4831 , n2062 );
and ( n4833 , n4828 , n4832 );
and ( n4834 , n2639 , n1972 );
and ( n4835 , n2556 , n1970 );
nor ( n4836 , n4834 , n4835 );
xnor ( n4837 , n4836 , n1980 );
and ( n4838 , n4832 , n4837 );
and ( n4839 , n4828 , n4837 );
or ( n4840 , n4833 , n4838 , n4839 );
and ( n4841 , n2024 , n2612 );
and ( n4842 , n2035 , n2610 );
nor ( n4843 , n4841 , n4842 );
xnor ( n4844 , n4843 , n2515 );
and ( n4845 , n3061 , n1993 );
and ( n4846 , n2919 , n1991 );
nor ( n4847 , n4845 , n4846 );
xnor ( n4848 , n4847 , n2001 );
and ( n4849 , n4844 , n4848 );
and ( n4850 , n3333 , n1893 );
and ( n4851 , n3222 , n1891 );
nor ( n4852 , n4850 , n4851 );
xnor ( n4853 , n4852 , n1901 );
and ( n4854 , n4848 , n4853 );
and ( n4855 , n4844 , n4853 );
or ( n4856 , n4849 , n4854 , n4855 );
and ( n4857 , n4840 , n4856 );
and ( n4858 , n1987 , n3803 );
and ( n4859 , n1996 , n3800 );
nor ( n4860 , n4858 , n4859 );
xnor ( n4861 , n4860 , n3289 );
and ( n4862 , n2065 , n2391 );
and ( n4863 , n2076 , n2389 );
nor ( n4864 , n4862 , n4863 );
xnor ( n4865 , n4864 , n1939 );
and ( n4866 , n4861 , n4865 );
and ( n4867 , n3522 , n1912 );
and ( n4868 , n3281 , n1910 );
nor ( n4869 , n4867 , n4868 );
xnor ( n4870 , n4869 , n1920 );
and ( n4871 , n4865 , n4870 );
and ( n4872 , n4861 , n4870 );
or ( n4873 , n4866 , n4871 , n4872 );
and ( n4874 , n4856 , n4873 );
and ( n4875 , n4840 , n4873 );
or ( n4876 , n4857 , n4874 , n4875 );
and ( n4877 , n1904 , n3154 );
and ( n4878 , n1915 , n3152 );
nor ( n4879 , n4877 , n4878 );
xnor ( n4880 , n4879 , n2978 );
and ( n4881 , n2085 , n1950 );
and ( n4882 , n2094 , n1948 );
nor ( n4883 , n4881 , n4882 );
xnor ( n4884 , n4883 , n1958 );
and ( n4885 , n4880 , n4884 );
and ( n4886 , n3813 , n2012 );
and ( n4887 , n3659 , n2010 );
nor ( n4888 , n4886 , n4887 );
xnor ( n4889 , n4888 , n2020 );
and ( n4890 , n4884 , n4889 );
and ( n4891 , n4880 , n4889 );
or ( n4892 , n4885 , n4890 , n4891 );
xor ( n4893 , n4706 , n4710 );
xor ( n4894 , n4893 , n4559 );
and ( n4895 , n4892 , n4894 );
xor ( n4896 , n4686 , n4690 );
xor ( n4897 , n4896 , n4695 );
and ( n4898 , n4894 , n4897 );
and ( n4899 , n4892 , n4897 );
or ( n4900 , n4895 , n4898 , n4899 );
and ( n4901 , n4876 , n4900 );
xor ( n4902 , n4665 , n4681 );
xor ( n4903 , n4902 , n4698 );
and ( n4904 , n4900 , n4903 );
and ( n4905 , n4876 , n4903 );
or ( n4906 , n4901 , n4904 , n4905 );
and ( n4907 , n4824 , n4906 );
xor ( n4908 , n4567 , n4569 );
xor ( n4909 , n4908 , n4572 );
and ( n4910 , n4906 , n4909 );
and ( n4911 , n4824 , n4909 );
or ( n4912 , n4907 , n4910 , n4911 );
xor ( n4913 , n4653 , n4657 );
xor ( n4914 , n4913 , n4662 );
xor ( n4915 , n4669 , n4673 );
xor ( n4916 , n4915 , n4678 );
and ( n4917 , n4914 , n4916 );
xor ( n4918 , n4804 , n4808 );
xor ( n4919 , n4918 , n4813 );
and ( n4920 , n4916 , n4919 );
and ( n4921 , n4914 , n4919 );
or ( n4922 , n4917 , n4920 , n4921 );
xor ( n4923 , n4730 , n4732 );
xor ( n4924 , n4923 , n4735 );
and ( n4925 , n4922 , n4924 );
xor ( n4926 , n4816 , n4818 );
xor ( n4927 , n4926 , n4821 );
and ( n4928 , n4924 , n4927 );
and ( n4929 , n4922 , n4927 );
or ( n4930 , n4925 , n4928 , n4929 );
xor ( n4931 , n4701 , n4722 );
xor ( n4932 , n4931 , n4725 );
and ( n4933 , n4930 , n4932 );
xor ( n4934 , n4738 , n4740 );
xor ( n4935 , n4934 , n4743 );
and ( n4936 , n4932 , n4935 );
and ( n4937 , n4930 , n4935 );
or ( n4938 , n4933 , n4936 , n4937 );
and ( n4939 , n4912 , n4938 );
xor ( n4940 , n4776 , n4778 );
xor ( n4941 , n4940 , n4781 );
and ( n4942 , n4938 , n4941 );
and ( n4943 , n4912 , n4941 );
or ( n4944 , n4939 , n4942 , n4943 );
and ( n4945 , n4796 , n4944 );
xor ( n4946 , n4796 , n4944 );
xor ( n4947 , n4912 , n4938 );
xor ( n4948 , n4947 , n4941 );
xor ( n4949 , n4800 , n4803 );
and ( n4950 , n1896 , n3803 );
and ( n4951 , n1987 , n3800 );
nor ( n4952 , n4950 , n4951 );
xnor ( n4953 , n4952 , n3289 );
and ( n4954 , n3222 , n1993 );
and ( n4955 , n3061 , n1991 );
nor ( n4956 , n4954 , n4955 );
xnor ( n4957 , n4956 , n2001 );
and ( n4958 , n4953 , n4957 );
and ( n4959 , n3281 , n1893 );
and ( n4960 , n3333 , n1891 );
nor ( n4961 , n4959 , n4960 );
xnor ( n4962 , n4961 , n1901 );
and ( n4963 , n4957 , n4962 );
and ( n4964 , n4953 , n4962 );
or ( n4965 , n4958 , n4963 , n4964 );
and ( n4966 , n4949 , n4965 );
and ( n4967 , n2076 , n2612 );
and ( n4968 , n2024 , n2610 );
nor ( n4969 , n4967 , n4968 );
xnor ( n4970 , n4969 , n2515 );
and ( n4971 , n2556 , n2054 );
and ( n4972 , n2401 , n2052 );
nor ( n4973 , n4971 , n4972 );
xnor ( n4974 , n4973 , n2062 );
and ( n4975 , n4970 , n4974 );
and ( n4976 , n2919 , n1972 );
and ( n4977 , n2639 , n1970 );
nor ( n4978 , n4976 , n4977 );
xnor ( n4979 , n4978 , n1980 );
and ( n4980 , n4974 , n4979 );
and ( n4981 , n4970 , n4979 );
or ( n4982 , n4975 , n4980 , n4981 );
and ( n4983 , n4965 , n4982 );
and ( n4984 , n4949 , n4982 );
or ( n4985 , n4966 , n4983 , n4984 );
xor ( n4986 , n4828 , n4832 );
xor ( n4987 , n4986 , n4837 );
xor ( n4988 , n4844 , n4848 );
xor ( n4989 , n4988 , n4853 );
and ( n4990 , n4987 , n4989 );
xor ( n4991 , n4861 , n4865 );
xor ( n4992 , n4991 , n4870 );
and ( n4993 , n4989 , n4992 );
and ( n4994 , n4987 , n4992 );
or ( n4995 , n4990 , n4993 , n4994 );
and ( n4996 , n4985 , n4995 );
and ( n4997 , n2015 , n3154 );
and ( n4998 , n1904 , n3152 );
nor ( n4999 , n4997 , n4998 );
xnor ( n5000 , n4999 , n2978 );
and ( n5001 , n2094 , n2391 );
and ( n5002 , n2065 , n2389 );
nor ( n5003 , n5001 , n5002 );
xnor ( n5004 , n5003 , n1939 );
and ( n5005 , n5000 , n5004 );
and ( n5006 , n3659 , n1912 );
and ( n5007 , n3522 , n1910 );
nor ( n5008 , n5006 , n5007 );
xnor ( n5009 , n5008 , n1920 );
and ( n5010 , n5004 , n5009 );
and ( n5011 , n5000 , n5009 );
or ( n5012 , n5005 , n5010 , n5011 );
and ( n5013 , n1915 , n3530 );
and ( n5014 , n1883 , n3528 );
nor ( n5015 , n5013 , n5014 );
xnor ( n5016 , n5015 , n3292 );
and ( n5017 , n2035 , n2872 );
and ( n5018 , n2004 , n2870 );
nor ( n5019 , n5017 , n5018 );
xnor ( n5020 , n5019 , n2811 );
and ( n5021 , n5016 , n5020 );
and ( n5022 , n5020 , n4801 );
and ( n5023 , n5016 , n4801 );
or ( n5024 , n5021 , n5022 , n5023 );
and ( n5025 , n5012 , n5024 );
xor ( n5026 , n4880 , n4884 );
xor ( n5027 , n5026 , n4889 );
and ( n5028 , n5024 , n5027 );
and ( n5029 , n5012 , n5027 );
or ( n5030 , n5025 , n5028 , n5029 );
and ( n5031 , n4995 , n5030 );
and ( n5032 , n4985 , n5030 );
or ( n5033 , n4996 , n5031 , n5032 );
xor ( n5034 , n4840 , n4856 );
xor ( n5035 , n5034 , n4873 );
xor ( n5036 , n4892 , n4894 );
xor ( n5037 , n5036 , n4897 );
and ( n5038 , n5035 , n5037 );
xor ( n5039 , n4914 , n4916 );
xor ( n5040 , n5039 , n4919 );
and ( n5041 , n5037 , n5040 );
and ( n5042 , n5035 , n5040 );
or ( n5043 , n5038 , n5041 , n5042 );
and ( n5044 , n5033 , n5043 );
xor ( n5045 , n4876 , n4900 );
xor ( n5046 , n5045 , n4903 );
and ( n5047 , n5043 , n5046 );
and ( n5048 , n5033 , n5046 );
or ( n5049 , n5044 , n5047 , n5048 );
xor ( n5050 , n4824 , n4906 );
xor ( n5051 , n5050 , n4909 );
and ( n5052 , n5049 , n5051 );
xor ( n5053 , n4930 , n4932 );
xor ( n5054 , n5053 , n4935 );
and ( n5055 , n5051 , n5054 );
and ( n5056 , n5049 , n5054 );
or ( n5057 , n5052 , n5055 , n5056 );
and ( n5058 , n4948 , n5057 );
xor ( n5059 , n4948 , n5057 );
xor ( n5060 , n5049 , n5051 );
xor ( n5061 , n5060 , n5054 );
and ( n5062 , n2024 , n2872 );
and ( n5063 , n2035 , n2870 );
nor ( n5064 , n5062 , n5063 );
xnor ( n5065 , n5064 , n2811 );
and ( n5066 , n2639 , n2054 );
and ( n5067 , n2556 , n2052 );
nor ( n5068 , n5066 , n5067 );
xnor ( n5069 , n5068 , n2062 );
and ( n5070 , n5065 , n5069 );
and ( n5071 , n3061 , n1972 );
and ( n5072 , n2919 , n1970 );
nor ( n5073 , n5071 , n5072 );
xnor ( n5074 , n5073 , n1980 );
and ( n5075 , n5069 , n5074 );
and ( n5076 , n5065 , n5074 );
or ( n5077 , n5070 , n5075 , n5076 );
and ( n5078 , n1883 , n3803 );
and ( n5079 , n1896 , n3800 );
nor ( n5080 , n5078 , n5079 );
xnor ( n5081 , n5080 , n3289 );
and ( n5082 , n2004 , n3154 );
and ( n5083 , n2015 , n3152 );
nor ( n5084 , n5082 , n5083 );
xnor ( n5085 , n5084 , n2978 );
and ( n5086 , n5081 , n5085 );
and ( n5087 , n3813 , n1912 );
and ( n5088 , n3659 , n1910 );
nor ( n5089 , n5087 , n5088 );
xnor ( n5090 , n5089 , n1920 );
and ( n5091 , n5085 , n5090 );
and ( n5092 , n5081 , n5090 );
or ( n5093 , n5086 , n5091 , n5092 );
and ( n5094 , n5077 , n5093 );
xor ( n5095 , n5000 , n5004 );
xor ( n5096 , n5095 , n5009 );
and ( n5097 , n5093 , n5096 );
and ( n5098 , n5077 , n5096 );
or ( n5099 , n5094 , n5097 , n5098 );
xor ( n5100 , n4949 , n4965 );
xor ( n5101 , n5100 , n4982 );
and ( n5102 , n5099 , n5101 );
xor ( n5103 , n4987 , n4989 );
xor ( n5104 , n5103 , n4992 );
and ( n5105 , n5101 , n5104 );
and ( n5106 , n5099 , n5104 );
or ( n5107 , n5102 , n5105 , n5106 );
and ( n5108 , n2065 , n2612 );
and ( n5109 , n2076 , n2610 );
nor ( n5110 , n5108 , n5109 );
xnor ( n5111 , n5110 , n2515 );
and ( n5112 , n3333 , n1993 );
and ( n5113 , n3222 , n1991 );
nor ( n5114 , n5112 , n5113 );
xnor ( n5115 , n5114 , n2001 );
and ( n5116 , n5111 , n5115 );
and ( n5117 , n3522 , n1893 );
and ( n5118 , n3281 , n1891 );
nor ( n5119 , n5117 , n5118 );
xnor ( n5120 , n5119 , n1901 );
and ( n5121 , n5115 , n5120 );
and ( n5122 , n5111 , n5120 );
or ( n5123 , n5116 , n5121 , n5122 );
and ( n5124 , n1904 , n3530 );
and ( n5125 , n1915 , n3528 );
nor ( n5126 , n5124 , n5125 );
xnor ( n5127 , n5126 , n3292 );
and ( n5128 , n3813 , n1910 );
not ( n5129 , n5128 );
and ( n5130 , n5129 , n1920 );
and ( n5131 , n5127 , n5130 );
and ( n5132 , n5123 , n5131 );
and ( n5133 , n1924 , n1950 );
and ( n5134 , n2085 , n1948 );
nor ( n5135 , n5133 , n5134 );
xnor ( n5136 , n5135 , n1958 );
and ( n5137 , n5131 , n5136 );
and ( n5138 , n5123 , n5136 );
or ( n5139 , n5132 , n5137 , n5138 );
xor ( n5140 , n4953 , n4957 );
xor ( n5141 , n5140 , n4962 );
xor ( n5142 , n5016 , n5020 );
xor ( n5143 , n5142 , n4801 );
and ( n5144 , n5141 , n5143 );
xor ( n5145 , n4970 , n4974 );
xor ( n5146 , n5145 , n4979 );
and ( n5147 , n5143 , n5146 );
and ( n5148 , n5141 , n5146 );
or ( n5149 , n5144 , n5147 , n5148 );
and ( n5150 , n5139 , n5149 );
xor ( n5151 , n5012 , n5024 );
xor ( n5152 , n5151 , n5027 );
and ( n5153 , n5149 , n5152 );
and ( n5154 , n5139 , n5152 );
or ( n5155 , n5150 , n5153 , n5154 );
and ( n5156 , n5107 , n5155 );
xor ( n5157 , n4985 , n4995 );
xor ( n5158 , n5157 , n5030 );
and ( n5159 , n5155 , n5158 );
and ( n5160 , n5107 , n5158 );
or ( n5161 , n5156 , n5159 , n5160 );
xor ( n5162 , n4922 , n4924 );
xor ( n5163 , n5162 , n4927 );
and ( n5164 , n5161 , n5163 );
xor ( n5165 , n5033 , n5043 );
xor ( n5166 , n5165 , n5046 );
and ( n5167 , n5163 , n5166 );
and ( n5168 , n5161 , n5166 );
or ( n5169 , n5164 , n5167 , n5168 );
and ( n5170 , n5061 , n5169 );
xor ( n5171 , n5061 , n5169 );
and ( n5172 , n2035 , n3154 );
and ( n5173 , n2004 , n3152 );
nor ( n5174 , n5172 , n5173 );
xnor ( n5175 , n5174 , n2978 );
and ( n5176 , n1924 , n2391 );
and ( n5177 , n2085 , n2389 );
nor ( n5178 , n5176 , n5177 );
xnor ( n5179 , n5178 , n1939 );
and ( n5180 , n5175 , n5179 );
and ( n5181 , n2556 , n1950 );
and ( n5182 , n2401 , n1948 );
nor ( n5183 , n5181 , n5182 );
xnor ( n5184 , n5183 , n1958 );
and ( n5185 , n5179 , n5184 );
and ( n5186 , n5175 , n5184 );
or ( n5187 , n5180 , n5185 , n5186 );
and ( n5188 , n1915 , n3803 );
and ( n5189 , n1883 , n3800 );
nor ( n5190 , n5188 , n5189 );
xnor ( n5191 , n5190 , n3289 );
and ( n5192 , n3281 , n1993 );
and ( n5193 , n3333 , n1991 );
nor ( n5194 , n5192 , n5193 );
xnor ( n5195 , n5194 , n2001 );
and ( n5196 , n5191 , n5195 );
and ( n5197 , n3659 , n1893 );
and ( n5198 , n3522 , n1891 );
nor ( n5199 , n5197 , n5198 );
xnor ( n5200 , n5199 , n1901 );
and ( n5201 , n5195 , n5200 );
and ( n5202 , n5191 , n5200 );
or ( n5203 , n5196 , n5201 , n5202 );
and ( n5204 , n5187 , n5203 );
and ( n5205 , n2015 , n3530 );
and ( n5206 , n1904 , n3528 );
nor ( n5207 , n5205 , n5206 );
xnor ( n5208 , n5207 , n3292 );
and ( n5209 , n2076 , n2872 );
and ( n5210 , n2024 , n2870 );
nor ( n5211 , n5209 , n5210 );
xnor ( n5212 , n5211 , n2811 );
and ( n5213 , n5208 , n5212 );
and ( n5214 , n5212 , n5128 );
and ( n5215 , n5208 , n5128 );
or ( n5216 , n5213 , n5214 , n5215 );
and ( n5217 , n5203 , n5216 );
and ( n5218 , n5187 , n5216 );
or ( n5219 , n5204 , n5217 , n5218 );
xor ( n5220 , n5127 , n5130 );
and ( n5221 , n2085 , n2391 );
and ( n5222 , n2094 , n2389 );
nor ( n5223 , n5221 , n5222 );
xnor ( n5224 , n5223 , n1939 );
and ( n5225 , n5220 , n5224 );
and ( n5226 , n2401 , n1950 );
and ( n5227 , n1924 , n1948 );
nor ( n5228 , n5226 , n5227 );
xnor ( n5229 , n5228 , n1958 );
and ( n5230 , n5224 , n5229 );
and ( n5231 , n5220 , n5229 );
or ( n5232 , n5225 , n5230 , n5231 );
and ( n5233 , n5219 , n5232 );
xor ( n5234 , n5123 , n5131 );
xor ( n5235 , n5234 , n5136 );
and ( n5236 , n5232 , n5235 );
and ( n5237 , n5219 , n5235 );
or ( n5238 , n5233 , n5236 , n5237 );
and ( n5239 , n2094 , n2612 );
and ( n5240 , n2065 , n2610 );
nor ( n5241 , n5239 , n5240 );
xnor ( n5242 , n5241 , n2515 );
and ( n5243 , n2919 , n2054 );
and ( n5244 , n2639 , n2052 );
nor ( n5245 , n5243 , n5244 );
xnor ( n5246 , n5245 , n2062 );
and ( n5247 , n5242 , n5246 );
and ( n5248 , n3222 , n1972 );
and ( n5249 , n3061 , n1970 );
nor ( n5250 , n5248 , n5249 );
xnor ( n5251 , n5250 , n1980 );
and ( n5252 , n5246 , n5251 );
and ( n5253 , n5242 , n5251 );
or ( n5254 , n5247 , n5252 , n5253 );
xor ( n5255 , n5081 , n5085 );
xor ( n5256 , n5255 , n5090 );
and ( n5257 , n5254 , n5256 );
xor ( n5258 , n5111 , n5115 );
xor ( n5259 , n5258 , n5120 );
and ( n5260 , n5256 , n5259 );
and ( n5261 , n5254 , n5259 );
or ( n5262 , n5257 , n5260 , n5261 );
xor ( n5263 , n5077 , n5093 );
xor ( n5264 , n5263 , n5096 );
and ( n5265 , n5262 , n5264 );
xor ( n5266 , n5141 , n5143 );
xor ( n5267 , n5266 , n5146 );
and ( n5268 , n5264 , n5267 );
and ( n5269 , n5262 , n5267 );
or ( n5270 , n5265 , n5268 , n5269 );
and ( n5271 , n5238 , n5270 );
xor ( n5272 , n5139 , n5149 );
xor ( n5273 , n5272 , n5152 );
and ( n5274 , n5270 , n5273 );
and ( n5275 , n5238 , n5273 );
or ( n5276 , n5271 , n5274 , n5275 );
xor ( n5277 , n5107 , n5155 );
xor ( n5278 , n5277 , n5158 );
and ( n5279 , n5276 , n5278 );
xor ( n5280 , n5035 , n5037 );
xor ( n5281 , n5280 , n5040 );
and ( n5282 , n5278 , n5281 );
and ( n5283 , n5276 , n5281 );
or ( n5284 , n5279 , n5282 , n5283 );
xor ( n5285 , n5161 , n5163 );
xor ( n5286 , n5285 , n5166 );
and ( n5287 , n5284 , n5286 );
xor ( n5288 , n5284 , n5286 );
xor ( n5289 , n5276 , n5278 );
xor ( n5290 , n5289 , n5281 );
and ( n5291 , n2085 , n2612 );
and ( n5292 , n2094 , n2610 );
nor ( n5293 , n5291 , n5292 );
xnor ( n5294 , n5293 , n2515 );
and ( n5295 , n3522 , n1993 );
and ( n5296 , n3281 , n1991 );
nor ( n5297 , n5295 , n5296 );
xnor ( n5298 , n5297 , n2001 );
and ( n5299 , n5294 , n5298 );
and ( n5300 , n3813 , n1893 );
and ( n5301 , n3659 , n1891 );
nor ( n5302 , n5300 , n5301 );
xnor ( n5303 , n5302 , n1901 );
and ( n5304 , n5298 , n5303 );
and ( n5305 , n5294 , n5303 );
or ( n5306 , n5299 , n5304 , n5305 );
and ( n5307 , n1904 , n3803 );
and ( n5308 , n1915 , n3800 );
nor ( n5309 , n5307 , n5308 );
xnor ( n5310 , n5309 , n3289 );
and ( n5311 , n2024 , n3154 );
and ( n5312 , n2035 , n3152 );
nor ( n5313 , n5311 , n5312 );
xnor ( n5314 , n5313 , n2978 );
and ( n5315 , n5310 , n5314 );
and ( n5316 , n2401 , n2391 );
and ( n5317 , n1924 , n2389 );
nor ( n5318 , n5316 , n5317 );
xnor ( n5319 , n5318 , n1939 );
and ( n5320 , n5314 , n5319 );
and ( n5321 , n5310 , n5319 );
or ( n5322 , n5315 , n5320 , n5321 );
and ( n5323 , n5306 , n5322 );
and ( n5324 , n2004 , n3530 );
and ( n5325 , n2015 , n3528 );
nor ( n5326 , n5324 , n5325 );
xnor ( n5327 , n5326 , n3292 );
and ( n5328 , n3813 , n1891 );
not ( n5329 , n5328 );
and ( n5330 , n5329 , n1901 );
and ( n5331 , n5327 , n5330 );
and ( n5332 , n5322 , n5331 );
and ( n5333 , n5306 , n5331 );
or ( n5334 , n5323 , n5332 , n5333 );
xor ( n5335 , n5065 , n5069 );
xor ( n5336 , n5335 , n5074 );
and ( n5337 , n5334 , n5336 );
xor ( n5338 , n5220 , n5224 );
xor ( n5339 , n5338 , n5229 );
and ( n5340 , n5336 , n5339 );
and ( n5341 , n5334 , n5339 );
or ( n5342 , n5337 , n5340 , n5341 );
and ( n5343 , n2065 , n2872 );
and ( n5344 , n2076 , n2870 );
nor ( n5345 , n5343 , n5344 );
xnor ( n5346 , n5345 , n2811 );
and ( n5347 , n3061 , n2054 );
and ( n5348 , n2919 , n2052 );
nor ( n5349 , n5347 , n5348 );
xnor ( n5350 , n5349 , n2062 );
and ( n5351 , n5346 , n5350 );
and ( n5352 , n3333 , n1972 );
and ( n5353 , n3222 , n1970 );
nor ( n5354 , n5352 , n5353 );
xnor ( n5355 , n5354 , n1980 );
and ( n5356 , n5350 , n5355 );
and ( n5357 , n5346 , n5355 );
or ( n5358 , n5351 , n5356 , n5357 );
xor ( n5359 , n5175 , n5179 );
xor ( n5360 , n5359 , n5184 );
and ( n5361 , n5358 , n5360 );
xor ( n5362 , n5242 , n5246 );
xor ( n5363 , n5362 , n5251 );
and ( n5364 , n5360 , n5363 );
and ( n5365 , n5358 , n5363 );
or ( n5366 , n5361 , n5364 , n5365 );
xor ( n5367 , n5187 , n5203 );
xor ( n5368 , n5367 , n5216 );
and ( n5369 , n5366 , n5368 );
xor ( n5370 , n5254 , n5256 );
xor ( n5371 , n5370 , n5259 );
and ( n5372 , n5368 , n5371 );
and ( n5373 , n5366 , n5371 );
or ( n5374 , n5369 , n5372 , n5373 );
and ( n5375 , n5342 , n5374 );
xor ( n5376 , n5219 , n5232 );
xor ( n5377 , n5376 , n5235 );
and ( n5378 , n5374 , n5377 );
and ( n5379 , n5342 , n5377 );
or ( n5380 , n5375 , n5378 , n5379 );
xor ( n5381 , n5099 , n5101 );
xor ( n5382 , n5381 , n5104 );
and ( n5383 , n5380 , n5382 );
xor ( n5384 , n5238 , n5270 );
xor ( n5385 , n5384 , n5273 );
and ( n5386 , n5382 , n5385 );
and ( n5387 , n5380 , n5385 );
or ( n5388 , n5383 , n5386 , n5387 );
and ( n5389 , n5290 , n5388 );
xor ( n5390 , n5290 , n5388 );
xor ( n5391 , n5380 , n5382 );
xor ( n5392 , n5391 , n5385 );
xor ( n5393 , n5327 , n5330 );
and ( n5394 , n2035 , n3530 );
and ( n5395 , n2004 , n3528 );
nor ( n5396 , n5394 , n5395 );
xnor ( n5397 , n5396 , n3292 );
and ( n5398 , n3222 , n2054 );
and ( n5399 , n3061 , n2052 );
nor ( n5400 , n5398 , n5399 );
xnor ( n5401 , n5400 , n2062 );
and ( n5402 , n5397 , n5401 );
and ( n5403 , n3281 , n1972 );
and ( n5404 , n3333 , n1970 );
nor ( n5405 , n5403 , n5404 );
xnor ( n5406 , n5405 , n1980 );
and ( n5407 , n5401 , n5406 );
and ( n5408 , n5397 , n5406 );
or ( n5409 , n5402 , n5407 , n5408 );
and ( n5410 , n5393 , n5409 );
and ( n5411 , n2639 , n1950 );
and ( n5412 , n2556 , n1948 );
nor ( n5413 , n5411 , n5412 );
xnor ( n5414 , n5413 , n1958 );
and ( n5415 , n5409 , n5414 );
and ( n5416 , n5393 , n5414 );
or ( n5417 , n5410 , n5415 , n5416 );
xor ( n5418 , n5191 , n5195 );
xor ( n5419 , n5418 , n5200 );
and ( n5420 , n5417 , n5419 );
xor ( n5421 , n5208 , n5212 );
xor ( n5422 , n5421 , n5128 );
and ( n5423 , n5419 , n5422 );
and ( n5424 , n5417 , n5422 );
or ( n5425 , n5420 , n5423 , n5424 );
xor ( n5426 , n5334 , n5336 );
xor ( n5427 , n5426 , n5339 );
and ( n5428 , n5425 , n5427 );
xor ( n5429 , n5366 , n5368 );
xor ( n5430 , n5429 , n5371 );
and ( n5431 , n5427 , n5430 );
and ( n5432 , n5425 , n5430 );
or ( n5433 , n5428 , n5431 , n5432 );
xor ( n5434 , n5262 , n5264 );
xor ( n5435 , n5434 , n5267 );
and ( n5436 , n5433 , n5435 );
xor ( n5437 , n5342 , n5374 );
xor ( n5438 , n5437 , n5377 );
and ( n5439 , n5435 , n5438 );
and ( n5440 , n5433 , n5438 );
or ( n5441 , n5436 , n5439 , n5440 );
and ( n5442 , n5392 , n5441 );
xor ( n5443 , n5392 , n5441 );
xor ( n5444 , n5433 , n5435 );
xor ( n5445 , n5444 , n5438 );
and ( n5446 , n2015 , n3803 );
and ( n5447 , n1904 , n3800 );
nor ( n5448 , n5446 , n5447 );
xnor ( n5449 , n5448 , n3289 );
and ( n5450 , n2094 , n2872 );
and ( n5451 , n2065 , n2870 );
nor ( n5452 , n5450 , n5451 );
xnor ( n5453 , n5452 , n2811 );
and ( n5454 , n5449 , n5453 );
and ( n5455 , n5453 , n5328 );
and ( n5456 , n5449 , n5328 );
or ( n5457 , n5454 , n5455 , n5456 );
and ( n5458 , n2076 , n3154 );
and ( n5459 , n2024 , n3152 );
nor ( n5460 , n5458 , n5459 );
xnor ( n5461 , n5460 , n2978 );
and ( n5462 , n1924 , n2612 );
and ( n5463 , n2085 , n2610 );
nor ( n5464 , n5462 , n5463 );
xnor ( n5465 , n5464 , n2515 );
and ( n5466 , n5461 , n5465 );
and ( n5467 , n3659 , n1993 );
and ( n5468 , n3522 , n1991 );
nor ( n5469 , n5467 , n5468 );
xnor ( n5470 , n5469 , n2001 );
and ( n5471 , n5465 , n5470 );
and ( n5472 , n5461 , n5470 );
or ( n5473 , n5466 , n5471 , n5472 );
and ( n5474 , n5457 , n5473 );
xor ( n5475 , n5310 , n5314 );
xor ( n5476 , n5475 , n5319 );
and ( n5477 , n5473 , n5476 );
and ( n5478 , n5457 , n5476 );
or ( n5479 , n5474 , n5477 , n5478 );
and ( n5480 , n2004 , n3803 );
and ( n5481 , n2015 , n3800 );
nor ( n5482 , n5480 , n5481 );
xnor ( n5483 , n5482 , n3289 );
and ( n5484 , n3813 , n1991 );
not ( n5485 , n5484 );
and ( n5486 , n5485 , n2001 );
and ( n5487 , n5483 , n5486 );
and ( n5488 , n2556 , n2391 );
and ( n5489 , n2401 , n2389 );
nor ( n5490 , n5488 , n5489 );
xnor ( n5491 , n5490 , n1939 );
and ( n5492 , n5487 , n5491 );
and ( n5493 , n2919 , n1950 );
and ( n5494 , n2639 , n1948 );
nor ( n5495 , n5493 , n5494 );
xnor ( n5496 , n5495 , n1958 );
and ( n5497 , n5491 , n5496 );
and ( n5498 , n5487 , n5496 );
or ( n5499 , n5492 , n5497 , n5498 );
xor ( n5500 , n5346 , n5350 );
xor ( n5501 , n5500 , n5355 );
and ( n5502 , n5499 , n5501 );
xor ( n5503 , n5294 , n5298 );
xor ( n5504 , n5503 , n5303 );
and ( n5505 , n5501 , n5504 );
and ( n5506 , n5499 , n5504 );
or ( n5507 , n5502 , n5505 , n5506 );
and ( n5508 , n5479 , n5507 );
xor ( n5509 , n5306 , n5322 );
xor ( n5510 , n5509 , n5331 );
and ( n5511 , n5507 , n5510 );
and ( n5512 , n5479 , n5510 );
or ( n5513 , n5508 , n5511 , n5512 );
and ( n5514 , n2024 , n3530 );
and ( n5515 , n2035 , n3528 );
nor ( n5516 , n5514 , n5515 );
xnor ( n5517 , n5516 , n3292 );
and ( n5518 , n2401 , n2612 );
and ( n5519 , n1924 , n2610 );
nor ( n5520 , n5518 , n5519 );
xnor ( n5521 , n5520 , n2515 );
and ( n5522 , n5517 , n5521 );
and ( n5523 , n3813 , n1993 );
and ( n5524 , n3659 , n1991 );
nor ( n5525 , n5523 , n5524 );
xnor ( n5526 , n5525 , n2001 );
and ( n5527 , n5521 , n5526 );
and ( n5528 , n5517 , n5526 );
or ( n5529 , n5522 , n5527 , n5528 );
and ( n5530 , n2065 , n3154 );
and ( n5531 , n2076 , n3152 );
nor ( n5532 , n5530 , n5531 );
xnor ( n5533 , n5532 , n2978 );
and ( n5534 , n2639 , n2391 );
and ( n5535 , n2556 , n2389 );
nor ( n5536 , n5534 , n5535 );
xnor ( n5537 , n5536 , n1939 );
and ( n5538 , n5533 , n5537 );
and ( n5539 , n3061 , n1950 );
and ( n5540 , n2919 , n1948 );
nor ( n5541 , n5539 , n5540 );
xnor ( n5542 , n5541 , n1958 );
and ( n5543 , n5537 , n5542 );
and ( n5544 , n5533 , n5542 );
or ( n5545 , n5538 , n5543 , n5544 );
and ( n5546 , n5529 , n5545 );
and ( n5547 , n2085 , n2872 );
and ( n5548 , n2094 , n2870 );
nor ( n5549 , n5547 , n5548 );
xnor ( n5550 , n5549 , n2811 );
and ( n5551 , n3333 , n2054 );
and ( n5552 , n3222 , n2052 );
nor ( n5553 , n5551 , n5552 );
xnor ( n5554 , n5553 , n2062 );
and ( n5555 , n5550 , n5554 );
and ( n5556 , n3522 , n1972 );
and ( n5557 , n3281 , n1970 );
nor ( n5558 , n5556 , n5557 );
xnor ( n5559 , n5558 , n1980 );
and ( n5560 , n5554 , n5559 );
and ( n5561 , n5550 , n5559 );
or ( n5562 , n5555 , n5560 , n5561 );
and ( n5563 , n5545 , n5562 );
and ( n5564 , n5529 , n5562 );
or ( n5565 , n5546 , n5563 , n5564 );
xor ( n5566 , n5393 , n5409 );
xor ( n5567 , n5566 , n5414 );
and ( n5568 , n5565 , n5567 );
xor ( n5569 , n5457 , n5473 );
xor ( n5570 , n5569 , n5476 );
and ( n5571 , n5567 , n5570 );
and ( n5572 , n5565 , n5570 );
or ( n5573 , n5568 , n5571 , n5572 );
xor ( n5574 , n5358 , n5360 );
xor ( n5575 , n5574 , n5363 );
and ( n5576 , n5573 , n5575 );
xor ( n5577 , n5417 , n5419 );
xor ( n5578 , n5577 , n5422 );
and ( n5579 , n5575 , n5578 );
and ( n5580 , n5573 , n5578 );
or ( n5581 , n5576 , n5579 , n5580 );
and ( n5582 , n5513 , n5581 );
xor ( n5583 , n5425 , n5427 );
xor ( n5584 , n5583 , n5430 );
and ( n5585 , n5581 , n5584 );
and ( n5586 , n5513 , n5584 );
or ( n5587 , n5582 , n5585 , n5586 );
and ( n5588 , n5445 , n5587 );
xor ( n5589 , n5445 , n5587 );
xor ( n5590 , n5513 , n5581 );
xor ( n5591 , n5590 , n5584 );
xor ( n5592 , n5449 , n5453 );
xor ( n5593 , n5592 , n5328 );
xor ( n5594 , n5397 , n5401 );
xor ( n5595 , n5594 , n5406 );
and ( n5596 , n5593 , n5595 );
xor ( n5597 , n5461 , n5465 );
xor ( n5598 , n5597 , n5470 );
and ( n5599 , n5595 , n5598 );
and ( n5600 , n5593 , n5598 );
or ( n5601 , n5596 , n5599 , n5600 );
xor ( n5602 , n5499 , n5501 );
xor ( n5603 , n5602 , n5504 );
and ( n5604 , n5601 , n5603 );
xor ( n5605 , n5565 , n5567 );
xor ( n5606 , n5605 , n5570 );
and ( n5607 , n5603 , n5606 );
and ( n5608 , n5601 , n5606 );
or ( n5609 , n5604 , n5607 , n5608 );
xor ( n5610 , n5479 , n5507 );
xor ( n5611 , n5610 , n5510 );
and ( n5612 , n5609 , n5611 );
xor ( n5613 , n5573 , n5575 );
xor ( n5614 , n5613 , n5578 );
and ( n5615 , n5611 , n5614 );
and ( n5616 , n5609 , n5614 );
or ( n5617 , n5612 , n5615 , n5616 );
and ( n5618 , n5591 , n5617 );
xor ( n5619 , n5591 , n5617 );
xor ( n5620 , n5609 , n5611 );
xor ( n5621 , n5620 , n5614 );
xor ( n5622 , n5483 , n5486 );
and ( n5623 , n2076 , n3530 );
and ( n5624 , n2024 , n3528 );
nor ( n5625 , n5623 , n5624 );
xnor ( n5626 , n5625 , n3292 );
and ( n5627 , n3281 , n2054 );
and ( n5628 , n3333 , n2052 );
nor ( n5629 , n5627 , n5628 );
xnor ( n5630 , n5629 , n2062 );
and ( n5631 , n5626 , n5630 );
and ( n5632 , n3659 , n1972 );
and ( n5633 , n3522 , n1970 );
nor ( n5634 , n5632 , n5633 );
xnor ( n5635 , n5634 , n1980 );
and ( n5636 , n5630 , n5635 );
and ( n5637 , n5626 , n5635 );
or ( n5638 , n5631 , n5636 , n5637 );
and ( n5639 , n5622 , n5638 );
and ( n5640 , n2035 , n3803 );
and ( n5641 , n2004 , n3800 );
nor ( n5642 , n5640 , n5641 );
xnor ( n5643 , n5642 , n3289 );
and ( n5644 , n1924 , n2872 );
and ( n5645 , n2085 , n2870 );
nor ( n5646 , n5644 , n5645 );
xnor ( n5647 , n5646 , n2811 );
and ( n5648 , n5643 , n5647 );
and ( n5649 , n5647 , n5484 );
and ( n5650 , n5643 , n5484 );
or ( n5651 , n5648 , n5649 , n5650 );
and ( n5652 , n5638 , n5651 );
and ( n5653 , n5622 , n5651 );
or ( n5654 , n5639 , n5652 , n5653 );
and ( n5655 , n2094 , n3154 );
and ( n5656 , n2065 , n3152 );
nor ( n5657 , n5655 , n5656 );
xnor ( n5658 , n5657 , n2978 );
and ( n5659 , n2556 , n2612 );
and ( n5660 , n2401 , n2610 );
nor ( n5661 , n5659 , n5660 );
xnor ( n5662 , n5661 , n2515 );
and ( n5663 , n5658 , n5662 );
and ( n5664 , n2919 , n2391 );
and ( n5665 , n2639 , n2389 );
nor ( n5666 , n5664 , n5665 );
xnor ( n5667 , n5666 , n1939 );
and ( n5668 , n5662 , n5667 );
and ( n5669 , n5658 , n5667 );
or ( n5670 , n5663 , n5668 , n5669 );
xor ( n5671 , n5533 , n5537 );
xor ( n5672 , n5671 , n5542 );
and ( n5673 , n5670 , n5672 );
xor ( n5674 , n5550 , n5554 );
xor ( n5675 , n5674 , n5559 );
and ( n5676 , n5672 , n5675 );
and ( n5677 , n5670 , n5675 );
or ( n5678 , n5673 , n5676 , n5677 );
and ( n5679 , n5654 , n5678 );
xor ( n5680 , n5487 , n5491 );
xor ( n5681 , n5680 , n5496 );
and ( n5682 , n5678 , n5681 );
and ( n5683 , n5654 , n5681 );
or ( n5684 , n5679 , n5682 , n5683 );
xor ( n5685 , n5529 , n5545 );
xor ( n5686 , n5685 , n5562 );
xor ( n5687 , n5593 , n5595 );
xor ( n5688 , n5687 , n5598 );
and ( n5689 , n5686 , n5688 );
xor ( n5690 , n5654 , n5678 );
xor ( n5691 , n5690 , n5681 );
and ( n5692 , n5688 , n5691 );
and ( n5693 , n5686 , n5691 );
or ( n5694 , n5689 , n5692 , n5693 );
and ( n5695 , n5684 , n5694 );
xor ( n5696 , n5601 , n5603 );
xor ( n5697 , n5696 , n5606 );
and ( n5698 , n5694 , n5697 );
and ( n5699 , n5684 , n5697 );
or ( n5700 , n5695 , n5698 , n5699 );
and ( n5701 , n5621 , n5700 );
xor ( n5702 , n5621 , n5700 );
xor ( n5703 , n5684 , n5694 );
xor ( n5704 , n5703 , n5697 );
and ( n5705 , n2401 , n2872 );
and ( n5706 , n1924 , n2870 );
nor ( n5707 , n5705 , n5706 );
xnor ( n5708 , n5707 , n2811 );
and ( n5709 , n3522 , n2054 );
and ( n5710 , n3281 , n2052 );
nor ( n5711 , n5709 , n5710 );
xnor ( n5712 , n5711 , n2062 );
and ( n5713 , n5708 , n5712 );
and ( n5714 , n3813 , n1972 );
and ( n5715 , n3659 , n1970 );
nor ( n5716 , n5714 , n5715 );
xnor ( n5717 , n5716 , n1980 );
and ( n5718 , n5712 , n5717 );
and ( n5719 , n5708 , n5717 );
or ( n5720 , n5713 , n5718 , n5719 );
and ( n5721 , n2024 , n3803 );
and ( n5722 , n2035 , n3800 );
nor ( n5723 , n5721 , n5722 );
xnor ( n5724 , n5723 , n3289 );
and ( n5725 , n3813 , n1970 );
not ( n5726 , n5725 );
and ( n5727 , n5726 , n1980 );
and ( n5728 , n5724 , n5727 );
and ( n5729 , n5720 , n5728 );
and ( n5730 , n3222 , n1950 );
and ( n5731 , n3061 , n1948 );
nor ( n5732 , n5730 , n5731 );
xnor ( n5733 , n5732 , n1958 );
and ( n5734 , n5728 , n5733 );
and ( n5735 , n5720 , n5733 );
or ( n5736 , n5729 , n5734 , n5735 );
xor ( n5737 , n5517 , n5521 );
xor ( n5738 , n5737 , n5526 );
and ( n5739 , n5736 , n5738 );
xor ( n5740 , n5622 , n5638 );
xor ( n5741 , n5740 , n5651 );
and ( n5742 , n5738 , n5741 );
and ( n5743 , n5736 , n5741 );
or ( n5744 , n5739 , n5742 , n5743 );
and ( n5745 , n2065 , n3530 );
and ( n5746 , n2076 , n3528 );
nor ( n5747 , n5745 , n5746 );
xnor ( n5748 , n5747 , n3292 );
and ( n5749 , n2085 , n3154 );
and ( n5750 , n2094 , n3152 );
nor ( n5751 , n5749 , n5750 );
xnor ( n5752 , n5751 , n2978 );
and ( n5753 , n5748 , n5752 );
and ( n5754 , n2639 , n2612 );
and ( n5755 , n2556 , n2610 );
nor ( n5756 , n5754 , n5755 );
xnor ( n5757 , n5756 , n2515 );
and ( n5758 , n5752 , n5757 );
and ( n5759 , n5748 , n5757 );
or ( n5760 , n5753 , n5758 , n5759 );
xor ( n5761 , n5658 , n5662 );
xor ( n5762 , n5761 , n5667 );
and ( n5763 , n5760 , n5762 );
xor ( n5764 , n5643 , n5647 );
xor ( n5765 , n5764 , n5484 );
and ( n5766 , n5762 , n5765 );
and ( n5767 , n5760 , n5765 );
or ( n5768 , n5763 , n5766 , n5767 );
xor ( n5769 , n5724 , n5727 );
and ( n5770 , n3061 , n2391 );
and ( n5771 , n2919 , n2389 );
nor ( n5772 , n5770 , n5771 );
xnor ( n5773 , n5772 , n1939 );
and ( n5774 , n5769 , n5773 );
and ( n5775 , n3333 , n1950 );
and ( n5776 , n3222 , n1948 );
nor ( n5777 , n5775 , n5776 );
xnor ( n5778 , n5777 , n1958 );
and ( n5779 , n5773 , n5778 );
and ( n5780 , n5769 , n5778 );
or ( n5781 , n5774 , n5779 , n5780 );
xor ( n5782 , n5626 , n5630 );
xor ( n5783 , n5782 , n5635 );
and ( n5784 , n5781 , n5783 );
xor ( n5785 , n5720 , n5728 );
xor ( n5786 , n5785 , n5733 );
and ( n5787 , n5783 , n5786 );
and ( n5788 , n5781 , n5786 );
or ( n5789 , n5784 , n5787 , n5788 );
and ( n5790 , n5768 , n5789 );
xor ( n5791 , n5670 , n5672 );
xor ( n5792 , n5791 , n5675 );
and ( n5793 , n5789 , n5792 );
and ( n5794 , n5768 , n5792 );
or ( n5795 , n5790 , n5793 , n5794 );
and ( n5796 , n5744 , n5795 );
xor ( n5797 , n5686 , n5688 );
xor ( n5798 , n5797 , n5691 );
and ( n5799 , n5795 , n5798 );
and ( n5800 , n5744 , n5798 );
or ( n5801 , n5796 , n5799 , n5800 );
and ( n5802 , n5704 , n5801 );
xor ( n5803 , n5704 , n5801 );
xor ( n5804 , n5744 , n5795 );
xor ( n5805 , n5804 , n5798 );
and ( n5806 , n1924 , n3154 );
and ( n5807 , n2085 , n3152 );
nor ( n5808 , n5806 , n5807 );
xnor ( n5809 , n5808 , n2978 );
and ( n5810 , n3222 , n2391 );
and ( n5811 , n3061 , n2389 );
nor ( n5812 , n5810 , n5811 );
xnor ( n5813 , n5812 , n1939 );
and ( n5814 , n5809 , n5813 );
and ( n5815 , n3281 , n1950 );
and ( n5816 , n3333 , n1948 );
nor ( n5817 , n5815 , n5816 );
xnor ( n5818 , n5817 , n1958 );
and ( n5819 , n5813 , n5818 );
and ( n5820 , n5809 , n5818 );
or ( n5821 , n5814 , n5819 , n5820 );
and ( n5822 , n2076 , n3803 );
and ( n5823 , n2024 , n3800 );
nor ( n5824 , n5822 , n5823 );
xnor ( n5825 , n5824 , n3289 );
and ( n5826 , n2094 , n3530 );
and ( n5827 , n2065 , n3528 );
nor ( n5828 , n5826 , n5827 );
xnor ( n5829 , n5828 , n3292 );
and ( n5830 , n5825 , n5829 );
and ( n5831 , n5829 , n5725 );
and ( n5832 , n5825 , n5725 );
or ( n5833 , n5830 , n5831 , n5832 );
and ( n5834 , n5821 , n5833 );
and ( n5835 , n2556 , n2872 );
and ( n5836 , n2401 , n2870 );
nor ( n5837 , n5835 , n5836 );
xnor ( n5838 , n5837 , n2811 );
and ( n5839 , n2919 , n2612 );
and ( n5840 , n2639 , n2610 );
nor ( n5841 , n5839 , n5840 );
xnor ( n5842 , n5841 , n2515 );
and ( n5843 , n5838 , n5842 );
and ( n5844 , n3659 , n2054 );
and ( n5845 , n3522 , n2052 );
nor ( n5846 , n5844 , n5845 );
xnor ( n5847 , n5846 , n2062 );
and ( n5848 , n5842 , n5847 );
and ( n5849 , n5838 , n5847 );
or ( n5850 , n5843 , n5848 , n5849 );
and ( n5851 , n5833 , n5850 );
and ( n5852 , n5821 , n5850 );
or ( n5853 , n5834 , n5851 , n5852 );
xor ( n5854 , n5708 , n5712 );
xor ( n5855 , n5854 , n5717 );
xor ( n5856 , n5748 , n5752 );
xor ( n5857 , n5856 , n5757 );
and ( n5858 , n5855 , n5857 );
xor ( n5859 , n5769 , n5773 );
xor ( n5860 , n5859 , n5778 );
and ( n5861 , n5857 , n5860 );
and ( n5862 , n5855 , n5860 );
or ( n5863 , n5858 , n5861 , n5862 );
and ( n5864 , n5853 , n5863 );
xor ( n5865 , n5760 , n5762 );
xor ( n5866 , n5865 , n5765 );
and ( n5867 , n5863 , n5866 );
and ( n5868 , n5853 , n5866 );
or ( n5869 , n5864 , n5867 , n5868 );
xor ( n5870 , n5736 , n5738 );
xor ( n5871 , n5870 , n5741 );
and ( n5872 , n5869 , n5871 );
xor ( n5873 , n5768 , n5789 );
xor ( n5874 , n5873 , n5792 );
and ( n5875 , n5871 , n5874 );
and ( n5876 , n5869 , n5874 );
or ( n5877 , n5872 , n5875 , n5876 );
and ( n5878 , n5805 , n5877 );
xor ( n5879 , n5805 , n5877 );
xor ( n5880 , n5869 , n5871 );
xor ( n5881 , n5880 , n5874 );
and ( n5882 , n2401 , n3154 );
and ( n5883 , n1924 , n3152 );
nor ( n5884 , n5882 , n5883 );
xnor ( n5885 , n5884 , n2978 );
and ( n5886 , n3061 , n2612 );
and ( n5887 , n2919 , n2610 );
nor ( n5888 , n5886 , n5887 );
xnor ( n5889 , n5888 , n2515 );
and ( n5890 , n5885 , n5889 );
and ( n5891 , n3333 , n2391 );
and ( n5892 , n3222 , n2389 );
nor ( n5893 , n5891 , n5892 );
xnor ( n5894 , n5893 , n1939 );
and ( n5895 , n5889 , n5894 );
and ( n5896 , n5885 , n5894 );
or ( n5897 , n5890 , n5895 , n5896 );
and ( n5898 , n2085 , n3530 );
and ( n5899 , n2094 , n3528 );
nor ( n5900 , n5898 , n5899 );
xnor ( n5901 , n5900 , n3292 );
and ( n5902 , n2639 , n2872 );
and ( n5903 , n2556 , n2870 );
nor ( n5904 , n5902 , n5903 );
xnor ( n5905 , n5904 , n2811 );
and ( n5906 , n5901 , n5905 );
and ( n5907 , n3813 , n2054 );
and ( n5908 , n3659 , n2052 );
nor ( n5909 , n5907 , n5908 );
xnor ( n5910 , n5909 , n2062 );
and ( n5911 , n5905 , n5910 );
and ( n5912 , n5901 , n5910 );
or ( n5913 , n5906 , n5911 , n5912 );
and ( n5914 , n5897 , n5913 );
and ( n5915 , n2065 , n3803 );
and ( n5916 , n2076 , n3800 );
nor ( n5917 , n5915 , n5916 );
xnor ( n5918 , n5917 , n3289 );
and ( n5919 , n3813 , n2052 );
not ( n5920 , n5919 );
and ( n5921 , n5920 , n2062 );
and ( n5922 , n5918 , n5921 );
and ( n5923 , n5913 , n5922 );
and ( n5924 , n5897 , n5922 );
or ( n5925 , n5914 , n5923 , n5924 );
xor ( n5926 , n5809 , n5813 );
xor ( n5927 , n5926 , n5818 );
xor ( n5928 , n5825 , n5829 );
xor ( n5929 , n5928 , n5725 );
and ( n5930 , n5927 , n5929 );
xor ( n5931 , n5838 , n5842 );
xor ( n5932 , n5931 , n5847 );
and ( n5933 , n5929 , n5932 );
and ( n5934 , n5927 , n5932 );
or ( n5935 , n5930 , n5933 , n5934 );
and ( n5936 , n5925 , n5935 );
xor ( n5937 , n5821 , n5833 );
xor ( n5938 , n5937 , n5850 );
and ( n5939 , n5935 , n5938 );
and ( n5940 , n5925 , n5938 );
or ( n5941 , n5936 , n5939 , n5940 );
xor ( n5942 , n5781 , n5783 );
xor ( n5943 , n5942 , n5786 );
and ( n5944 , n5941 , n5943 );
xor ( n5945 , n5853 , n5863 );
xor ( n5946 , n5945 , n5866 );
and ( n5947 , n5943 , n5946 );
and ( n5948 , n5941 , n5946 );
or ( n5949 , n5944 , n5947 , n5948 );
and ( n5950 , n5881 , n5949 );
xor ( n5951 , n5881 , n5949 );
xor ( n5952 , n5918 , n5921 );
and ( n5953 , n2094 , n3803 );
and ( n5954 , n2065 , n3800 );
nor ( n5955 , n5953 , n5954 );
xnor ( n5956 , n5955 , n3289 );
and ( n5957 , n1924 , n3530 );
and ( n5958 , n2085 , n3528 );
nor ( n5959 , n5957 , n5958 );
xnor ( n5960 , n5959 , n3292 );
and ( n5961 , n5956 , n5960 );
and ( n5962 , n5960 , n5919 );
and ( n5963 , n5956 , n5919 );
or ( n5964 , n5961 , n5962 , n5963 );
and ( n5965 , n5952 , n5964 );
and ( n5966 , n3522 , n1950 );
and ( n5967 , n3281 , n1948 );
nor ( n5968 , n5966 , n5967 );
xnor ( n5969 , n5968 , n1958 );
and ( n5970 , n5964 , n5969 );
and ( n5971 , n5952 , n5969 );
or ( n5972 , n5965 , n5970 , n5971 );
and ( n5973 , n2556 , n3154 );
and ( n5974 , n2401 , n3152 );
nor ( n5975 , n5973 , n5974 );
xnor ( n5976 , n5975 , n2978 );
and ( n5977 , n2919 , n2872 );
and ( n5978 , n2639 , n2870 );
nor ( n5979 , n5977 , n5978 );
xnor ( n5980 , n5979 , n2811 );
and ( n5981 , n5976 , n5980 );
and ( n5982 , n3222 , n2612 );
and ( n5983 , n3061 , n2610 );
nor ( n5984 , n5982 , n5983 );
xnor ( n5985 , n5984 , n2515 );
and ( n5986 , n5980 , n5985 );
and ( n5987 , n5976 , n5985 );
or ( n5988 , n5981 , n5986 , n5987 );
xor ( n5989 , n5885 , n5889 );
xor ( n5990 , n5989 , n5894 );
and ( n5991 , n5988 , n5990 );
xor ( n5992 , n5901 , n5905 );
xor ( n5993 , n5992 , n5910 );
and ( n5994 , n5990 , n5993 );
and ( n5995 , n5988 , n5993 );
or ( n5996 , n5991 , n5994 , n5995 );
and ( n5997 , n5972 , n5996 );
xor ( n5998 , n5897 , n5913 );
xor ( n5999 , n5998 , n5922 );
and ( n6000 , n5996 , n5999 );
and ( n6001 , n5972 , n5999 );
or ( n6002 , n5997 , n6000 , n6001 );
xor ( n6003 , n5855 , n5857 );
xor ( n6004 , n6003 , n5860 );
and ( n6005 , n6002 , n6004 );
xor ( n6006 , n5925 , n5935 );
xor ( n6007 , n6006 , n5938 );
and ( n6008 , n6004 , n6007 );
and ( n6009 , n6002 , n6007 );
or ( n6010 , n6005 , n6008 , n6009 );
xor ( n6011 , n5941 , n5943 );
xor ( n6012 , n6011 , n5946 );
and ( n6013 , n6010 , n6012 );
xor ( n6014 , n6010 , n6012 );
xor ( n6015 , n6002 , n6004 );
xor ( n6016 , n6015 , n6007 );
and ( n6017 , n2085 , n3803 );
and ( n6018 , n2094 , n3800 );
nor ( n6019 , n6017 , n6018 );
xnor ( n6020 , n6019 , n3289 );
and ( n6021 , n3813 , n1948 );
not ( n6022 , n6021 );
and ( n6023 , n6022 , n1958 );
and ( n6024 , n6020 , n6023 );
and ( n6025 , n3281 , n2391 );
and ( n6026 , n3333 , n2389 );
nor ( n6027 , n6025 , n6026 );
xnor ( n6028 , n6027 , n1939 );
and ( n6029 , n6024 , n6028 );
and ( n6030 , n3659 , n1950 );
and ( n6031 , n3522 , n1948 );
nor ( n6032 , n6030 , n6031 );
xnor ( n6033 , n6032 , n1958 );
and ( n6034 , n6028 , n6033 );
and ( n6035 , n6024 , n6033 );
or ( n6036 , n6029 , n6034 , n6035 );
and ( n6037 , n2639 , n3154 );
and ( n6038 , n2556 , n3152 );
nor ( n6039 , n6037 , n6038 );
xnor ( n6040 , n6039 , n2978 );
and ( n6041 , n3522 , n2391 );
and ( n6042 , n3281 , n2389 );
nor ( n6043 , n6041 , n6042 );
xnor ( n6044 , n6043 , n1939 );
and ( n6045 , n6040 , n6044 );
and ( n6046 , n3813 , n1950 );
and ( n6047 , n3659 , n1948 );
nor ( n6048 , n6046 , n6047 );
xnor ( n6049 , n6048 , n1958 );
and ( n6050 , n6044 , n6049 );
and ( n6051 , n6040 , n6049 );
or ( n6052 , n6045 , n6050 , n6051 );
and ( n6053 , n2401 , n3530 );
and ( n6054 , n1924 , n3528 );
nor ( n6055 , n6053 , n6054 );
xnor ( n6056 , n6055 , n3292 );
and ( n6057 , n3061 , n2872 );
and ( n6058 , n2919 , n2870 );
nor ( n6059 , n6057 , n6058 );
xnor ( n6060 , n6059 , n2811 );
and ( n6061 , n6056 , n6060 );
and ( n6062 , n3333 , n2612 );
and ( n6063 , n3222 , n2610 );
nor ( n6064 , n6062 , n6063 );
xnor ( n6065 , n6064 , n2515 );
and ( n6066 , n6060 , n6065 );
and ( n6067 , n6056 , n6065 );
or ( n6068 , n6061 , n6066 , n6067 );
and ( n6069 , n6052 , n6068 );
xor ( n6070 , n5956 , n5960 );
xor ( n6071 , n6070 , n5919 );
and ( n6072 , n6068 , n6071 );
and ( n6073 , n6052 , n6071 );
or ( n6074 , n6069 , n6072 , n6073 );
and ( n6075 , n6036 , n6074 );
xor ( n6076 , n5952 , n5964 );
xor ( n6077 , n6076 , n5969 );
and ( n6078 , n6074 , n6077 );
and ( n6079 , n6036 , n6077 );
or ( n6080 , n6075 , n6078 , n6079 );
xor ( n6081 , n5927 , n5929 );
xor ( n6082 , n6081 , n5932 );
and ( n6083 , n6080 , n6082 );
xor ( n6084 , n5972 , n5996 );
xor ( n6085 , n6084 , n5999 );
and ( n6086 , n6082 , n6085 );
and ( n6087 , n6080 , n6085 );
or ( n6088 , n6083 , n6086 , n6087 );
and ( n6089 , n6016 , n6088 );
xor ( n6090 , n6016 , n6088 );
xor ( n6091 , n6080 , n6082 );
xor ( n6092 , n6091 , n6085 );
xor ( n6093 , n6020 , n6023 );
and ( n6094 , n1924 , n3803 );
and ( n6095 , n2085 , n3800 );
nor ( n6096 , n6094 , n6095 );
xnor ( n6097 , n6096 , n3289 );
and ( n6098 , n3281 , n2612 );
and ( n6099 , n3333 , n2610 );
nor ( n6100 , n6098 , n6099 );
xnor ( n6101 , n6100 , n2515 );
and ( n6102 , n6097 , n6101 );
and ( n6103 , n3659 , n2391 );
and ( n6104 , n3522 , n2389 );
nor ( n6105 , n6103 , n6104 );
xnor ( n6106 , n6105 , n1939 );
and ( n6107 , n6101 , n6106 );
and ( n6108 , n6097 , n6106 );
or ( n6109 , n6102 , n6107 , n6108 );
and ( n6110 , n6093 , n6109 );
and ( n6111 , n2556 , n3530 );
and ( n6112 , n2401 , n3528 );
nor ( n6113 , n6111 , n6112 );
xnor ( n6114 , n6113 , n3292 );
and ( n6115 , n3222 , n2872 );
and ( n6116 , n3061 , n2870 );
nor ( n6117 , n6115 , n6116 );
xnor ( n6118 , n6117 , n2811 );
and ( n6119 , n6114 , n6118 );
and ( n6120 , n6118 , n6021 );
and ( n6121 , n6114 , n6021 );
or ( n6122 , n6119 , n6120 , n6121 );
and ( n6123 , n6109 , n6122 );
and ( n6124 , n6093 , n6122 );
or ( n6125 , n6110 , n6123 , n6124 );
xor ( n6126 , n5976 , n5980 );
xor ( n6127 , n6126 , n5985 );
and ( n6128 , n6125 , n6127 );
xor ( n6129 , n6024 , n6028 );
xor ( n6130 , n6129 , n6033 );
and ( n6131 , n6127 , n6130 );
and ( n6132 , n6125 , n6130 );
or ( n6133 , n6128 , n6131 , n6132 );
xor ( n6134 , n5988 , n5990 );
xor ( n6135 , n6134 , n5993 );
and ( n6136 , n6133 , n6135 );
xor ( n6137 , n6036 , n6074 );
xor ( n6138 , n6137 , n6077 );
and ( n6139 , n6135 , n6138 );
and ( n6140 , n6133 , n6138 );
or ( n6141 , n6136 , n6139 , n6140 );
and ( n6142 , n6092 , n6141 );
xor ( n6143 , n6092 , n6141 );
xor ( n6144 , n6133 , n6135 );
xor ( n6145 , n6144 , n6138 );
and ( n6146 , n2401 , n3803 );
and ( n6147 , n1924 , n3800 );
nor ( n6148 , n6146 , n6147 );
xnor ( n6149 , n6148 , n3289 );
and ( n6150 , n3333 , n2872 );
and ( n6151 , n3222 , n2870 );
nor ( n6152 , n6150 , n6151 );
xnor ( n6153 , n6152 , n2811 );
and ( n6154 , n6149 , n6153 );
and ( n6155 , n3522 , n2612 );
and ( n6156 , n3281 , n2610 );
nor ( n6157 , n6155 , n6156 );
xnor ( n6158 , n6157 , n2515 );
and ( n6159 , n6153 , n6158 );
and ( n6160 , n6149 , n6158 );
or ( n6161 , n6154 , n6159 , n6160 );
and ( n6162 , n2639 , n3530 );
and ( n6163 , n2556 , n3528 );
nor ( n6164 , n6162 , n6163 );
xnor ( n6165 , n6164 , n3292 );
and ( n6166 , n3813 , n2389 );
not ( n6167 , n6166 );
and ( n6168 , n6167 , n1939 );
and ( n6169 , n6165 , n6168 );
and ( n6170 , n6161 , n6169 );
and ( n6171 , n2919 , n3154 );
and ( n6172 , n2639 , n3152 );
nor ( n6173 , n6171 , n6172 );
xnor ( n6174 , n6173 , n2978 );
and ( n6175 , n6169 , n6174 );
and ( n6176 , n6161 , n6174 );
or ( n6177 , n6170 , n6175 , n6176 );
xor ( n6178 , n6040 , n6044 );
xor ( n6179 , n6178 , n6049 );
and ( n6180 , n6177 , n6179 );
xor ( n6181 , n6056 , n6060 );
xor ( n6182 , n6181 , n6065 );
and ( n6183 , n6179 , n6182 );
and ( n6184 , n6177 , n6182 );
or ( n6185 , n6180 , n6183 , n6184 );
xor ( n6186 , n6052 , n6068 );
xor ( n6187 , n6186 , n6071 );
and ( n6188 , n6185 , n6187 );
xor ( n6189 , n6125 , n6127 );
xor ( n6190 , n6189 , n6130 );
and ( n6191 , n6187 , n6190 );
and ( n6192 , n6185 , n6190 );
or ( n6193 , n6188 , n6191 , n6192 );
and ( n6194 , n6145 , n6193 );
xor ( n6195 , n6145 , n6193 );
xor ( n6196 , n6185 , n6187 );
xor ( n6197 , n6196 , n6190 );
xor ( n6198 , n6165 , n6168 );
and ( n6199 , n3061 , n3154 );
and ( n6200 , n2919 , n3152 );
nor ( n6201 , n6199 , n6200 );
xnor ( n6202 , n6201 , n2978 );
and ( n6203 , n6198 , n6202 );
and ( n6204 , n3813 , n2391 );
and ( n6205 , n3659 , n2389 );
nor ( n6206 , n6204 , n6205 );
xnor ( n6207 , n6206 , n1939 );
and ( n6208 , n6202 , n6207 );
and ( n6209 , n6198 , n6207 );
or ( n6210 , n6203 , n6208 , n6209 );
xor ( n6211 , n6097 , n6101 );
xor ( n6212 , n6211 , n6106 );
and ( n6213 , n6210 , n6212 );
xor ( n6214 , n6114 , n6118 );
xor ( n6215 , n6214 , n6021 );
and ( n6216 , n6212 , n6215 );
and ( n6217 , n6210 , n6215 );
or ( n6218 , n6213 , n6216 , n6217 );
xor ( n6219 , n6093 , n6109 );
xor ( n6220 , n6219 , n6122 );
and ( n6221 , n6218 , n6220 );
xor ( n6222 , n6177 , n6179 );
xor ( n6223 , n6222 , n6182 );
and ( n6224 , n6220 , n6223 );
and ( n6225 , n6218 , n6223 );
or ( n6226 , n6221 , n6224 , n6225 );
and ( n6227 , n6197 , n6226 );
xor ( n6228 , n6197 , n6226 );
xor ( n6229 , n6218 , n6220 );
xor ( n6230 , n6229 , n6223 );
and ( n6231 , n2556 , n3803 );
and ( n6232 , n2401 , n3800 );
nor ( n6233 , n6231 , n6232 );
xnor ( n6234 , n6233 , n3289 );
and ( n6235 , n3222 , n3154 );
and ( n6236 , n3061 , n3152 );
nor ( n6237 , n6235 , n6236 );
xnor ( n6238 , n6237 , n2978 );
and ( n6239 , n6234 , n6238 );
and ( n6240 , n3659 , n2612 );
and ( n6241 , n3522 , n2610 );
nor ( n6242 , n6240 , n6241 );
xnor ( n6243 , n6242 , n2515 );
and ( n6244 , n6238 , n6243 );
and ( n6245 , n6234 , n6243 );
or ( n6246 , n6239 , n6244 , n6245 );
and ( n6247 , n2919 , n3530 );
and ( n6248 , n2639 , n3528 );
nor ( n6249 , n6247 , n6248 );
xnor ( n6250 , n6249 , n3292 );
and ( n6251 , n3281 , n2872 );
and ( n6252 , n3333 , n2870 );
nor ( n6253 , n6251 , n6252 );
xnor ( n6254 , n6253 , n2811 );
and ( n6255 , n6250 , n6254 );
and ( n6256 , n6254 , n6166 );
and ( n6257 , n6250 , n6166 );
or ( n6258 , n6255 , n6256 , n6257 );
and ( n6259 , n6246 , n6258 );
xor ( n6260 , n6149 , n6153 );
xor ( n6261 , n6260 , n6158 );
and ( n6262 , n6258 , n6261 );
and ( n6263 , n6246 , n6261 );
or ( n6264 , n6259 , n6262 , n6263 );
xor ( n6265 , n6161 , n6169 );
xor ( n6266 , n6265 , n6174 );
and ( n6267 , n6264 , n6266 );
xor ( n6268 , n6210 , n6212 );
xor ( n6269 , n6268 , n6215 );
and ( n6270 , n6266 , n6269 );
and ( n6271 , n6264 , n6269 );
or ( n6272 , n6267 , n6270 , n6271 );
and ( n6273 , n6230 , n6272 );
xor ( n6274 , n6230 , n6272 );
and ( n6275 , n2639 , n3803 );
and ( n6276 , n2556 , n3800 );
nor ( n6277 , n6275 , n6276 );
xnor ( n6278 , n6277 , n3289 );
and ( n6279 , n3522 , n2872 );
and ( n6280 , n3281 , n2870 );
nor ( n6281 , n6279 , n6280 );
xnor ( n6282 , n6281 , n2811 );
and ( n6283 , n6278 , n6282 );
and ( n6284 , n3813 , n2612 );
and ( n6285 , n3659 , n2610 );
nor ( n6286 , n6284 , n6285 );
xnor ( n6287 , n6286 , n2515 );
and ( n6288 , n6282 , n6287 );
and ( n6289 , n6278 , n6287 );
or ( n6290 , n6283 , n6288 , n6289 );
and ( n6291 , n3061 , n3530 );
and ( n6292 , n2919 , n3528 );
nor ( n6293 , n6291 , n6292 );
xnor ( n6294 , n6293 , n3292 );
and ( n6295 , n3813 , n2610 );
not ( n6296 , n6295 );
and ( n6297 , n6296 , n2515 );
and ( n6298 , n6294 , n6297 );
and ( n6299 , n6290 , n6298 );
xor ( n6300 , n6250 , n6254 );
xor ( n6301 , n6300 , n6166 );
and ( n6302 , n6298 , n6301 );
and ( n6303 , n6290 , n6301 );
or ( n6304 , n6299 , n6302 , n6303 );
xor ( n6305 , n6198 , n6202 );
xor ( n6306 , n6305 , n6207 );
and ( n6307 , n6304 , n6306 );
xor ( n6308 , n6246 , n6258 );
xor ( n6309 , n6308 , n6261 );
and ( n6310 , n6306 , n6309 );
and ( n6311 , n6304 , n6309 );
or ( n6312 , n6307 , n6310 , n6311 );
xor ( n6313 , n6264 , n6266 );
xor ( n6314 , n6313 , n6269 );
and ( n6315 , n6312 , n6314 );
xor ( n6316 , n6312 , n6314 );
xor ( n6317 , n6304 , n6306 );
xor ( n6318 , n6317 , n6309 );
xor ( n6319 , n6294 , n6297 );
and ( n6320 , n2919 , n3803 );
and ( n6321 , n2639 , n3800 );
nor ( n6322 , n6320 , n6321 );
xnor ( n6323 , n6322 , n3289 );
and ( n6324 , n3659 , n2872 );
and ( n6325 , n3522 , n2870 );
nor ( n6326 , n6324 , n6325 );
xnor ( n6327 , n6326 , n2811 );
and ( n6328 , n6323 , n6327 );
and ( n6329 , n6327 , n6295 );
and ( n6330 , n6323 , n6295 );
or ( n6331 , n6328 , n6329 , n6330 );
and ( n6332 , n6319 , n6331 );
and ( n6333 , n3333 , n3154 );
and ( n6334 , n3222 , n3152 );
nor ( n6335 , n6333 , n6334 );
xnor ( n6336 , n6335 , n2978 );
and ( n6337 , n6331 , n6336 );
and ( n6338 , n6319 , n6336 );
or ( n6339 , n6332 , n6337 , n6338 );
xor ( n6340 , n6234 , n6238 );
xor ( n6341 , n6340 , n6243 );
and ( n6342 , n6339 , n6341 );
xor ( n6343 , n6290 , n6298 );
xor ( n6344 , n6343 , n6301 );
and ( n6345 , n6341 , n6344 );
and ( n6346 , n6339 , n6344 );
or ( n6347 , n6342 , n6345 , n6346 );
and ( n6348 , n6318 , n6347 );
xor ( n6349 , n6318 , n6347 );
xor ( n6350 , n6339 , n6341 );
xor ( n6351 , n6350 , n6344 );
and ( n6352 , n3061 , n3803 );
and ( n6353 , n2919 , n3800 );
nor ( n6354 , n6352 , n6353 );
xnor ( n6355 , n6354 , n3289 );
and ( n6356 , n3813 , n2870 );
not ( n6357 , n6356 );
and ( n6358 , n6357 , n2811 );
and ( n6359 , n6355 , n6358 );
and ( n6360 , n3222 , n3530 );
and ( n6361 , n3061 , n3528 );
nor ( n6362 , n6360 , n6361 );
xnor ( n6363 , n6362 , n3292 );
and ( n6364 , n6359 , n6363 );
and ( n6365 , n3281 , n3154 );
and ( n6366 , n3333 , n3152 );
nor ( n6367 , n6365 , n6366 );
xnor ( n6368 , n6367 , n2978 );
and ( n6369 , n6363 , n6368 );
and ( n6370 , n6359 , n6368 );
or ( n6371 , n6364 , n6369 , n6370 );
xor ( n6372 , n6278 , n6282 );
xor ( n6373 , n6372 , n6287 );
and ( n6374 , n6371 , n6373 );
xor ( n6375 , n6319 , n6331 );
xor ( n6376 , n6375 , n6336 );
and ( n6377 , n6373 , n6376 );
and ( n6378 , n6371 , n6376 );
or ( n6379 , n6374 , n6377 , n6378 );
and ( n6380 , n6351 , n6379 );
xor ( n6381 , n6351 , n6379 );
xor ( n6382 , n6371 , n6373 );
xor ( n6383 , n6382 , n6376 );
and ( n6384 , n3333 , n3530 );
and ( n6385 , n3222 , n3528 );
nor ( n6386 , n6384 , n6385 );
xnor ( n6387 , n6386 , n3292 );
and ( n6388 , n3522 , n3154 );
and ( n6389 , n3281 , n3152 );
nor ( n6390 , n6388 , n6389 );
xnor ( n6391 , n6390 , n2978 );
and ( n6392 , n6387 , n6391 );
and ( n6393 , n3813 , n2872 );
and ( n6394 , n3659 , n2870 );
nor ( n6395 , n6393 , n6394 );
xnor ( n6396 , n6395 , n2811 );
and ( n6397 , n6391 , n6396 );
and ( n6398 , n6387 , n6396 );
or ( n6399 , n6392 , n6397 , n6398 );
xor ( n6400 , n6323 , n6327 );
xor ( n6401 , n6400 , n6295 );
and ( n6402 , n6399 , n6401 );
xor ( n6403 , n6359 , n6363 );
xor ( n6404 , n6403 , n6368 );
and ( n6405 , n6401 , n6404 );
and ( n6406 , n6399 , n6404 );
or ( n6407 , n6402 , n6405 , n6406 );
and ( n6408 , n6383 , n6407 );
xor ( n6409 , n6383 , n6407 );
xor ( n6410 , n6355 , n6358 );
and ( n6411 , n3222 , n3803 );
and ( n6412 , n3061 , n3800 );
nor ( n6413 , n6411 , n6412 );
xnor ( n6414 , n6413 , n3289 );
and ( n6415 , n3281 , n3530 );
and ( n6416 , n3333 , n3528 );
nor ( n6417 , n6415 , n6416 );
xnor ( n6418 , n6417 , n3292 );
and ( n6419 , n6414 , n6418 );
and ( n6420 , n6418 , n6356 );
and ( n6421 , n6414 , n6356 );
or ( n6422 , n6419 , n6420 , n6421 );
and ( n6423 , n6410 , n6422 );
xor ( n6424 , n6387 , n6391 );
xor ( n6425 , n6424 , n6396 );
and ( n6426 , n6422 , n6425 );
and ( n6427 , n6410 , n6425 );
or ( n6428 , n6423 , n6426 , n6427 );
xor ( n6429 , n6399 , n6401 );
xor ( n6430 , n6429 , n6404 );
and ( n6431 , n6428 , n6430 );
xor ( n6432 , n6428 , n6430 );
xor ( n6433 , n6410 , n6422 );
xor ( n6434 , n6433 , n6425 );
and ( n6435 , n3333 , n3803 );
and ( n6436 , n3222 , n3800 );
nor ( n6437 , n6435 , n6436 );
xnor ( n6438 , n6437 , n3289 );
and ( n6439 , n3813 , n3152 );
not ( n6440 , n6439 );
and ( n6441 , n6440 , n2978 );
and ( n6442 , n6438 , n6441 );
and ( n6443 , n3659 , n3154 );
and ( n6444 , n3522 , n3152 );
nor ( n6445 , n6443 , n6444 );
xnor ( n6446 , n6445 , n2978 );
and ( n6447 , n6442 , n6446 );
xor ( n6448 , n6414 , n6418 );
xor ( n6449 , n6448 , n6356 );
and ( n6450 , n6446 , n6449 );
and ( n6451 , n6442 , n6449 );
or ( n6452 , n6447 , n6450 , n6451 );
and ( n6453 , n6434 , n6452 );
xor ( n6454 , n6434 , n6452 );
xor ( n6455 , n6442 , n6446 );
xor ( n6456 , n6455 , n6449 );
xor ( n6457 , n6438 , n6441 );
and ( n6458 , n3522 , n3530 );
and ( n6459 , n3281 , n3528 );
nor ( n6460 , n6458 , n6459 );
xnor ( n6461 , n6460 , n3292 );
and ( n6462 , n6457 , n6461 );
and ( n6463 , n3813 , n3154 );
and ( n6464 , n3659 , n3152 );
nor ( n6465 , n6463 , n6464 );
xnor ( n6466 , n6465 , n2978 );
and ( n6467 , n6461 , n6466 );
and ( n6468 , n6457 , n6466 );
or ( n6469 , n6462 , n6467 , n6468 );
and ( n6470 , n6456 , n6469 );
xor ( n6471 , n6456 , n6469 );
and ( n6472 , n3281 , n3803 );
and ( n6473 , n3333 , n3800 );
nor ( n6474 , n6472 , n6473 );
xnor ( n6475 , n6474 , n3289 );
and ( n6476 , n3659 , n3530 );
and ( n6477 , n3522 , n3528 );
nor ( n6478 , n6476 , n6477 );
xnor ( n6479 , n6478 , n3292 );
and ( n6480 , n6475 , n6479 );
and ( n6481 , n6479 , n6439 );
and ( n6482 , n6475 , n6439 );
or ( n6483 , n6480 , n6481 , n6482 );
xor ( n6484 , n6457 , n6461 );
xor ( n6485 , n6484 , n6466 );
and ( n6486 , n6483 , n6485 );
xor ( n6487 , n6483 , n6485 );
xor ( n6488 , n6475 , n6479 );
xor ( n6489 , n6488 , n6439 );
and ( n6490 , n3522 , n3803 );
and ( n6491 , n3281 , n3800 );
nor ( n6492 , n6490 , n6491 );
xnor ( n6493 , n6492 , n3289 );
and ( n6494 , n3813 , n3528 );
not ( n6495 , n6494 );
and ( n6496 , n6495 , n3292 );
and ( n6497 , n6493 , n6496 );
and ( n6498 , n6489 , n6497 );
xor ( n6499 , n6489 , n6497 );
and ( n6500 , n3813 , n3530 );
and ( n6501 , n3659 , n3528 );
nor ( n6502 , n6500 , n6501 );
xnor ( n6503 , n6502 , n3292 );
xor ( n6504 , n6493 , n6496 );
and ( n6505 , n6503 , n6504 );
xor ( n6506 , n6503 , n6504 );
and ( n6507 , n3659 , n3803 );
and ( n6508 , n3522 , n3800 );
nor ( n6509 , n6507 , n6508 );
xnor ( n6510 , n6509 , n3289 );
and ( n6511 , n6510 , n6494 );
xor ( n6512 , n6510 , n6494 );
and ( n6513 , n3813 , n3803 );
and ( n6514 , n3659 , n3800 );
nor ( n6515 , n6513 , n6514 );
xnor ( n6516 , n6515 , n3289 );
and ( n6517 , n3813 , n3800 );
not ( n6518 , n6517 );
and ( n6519 , n6518 , n3289 );
and ( n6520 , n6516 , n6519 );
and ( n6521 , n6512 , n6520 );
or ( n6522 , n6511 , n6521 );
and ( n6523 , n6506 , n6522 );
or ( n6524 , n6505 , n6523 );
and ( n6525 , n6499 , n6524 );
or ( n6526 , n6498 , n6525 );
and ( n6527 , n6487 , n6526 );
or ( n6528 , n6486 , n6527 );
and ( n6529 , n6471 , n6528 );
or ( n6530 , n6470 , n6529 );
and ( n6531 , n6454 , n6530 );
or ( n6532 , n6453 , n6531 );
and ( n6533 , n6432 , n6532 );
or ( n6534 , n6431 , n6533 );
and ( n6535 , n6409 , n6534 );
or ( n6536 , n6408 , n6535 );
and ( n6537 , n6381 , n6536 );
or ( n6538 , n6380 , n6537 );
and ( n6539 , n6349 , n6538 );
or ( n6540 , n6348 , n6539 );
and ( n6541 , n6316 , n6540 );
or ( n6542 , n6315 , n6541 );
and ( n6543 , n6274 , n6542 );
or ( n6544 , n6273 , n6543 );
and ( n6545 , n6228 , n6544 );
or ( n6546 , n6227 , n6545 );
and ( n6547 , n6195 , n6546 );
or ( n6548 , n6194 , n6547 );
and ( n6549 , n6143 , n6548 );
or ( n6550 , n6142 , n6549 );
and ( n6551 , n6090 , n6550 );
or ( n6552 , n6089 , n6551 );
and ( n6553 , n6014 , n6552 );
or ( n6554 , n6013 , n6553 );
and ( n6555 , n5951 , n6554 );
or ( n6556 , n5950 , n6555 );
and ( n6557 , n5879 , n6556 );
or ( n6558 , n5878 , n6557 );
and ( n6559 , n5803 , n6558 );
or ( n6560 , n5802 , n6559 );
and ( n6561 , n5702 , n6560 );
or ( n6562 , n5701 , n6561 );
and ( n6563 , n5619 , n6562 );
or ( n6564 , n5618 , n6563 );
and ( n6565 , n5589 , n6564 );
or ( n6566 , n5588 , n6565 );
and ( n6567 , n5443 , n6566 );
or ( n6568 , n5442 , n6567 );
and ( n6569 , n5390 , n6568 );
or ( n6570 , n5389 , n6569 );
and ( n6571 , n5288 , n6570 );
or ( n6572 , n5287 , n6571 );
and ( n6573 , n5171 , n6572 );
or ( n6574 , n5170 , n6573 );
and ( n6575 , n5059 , n6574 );
or ( n6576 , n5058 , n6575 );
and ( n6577 , n4946 , n6576 );
or ( n6578 , n4945 , n6577 );
and ( n6579 , n4794 , n6578 );
or ( n6580 , n4793 , n6579 );
and ( n6581 , n4772 , n6580 );
or ( n6582 , n4771 , n6581 );
and ( n6583 , n4649 , n6582 );
or ( n6584 , n4648 , n6583 );
and ( n6585 , n4403 , n6584 );
or ( n6586 , n4402 , n6585 );
and ( n6587 , n4381 , n6586 );
or ( n6588 , n4380 , n6587 );
and ( n6589 , n4212 , n6588 );
or ( n6590 , n4211 , n6589 );
and ( n6591 , n4069 , n6590 );
or ( n6592 , n4068 , n6591 );
and ( n6593 , n3903 , n6592 );
or ( n6594 , n3902 , n6593 );
and ( n6595 , n3744 , n6594 );
or ( n6596 , n3743 , n6595 );
and ( n6597 , n3457 , n6596 );
or ( n6598 , n3456 , n6597 );
and ( n6599 , n3367 , n6598 );
or ( n6600 , n3366 , n6599 );
and ( n6601 , n3258 , n6600 );
or ( n6602 , n3257 , n6601 );
and ( n6603 , n3105 , n6602 );
or ( n6604 , n3104 , n6603 );
and ( n6605 , n2953 , n6604 );
or ( n6606 , n2952 , n6605 );
and ( n6607 , n2792 , n6606 );
or ( n6608 , n2791 , n6607 );
and ( n6609 , n2676 , n6608 );
or ( n6610 , n2675 , n6609 );
xor ( n6611 , n2455 , n6610 );
buf ( n533872 , n6611 );
buf ( n533873 , n533872 );
buf ( n6614 , n533873 );
buf ( n533875 , n1133 );
buf ( n533876 , n1106 );
xor ( n6617 , n533875 , n533876 );
buf ( n533878 , n1134 );
buf ( n533879 , n1107 );
and ( n6620 , n533878 , n533879 );
buf ( n533881 , n1135 );
buf ( n533882 , n1108 );
and ( n6623 , n533881 , n533882 );
buf ( n533884 , n1136 );
buf ( n533885 , n1109 );
and ( n6626 , n533884 , n533885 );
buf ( n533887 , n1137 );
buf ( n533888 , n1110 );
and ( n6629 , n533887 , n533888 );
buf ( n533890 , n1138 );
buf ( n533891 , n1111 );
and ( n6632 , n533890 , n533891 );
buf ( n533893 , n1139 );
buf ( n533894 , n1112 );
and ( n6635 , n533893 , n533894 );
buf ( n533896 , n1140 );
buf ( n533897 , n1113 );
and ( n6638 , n533896 , n533897 );
buf ( n533899 , n1141 );
buf ( n533900 , n1114 );
and ( n6641 , n533899 , n533900 );
buf ( n533902 , n1142 );
buf ( n533903 , n1115 );
and ( n6644 , n533902 , n533903 );
buf ( n533905 , n1143 );
buf ( n533906 , n1116 );
and ( n6647 , n533905 , n533906 );
buf ( n533908 , n1144 );
buf ( n533909 , n1117 );
and ( n6650 , n533908 , n533909 );
buf ( n533911 , n1145 );
buf ( n533912 , n1118 );
and ( n6653 , n533911 , n533912 );
buf ( n533914 , n1146 );
buf ( n533915 , n1119 );
and ( n6656 , n533914 , n533915 );
buf ( n533917 , n1147 );
buf ( n533918 , n1120 );
and ( n6659 , n533917 , n533918 );
buf ( n533920 , n1148 );
buf ( n533921 , n1121 );
and ( n6662 , n533920 , n533921 );
and ( n6663 , n533918 , n6662 );
and ( n6664 , n533917 , n6662 );
or ( n6665 , n6659 , n6663 , n6664 );
and ( n6666 , n533915 , n6665 );
and ( n6667 , n533914 , n6665 );
or ( n6668 , n6656 , n6666 , n6667 );
and ( n6669 , n533912 , n6668 );
and ( n6670 , n533911 , n6668 );
or ( n6671 , n6653 , n6669 , n6670 );
and ( n6672 , n533909 , n6671 );
and ( n6673 , n533908 , n6671 );
or ( n6674 , n6650 , n6672 , n6673 );
and ( n6675 , n533906 , n6674 );
and ( n6676 , n533905 , n6674 );
or ( n6677 , n6647 , n6675 , n6676 );
and ( n6678 , n533903 , n6677 );
and ( n6679 , n533902 , n6677 );
or ( n6680 , n6644 , n6678 , n6679 );
and ( n6681 , n533900 , n6680 );
and ( n6682 , n533899 , n6680 );
or ( n6683 , n6641 , n6681 , n6682 );
and ( n6684 , n533897 , n6683 );
and ( n6685 , n533896 , n6683 );
or ( n6686 , n6638 , n6684 , n6685 );
and ( n6687 , n533894 , n6686 );
and ( n6688 , n533893 , n6686 );
or ( n6689 , n6635 , n6687 , n6688 );
and ( n6690 , n533891 , n6689 );
and ( n6691 , n533890 , n6689 );
or ( n6692 , n6632 , n6690 , n6691 );
and ( n6693 , n533888 , n6692 );
and ( n6694 , n533887 , n6692 );
or ( n6695 , n6629 , n6693 , n6694 );
and ( n6696 , n533885 , n6695 );
and ( n6697 , n533884 , n6695 );
or ( n6698 , n6626 , n6696 , n6697 );
and ( n6699 , n533882 , n6698 );
and ( n6700 , n533881 , n6698 );
or ( n6701 , n6623 , n6699 , n6700 );
and ( n6702 , n533879 , n6701 );
and ( n6703 , n533878 , n6701 );
or ( n6704 , n6620 , n6702 , n6703 );
xor ( n6705 , n6617 , n6704 );
buf ( n533966 , n6705 );
buf ( n533967 , n533966 );
buf ( n6708 , n533967 );
xor ( n6709 , n533878 , n533879 );
xor ( n6710 , n6709 , n6701 );
buf ( n533971 , n6710 );
buf ( n533972 , n533971 );
buf ( n6713 , n533972 );
xor ( n6714 , n6708 , n6713 );
xor ( n6715 , n533881 , n533882 );
xor ( n6716 , n6715 , n6698 );
buf ( n533977 , n6716 );
buf ( n533978 , n533977 );
buf ( n6719 , n533978 );
xor ( n6720 , n6713 , n6719 );
not ( n6721 , n6720 );
and ( n6722 , n6714 , n6721 );
and ( n6723 , n6614 , n6722 );
and ( n6724 , n2334 , n2346 );
and ( n6725 , n2346 , n2385 );
and ( n6726 , n2334 , n2385 );
or ( n6727 , n6724 , n6725 , n6726 );
and ( n6728 , n2377 , n2378 );
and ( n6729 , n2378 , n2383 );
and ( n6730 , n2377 , n2383 );
or ( n6731 , n6728 , n6729 , n6730 );
and ( n6732 , n2311 , n2315 );
and ( n6733 , n2315 , n2327 );
and ( n6734 , n2311 , n2327 );
or ( n6735 , n6732 , n6733 , n6734 );
xor ( n6736 , n6731 , n6735 );
and ( n6737 , n2320 , n2324 );
and ( n6738 , n2324 , n2326 );
and ( n6739 , n2320 , n2326 );
or ( n6740 , n6737 , n6738 , n6739 );
and ( n6741 , n2348 , n2352 );
and ( n6742 , n2352 , n2357 );
and ( n6743 , n2348 , n2357 );
or ( n6744 , n6741 , n6742 , n6743 );
xor ( n6745 , n6740 , n6744 );
and ( n6746 , n2362 , n2366 );
and ( n6747 , n2366 , n2371 );
and ( n6748 , n2362 , n2371 );
or ( n6749 , n6746 , n6747 , n6748 );
xor ( n6750 , n6745 , n6749 );
xor ( n6751 , n6736 , n6750 );
xor ( n6752 , n6727 , n6751 );
and ( n6753 , n2358 , n2372 );
and ( n6754 , n2372 , n2384 );
and ( n6755 , n2358 , n2384 );
or ( n6756 , n6753 , n6754 , n6755 );
and ( n6757 , n2273 , n2306 );
and ( n6758 , n2306 , n2328 );
and ( n6759 , n2273 , n2328 );
or ( n6760 , n6757 , n6758 , n6759 );
xor ( n6761 , n6756 , n6760 );
and ( n6762 , n1996 , n1912 );
and ( n6763 , n1962 , n1910 );
nor ( n6764 , n6762 , n6763 );
xnor ( n6765 , n6764 , n1920 );
and ( n6766 , n2035 , n2091 );
and ( n6767 , n2004 , n2089 );
nor ( n6768 , n6766 , n6767 );
xnor ( n6769 , n6768 , n2099 );
xor ( n6770 , n6765 , n6769 );
and ( n6771 , n2024 , n1926 );
xor ( n6772 , n6770 , n6771 );
and ( n6773 , n2057 , n1993 );
and ( n6774 , n1942 , n1991 );
nor ( n6775 , n6773 , n6774 );
xnor ( n6776 , n6775 , n2001 );
and ( n6777 , n1975 , n1893 );
and ( n6778 , n2049 , n1891 );
nor ( n6779 , n6777 , n6778 );
xnor ( n6780 , n6779 , n1901 );
xor ( n6781 , n6776 , n6780 );
and ( n6782 , n1896 , n2012 );
and ( n6783 , n1987 , n2010 );
nor ( n6784 , n6782 , n6783 );
xnor ( n6785 , n6784 , n2020 );
xor ( n6786 , n6781 , n6785 );
xor ( n6787 , n6772 , n6786 );
and ( n6788 , n1953 , n1972 );
not ( n6789 , n6788 );
xnor ( n6790 , n6789 , n1980 );
not ( n6791 , n6790 );
and ( n6792 , n1915 , n2032 );
and ( n6793 , n1883 , n2030 );
nor ( n6794 , n6792 , n6793 );
xnor ( n6795 , n6794 , n2040 );
xor ( n6796 , n6791 , n6795 );
and ( n6797 , n2015 , n2073 );
and ( n6798 , n1904 , n2071 );
nor ( n6799 , n6797 , n6798 );
xnor ( n6800 , n6799 , n2081 );
xor ( n6801 , n6796 , n6800 );
xor ( n6802 , n6787 , n6801 );
xor ( n6803 , n6761 , n6802 );
xor ( n6804 , n6752 , n6803 );
and ( n6805 , n2257 , n2329 );
and ( n6806 , n2329 , n2386 );
and ( n6807 , n2257 , n2386 );
or ( n6808 , n6805 , n6806 , n6807 );
xor ( n6809 , n6804 , n6808 );
and ( n6810 , n2387 , n2454 );
and ( n6811 , n2455 , n6610 );
or ( n6812 , n6810 , n6811 );
xor ( n6813 , n6809 , n6812 );
buf ( n534074 , n6813 );
buf ( n534075 , n534074 );
buf ( n6816 , n534075 );
and ( n6817 , n6816 , n6720 );
nor ( n6818 , n6723 , n6817 );
and ( n6819 , n6713 , n6719 );
not ( n6820 , n6819 );
and ( n6821 , n6708 , n6820 );
xnor ( n6822 , n6818 , n6821 );
xor ( n6823 , n2792 , n6606 );
buf ( n534084 , n6823 );
buf ( n534085 , n534084 );
buf ( n6826 , n534085 );
buf ( n534087 , n1131 );
buf ( n534088 , n1104 );
xor ( n6829 , n534087 , n534088 );
buf ( n534090 , n1132 );
buf ( n534091 , n1105 );
and ( n6832 , n534090 , n534091 );
and ( n6833 , n533875 , n533876 );
and ( n6834 , n533876 , n6704 );
and ( n6835 , n533875 , n6704 );
or ( n6836 , n6833 , n6834 , n6835 );
and ( n6837 , n534091 , n6836 );
and ( n6838 , n534090 , n6836 );
or ( n6839 , n6832 , n6837 , n6838 );
xor ( n6840 , n6829 , n6839 );
buf ( n534101 , n6840 );
buf ( n534102 , n534101 );
buf ( n6843 , n534102 );
xor ( n6844 , n534090 , n534091 );
xor ( n6845 , n6844 , n6836 );
buf ( n534106 , n6845 );
buf ( n534107 , n534106 );
buf ( n6848 , n534107 );
xor ( n6849 , n6843 , n6848 );
xor ( n6850 , n6848 , n6708 );
not ( n6851 , n6850 );
and ( n6852 , n6849 , n6851 );
and ( n6853 , n6826 , n6852 );
xor ( n6854 , n2676 , n6608 );
buf ( n534115 , n6854 );
buf ( n534116 , n534115 );
buf ( n6857 , n534116 );
and ( n6858 , n6857 , n6850 );
nor ( n6859 , n6853 , n6858 );
and ( n6860 , n6848 , n6708 );
not ( n6861 , n6860 );
and ( n6862 , n6843 , n6861 );
xnor ( n6863 , n6859 , n6862 );
xor ( n6864 , n6822 , n6863 );
xor ( n6865 , n3744 , n6594 );
buf ( n534126 , n6865 );
buf ( n534127 , n534126 );
buf ( n6868 , n534127 );
buf ( n534129 , n1125 );
buf ( n534130 , n1098 );
xor ( n6871 , n534129 , n534130 );
buf ( n534132 , n1126 );
buf ( n534133 , n1099 );
and ( n6874 , n534132 , n534133 );
buf ( n534135 , n1127 );
buf ( n534136 , n1100 );
and ( n6877 , n534135 , n534136 );
buf ( n534138 , n1128 );
buf ( n534139 , n1101 );
and ( n6880 , n534138 , n534139 );
buf ( n534141 , n1129 );
buf ( n534142 , n1102 );
and ( n6883 , n534141 , n534142 );
buf ( n534144 , n1130 );
buf ( n534145 , n1103 );
and ( n6886 , n534144 , n534145 );
and ( n6887 , n534087 , n534088 );
and ( n6888 , n534088 , n6839 );
and ( n6889 , n534087 , n6839 );
or ( n6890 , n6887 , n6888 , n6889 );
and ( n6891 , n534145 , n6890 );
and ( n6892 , n534144 , n6890 );
or ( n6893 , n6886 , n6891 , n6892 );
and ( n6894 , n534142 , n6893 );
and ( n6895 , n534141 , n6893 );
or ( n6896 , n6883 , n6894 , n6895 );
and ( n6897 , n534139 , n6896 );
and ( n6898 , n534138 , n6896 );
or ( n6899 , n6880 , n6897 , n6898 );
and ( n6900 , n534136 , n6899 );
and ( n6901 , n534135 , n6899 );
or ( n6902 , n6877 , n6900 , n6901 );
and ( n6903 , n534133 , n6902 );
and ( n6904 , n534132 , n6902 );
or ( n6905 , n6874 , n6903 , n6904 );
xor ( n6906 , n6871 , n6905 );
buf ( n534167 , n6906 );
buf ( n534168 , n534167 );
buf ( n6909 , n534168 );
xor ( n6910 , n534132 , n534133 );
xor ( n6911 , n6910 , n6902 );
buf ( n534172 , n6911 );
buf ( n534173 , n534172 );
buf ( n6914 , n534173 );
xor ( n6915 , n6909 , n6914 );
xor ( n6916 , n534135 , n534136 );
xor ( n6917 , n6916 , n6899 );
buf ( n534178 , n6917 );
buf ( n534179 , n534178 );
buf ( n6920 , n534179 );
xor ( n6921 , n6914 , n6920 );
not ( n6922 , n6921 );
and ( n6923 , n6915 , n6922 );
and ( n6924 , n6868 , n6923 );
xor ( n6925 , n3457 , n6596 );
buf ( n534186 , n6925 );
buf ( n534187 , n534186 );
buf ( n6928 , n534187 );
and ( n6929 , n6928 , n6921 );
nor ( n6930 , n6924 , n6929 );
and ( n6931 , n6914 , n6920 );
not ( n6932 , n6931 );
and ( n6933 , n6909 , n6932 );
xnor ( n6934 , n6930 , n6933 );
xor ( n6935 , n6864 , n6934 );
and ( n6936 , n6756 , n6760 );
and ( n6937 , n6760 , n6802 );
and ( n6938 , n6756 , n6802 );
or ( n6939 , n6936 , n6937 , n6938 );
and ( n6940 , n6740 , n6744 );
and ( n6941 , n6744 , n6749 );
and ( n6942 , n6740 , n6749 );
or ( n6943 , n6940 , n6941 , n6942 );
and ( n6944 , n6791 , n6795 );
and ( n6945 , n6795 , n6800 );
and ( n6946 , n6791 , n6800 );
or ( n6947 , n6944 , n6945 , n6946 );
xor ( n6948 , n6943 , n6947 );
and ( n6949 , n6765 , n6769 );
and ( n6950 , n6769 , n6771 );
and ( n6951 , n6765 , n6771 );
or ( n6952 , n6949 , n6950 , n6951 );
and ( n6953 , n6776 , n6780 );
and ( n6954 , n6780 , n6785 );
and ( n6955 , n6776 , n6785 );
or ( n6956 , n6953 , n6954 , n6955 );
xor ( n6957 , n6952 , n6956 );
buf ( n6958 , n6790 );
xor ( n6959 , n6957 , n6958 );
xor ( n6960 , n6948 , n6959 );
xor ( n6961 , n6939 , n6960 );
and ( n6962 , n6772 , n6786 );
and ( n6963 , n6786 , n6801 );
and ( n6964 , n6772 , n6801 );
or ( n6965 , n6962 , n6963 , n6964 );
and ( n6966 , n6731 , n6735 );
and ( n6967 , n6735 , n6750 );
and ( n6968 , n6731 , n6750 );
or ( n6969 , n6966 , n6967 , n6968 );
xor ( n6970 , n6965 , n6969 );
not ( n6971 , n1980 );
and ( n6972 , n1942 , n1993 );
and ( n6973 , n1953 , n1991 );
nor ( n6974 , n6972 , n6973 );
xnor ( n6975 , n6974 , n2001 );
xor ( n6976 , n6971 , n6975 );
and ( n6977 , n1962 , n1912 );
and ( n6978 , n1975 , n1910 );
nor ( n6979 , n6977 , n6978 );
xnor ( n6980 , n6979 , n1920 );
xor ( n6981 , n6976 , n6980 );
and ( n6982 , n2049 , n1893 );
and ( n6983 , n2057 , n1891 );
nor ( n6984 , n6982 , n6983 );
xnor ( n6985 , n6984 , n1901 );
and ( n6986 , n1883 , n2032 );
and ( n6987 , n1896 , n2030 );
nor ( n6988 , n6986 , n6987 );
xnor ( n6989 , n6988 , n2040 );
xor ( n6990 , n6985 , n6989 );
and ( n6991 , n1904 , n2073 );
and ( n6992 , n1915 , n2071 );
nor ( n6993 , n6991 , n6992 );
xnor ( n6994 , n6993 , n2081 );
xor ( n6995 , n6990 , n6994 );
xor ( n6996 , n6981 , n6995 );
and ( n6997 , n1987 , n2012 );
and ( n6998 , n1996 , n2010 );
nor ( n6999 , n6997 , n6998 );
xnor ( n7000 , n6999 , n2020 );
and ( n7001 , n2004 , n2091 );
and ( n7002 , n2015 , n2089 );
nor ( n7003 , n7001 , n7002 );
xnor ( n7004 , n7003 , n2099 );
xor ( n7005 , n7000 , n7004 );
and ( n7006 , n2035 , n1926 );
xor ( n7007 , n7005 , n7006 );
xor ( n7008 , n6996 , n7007 );
xor ( n7009 , n6970 , n7008 );
xor ( n7010 , n6961 , n7009 );
and ( n7011 , n6727 , n6751 );
and ( n7012 , n6751 , n6803 );
and ( n7013 , n6727 , n6803 );
or ( n7014 , n7011 , n7012 , n7013 );
xor ( n7015 , n7010 , n7014 );
and ( n7016 , n6804 , n6808 );
and ( n7017 , n6809 , n6812 );
or ( n7018 , n7016 , n7017 );
xor ( n7019 , n7015 , n7018 );
buf ( n534280 , n7019 );
buf ( n534281 , n534280 );
buf ( n7022 , n534281 );
xor ( n7023 , n533884 , n533885 );
xor ( n7024 , n7023 , n6695 );
buf ( n534285 , n7024 );
buf ( n534286 , n534285 );
buf ( n7027 , n534286 );
xor ( n7028 , n6719 , n7027 );
xor ( n7029 , n533887 , n533888 );
xor ( n7030 , n7029 , n6692 );
buf ( n534291 , n7030 );
buf ( n534292 , n534291 );
buf ( n7033 , n534292 );
xor ( n7034 , n7027 , n7033 );
not ( n7035 , n7034 );
and ( n7036 , n7028 , n7035 );
and ( n7037 , n7022 , n7036 );
and ( n7038 , n6943 , n6947 );
and ( n7039 , n6947 , n6959 );
and ( n7040 , n6943 , n6959 );
or ( n7041 , n7038 , n7039 , n7040 );
and ( n7042 , n6965 , n6969 );
and ( n7043 , n6969 , n7008 );
and ( n7044 , n6965 , n7008 );
or ( n7045 , n7042 , n7043 , n7044 );
xor ( n7046 , n7041 , n7045 );
and ( n7047 , n6981 , n6995 );
and ( n7048 , n6995 , n7007 );
and ( n7049 , n6981 , n7007 );
or ( n7050 , n7047 , n7048 , n7049 );
and ( n7051 , n6985 , n6989 );
and ( n7052 , n6989 , n6994 );
and ( n7053 , n6985 , n6994 );
or ( n7054 , n7051 , n7052 , n7053 );
and ( n7055 , n7000 , n7004 );
and ( n7056 , n7004 , n7006 );
and ( n7057 , n7000 , n7006 );
or ( n7058 , n7055 , n7056 , n7057 );
xor ( n7059 , n7054 , n7058 );
and ( n7060 , n1975 , n1912 );
and ( n7061 , n2049 , n1910 );
nor ( n7062 , n7060 , n7061 );
xnor ( n7063 , n7062 , n1920 );
and ( n7064 , n1896 , n2032 );
and ( n7065 , n1987 , n2030 );
nor ( n7066 , n7064 , n7065 );
xnor ( n7067 , n7066 , n2040 );
xor ( n7068 , n7063 , n7067 );
and ( n7069 , n1915 , n2073 );
and ( n7070 , n1883 , n2071 );
nor ( n7071 , n7069 , n7070 );
xnor ( n7072 , n7071 , n2081 );
xor ( n7073 , n7068 , n7072 );
xor ( n7074 , n7059 , n7073 );
xor ( n7075 , n7050 , n7074 );
and ( n7076 , n6952 , n6956 );
and ( n7077 , n6956 , n6958 );
and ( n7078 , n6952 , n6958 );
or ( n7079 , n7076 , n7077 , n7078 );
and ( n7080 , n2057 , n1893 );
and ( n7081 , n1942 , n1891 );
nor ( n7082 , n7080 , n7081 );
xnor ( n7083 , n7082 , n1901 );
and ( n7084 , n1996 , n2012 );
and ( n7085 , n1962 , n2010 );
nor ( n7086 , n7084 , n7085 );
xnor ( n7087 , n7086 , n2020 );
xor ( n7088 , n7083 , n7087 );
and ( n7089 , n2004 , n1926 );
xor ( n7090 , n7088 , n7089 );
xor ( n7091 , n7079 , n7090 );
and ( n7092 , n6971 , n6975 );
and ( n7093 , n6975 , n6980 );
and ( n7094 , n6971 , n6980 );
or ( n7095 , n7092 , n7093 , n7094 );
and ( n7096 , n1953 , n1993 );
not ( n7097 , n7096 );
xnor ( n7098 , n7097 , n2001 );
not ( n7099 , n7098 );
xor ( n7100 , n7095 , n7099 );
and ( n7101 , n2015 , n2091 );
and ( n7102 , n1904 , n2089 );
nor ( n7103 , n7101 , n7102 );
xnor ( n7104 , n7103 , n2099 );
xor ( n7105 , n7100 , n7104 );
xor ( n7106 , n7091 , n7105 );
xor ( n7107 , n7075 , n7106 );
xor ( n7108 , n7046 , n7107 );
and ( n7109 , n6939 , n6960 );
and ( n7110 , n6960 , n7009 );
and ( n7111 , n6939 , n7009 );
or ( n7112 , n7109 , n7110 , n7111 );
xor ( n7113 , n7108 , n7112 );
and ( n7114 , n7010 , n7014 );
and ( n7115 , n7015 , n7018 );
or ( n7116 , n7114 , n7115 );
xor ( n7117 , n7113 , n7116 );
buf ( n534378 , n7117 );
buf ( n534379 , n534378 );
buf ( n7120 , n534379 );
and ( n7121 , n7120 , n7034 );
nor ( n7122 , n7037 , n7121 );
and ( n7123 , n7027 , n7033 );
not ( n7124 , n7123 );
and ( n7125 , n6719 , n7124 );
xnor ( n7126 , n7122 , n7125 );
xor ( n7127 , n3367 , n6598 );
buf ( n534388 , n7127 );
buf ( n534389 , n534388 );
buf ( n7130 , n534389 );
xor ( n7131 , n534138 , n534139 );
xor ( n7132 , n7131 , n6896 );
buf ( n534393 , n7132 );
buf ( n534394 , n534393 );
buf ( n7135 , n534394 );
xor ( n7136 , n6920 , n7135 );
xor ( n7137 , n534141 , n534142 );
xor ( n7138 , n7137 , n6893 );
buf ( n534399 , n7138 );
buf ( n534400 , n534399 );
buf ( n7141 , n534400 );
xor ( n7142 , n7135 , n7141 );
not ( n7143 , n7142 );
and ( n7144 , n7136 , n7143 );
and ( n7145 , n7130 , n7144 );
xor ( n7146 , n3258 , n6600 );
buf ( n534407 , n7146 );
buf ( n534408 , n534407 );
buf ( n7149 , n534408 );
and ( n7150 , n7149 , n7142 );
nor ( n7151 , n7145 , n7150 );
and ( n7152 , n7135 , n7141 );
not ( n7153 , n7152 );
and ( n7154 , n6920 , n7153 );
xnor ( n7155 , n7151 , n7154 );
xor ( n7156 , n7126 , n7155 );
and ( n7157 , n6935 , n7156 );
not ( n7158 , n2040 );
and ( n7159 , n1942 , n2073 );
and ( n7160 , n1953 , n2071 );
nor ( n7161 , n7159 , n7160 );
xnor ( n7162 , n7161 , n2081 );
and ( n7163 , n7158 , n7162 );
and ( n7164 , n1975 , n1926 );
and ( n7165 , n7162 , n7164 );
and ( n7166 , n7158 , n7164 );
or ( n7167 , n7163 , n7165 , n7166 );
and ( n7168 , n2057 , n2073 );
and ( n7169 , n1942 , n2071 );
nor ( n7170 , n7168 , n7169 );
xnor ( n7171 , n7170 , n2081 );
and ( n7172 , n1975 , n2091 );
and ( n7173 , n2049 , n2089 );
nor ( n7174 , n7172 , n7173 );
xnor ( n7175 , n7174 , n2099 );
and ( n7176 , n7171 , n7175 );
and ( n7177 , n1962 , n1926 );
and ( n7178 , n7175 , n7177 );
and ( n7179 , n7171 , n7177 );
or ( n7180 , n7176 , n7178 , n7179 );
and ( n7181 , n1953 , n2032 );
not ( n7182 , n7181 );
xnor ( n7183 , n7182 , n2040 );
buf ( n7184 , n7183 );
and ( n7185 , n7180 , n7184 );
and ( n7186 , n2049 , n2091 );
and ( n7187 , n2057 , n2089 );
nor ( n7188 , n7186 , n7187 );
xnor ( n7189 , n7188 , n2099 );
and ( n7190 , n7184 , n7189 );
and ( n7191 , n7180 , n7189 );
or ( n7192 , n7185 , n7190 , n7191 );
xor ( n7193 , n7167 , n7192 );
and ( n7194 , n1953 , n2073 );
not ( n7195 , n7194 );
xnor ( n7196 , n7195 , n2081 );
not ( n7197 , n7196 );
and ( n7198 , n2057 , n2091 );
and ( n7199 , n1942 , n2089 );
nor ( n7200 , n7198 , n7199 );
xnor ( n7201 , n7200 , n2099 );
xor ( n7202 , n7197 , n7201 );
and ( n7203 , n2049 , n1926 );
xor ( n7204 , n7202 , n7203 );
xor ( n7205 , n7193 , n7204 );
not ( n7206 , n2020 );
and ( n7207 , n1942 , n2032 );
and ( n7208 , n1953 , n2030 );
nor ( n7209 , n7207 , n7208 );
xnor ( n7210 , n7209 , n2040 );
and ( n7211 , n7206 , n7210 );
and ( n7212 , n1962 , n2091 );
and ( n7213 , n1975 , n2089 );
nor ( n7214 , n7212 , n7213 );
xnor ( n7215 , n7214 , n2099 );
and ( n7216 , n7210 , n7215 );
and ( n7217 , n7206 , n7215 );
or ( n7218 , n7211 , n7216 , n7217 );
not ( n7219 , n7183 );
and ( n7220 , n7218 , n7219 );
xor ( n7221 , n7171 , n7175 );
xor ( n7222 , n7221 , n7177 );
and ( n7223 , n7219 , n7222 );
and ( n7224 , n7218 , n7222 );
or ( n7225 , n7220 , n7223 , n7224 );
xor ( n7226 , n7158 , n7162 );
xor ( n7227 , n7226 , n7164 );
and ( n7228 , n7225 , n7227 );
xor ( n7229 , n7180 , n7184 );
xor ( n7230 , n7229 , n7189 );
and ( n7231 , n7227 , n7230 );
and ( n7232 , n7225 , n7230 );
or ( n7233 , n7228 , n7231 , n7232 );
xor ( n7234 , n7205 , n7233 );
xor ( n7235 , n7225 , n7227 );
xor ( n7236 , n7235 , n7230 );
and ( n7237 , n2057 , n2032 );
and ( n7238 , n1942 , n2030 );
nor ( n7239 , n7237 , n7238 );
xnor ( n7240 , n7239 , n2040 );
buf ( n7241 , n7240 );
and ( n7242 , n2049 , n2073 );
and ( n7243 , n2057 , n2071 );
nor ( n7244 , n7242 , n7243 );
xnor ( n7245 , n7244 , n2081 );
and ( n7246 , n7241 , n7245 );
and ( n7247 , n1996 , n1926 );
and ( n7248 , n7245 , n7247 );
and ( n7249 , n7241 , n7247 );
or ( n7250 , n7246 , n7248 , n7249 );
and ( n7251 , n1953 , n2012 );
not ( n7252 , n7251 );
xnor ( n7253 , n7252 , n2020 );
and ( n7254 , n1996 , n2091 );
and ( n7255 , n1962 , n2089 );
nor ( n7256 , n7254 , n7255 );
xnor ( n7257 , n7256 , n2099 );
and ( n7258 , n7253 , n7257 );
and ( n7259 , n1987 , n1926 );
and ( n7260 , n7257 , n7259 );
and ( n7261 , n7253 , n7259 );
or ( n7262 , n7258 , n7260 , n7261 );
xor ( n7263 , n7206 , n7210 );
xor ( n7264 , n7263 , n7215 );
and ( n7265 , n7262 , n7264 );
xor ( n7266 , n7241 , n7245 );
xor ( n7267 , n7266 , n7247 );
and ( n7268 , n7264 , n7267 );
and ( n7269 , n7262 , n7267 );
or ( n7270 , n7265 , n7268 , n7269 );
and ( n7271 , n7250 , n7270 );
xor ( n7272 , n7218 , n7219 );
xor ( n7273 , n7272 , n7222 );
and ( n7274 , n7270 , n7273 );
and ( n7275 , n7250 , n7273 );
or ( n7276 , n7271 , n7274 , n7275 );
and ( n7277 , n7236 , n7276 );
xor ( n7278 , n7236 , n7276 );
xor ( n7279 , n7250 , n7270 );
xor ( n7280 , n7279 , n7273 );
and ( n7281 , n2049 , n2032 );
and ( n7282 , n2057 , n2030 );
nor ( n7283 , n7281 , n7282 );
xnor ( n7284 , n7283 , n2040 );
and ( n7285 , n1987 , n2091 );
and ( n7286 , n1996 , n2089 );
nor ( n7287 , n7285 , n7286 );
xnor ( n7288 , n7287 , n2099 );
and ( n7289 , n7284 , n7288 );
and ( n7290 , n1896 , n1926 );
and ( n7291 , n7288 , n7290 );
and ( n7292 , n7284 , n7290 );
or ( n7293 , n7289 , n7291 , n7292 );
not ( n7294 , n7240 );
and ( n7295 , n7293 , n7294 );
and ( n7296 , n1975 , n2073 );
and ( n7297 , n2049 , n2071 );
nor ( n7298 , n7296 , n7297 );
xnor ( n7299 , n7298 , n2081 );
and ( n7300 , n7294 , n7299 );
and ( n7301 , n7293 , n7299 );
or ( n7302 , n7295 , n7300 , n7301 );
not ( n7303 , n1920 );
and ( n7304 , n1942 , n2012 );
and ( n7305 , n1953 , n2010 );
nor ( n7306 , n7304 , n7305 );
xnor ( n7307 , n7306 , n2020 );
and ( n7308 , n7303 , n7307 );
and ( n7309 , n1962 , n2073 );
and ( n7310 , n1975 , n2071 );
nor ( n7311 , n7309 , n7310 );
xnor ( n7312 , n7311 , n2081 );
and ( n7313 , n7307 , n7312 );
and ( n7314 , n7303 , n7312 );
or ( n7315 , n7308 , n7313 , n7314 );
xor ( n7316 , n7253 , n7257 );
xor ( n7317 , n7316 , n7259 );
and ( n7318 , n7315 , n7317 );
xor ( n7319 , n7293 , n7294 );
xor ( n7320 , n7319 , n7299 );
and ( n7321 , n7317 , n7320 );
and ( n7322 , n7315 , n7320 );
or ( n7323 , n7318 , n7321 , n7322 );
and ( n7324 , n7302 , n7323 );
xor ( n7325 , n7262 , n7264 );
xor ( n7326 , n7325 , n7267 );
and ( n7327 , n7323 , n7326 );
and ( n7328 , n7302 , n7326 );
or ( n7329 , n7324 , n7327 , n7328 );
and ( n7330 , n7280 , n7329 );
xor ( n7331 , n7280 , n7329 );
and ( n7332 , n1953 , n1912 );
not ( n7333 , n7332 );
xnor ( n7334 , n7333 , n1920 );
and ( n7335 , n1996 , n2073 );
and ( n7336 , n1962 , n2071 );
nor ( n7337 , n7335 , n7336 );
xnor ( n7338 , n7337 , n2081 );
and ( n7339 , n7334 , n7338 );
and ( n7340 , n1896 , n2091 );
and ( n7341 , n1987 , n2089 );
nor ( n7342 , n7340 , n7341 );
xnor ( n7343 , n7342 , n2099 );
and ( n7344 , n7338 , n7343 );
and ( n7345 , n7334 , n7343 );
or ( n7346 , n7339 , n7344 , n7345 );
and ( n7347 , n2057 , n2012 );
and ( n7348 , n1942 , n2010 );
nor ( n7349 , n7347 , n7348 );
xnor ( n7350 , n7349 , n2020 );
buf ( n7351 , n7350 );
and ( n7352 , n7346 , n7351 );
xor ( n7353 , n7284 , n7288 );
xor ( n7354 , n7353 , n7290 );
and ( n7355 , n7351 , n7354 );
and ( n7356 , n7346 , n7354 );
or ( n7357 , n7352 , n7355 , n7356 );
not ( n7358 , n7350 );
and ( n7359 , n1975 , n2032 );
and ( n7360 , n2049 , n2030 );
nor ( n7361 , n7359 , n7360 );
xnor ( n7362 , n7361 , n2040 );
and ( n7363 , n7358 , n7362 );
and ( n7364 , n1883 , n1926 );
and ( n7365 , n7362 , n7364 );
and ( n7366 , n7358 , n7364 );
or ( n7367 , n7363 , n7365 , n7366 );
xor ( n7368 , n7303 , n7307 );
xor ( n7369 , n7368 , n7312 );
and ( n7370 , n7367 , n7369 );
xor ( n7371 , n7346 , n7351 );
xor ( n7372 , n7371 , n7354 );
and ( n7373 , n7369 , n7372 );
and ( n7374 , n7367 , n7372 );
or ( n7375 , n7370 , n7373 , n7374 );
and ( n7376 , n7357 , n7375 );
xor ( n7377 , n7315 , n7317 );
xor ( n7378 , n7377 , n7320 );
and ( n7379 , n7375 , n7378 );
and ( n7380 , n7357 , n7378 );
or ( n7381 , n7376 , n7379 , n7380 );
xor ( n7382 , n7302 , n7323 );
xor ( n7383 , n7382 , n7326 );
and ( n7384 , n7381 , n7383 );
xor ( n7385 , n7381 , n7383 );
xor ( n7386 , n7357 , n7375 );
xor ( n7387 , n7386 , n7378 );
and ( n7388 , n2049 , n2012 );
and ( n7389 , n2057 , n2010 );
nor ( n7390 , n7388 , n7389 );
xnor ( n7391 , n7390 , n2020 );
and ( n7392 , n1987 , n2073 );
and ( n7393 , n1996 , n2071 );
nor ( n7394 , n7392 , n7393 );
xnor ( n7395 , n7394 , n2081 );
and ( n7396 , n7391 , n7395 );
and ( n7397 , n1883 , n2091 );
and ( n7398 , n1896 , n2089 );
nor ( n7399 , n7397 , n7398 );
xnor ( n7400 , n7399 , n2099 );
and ( n7401 , n7395 , n7400 );
and ( n7402 , n7391 , n7400 );
or ( n7403 , n7396 , n7401 , n7402 );
not ( n7404 , n1901 );
and ( n7405 , n1942 , n1912 );
and ( n7406 , n1953 , n1910 );
nor ( n7407 , n7405 , n7406 );
xnor ( n7408 , n7407 , n1920 );
and ( n7409 , n7404 , n7408 );
and ( n7410 , n1962 , n2032 );
and ( n7411 , n1975 , n2030 );
nor ( n7412 , n7410 , n7411 );
xnor ( n7413 , n7412 , n2040 );
and ( n7414 , n7408 , n7413 );
and ( n7415 , n7404 , n7413 );
or ( n7416 , n7409 , n7414 , n7415 );
and ( n7417 , n7403 , n7416 );
xor ( n7418 , n7334 , n7338 );
xor ( n7419 , n7418 , n7343 );
and ( n7420 , n7416 , n7419 );
and ( n7421 , n7403 , n7419 );
or ( n7422 , n7417 , n7420 , n7421 );
and ( n7423 , n2057 , n1912 );
and ( n7424 , n1942 , n1910 );
nor ( n7425 , n7423 , n7424 );
xnor ( n7426 , n7425 , n1920 );
and ( n7427 , n1996 , n2032 );
and ( n7428 , n1962 , n2030 );
nor ( n7429 , n7427 , n7428 );
xnor ( n7430 , n7429 , n2040 );
and ( n7431 , n7426 , n7430 );
and ( n7432 , n1896 , n2073 );
and ( n7433 , n1987 , n2071 );
nor ( n7434 , n7432 , n7433 );
xnor ( n7435 , n7434 , n2081 );
and ( n7436 , n7430 , n7435 );
and ( n7437 , n7426 , n7435 );
or ( n7438 , n7431 , n7436 , n7437 );
and ( n7439 , n1953 , n1893 );
not ( n7440 , n7439 );
xnor ( n7441 , n7440 , n1901 );
buf ( n7442 , n7441 );
and ( n7443 , n7438 , n7442 );
and ( n7444 , n1915 , n1926 );
and ( n7445 , n7442 , n7444 );
and ( n7446 , n7438 , n7444 );
or ( n7447 , n7443 , n7445 , n7446 );
and ( n7448 , n1975 , n2012 );
and ( n7449 , n2049 , n2010 );
nor ( n7450 , n7448 , n7449 );
xnor ( n7451 , n7450 , n2020 );
and ( n7452 , n1915 , n2091 );
and ( n7453 , n1883 , n2089 );
nor ( n7454 , n7452 , n7453 );
xnor ( n7455 , n7454 , n2099 );
and ( n7456 , n7451 , n7455 );
and ( n7457 , n1904 , n1926 );
and ( n7458 , n7455 , n7457 );
and ( n7459 , n7451 , n7457 );
or ( n7460 , n7456 , n7458 , n7459 );
xor ( n7461 , n7391 , n7395 );
xor ( n7462 , n7461 , n7400 );
and ( n7463 , n7460 , n7462 );
xor ( n7464 , n7404 , n7408 );
xor ( n7465 , n7464 , n7413 );
and ( n7466 , n7462 , n7465 );
and ( n7467 , n7460 , n7465 );
or ( n7468 , n7463 , n7466 , n7467 );
and ( n7469 , n7447 , n7468 );
xor ( n7470 , n7358 , n7362 );
xor ( n7471 , n7470 , n7364 );
and ( n7472 , n7468 , n7471 );
and ( n7473 , n7447 , n7471 );
or ( n7474 , n7469 , n7472 , n7473 );
and ( n7475 , n7422 , n7474 );
xor ( n7476 , n7367 , n7369 );
xor ( n7477 , n7476 , n7372 );
and ( n7478 , n7474 , n7477 );
and ( n7479 , n7422 , n7477 );
or ( n7480 , n7475 , n7478 , n7479 );
and ( n7481 , n7387 , n7480 );
xor ( n7482 , n7387 , n7480 );
xor ( n7483 , n7422 , n7474 );
xor ( n7484 , n7483 , n7477 );
and ( n7485 , n2049 , n1912 );
and ( n7486 , n2057 , n1910 );
nor ( n7487 , n7485 , n7486 );
xnor ( n7488 , n7487 , n1920 );
and ( n7489 , n1987 , n2032 );
and ( n7490 , n1996 , n2030 );
nor ( n7491 , n7489 , n7490 );
xnor ( n7492 , n7491 , n2040 );
and ( n7493 , n7488 , n7492 );
and ( n7494 , n2015 , n1926 );
and ( n7495 , n7492 , n7494 );
and ( n7496 , n7488 , n7494 );
or ( n7497 , n7493 , n7495 , n7496 );
not ( n7498 , n2001 );
and ( n7499 , n1942 , n1893 );
and ( n7500 , n1953 , n1891 );
nor ( n7501 , n7499 , n7500 );
xnor ( n7502 , n7501 , n1901 );
and ( n7503 , n7498 , n7502 );
and ( n7504 , n1962 , n2012 );
and ( n7505 , n1975 , n2010 );
nor ( n7506 , n7504 , n7505 );
xnor ( n7507 , n7506 , n2020 );
and ( n7508 , n7502 , n7507 );
and ( n7509 , n7498 , n7507 );
or ( n7510 , n7503 , n7508 , n7509 );
and ( n7511 , n7497 , n7510 );
not ( n7512 , n7441 );
and ( n7513 , n7510 , n7512 );
and ( n7514 , n7497 , n7512 );
or ( n7515 , n7511 , n7513 , n7514 );
buf ( n7516 , n7098 );
and ( n7517 , n1883 , n2073 );
and ( n7518 , n1896 , n2071 );
nor ( n7519 , n7517 , n7518 );
xnor ( n7520 , n7519 , n2081 );
and ( n7521 , n7516 , n7520 );
and ( n7522 , n1904 , n2091 );
and ( n7523 , n1915 , n2089 );
nor ( n7524 , n7522 , n7523 );
xnor ( n7525 , n7524 , n2099 );
and ( n7526 , n7520 , n7525 );
and ( n7527 , n7516 , n7525 );
or ( n7528 , n7521 , n7526 , n7527 );
xor ( n7529 , n7451 , n7455 );
xor ( n7530 , n7529 , n7457 );
and ( n7531 , n7528 , n7530 );
xor ( n7532 , n7426 , n7430 );
xor ( n7533 , n7532 , n7435 );
and ( n7534 , n7530 , n7533 );
and ( n7535 , n7528 , n7533 );
or ( n7536 , n7531 , n7534 , n7535 );
and ( n7537 , n7515 , n7536 );
xor ( n7538 , n7438 , n7442 );
xor ( n7539 , n7538 , n7444 );
and ( n7540 , n7536 , n7539 );
and ( n7541 , n7515 , n7539 );
or ( n7542 , n7537 , n7540 , n7541 );
xor ( n7543 , n7403 , n7416 );
xor ( n7544 , n7543 , n7419 );
and ( n7545 , n7542 , n7544 );
xor ( n7546 , n7447 , n7468 );
xor ( n7547 , n7546 , n7471 );
and ( n7548 , n7544 , n7547 );
and ( n7549 , n7542 , n7547 );
or ( n7550 , n7545 , n7548 , n7549 );
and ( n7551 , n7484 , n7550 );
xor ( n7552 , n7484 , n7550 );
xor ( n7553 , n7542 , n7544 );
xor ( n7554 , n7553 , n7547 );
and ( n7555 , n7063 , n7067 );
and ( n7556 , n7067 , n7072 );
and ( n7557 , n7063 , n7072 );
or ( n7558 , n7555 , n7556 , n7557 );
and ( n7559 , n7083 , n7087 );
and ( n7560 , n7087 , n7089 );
and ( n7561 , n7083 , n7089 );
or ( n7562 , n7559 , n7560 , n7561 );
and ( n7563 , n7558 , n7562 );
xor ( n7564 , n7498 , n7502 );
xor ( n7565 , n7564 , n7507 );
and ( n7566 , n7562 , n7565 );
and ( n7567 , n7558 , n7565 );
or ( n7568 , n7563 , n7566 , n7567 );
xor ( n7569 , n7497 , n7510 );
xor ( n7570 , n7569 , n7512 );
and ( n7571 , n7568 , n7570 );
xor ( n7572 , n7528 , n7530 );
xor ( n7573 , n7572 , n7533 );
and ( n7574 , n7570 , n7573 );
and ( n7575 , n7568 , n7573 );
or ( n7576 , n7571 , n7574 , n7575 );
xor ( n7577 , n7460 , n7462 );
xor ( n7578 , n7577 , n7465 );
and ( n7579 , n7576 , n7578 );
xor ( n7580 , n7515 , n7536 );
xor ( n7581 , n7580 , n7539 );
and ( n7582 , n7578 , n7581 );
and ( n7583 , n7576 , n7581 );
or ( n7584 , n7579 , n7582 , n7583 );
and ( n7585 , n7554 , n7584 );
xor ( n7586 , n7554 , n7584 );
xor ( n7587 , n7576 , n7578 );
xor ( n7588 , n7587 , n7581 );
and ( n7589 , n7095 , n7099 );
and ( n7590 , n7099 , n7104 );
and ( n7591 , n7095 , n7104 );
or ( n7592 , n7589 , n7590 , n7591 );
xor ( n7593 , n7488 , n7492 );
xor ( n7594 , n7593 , n7494 );
and ( n7595 , n7592 , n7594 );
xor ( n7596 , n7516 , n7520 );
xor ( n7597 , n7596 , n7525 );
and ( n7598 , n7594 , n7597 );
and ( n7599 , n7592 , n7597 );
or ( n7600 , n7595 , n7598 , n7599 );
and ( n7601 , n7054 , n7058 );
and ( n7602 , n7058 , n7073 );
and ( n7603 , n7054 , n7073 );
or ( n7604 , n7601 , n7602 , n7603 );
and ( n7605 , n7079 , n7090 );
and ( n7606 , n7090 , n7105 );
and ( n7607 , n7079 , n7105 );
or ( n7608 , n7605 , n7606 , n7607 );
and ( n7609 , n7604 , n7608 );
xor ( n7610 , n7558 , n7562 );
xor ( n7611 , n7610 , n7565 );
and ( n7612 , n7608 , n7611 );
and ( n7613 , n7604 , n7611 );
or ( n7614 , n7609 , n7612 , n7613 );
and ( n7615 , n7600 , n7614 );
xor ( n7616 , n7568 , n7570 );
xor ( n7617 , n7616 , n7573 );
and ( n7618 , n7614 , n7617 );
and ( n7619 , n7600 , n7617 );
or ( n7620 , n7615 , n7618 , n7619 );
and ( n7621 , n7588 , n7620 );
xor ( n7622 , n7588 , n7620 );
and ( n7623 , n7050 , n7074 );
and ( n7624 , n7074 , n7106 );
and ( n7625 , n7050 , n7106 );
or ( n7626 , n7623 , n7624 , n7625 );
xor ( n7627 , n7592 , n7594 );
xor ( n7628 , n7627 , n7597 );
and ( n7629 , n7626 , n7628 );
xor ( n7630 , n7604 , n7608 );
xor ( n7631 , n7630 , n7611 );
and ( n7632 , n7628 , n7631 );
and ( n7633 , n7626 , n7631 );
or ( n7634 , n7629 , n7632 , n7633 );
xor ( n7635 , n7600 , n7614 );
xor ( n7636 , n7635 , n7617 );
and ( n7637 , n7634 , n7636 );
xor ( n7638 , n7634 , n7636 );
xor ( n7639 , n7626 , n7628 );
xor ( n7640 , n7639 , n7631 );
and ( n7641 , n7041 , n7045 );
and ( n7642 , n7045 , n7107 );
and ( n7643 , n7041 , n7107 );
or ( n7644 , n7641 , n7642 , n7643 );
and ( n7645 , n7640 , n7644 );
xor ( n7646 , n7640 , n7644 );
and ( n7647 , n7108 , n7112 );
and ( n7648 , n7113 , n7116 );
or ( n7649 , n7647 , n7648 );
and ( n7650 , n7646 , n7649 );
or ( n7651 , n7645 , n7650 );
and ( n7652 , n7638 , n7651 );
or ( n7653 , n7637 , n7652 );
and ( n7654 , n7622 , n7653 );
or ( n7655 , n7621 , n7654 );
and ( n7656 , n7586 , n7655 );
or ( n7657 , n7585 , n7656 );
and ( n7658 , n7552 , n7657 );
or ( n7659 , n7551 , n7658 );
and ( n7660 , n7482 , n7659 );
or ( n7661 , n7481 , n7660 );
and ( n7662 , n7385 , n7661 );
or ( n7663 , n7384 , n7662 );
and ( n7664 , n7331 , n7663 );
or ( n7665 , n7330 , n7664 );
and ( n7666 , n7278 , n7665 );
or ( n7667 , n7277 , n7666 );
xor ( n7668 , n7234 , n7667 );
buf ( n534929 , n7668 );
buf ( n534930 , n534929 );
buf ( n7671 , n534930 );
xor ( n7672 , n533917 , n533918 );
xor ( n7673 , n7672 , n6662 );
buf ( n534934 , n7673 );
buf ( n534935 , n534934 );
buf ( n7676 , n534935 );
xor ( n7677 , n533920 , n533921 );
buf ( n534938 , n7677 );
buf ( n534939 , n534938 );
buf ( n7680 , n534939 );
xor ( n7681 , n7676 , n7680 );
not ( n7682 , n7680 );
and ( n7683 , n7681 , n7682 );
and ( n7684 , n7671 , n7683 );
and ( n7685 , n7197 , n7201 );
and ( n7686 , n7201 , n7203 );
and ( n7687 , n7197 , n7203 );
or ( n7688 , n7685 , n7686 , n7687 );
buf ( n7689 , n7196 );
xor ( n7690 , n7688 , n7689 );
not ( n7691 , n2081 );
and ( n7692 , n1942 , n2091 );
and ( n7693 , n1953 , n2089 );
nor ( n7694 , n7692 , n7693 );
xnor ( n7695 , n7694 , n2099 );
xor ( n7696 , n7691 , n7695 );
and ( n7697 , n2057 , n1926 );
xor ( n7698 , n7696 , n7697 );
xor ( n7699 , n7690 , n7698 );
and ( n7700 , n7167 , n7192 );
and ( n7701 , n7192 , n7204 );
and ( n7702 , n7167 , n7204 );
or ( n7703 , n7700 , n7701 , n7702 );
xor ( n7704 , n7699 , n7703 );
and ( n7705 , n7205 , n7233 );
and ( n7706 , n7234 , n7667 );
or ( n7707 , n7705 , n7706 );
xor ( n7708 , n7704 , n7707 );
buf ( n534969 , n7708 );
buf ( n534970 , n534969 );
buf ( n7711 , n534970 );
and ( n7712 , n7711 , n7680 );
nor ( n7713 , n7684 , n7712 );
xnor ( n7714 , n7713 , n7676 );
xor ( n7715 , n7331 , n7663 );
buf ( n534976 , n7715 );
buf ( n534977 , n534976 );
buf ( n7718 , n534977 );
xor ( n7719 , n533911 , n533912 );
xor ( n7720 , n7719 , n6668 );
buf ( n534981 , n7720 );
buf ( n534982 , n534981 );
buf ( n7723 , n534982 );
xor ( n7724 , n533914 , n533915 );
xor ( n7725 , n7724 , n6665 );
buf ( n534986 , n7725 );
buf ( n534987 , n534986 );
buf ( n7728 , n534987 );
xor ( n7729 , n7723 , n7728 );
xor ( n7730 , n7728 , n7676 );
not ( n7731 , n7730 );
and ( n7732 , n7729 , n7731 );
and ( n7733 , n7718 , n7732 );
xor ( n7734 , n7278 , n7665 );
buf ( n534995 , n7734 );
buf ( n534996 , n534995 );
buf ( n7737 , n534996 );
and ( n7738 , n7737 , n7730 );
nor ( n7739 , n7733 , n7738 );
and ( n7740 , n7728 , n7676 );
not ( n7741 , n7740 );
and ( n7742 , n7723 , n7741 );
xnor ( n7743 , n7739 , n7742 );
and ( n7744 , n7714 , n7743 );
xor ( n7745 , n7482 , n7659 );
buf ( n535006 , n7745 );
buf ( n535007 , n535006 );
buf ( n7748 , n535007 );
xor ( n7749 , n533905 , n533906 );
xor ( n7750 , n7749 , n6674 );
buf ( n535011 , n7750 );
buf ( n535012 , n535011 );
buf ( n7753 , n535012 );
xor ( n7754 , n533908 , n533909 );
xor ( n7755 , n7754 , n6671 );
buf ( n535016 , n7755 );
buf ( n535017 , n535016 );
buf ( n7758 , n535017 );
xor ( n7759 , n7753 , n7758 );
xor ( n7760 , n7758 , n7723 );
not ( n7761 , n7760 );
and ( n7762 , n7759 , n7761 );
and ( n7763 , n7748 , n7762 );
xor ( n7764 , n7385 , n7661 );
buf ( n535025 , n7764 );
buf ( n535026 , n535025 );
buf ( n7767 , n535026 );
and ( n7768 , n7767 , n7760 );
nor ( n7769 , n7763 , n7768 );
and ( n7770 , n7758 , n7723 );
not ( n7771 , n7770 );
and ( n7772 , n7753 , n7771 );
xnor ( n7773 , n7769 , n7772 );
and ( n7774 , n7743 , n7773 );
and ( n7775 , n7714 , n7773 );
or ( n7776 , n7744 , n7774 , n7775 );
and ( n7777 , n7156 , n7776 );
and ( n7778 , n6935 , n7776 );
or ( n7779 , n7157 , n7777 , n7778 );
xor ( n7780 , n7586 , n7655 );
buf ( n535041 , n7780 );
buf ( n535042 , n535041 );
buf ( n7783 , n535042 );
xor ( n7784 , n533899 , n533900 );
xor ( n7785 , n7784 , n6680 );
buf ( n535046 , n7785 );
buf ( n535047 , n535046 );
buf ( n7788 , n535047 );
xor ( n7789 , n533902 , n533903 );
xor ( n7790 , n7789 , n6677 );
buf ( n535051 , n7790 );
buf ( n535052 , n535051 );
buf ( n7793 , n535052 );
xor ( n7794 , n7788 , n7793 );
xor ( n7795 , n7793 , n7753 );
not ( n7796 , n7795 );
and ( n7797 , n7794 , n7796 );
and ( n7798 , n7783 , n7797 );
xor ( n7799 , n7552 , n7657 );
buf ( n535060 , n7799 );
buf ( n535061 , n535060 );
buf ( n7802 , n535061 );
and ( n7803 , n7802 , n7795 );
nor ( n7804 , n7798 , n7803 );
and ( n7805 , n7793 , n7753 );
not ( n7806 , n7805 );
and ( n7807 , n7788 , n7806 );
xnor ( n7808 , n7804 , n7807 );
xor ( n7809 , n7638 , n7651 );
buf ( n535070 , n7809 );
buf ( n535071 , n535070 );
buf ( n7812 , n535071 );
xor ( n7813 , n533893 , n533894 );
xor ( n7814 , n7813 , n6686 );
buf ( n535075 , n7814 );
buf ( n535076 , n535075 );
buf ( n7817 , n535076 );
xor ( n7818 , n533896 , n533897 );
xor ( n7819 , n7818 , n6683 );
buf ( n535080 , n7819 );
buf ( n535081 , n535080 );
buf ( n7822 , n535081 );
xor ( n7823 , n7817 , n7822 );
xor ( n7824 , n7822 , n7788 );
not ( n7825 , n7824 );
and ( n7826 , n7823 , n7825 );
and ( n7827 , n7812 , n7826 );
xor ( n7828 , n7622 , n7653 );
buf ( n535089 , n7828 );
buf ( n535090 , n535089 );
buf ( n7831 , n535090 );
and ( n7832 , n7831 , n7824 );
nor ( n7833 , n7827 , n7832 );
and ( n7834 , n7822 , n7788 );
not ( n7835 , n7834 );
and ( n7836 , n7817 , n7835 );
xnor ( n7837 , n7833 , n7836 );
and ( n7838 , n7808 , n7837 );
xor ( n7839 , n533890 , n533891 );
xor ( n7840 , n7839 , n6689 );
buf ( n535101 , n7840 );
buf ( n535102 , n535101 );
buf ( n7843 , n535102 );
xor ( n7844 , n7033 , n7843 );
xor ( n7845 , n7843 , n7817 );
not ( n7846 , n7845 );
and ( n7847 , n7844 , n7846 );
and ( n7848 , n7120 , n7847 );
xor ( n7849 , n7646 , n7649 );
buf ( n535110 , n7849 );
buf ( n535111 , n535110 );
buf ( n7852 , n535111 );
and ( n7853 , n7852 , n7845 );
nor ( n7854 , n7848 , n7853 );
and ( n7855 , n7843 , n7817 );
not ( n7856 , n7855 );
and ( n7857 , n7033 , n7856 );
xnor ( n7858 , n7854 , n7857 );
and ( n7859 , n7837 , n7858 );
and ( n7860 , n7808 , n7858 );
or ( n7861 , n7838 , n7859 , n7860 );
and ( n7862 , n6857 , n6722 );
and ( n7863 , n6614 , n6720 );
nor ( n7864 , n7862 , n7863 );
xnor ( n7865 , n7864 , n6821 );
xor ( n7866 , n534144 , n534145 );
xor ( n7867 , n7866 , n6890 );
buf ( n535128 , n7867 );
buf ( n535129 , n535128 );
buf ( n7870 , n535129 );
xor ( n7871 , n7141 , n7870 );
xor ( n7872 , n7870 , n6843 );
not ( n7873 , n7872 );
and ( n7874 , n7871 , n7873 );
and ( n7875 , n7149 , n7874 );
xor ( n7876 , n3105 , n6602 );
buf ( n535137 , n7876 );
buf ( n535138 , n535137 );
buf ( n7879 , n535138 );
and ( n7880 , n7879 , n7872 );
nor ( n7881 , n7875 , n7880 );
and ( n7882 , n7870 , n6843 );
not ( n7883 , n7882 );
and ( n7884 , n7141 , n7883 );
xnor ( n7885 , n7881 , n7884 );
and ( n7886 , n7865 , n7885 );
and ( n7887 , n6928 , n7144 );
and ( n7888 , n7130 , n7142 );
nor ( n7889 , n7887 , n7888 );
xnor ( n7890 , n7889 , n7154 );
and ( n7891 , n7885 , n7890 );
and ( n7892 , n7865 , n7890 );
or ( n7893 , n7886 , n7891 , n7892 );
and ( n7894 , n7861 , n7893 );
xor ( n7895 , n4212 , n6588 );
buf ( n535156 , n7895 );
buf ( n535157 , n535156 );
buf ( n7898 , n535157 );
buf ( n535159 , n1123 );
buf ( n535160 , n1096 );
xor ( n7901 , n535159 , n535160 );
buf ( n535162 , n1124 );
buf ( n535163 , n1097 );
and ( n7904 , n535162 , n535163 );
and ( n7905 , n534129 , n534130 );
and ( n7906 , n534130 , n6905 );
and ( n7907 , n534129 , n6905 );
or ( n7908 , n7905 , n7906 , n7907 );
and ( n7909 , n535163 , n7908 );
and ( n7910 , n535162 , n7908 );
or ( n7911 , n7904 , n7909 , n7910 );
xor ( n7912 , n7901 , n7911 );
buf ( n535173 , n7912 );
buf ( n535174 , n535173 );
buf ( n7915 , n535174 );
xor ( n7916 , n535162 , n535163 );
xor ( n7917 , n7916 , n7908 );
buf ( n535178 , n7917 );
buf ( n535179 , n535178 );
buf ( n7920 , n535179 );
xor ( n7921 , n7915 , n7920 );
xor ( n7922 , n7920 , n6909 );
not ( n7923 , n7922 );
and ( n7924 , n7921 , n7923 );
and ( n7925 , n7898 , n7924 );
xor ( n7926 , n4069 , n6590 );
buf ( n535187 , n7926 );
buf ( n535188 , n535187 );
buf ( n7929 , n535188 );
and ( n7930 , n7929 , n7922 );
nor ( n7931 , n7925 , n7930 );
and ( n7932 , n7920 , n6909 );
not ( n7933 , n7932 );
and ( n7934 , n7915 , n7933 );
xnor ( n7935 , n7931 , n7934 );
xor ( n7936 , n4403 , n6584 );
buf ( n535197 , n7936 );
buf ( n535198 , n535197 );
buf ( n7939 , n535198 );
buf ( n535200 , n1094 );
buf ( n535201 , n1122 );
buf ( n535202 , n1095 );
and ( n7943 , n535201 , n535202 );
and ( n7944 , n535159 , n535160 );
and ( n7945 , n535160 , n7911 );
and ( n7946 , n535159 , n7911 );
or ( n7947 , n7944 , n7945 , n7946 );
and ( n7948 , n535202 , n7947 );
and ( n7949 , n535201 , n7947 );
or ( n7950 , n7943 , n7948 , n7949 );
xor ( n7951 , n535200 , n7950 );
buf ( n535212 , n7951 );
buf ( n535213 , n535212 );
buf ( n7954 , n535213 );
xor ( n7955 , n535201 , n535202 );
xor ( n7956 , n7955 , n7947 );
buf ( n535217 , n7956 );
buf ( n535218 , n535217 );
buf ( n7959 , n535218 );
xor ( n7960 , n7954 , n7959 );
xor ( n7961 , n7959 , n7915 );
not ( n7962 , n7961 );
and ( n7963 , n7960 , n7962 );
and ( n7964 , n7939 , n7963 );
xor ( n7965 , n4381 , n6586 );
buf ( n535226 , n7965 );
buf ( n535227 , n535226 );
buf ( n7968 , n535227 );
and ( n7969 , n7968 , n7961 );
nor ( n7970 , n7964 , n7969 );
and ( n7971 , n7959 , n7915 );
not ( n7972 , n7971 );
and ( n7973 , n7954 , n7972 );
xnor ( n7974 , n7970 , n7973 );
and ( n7975 , n7935 , n7974 );
xor ( n7976 , n4772 , n6580 );
buf ( n535237 , n7976 );
buf ( n535238 , n535237 );
buf ( n7979 , n535238 );
buf ( n535240 , n1092 );
buf ( n535241 , n1093 );
and ( n7982 , n535200 , n7950 );
and ( n7983 , n535241 , n7982 );
xor ( n7984 , n535240 , n7983 );
buf ( n535245 , n7984 );
buf ( n535246 , n535245 );
buf ( n7987 , n535246 );
xor ( n7988 , n535241 , n7982 );
buf ( n535249 , n7988 );
buf ( n535250 , n535249 );
buf ( n7991 , n535250 );
xor ( n7992 , n7987 , n7991 );
xor ( n7993 , n7991 , n7954 );
not ( n7994 , n7993 );
and ( n7995 , n7992 , n7994 );
and ( n7996 , n7979 , n7995 );
xor ( n7997 , n4649 , n6582 );
buf ( n535258 , n7997 );
buf ( n535259 , n535258 );
buf ( n8000 , n535259 );
and ( n8001 , n8000 , n7993 );
nor ( n8002 , n7996 , n8001 );
and ( n8003 , n7991 , n7954 );
not ( n8004 , n8003 );
and ( n8005 , n7987 , n8004 );
xnor ( n8006 , n8002 , n8005 );
and ( n8007 , n7974 , n8006 );
and ( n8008 , n7935 , n8006 );
or ( n8009 , n7975 , n8007 , n8008 );
and ( n8010 , n7893 , n8009 );
and ( n8011 , n7861 , n8009 );
or ( n8012 , n7894 , n8010 , n8011 );
xor ( n8013 , n7779 , n8012 );
and ( n8014 , n6857 , n6852 );
and ( n8015 , n6614 , n6850 );
nor ( n8016 , n8014 , n8015 );
xnor ( n8017 , n8016 , n6862 );
xor ( n8018 , n2953 , n6604 );
buf ( n535279 , n8018 );
buf ( n535280 , n535279 );
buf ( n8021 , n535280 );
and ( n8022 , n8021 , n7874 );
and ( n8023 , n6826 , n7872 );
nor ( n8024 , n8022 , n8023 );
xnor ( n8025 , n8024 , n7884 );
xor ( n8026 , n8017 , n8025 );
and ( n8027 , n7149 , n7144 );
and ( n8028 , n7879 , n7142 );
nor ( n8029 , n8027 , n8028 );
xnor ( n8030 , n8029 , n7154 );
xor ( n8031 , n8026 , n8030 );
and ( n8032 , n6928 , n6923 );
and ( n8033 , n7130 , n6921 );
nor ( n8034 , n8032 , n8033 );
xnor ( n8035 , n8034 , n6933 );
xor ( n8036 , n3903 , n6592 );
buf ( n535297 , n8036 );
buf ( n535298 , n535297 );
buf ( n8039 , n535298 );
and ( n8040 , n8039 , n7924 );
and ( n8041 , n6868 , n7922 );
nor ( n8042 , n8040 , n8041 );
xnor ( n8043 , n8042 , n7934 );
xor ( n8044 , n8035 , n8043 );
and ( n8045 , n7898 , n7963 );
and ( n8046 , n7929 , n7961 );
nor ( n8047 , n8045 , n8046 );
xnor ( n8048 , n8047 , n7973 );
xor ( n8049 , n8044 , n8048 );
xor ( n8050 , n8031 , n8049 );
and ( n8051 , n6822 , n6863 );
and ( n8052 , n6863 , n6934 );
and ( n8053 , n6822 , n6934 );
or ( n8054 , n8051 , n8052 , n8053 );
xor ( n8055 , n8050 , n8054 );
xor ( n8056 , n8013 , n8055 );
xor ( n8057 , n7861 , n7893 );
xor ( n8058 , n8057 , n8009 );
and ( n8059 , n8039 , n7144 );
and ( n8060 , n6868 , n7142 );
nor ( n8061 , n8059 , n8060 );
xnor ( n8062 , n8061 , n7154 );
and ( n8063 , n7939 , n7924 );
and ( n8064 , n7968 , n7922 );
nor ( n8065 , n8063 , n8064 );
xnor ( n8066 , n8065 , n7934 );
and ( n8067 , n8062 , n8066 );
xor ( n8068 , n4946 , n6576 );
buf ( n535329 , n8068 );
buf ( n535330 , n535329 );
buf ( n8071 , n535330 );
and ( n8072 , n8071 , n7995 );
xor ( n8073 , n4794 , n6578 );
buf ( n535334 , n8073 );
buf ( n535335 , n535334 );
buf ( n8076 , n535335 );
and ( n8077 , n8076 , n7993 );
nor ( n8078 , n8072 , n8077 );
xnor ( n8079 , n8078 , n8005 );
and ( n8080 , n8066 , n8079 );
and ( n8081 , n8062 , n8079 );
or ( n8082 , n8067 , n8080 , n8081 );
and ( n8083 , n7831 , n7797 );
and ( n8084 , n7783 , n7795 );
nor ( n8085 , n8083 , n8084 );
xnor ( n8086 , n8085 , n7807 );
and ( n8087 , n8082 , n8086 );
xor ( n8088 , n5288 , n6570 );
buf ( n535349 , n8088 );
buf ( n535350 , n535349 );
buf ( n8091 , n535350 );
buf ( n535352 , n1090 );
buf ( n535353 , n1091 );
and ( n8094 , n535240 , n7983 );
and ( n8095 , n535353 , n8094 );
and ( n8096 , n535352 , n8095 );
buf ( n535357 , n8096 );
buf ( n535358 , n535357 );
buf ( n8099 , n535358 );
xor ( n8100 , n535352 , n8095 );
buf ( n535361 , n8100 );
buf ( n535362 , n535361 );
buf ( n8103 , n535362 );
xor ( n8104 , n8099 , n8103 );
not ( n8105 , n8104 );
and ( n8106 , n8099 , n8105 );
and ( n8107 , n8091 , n8106 );
xor ( n8108 , n5171 , n6572 );
buf ( n535369 , n8108 );
buf ( n535370 , n535369 );
buf ( n8111 , n535370 );
and ( n8112 , n8111 , n8104 );
nor ( n8113 , n8107 , n8112 );
not ( n8114 , n8113 );
and ( n8115 , n6614 , n7036 );
and ( n8116 , n6816 , n7034 );
nor ( n8117 , n8115 , n8116 );
xnor ( n8118 , n8117 , n7125 );
and ( n8119 , n6868 , n7144 );
and ( n8120 , n6928 , n7142 );
nor ( n8121 , n8119 , n8120 );
xnor ( n8122 , n8121 , n7154 );
xor ( n8123 , n8118 , n8122 );
and ( n8124 , n7929 , n6923 );
and ( n8125 , n8039 , n6921 );
nor ( n8126 , n8124 , n8125 );
xnor ( n8127 , n8126 , n6933 );
xor ( n8128 , n8123 , n8127 );
and ( n8129 , n8114 , n8128 );
and ( n8130 , n7149 , n6852 );
and ( n8131 , n7879 , n6850 );
nor ( n8132 , n8130 , n8131 );
xnor ( n8133 , n8132 , n6862 );
and ( n8134 , n6928 , n7874 );
and ( n8135 , n7130 , n7872 );
nor ( n8136 , n8134 , n8135 );
xnor ( n8137 , n8136 , n7884 );
and ( n8138 , n8133 , n8137 );
and ( n8139 , n7898 , n6923 );
and ( n8140 , n7929 , n6921 );
nor ( n8141 , n8139 , n8140 );
xnor ( n8142 , n8141 , n6933 );
and ( n8143 , n8137 , n8142 );
and ( n8144 , n8133 , n8142 );
or ( n8145 , n8138 , n8143 , n8144 );
and ( n8146 , n8128 , n8145 );
and ( n8147 , n8114 , n8145 );
or ( n8148 , n8129 , n8146 , n8147 );
and ( n8149 , n8087 , n8148 );
and ( n8150 , n7748 , n7732 );
and ( n8151 , n7767 , n7730 );
nor ( n8152 , n8150 , n8151 );
xnor ( n8153 , n8152 , n7742 );
and ( n8154 , n7783 , n7762 );
and ( n8155 , n7802 , n7760 );
nor ( n8156 , n8154 , n8155 );
xnor ( n8157 , n8156 , n7772 );
and ( n8158 , n8153 , n8157 );
and ( n8159 , n7812 , n7797 );
and ( n8160 , n7831 , n7795 );
nor ( n8161 , n8159 , n8160 );
xnor ( n8162 , n8161 , n7807 );
and ( n8163 , n8157 , n8162 );
and ( n8164 , n8153 , n8162 );
or ( n8165 , n8158 , n8163 , n8164 );
and ( n8166 , n6816 , n7847 );
and ( n8167 , n7022 , n7845 );
nor ( n8168 , n8166 , n8167 );
xnor ( n8169 , n8168 , n7857 );
and ( n8170 , n8021 , n6722 );
and ( n8171 , n6826 , n6720 );
nor ( n8172 , n8170 , n8171 );
xnor ( n8173 , n8172 , n6821 );
and ( n8174 , n8169 , n8173 );
and ( n8175 , n7979 , n7963 );
and ( n8176 , n8000 , n7961 );
nor ( n8177 , n8175 , n8176 );
xnor ( n8178 , n8177 , n7973 );
and ( n8179 , n8173 , n8178 );
and ( n8180 , n8169 , n8178 );
or ( n8181 , n8174 , n8179 , n8180 );
and ( n8182 , n8165 , n8181 );
and ( n8183 , n7737 , n7683 );
and ( n8184 , n7671 , n7680 );
nor ( n8185 , n8183 , n8184 );
xnor ( n8186 , n8185 , n7676 );
and ( n8187 , n7767 , n7732 );
and ( n8188 , n7718 , n7730 );
nor ( n8189 , n8187 , n8188 );
xnor ( n8190 , n8189 , n7742 );
xor ( n8191 , n8186 , n8190 );
and ( n8192 , n7802 , n7762 );
and ( n8193 , n7748 , n7760 );
nor ( n8194 , n8192 , n8193 );
xnor ( n8195 , n8194 , n7772 );
xor ( n8196 , n8191 , n8195 );
and ( n8197 , n8181 , n8196 );
and ( n8198 , n8165 , n8196 );
or ( n8199 , n8182 , n8197 , n8198 );
and ( n8200 , n8148 , n8199 );
and ( n8201 , n8087 , n8199 );
or ( n8202 , n8149 , n8200 , n8201 );
and ( n8203 , n8058 , n8202 );
and ( n8204 , n7852 , n7826 );
and ( n8205 , n7812 , n7824 );
nor ( n8206 , n8204 , n8205 );
xnor ( n8207 , n8206 , n7836 );
and ( n8208 , n7022 , n7847 );
and ( n8209 , n7120 , n7845 );
nor ( n8210 , n8208 , n8209 );
xnor ( n8211 , n8210 , n7857 );
xor ( n8212 , n8207 , n8211 );
and ( n8213 , n6826 , n6722 );
and ( n8214 , n6857 , n6720 );
nor ( n8215 , n8213 , n8214 );
xnor ( n8216 , n8215 , n6821 );
xor ( n8217 , n8212 , n8216 );
and ( n8218 , n7879 , n6852 );
and ( n8219 , n8021 , n6850 );
nor ( n8220 , n8218 , n8219 );
xnor ( n8221 , n8220 , n6862 );
and ( n8222 , n7130 , n7874 );
and ( n8223 , n7149 , n7872 );
nor ( n8224 , n8222 , n8223 );
xnor ( n8225 , n8224 , n7884 );
xor ( n8226 , n8221 , n8225 );
and ( n8227 , n7968 , n7924 );
and ( n8228 , n7898 , n7922 );
nor ( n8229 , n8227 , n8228 );
xnor ( n8230 , n8229 , n7934 );
xor ( n8231 , n8226 , n8230 );
and ( n8232 , n8217 , n8231 );
and ( n8233 , n8000 , n7963 );
and ( n8234 , n7939 , n7961 );
nor ( n8235 , n8233 , n8234 );
xnor ( n8236 , n8235 , n7973 );
and ( n8237 , n8076 , n7995 );
and ( n8238 , n7979 , n7993 );
nor ( n8239 , n8237 , n8238 );
xnor ( n8240 , n8239 , n8005 );
xor ( n8241 , n8236 , n8240 );
xor ( n8242 , n5059 , n6574 );
buf ( n535503 , n8242 );
buf ( n535504 , n535503 );
buf ( n8245 , n535504 );
xor ( n8246 , n535353 , n8094 );
buf ( n535507 , n8246 );
buf ( n535508 , n535507 );
buf ( n8249 , n535508 );
xor ( n8250 , n8103 , n8249 );
xor ( n8251 , n8249 , n7987 );
not ( n8252 , n8251 );
and ( n8253 , n8250 , n8252 );
and ( n8254 , n8245 , n8253 );
and ( n8255 , n8071 , n8251 );
nor ( n8256 , n8254 , n8255 );
and ( n8257 , n8249 , n7987 );
not ( n8258 , n8257 );
and ( n8259 , n8103 , n8258 );
xnor ( n8260 , n8256 , n8259 );
xor ( n8261 , n8241 , n8260 );
and ( n8262 , n8231 , n8261 );
and ( n8263 , n8217 , n8261 );
or ( n8264 , n8232 , n8262 , n8263 );
and ( n8265 , n8071 , n8253 );
and ( n8266 , n8076 , n8251 );
nor ( n8267 , n8265 , n8266 );
xnor ( n8268 , n8267 , n8259 );
and ( n8269 , n8111 , n8106 );
and ( n8270 , n8245 , n8104 );
nor ( n8271 , n8269 , n8270 );
not ( n8272 , n8271 );
xor ( n8273 , n8268 , n8272 );
and ( n8274 , n6816 , n7036 );
and ( n8275 , n7022 , n7034 );
nor ( n8276 , n8274 , n8275 );
xnor ( n8277 , n8276 , n7125 );
and ( n8278 , n8021 , n6852 );
and ( n8279 , n6826 , n6850 );
nor ( n8280 , n8278 , n8279 );
xnor ( n8281 , n8280 , n6862 );
xor ( n8282 , n8277 , n8281 );
and ( n8283 , n8039 , n6923 );
and ( n8284 , n6868 , n6921 );
nor ( n8285 , n8283 , n8284 );
xnor ( n8286 , n8285 , n6933 );
xor ( n8287 , n8282 , n8286 );
xor ( n8288 , n8273 , n8287 );
and ( n8289 , n8264 , n8288 );
and ( n8290 , n8118 , n8122 );
and ( n8291 , n8122 , n8127 );
and ( n8292 , n8118 , n8127 );
or ( n8293 , n8290 , n8291 , n8292 );
and ( n8294 , n8186 , n8190 );
and ( n8295 , n8190 , n8195 );
and ( n8296 , n8186 , n8195 );
or ( n8297 , n8294 , n8295 , n8296 );
xor ( n8298 , n8293 , n8297 );
and ( n8299 , n8207 , n8211 );
and ( n8300 , n8211 , n8216 );
and ( n8301 , n8207 , n8216 );
or ( n8302 , n8299 , n8300 , n8301 );
xor ( n8303 , n8298 , n8302 );
and ( n8304 , n8288 , n8303 );
and ( n8305 , n8264 , n8303 );
or ( n8306 , n8289 , n8304 , n8305 );
and ( n8307 , n8202 , n8306 );
and ( n8308 , n8058 , n8306 );
or ( n8309 , n8203 , n8307 , n8308 );
xor ( n8310 , n8056 , n8309 );
and ( n8311 , n7711 , n7683 );
and ( n8312 , n7691 , n7695 );
and ( n8313 , n7695 , n7697 );
and ( n8314 , n7691 , n7697 );
or ( n8315 , n8312 , n8313 , n8314 );
and ( n8316 , n1953 , n2091 );
not ( n8317 , n8316 );
xnor ( n8318 , n8317 , n2099 );
xor ( n8319 , n8315 , n8318 );
and ( n8320 , n1942 , n1926 );
not ( n8321 , n8320 );
xor ( n8322 , n8319 , n8321 );
and ( n8323 , n7688 , n7689 );
and ( n8324 , n7689 , n7698 );
and ( n8325 , n7688 , n7698 );
or ( n8326 , n8323 , n8324 , n8325 );
xor ( n8327 , n8322 , n8326 );
and ( n8328 , n7699 , n7703 );
and ( n8329 , n7704 , n7707 );
or ( n8330 , n8328 , n8329 );
xor ( n8331 , n8327 , n8330 );
buf ( n535592 , n8331 );
buf ( n535593 , n535592 );
buf ( n8334 , n535593 );
and ( n8335 , n8334 , n7680 );
nor ( n8336 , n8311 , n8335 );
xnor ( n8337 , n8336 , n7676 );
and ( n8338 , n7737 , n7732 );
and ( n8339 , n7671 , n7730 );
nor ( n8340 , n8338 , n8339 );
xnor ( n8341 , n8340 , n7742 );
xor ( n8342 , n8337 , n8341 );
and ( n8343 , n7767 , n7762 );
and ( n8344 , n7718 , n7760 );
nor ( n8345 , n8343 , n8344 );
xnor ( n8346 , n8345 , n7772 );
xor ( n8347 , n8342 , n8346 );
and ( n8348 , n7802 , n7797 );
and ( n8349 , n7748 , n7795 );
nor ( n8350 , n8348 , n8349 );
xnor ( n8351 , n8350 , n7807 );
and ( n8352 , n7831 , n7826 );
and ( n8353 , n7783 , n7824 );
nor ( n8354 , n8352 , n8353 );
xnor ( n8355 , n8354 , n7836 );
xor ( n8356 , n8351 , n8355 );
and ( n8357 , n7929 , n7924 );
and ( n8358 , n8039 , n7922 );
nor ( n8359 , n8357 , n8358 );
xnor ( n8360 , n8359 , n7934 );
xor ( n8361 , n8356 , n8360 );
xor ( n8362 , n8347 , n8361 );
and ( n8363 , n8277 , n8281 );
and ( n8364 , n8281 , n8286 );
and ( n8365 , n8277 , n8286 );
or ( n8366 , n8363 , n8364 , n8365 );
and ( n8367 , n7852 , n7847 );
and ( n8368 , n7812 , n7845 );
nor ( n8369 , n8367 , n8368 );
xnor ( n8370 , n8369 , n7857 );
xor ( n8371 , n8366 , n8370 );
xor ( n8372 , n8362 , n8371 );
and ( n8373 , n8268 , n8272 );
and ( n8374 , n8272 , n8287 );
and ( n8375 , n8268 , n8287 );
or ( n8376 , n8373 , n8374 , n8375 );
and ( n8377 , n8293 , n8297 );
and ( n8378 , n8297 , n8302 );
and ( n8379 , n8293 , n8302 );
or ( n8380 , n8377 , n8378 , n8379 );
xor ( n8381 , n8376 , n8380 );
and ( n8382 , n8221 , n8225 );
and ( n8383 , n8225 , n8230 );
and ( n8384 , n8221 , n8230 );
or ( n8385 , n8382 , n8383 , n8384 );
and ( n8386 , n8236 , n8240 );
and ( n8387 , n8240 , n8260 );
and ( n8388 , n8236 , n8260 );
or ( n8389 , n8386 , n8387 , n8388 );
and ( n8390 , n8385 , n8389 );
xor ( n8391 , n7714 , n7743 );
xor ( n8392 , n8391 , n7773 );
and ( n8393 , n8389 , n8392 );
and ( n8394 , n8385 , n8392 );
or ( n8395 , n8390 , n8393 , n8394 );
xor ( n8396 , n8381 , n8395 );
and ( n8397 , n8372 , n8396 );
xor ( n8398 , n7808 , n7837 );
xor ( n8399 , n8398 , n7858 );
xor ( n8400 , n7865 , n7885 );
xor ( n8401 , n8400 , n7890 );
and ( n8402 , n8399 , n8401 );
xor ( n8403 , n7935 , n7974 );
xor ( n8404 , n8403 , n8006 );
and ( n8405 , n8401 , n8404 );
and ( n8406 , n8399 , n8404 );
or ( n8407 , n8402 , n8405 , n8406 );
and ( n8408 , n8000 , n7995 );
and ( n8409 , n7939 , n7993 );
nor ( n8410 , n8408 , n8409 );
xnor ( n8411 , n8410 , n8005 );
and ( n8412 , n8245 , n8106 );
and ( n8413 , n8071 , n8104 );
nor ( n8414 , n8412 , n8413 );
not ( n8415 , n8414 );
xor ( n8416 , n8411 , n8415 );
and ( n8417 , n7879 , n7874 );
and ( n8418 , n8021 , n7872 );
nor ( n8419 , n8417 , n8418 );
xnor ( n8420 , n8419 , n7884 );
and ( n8421 , n7968 , n7963 );
and ( n8422 , n7898 , n7961 );
nor ( n8423 , n8421 , n8422 );
xnor ( n8424 , n8423 , n7973 );
xor ( n8425 , n8420 , n8424 );
and ( n8426 , n8076 , n8253 );
and ( n8427 , n7979 , n8251 );
nor ( n8428 , n8426 , n8427 );
xnor ( n8429 , n8428 , n8259 );
xor ( n8430 , n8425 , n8429 );
xor ( n8431 , n8416 , n8430 );
xor ( n8432 , n8407 , n8431 );
xor ( n8433 , n6935 , n7156 );
xor ( n8434 , n8433 , n7776 );
xor ( n8435 , n8432 , n8434 );
and ( n8436 , n8396 , n8435 );
and ( n8437 , n8372 , n8435 );
or ( n8438 , n8397 , n8436 , n8437 );
xor ( n8439 , n8310 , n8438 );
xor ( n8440 , n8372 , n8396 );
xor ( n8441 , n8440 , n8435 );
xor ( n8442 , n8264 , n8288 );
xor ( n8443 , n8442 , n8303 );
and ( n8444 , n6816 , n7826 );
and ( n8445 , n7022 , n7824 );
nor ( n8446 , n8444 , n8445 );
xnor ( n8447 , n8446 , n7836 );
and ( n8448 , n6857 , n7847 );
and ( n8449 , n6614 , n7845 );
nor ( n8450 , n8448 , n8449 );
xnor ( n8451 , n8450 , n7857 );
and ( n8452 , n8447 , n8451 );
and ( n8453 , n8021 , n7036 );
and ( n8454 , n6826 , n7034 );
nor ( n8455 , n8453 , n8454 );
xnor ( n8456 , n8455 , n7125 );
and ( n8457 , n8451 , n8456 );
and ( n8458 , n8447 , n8456 );
or ( n8459 , n8452 , n8457 , n8458 );
and ( n8460 , n8039 , n7874 );
and ( n8461 , n6868 , n7872 );
nor ( n8462 , n8460 , n8461 );
xnor ( n8463 , n8462 , n7884 );
and ( n8464 , n7898 , n7144 );
and ( n8465 , n7929 , n7142 );
nor ( n8466 , n8464 , n8465 );
xnor ( n8467 , n8466 , n7154 );
and ( n8468 , n8463 , n8467 );
and ( n8469 , n7939 , n6923 );
and ( n8470 , n7968 , n6921 );
nor ( n8471 , n8469 , n8470 );
xnor ( n8472 , n8471 , n6933 );
and ( n8473 , n8467 , n8472 );
and ( n8474 , n8463 , n8472 );
or ( n8475 , n8468 , n8473 , n8474 );
and ( n8476 , n8459 , n8475 );
and ( n8477 , n7852 , n7797 );
and ( n8478 , n7812 , n7795 );
nor ( n8479 , n8477 , n8478 );
xnor ( n8480 , n8479 , n7807 );
and ( n8481 , n8475 , n8480 );
and ( n8482 , n8459 , n8480 );
or ( n8483 , n8476 , n8481 , n8482 );
and ( n8484 , n7718 , n7683 );
and ( n8485 , n7737 , n7680 );
nor ( n8486 , n8484 , n8485 );
xnor ( n8487 , n8486 , n7676 );
and ( n8488 , n8483 , n8487 );
and ( n8489 , n7879 , n6722 );
and ( n8490 , n8021 , n6720 );
nor ( n8491 , n8489 , n8490 );
xnor ( n8492 , n8491 , n6821 );
and ( n8493 , n6868 , n7874 );
and ( n8494 , n6928 , n7872 );
nor ( n8495 , n8493 , n8494 );
xnor ( n8496 , n8495 , n7884 );
and ( n8497 , n8492 , n8496 );
and ( n8498 , n7929 , n7144 );
and ( n8499 , n8039 , n7142 );
nor ( n8500 , n8498 , n8499 );
xnor ( n8501 , n8500 , n7154 );
and ( n8502 , n8496 , n8501 );
and ( n8503 , n8492 , n8501 );
or ( n8504 , n8497 , n8502 , n8503 );
and ( n8505 , n7120 , n7826 );
and ( n8506 , n7852 , n7824 );
nor ( n8507 , n8505 , n8506 );
xnor ( n8508 , n8507 , n7836 );
xor ( n8509 , n8504 , n8508 );
xor ( n8510 , n8062 , n8066 );
xor ( n8511 , n8510 , n8079 );
xor ( n8512 , n8509 , n8511 );
and ( n8513 , n8487 , n8512 );
and ( n8514 , n8483 , n8512 );
or ( n8515 , n8488 , n8513 , n8514 );
and ( n8516 , n7968 , n6923 );
and ( n8517 , n7898 , n6921 );
nor ( n8518 , n8516 , n8517 );
xnor ( n8519 , n8518 , n6933 );
and ( n8520 , n8000 , n7924 );
and ( n8521 , n7939 , n7922 );
nor ( n8522 , n8520 , n8521 );
xnor ( n8523 , n8522 , n7934 );
and ( n8524 , n8519 , n8523 );
and ( n8525 , n8076 , n7963 );
and ( n8526 , n7979 , n7961 );
nor ( n8527 , n8525 , n8526 );
xnor ( n8528 , n8527 , n7973 );
and ( n8529 , n8523 , n8528 );
and ( n8530 , n8519 , n8528 );
or ( n8531 , n8524 , n8529 , n8530 );
and ( n8532 , n6857 , n7036 );
and ( n8533 , n6614 , n7034 );
nor ( n8534 , n8532 , n8533 );
xnor ( n8535 , n8534 , n7125 );
xor ( n8536 , n8531 , n8535 );
xor ( n8537 , n8519 , n8523 );
xor ( n8538 , n8537 , n8528 );
and ( n8539 , n6614 , n7847 );
and ( n8540 , n6816 , n7845 );
nor ( n8541 , n8539 , n8540 );
xnor ( n8542 , n8541 , n7857 );
and ( n8543 , n7130 , n6852 );
and ( n8544 , n7149 , n6850 );
nor ( n8545 , n8543 , n8544 );
xnor ( n8546 , n8545 , n6862 );
xor ( n8547 , n8542 , n8546 );
and ( n8548 , n8538 , n8547 );
and ( n8549 , n7022 , n7826 );
and ( n8550 , n7120 , n7824 );
nor ( n8551 , n8549 , n8550 );
xnor ( n8552 , n8551 , n7836 );
and ( n8553 , n6826 , n7036 );
and ( n8554 , n6857 , n7034 );
nor ( n8555 , n8553 , n8554 );
xnor ( n8556 , n8555 , n7125 );
xor ( n8557 , n8552 , n8556 );
and ( n8558 , n8547 , n8557 );
and ( n8559 , n8538 , n8557 );
or ( n8560 , n8548 , n8558 , n8559 );
and ( n8561 , n8536 , n8560 );
and ( n8562 , n7979 , n7924 );
and ( n8563 , n8000 , n7922 );
nor ( n8564 , n8562 , n8563 );
xnor ( n8565 , n8564 , n7934 );
and ( n8566 , n8071 , n7963 );
and ( n8567 , n8076 , n7961 );
nor ( n8568 , n8566 , n8567 );
xnor ( n8569 , n8568 , n7973 );
and ( n8570 , n8565 , n8569 );
and ( n8571 , n7783 , n7732 );
and ( n8572 , n7802 , n7730 );
nor ( n8573 , n8571 , n8572 );
xnor ( n8574 , n8573 , n7742 );
and ( n8575 , n7812 , n7762 );
and ( n8576 , n7831 , n7760 );
nor ( n8577 , n8575 , n8576 );
xnor ( n8578 , n8577 , n7772 );
and ( n8579 , n8574 , n8578 );
and ( n8580 , n7120 , n7797 );
and ( n8581 , n7852 , n7795 );
nor ( n8582 , n8580 , n8581 );
xnor ( n8583 , n8582 , n7807 );
and ( n8584 , n8578 , n8583 );
and ( n8585 , n8574 , n8583 );
or ( n8586 , n8579 , n8584 , n8585 );
and ( n8587 , n8570 , n8586 );
and ( n8588 , n8111 , n7995 );
and ( n8589 , n8245 , n7993 );
nor ( n8590 , n8588 , n8589 );
xnor ( n8591 , n8590 , n8005 );
xor ( n8592 , n5390 , n6568 );
buf ( n535853 , n8592 );
buf ( n535854 , n535853 );
buf ( n8595 , n535854 );
and ( n8596 , n8595 , n8253 );
and ( n8597 , n8091 , n8251 );
nor ( n8598 , n8596 , n8597 );
xnor ( n8599 , n8598 , n8259 );
and ( n8600 , n8591 , n8599 );
xor ( n8601 , n5589 , n6564 );
buf ( n535862 , n8601 );
buf ( n535863 , n535862 );
buf ( n8604 , n535863 );
and ( n8605 , n8604 , n8106 );
xor ( n8606 , n5443 , n6566 );
buf ( n535867 , n8606 );
buf ( n535868 , n535867 );
buf ( n8609 , n535868 );
and ( n8610 , n8609 , n8104 );
nor ( n8611 , n8605 , n8610 );
not ( n8612 , n8611 );
and ( n8613 , n8599 , n8612 );
and ( n8614 , n8591 , n8612 );
or ( n8615 , n8600 , n8613 , n8614 );
and ( n8616 , n8586 , n8615 );
and ( n8617 , n8570 , n8615 );
or ( n8618 , n8587 , n8616 , n8617 );
and ( n8619 , n8560 , n8618 );
and ( n8620 , n8536 , n8618 );
or ( n8621 , n8561 , n8619 , n8620 );
and ( n8622 , n8515 , n8621 );
and ( n8623 , n8111 , n8253 );
and ( n8624 , n8245 , n8251 );
nor ( n8625 , n8623 , n8624 );
xnor ( n8626 , n8625 , n8259 );
and ( n8627 , n8595 , n8106 );
and ( n8628 , n8091 , n8104 );
nor ( n8629 , n8627 , n8628 );
not ( n8630 , n8629 );
xor ( n8631 , n8626 , n8630 );
xor ( n8632 , n8133 , n8137 );
xor ( n8633 , n8632 , n8142 );
xor ( n8634 , n8631 , n8633 );
and ( n8635 , n8542 , n8546 );
and ( n8636 , n8552 , n8556 );
xor ( n8637 , n8635 , n8636 );
and ( n8638 , n7767 , n7683 );
and ( n8639 , n7718 , n7680 );
nor ( n8640 , n8638 , n8639 );
xnor ( n8641 , n8640 , n7676 );
and ( n8642 , n7802 , n7732 );
and ( n8643 , n7748 , n7730 );
nor ( n8644 , n8642 , n8643 );
xnor ( n8645 , n8644 , n7742 );
and ( n8646 , n8641 , n8645 );
and ( n8647 , n7831 , n7762 );
and ( n8648 , n7783 , n7760 );
nor ( n8649 , n8647 , n8648 );
xnor ( n8650 , n8649 , n7772 );
and ( n8651 , n8645 , n8650 );
and ( n8652 , n8641 , n8650 );
or ( n8653 , n8646 , n8651 , n8652 );
xor ( n8654 , n8637 , n8653 );
and ( n8655 , n8634 , n8654 );
and ( n8656 , n8245 , n7995 );
and ( n8657 , n8071 , n7993 );
nor ( n8658 , n8656 , n8657 );
xnor ( n8659 , n8658 , n8005 );
and ( n8660 , n8091 , n8253 );
and ( n8661 , n8111 , n8251 );
nor ( n8662 , n8660 , n8661 );
xnor ( n8663 , n8662 , n8259 );
and ( n8664 , n8659 , n8663 );
and ( n8665 , n8609 , n8106 );
and ( n8666 , n8595 , n8104 );
nor ( n8667 , n8665 , n8666 );
not ( n8668 , n8667 );
and ( n8669 , n8663 , n8668 );
and ( n8670 , n8659 , n8668 );
or ( n8671 , n8664 , n8669 , n8670 );
xor ( n8672 , n8153 , n8157 );
xor ( n8673 , n8672 , n8162 );
xor ( n8674 , n8671 , n8673 );
xor ( n8675 , n8169 , n8173 );
xor ( n8676 , n8675 , n8178 );
xor ( n8677 , n8674 , n8676 );
and ( n8678 , n8654 , n8677 );
and ( n8679 , n8634 , n8677 );
or ( n8680 , n8655 , n8678 , n8679 );
and ( n8681 , n8621 , n8680 );
and ( n8682 , n8515 , n8680 );
or ( n8683 , n8622 , n8681 , n8682 );
and ( n8684 , n8443 , n8683 );
xor ( n8685 , n8082 , n8086 );
and ( n8686 , n8504 , n8508 );
and ( n8687 , n8508 , n8511 );
and ( n8688 , n8504 , n8511 );
or ( n8689 , n8686 , n8687 , n8688 );
xor ( n8690 , n8685 , n8689 );
and ( n8691 , n8531 , n8535 );
xor ( n8692 , n8690 , n8691 );
and ( n8693 , n8626 , n8630 );
and ( n8694 , n8630 , n8633 );
and ( n8695 , n8626 , n8633 );
or ( n8696 , n8693 , n8694 , n8695 );
and ( n8697 , n8635 , n8636 );
and ( n8698 , n8636 , n8653 );
and ( n8699 , n8635 , n8653 );
or ( n8700 , n8697 , n8698 , n8699 );
xor ( n8701 , n8696 , n8700 );
and ( n8702 , n8671 , n8673 );
and ( n8703 , n8673 , n8676 );
and ( n8704 , n8671 , n8676 );
or ( n8705 , n8702 , n8703 , n8704 );
xor ( n8706 , n8701 , n8705 );
and ( n8707 , n8692 , n8706 );
xor ( n8708 , n8114 , n8128 );
xor ( n8709 , n8708 , n8145 );
xor ( n8710 , n8165 , n8181 );
xor ( n8711 , n8710 , n8196 );
xor ( n8712 , n8709 , n8711 );
xor ( n8713 , n8217 , n8231 );
xor ( n8714 , n8713 , n8261 );
xor ( n8715 , n8712 , n8714 );
and ( n8716 , n8706 , n8715 );
and ( n8717 , n8692 , n8715 );
or ( n8718 , n8707 , n8716 , n8717 );
and ( n8719 , n8683 , n8718 );
and ( n8720 , n8443 , n8718 );
or ( n8721 , n8684 , n8719 , n8720 );
and ( n8722 , n8441 , n8721 );
xor ( n8723 , n8385 , n8389 );
xor ( n8724 , n8723 , n8392 );
xor ( n8725 , n8399 , n8401 );
xor ( n8726 , n8725 , n8404 );
and ( n8727 , n8724 , n8726 );
and ( n8728 , n8685 , n8689 );
and ( n8729 , n8689 , n8691 );
and ( n8730 , n8685 , n8691 );
or ( n8731 , n8728 , n8729 , n8730 );
and ( n8732 , n8726 , n8731 );
and ( n8733 , n8724 , n8731 );
or ( n8734 , n8727 , n8732 , n8733 );
and ( n8735 , n8696 , n8700 );
and ( n8736 , n8700 , n8705 );
and ( n8737 , n8696 , n8705 );
or ( n8738 , n8735 , n8736 , n8737 );
and ( n8739 , n8709 , n8711 );
and ( n8740 , n8711 , n8714 );
and ( n8741 , n8709 , n8714 );
or ( n8742 , n8739 , n8740 , n8741 );
and ( n8743 , n8738 , n8742 );
xor ( n8744 , n8087 , n8148 );
xor ( n8745 , n8744 , n8199 );
and ( n8746 , n8742 , n8745 );
and ( n8747 , n8738 , n8745 );
or ( n8748 , n8743 , n8746 , n8747 );
xor ( n8749 , n8734 , n8748 );
xor ( n8750 , n8058 , n8202 );
xor ( n8751 , n8750 , n8306 );
xor ( n8752 , n8749 , n8751 );
and ( n8753 , n8721 , n8752 );
and ( n8754 , n8441 , n8752 );
or ( n8755 , n8722 , n8753 , n8754 );
xor ( n8756 , n8439 , n8755 );
and ( n8757 , n7126 , n7155 );
and ( n8758 , n8337 , n8341 );
and ( n8759 , n8341 , n8346 );
and ( n8760 , n8337 , n8346 );
or ( n8761 , n8758 , n8759 , n8760 );
xor ( n8762 , n8757 , n8761 );
and ( n8763 , n8351 , n8355 );
and ( n8764 , n8355 , n8360 );
and ( n8765 , n8351 , n8360 );
or ( n8766 , n8763 , n8764 , n8765 );
xor ( n8767 , n8762 , n8766 );
and ( n8768 , n8334 , n7683 );
and ( n8769 , n8315 , n8318 );
and ( n8770 , n8318 , n8321 );
and ( n8771 , n8315 , n8321 );
or ( n8772 , n8769 , n8770 , n8771 );
buf ( n8773 , n8320 );
not ( n8774 , n2099 );
xor ( n8775 , n8773 , n8774 );
and ( n8776 , n1953 , n1926 );
xor ( n8777 , n8775 , n8776 );
xor ( n8778 , n8772 , n8777 );
and ( n8779 , n8322 , n8326 );
and ( n8780 , n8327 , n8330 );
or ( n8781 , n8779 , n8780 );
xor ( n8782 , n8778 , n8781 );
buf ( n536043 , n8782 );
buf ( n536044 , n536043 );
buf ( n8785 , n536044 );
and ( n8786 , n8785 , n7680 );
nor ( n8787 , n8768 , n8786 );
xnor ( n8788 , n8787 , n7676 );
and ( n8789 , n7671 , n7732 );
and ( n8790 , n7711 , n7730 );
nor ( n8791 , n8789 , n8790 );
xnor ( n8792 , n8791 , n7742 );
xor ( n8793 , n8788 , n8792 );
and ( n8794 , n7718 , n7762 );
and ( n8795 , n7737 , n7760 );
nor ( n8796 , n8794 , n8795 );
xnor ( n8797 , n8796 , n7772 );
xor ( n8798 , n8793 , n8797 );
and ( n8799 , n7748 , n7797 );
and ( n8800 , n7767 , n7795 );
nor ( n8801 , n8799 , n8800 );
xnor ( n8802 , n8801 , n7807 );
and ( n8803 , n7783 , n7826 );
and ( n8804 , n7802 , n7824 );
nor ( n8805 , n8803 , n8804 );
xnor ( n8806 , n8805 , n7836 );
xor ( n8807 , n8802 , n8806 );
and ( n8808 , n7120 , n7036 );
and ( n8809 , n7852 , n7034 );
nor ( n8810 , n8808 , n8809 );
xnor ( n8811 , n8810 , n7125 );
xor ( n8812 , n8807 , n8811 );
xor ( n8813 , n8798 , n8812 );
and ( n8814 , n7939 , n7995 );
and ( n8815 , n7968 , n7993 );
nor ( n8816 , n8814 , n8815 );
xnor ( n8817 , n8816 , n8005 );
and ( n8818 , n7979 , n8253 );
and ( n8819 , n8000 , n8251 );
nor ( n8820 , n8818 , n8819 );
xnor ( n8821 , n8820 , n8259 );
xor ( n8822 , n8817 , n8821 );
and ( n8823 , n8071 , n8106 );
and ( n8824 , n8076 , n8104 );
nor ( n8825 , n8823 , n8824 );
not ( n8826 , n8825 );
xor ( n8827 , n8822 , n8826 );
xor ( n8828 , n8813 , n8827 );
xor ( n8829 , n8767 , n8828 );
and ( n8830 , n8347 , n8361 );
and ( n8831 , n8361 , n8371 );
and ( n8832 , n8347 , n8371 );
or ( n8833 , n8830 , n8831 , n8832 );
xor ( n8834 , n8829 , n8833 );
and ( n8835 , n8376 , n8380 );
and ( n8836 , n8380 , n8395 );
and ( n8837 , n8376 , n8395 );
or ( n8838 , n8835 , n8836 , n8837 );
and ( n8839 , n8407 , n8431 );
and ( n8840 , n8431 , n8434 );
and ( n8841 , n8407 , n8434 );
or ( n8842 , n8839 , n8840 , n8841 );
xor ( n8843 , n8838 , n8842 );
and ( n8844 , n8420 , n8424 );
and ( n8845 , n8424 , n8429 );
and ( n8846 , n8420 , n8429 );
or ( n8847 , n8844 , n8845 , n8846 );
and ( n8848 , n7812 , n7847 );
and ( n8849 , n7831 , n7845 );
nor ( n8850 , n8848 , n8849 );
xnor ( n8851 , n8850 , n7857 );
xor ( n8852 , n8847 , n8851 );
and ( n8853 , n6816 , n6722 );
and ( n8854 , n7022 , n6720 );
nor ( n8855 , n8853 , n8854 );
xnor ( n8856 , n8855 , n6821 );
xor ( n8857 , n8852 , n8856 );
and ( n8858 , n8366 , n8370 );
xor ( n8859 , n8857 , n8858 );
and ( n8860 , n8411 , n8415 );
and ( n8861 , n8415 , n8430 );
and ( n8862 , n8411 , n8430 );
or ( n8863 , n8860 , n8861 , n8862 );
xor ( n8864 , n8859 , n8863 );
xor ( n8865 , n8843 , n8864 );
xor ( n8866 , n8834 , n8865 );
and ( n8867 , n8734 , n8748 );
and ( n8868 , n8748 , n8751 );
and ( n8869 , n8734 , n8751 );
or ( n8870 , n8867 , n8868 , n8869 );
xor ( n8871 , n8866 , n8870 );
xor ( n8872 , n8756 , n8871 );
xor ( n8873 , n8724 , n8726 );
xor ( n8874 , n8873 , n8731 );
xor ( n8875 , n8738 , n8742 );
xor ( n8876 , n8875 , n8745 );
and ( n8877 , n8874 , n8876 );
xor ( n8878 , n8483 , n8487 );
xor ( n8879 , n8878 , n8512 );
and ( n8880 , n8000 , n6923 );
and ( n8881 , n7939 , n6921 );
nor ( n8882 , n8880 , n8881 );
xnor ( n8883 , n8882 , n6933 );
and ( n8884 , n8076 , n7924 );
and ( n8885 , n7979 , n7922 );
nor ( n8886 , n8884 , n8885 );
xnor ( n8887 , n8886 , n7934 );
and ( n8888 , n8883 , n8887 );
and ( n8889 , n8245 , n7963 );
and ( n8890 , n8071 , n7961 );
nor ( n8891 , n8889 , n8890 );
xnor ( n8892 , n8891 , n7973 );
and ( n8893 , n8887 , n8892 );
and ( n8894 , n8883 , n8892 );
or ( n8895 , n8888 , n8893 , n8894 );
and ( n8896 , n7149 , n6722 );
and ( n8897 , n7879 , n6720 );
nor ( n8898 , n8896 , n8897 );
xnor ( n8899 , n8898 , n6821 );
and ( n8900 , n8895 , n8899 );
and ( n8901 , n6928 , n6852 );
and ( n8902 , n7130 , n6850 );
nor ( n8903 , n8901 , n8902 );
xnor ( n8904 , n8903 , n6862 );
and ( n8905 , n8899 , n8904 );
and ( n8906 , n8895 , n8904 );
or ( n8907 , n8900 , n8905 , n8906 );
xor ( n8908 , n8492 , n8496 );
xor ( n8909 , n8908 , n8501 );
and ( n8910 , n8907 , n8909 );
and ( n8911 , n8879 , n8910 );
xor ( n8912 , n8641 , n8645 );
xor ( n8913 , n8912 , n8650 );
xor ( n8914 , n8659 , n8663 );
xor ( n8915 , n8914 , n8668 );
and ( n8916 , n8913 , n8915 );
xor ( n8917 , n8463 , n8467 );
xor ( n8918 , n8917 , n8472 );
xor ( n8919 , n8565 , n8569 );
and ( n8920 , n8918 , n8919 );
and ( n8921 , n7879 , n7036 );
and ( n8922 , n8021 , n7034 );
nor ( n8923 , n8921 , n8922 );
xnor ( n8924 , n8923 , n7125 );
and ( n8925 , n6868 , n6852 );
and ( n8926 , n6928 , n6850 );
nor ( n8927 , n8925 , n8926 );
xnor ( n8928 , n8927 , n6862 );
and ( n8929 , n8924 , n8928 );
and ( n8930 , n7929 , n7874 );
and ( n8931 , n8039 , n7872 );
nor ( n8932 , n8930 , n8931 );
xnor ( n8933 , n8932 , n7884 );
and ( n8934 , n8928 , n8933 );
and ( n8935 , n8924 , n8933 );
or ( n8936 , n8929 , n8934 , n8935 );
and ( n8937 , n8919 , n8936 );
and ( n8938 , n8918 , n8936 );
or ( n8939 , n8920 , n8937 , n8938 );
and ( n8940 , n8915 , n8939 );
and ( n8941 , n8913 , n8939 );
or ( n8942 , n8916 , n8940 , n8941 );
and ( n8943 , n8910 , n8942 );
and ( n8944 , n8879 , n8942 );
or ( n8945 , n8911 , n8943 , n8944 );
and ( n8946 , n7802 , n7683 );
and ( n8947 , n7748 , n7680 );
nor ( n8948 , n8946 , n8947 );
xnor ( n8949 , n8948 , n7676 );
and ( n8950 , n7831 , n7732 );
and ( n8951 , n7783 , n7730 );
nor ( n8952 , n8950 , n8951 );
xnor ( n8953 , n8952 , n7742 );
and ( n8954 , n8949 , n8953 );
and ( n8955 , n7852 , n7762 );
and ( n8956 , n7812 , n7760 );
nor ( n8957 , n8955 , n8956 );
xnor ( n8958 , n8957 , n7772 );
and ( n8959 , n8953 , n8958 );
and ( n8960 , n8949 , n8958 );
or ( n8961 , n8954 , n8959 , n8960 );
and ( n8962 , n7022 , n7797 );
and ( n8963 , n7120 , n7795 );
nor ( n8964 , n8962 , n8963 );
xnor ( n8965 , n8964 , n7807 );
and ( n8966 , n6614 , n7826 );
and ( n8967 , n6816 , n7824 );
nor ( n8968 , n8966 , n8967 );
xnor ( n8969 , n8968 , n7836 );
and ( n8970 , n8965 , n8969 );
and ( n8971 , n7130 , n6722 );
and ( n8972 , n7149 , n6720 );
nor ( n8973 , n8971 , n8972 );
xnor ( n8974 , n8973 , n6821 );
and ( n8975 , n8969 , n8974 );
and ( n8976 , n8965 , n8974 );
or ( n8977 , n8970 , n8975 , n8976 );
and ( n8978 , n8961 , n8977 );
and ( n8979 , n7968 , n7144 );
and ( n8980 , n7898 , n7142 );
nor ( n8981 , n8979 , n8980 );
xnor ( n8982 , n8981 , n7154 );
and ( n8983 , n8091 , n7995 );
and ( n8984 , n8111 , n7993 );
nor ( n8985 , n8983 , n8984 );
xnor ( n8986 , n8985 , n8005 );
and ( n8987 , n8982 , n8986 );
and ( n8988 , n8609 , n8253 );
and ( n8989 , n8595 , n8251 );
nor ( n8990 , n8988 , n8989 );
xnor ( n8991 , n8990 , n8259 );
and ( n8992 , n8986 , n8991 );
and ( n8993 , n8982 , n8991 );
or ( n8994 , n8987 , n8992 , n8993 );
and ( n8995 , n8977 , n8994 );
and ( n8996 , n8961 , n8994 );
or ( n8997 , n8978 , n8995 , n8996 );
xor ( n8998 , n8538 , n8547 );
xor ( n8999 , n8998 , n8557 );
and ( n9000 , n8997 , n8999 );
xor ( n9001 , n8570 , n8586 );
xor ( n9002 , n9001 , n8615 );
and ( n9003 , n8999 , n9002 );
and ( n9004 , n8997 , n9002 );
or ( n9005 , n9000 , n9003 , n9004 );
xor ( n9006 , n8536 , n8560 );
xor ( n9007 , n9006 , n8618 );
and ( n9008 , n9005 , n9007 );
xor ( n9009 , n8634 , n8654 );
xor ( n9010 , n9009 , n8677 );
and ( n9011 , n9007 , n9010 );
and ( n9012 , n9005 , n9010 );
or ( n9013 , n9008 , n9011 , n9012 );
and ( n9014 , n8945 , n9013 );
xor ( n9015 , n8515 , n8621 );
xor ( n9016 , n9015 , n8680 );
and ( n9017 , n9013 , n9016 );
and ( n9018 , n8945 , n9016 );
or ( n9019 , n9014 , n9017 , n9018 );
and ( n9020 , n8876 , n9019 );
and ( n9021 , n8874 , n9019 );
or ( n9022 , n8877 , n9020 , n9021 );
xor ( n9023 , n8441 , n8721 );
xor ( n9024 , n9023 , n8752 );
and ( n9025 , n9022 , n9024 );
xor ( n9026 , n8443 , n8683 );
xor ( n9027 , n9026 , n8718 );
xor ( n9028 , n8692 , n8706 );
xor ( n9029 , n9028 , n8715 );
and ( n9030 , n7979 , n6923 );
and ( n9031 , n8000 , n6921 );
nor ( n9032 , n9030 , n9031 );
xnor ( n9033 , n9032 , n6933 );
and ( n9034 , n8071 , n7924 );
and ( n9035 , n8076 , n7922 );
nor ( n9036 , n9034 , n9035 );
xnor ( n9037 , n9036 , n7934 );
and ( n9038 , n9033 , n9037 );
and ( n9039 , n8595 , n7995 );
and ( n9040 , n8091 , n7993 );
nor ( n9041 , n9039 , n9040 );
xnor ( n9042 , n9041 , n8005 );
and ( n9043 , n9037 , n9042 );
and ( n9044 , n9033 , n9042 );
or ( n9045 , n9038 , n9043 , n9044 );
and ( n9046 , n6826 , n7847 );
and ( n9047 , n6857 , n7845 );
nor ( n9048 , n9046 , n9047 );
xnor ( n9049 , n9048 , n7857 );
and ( n9050 , n9045 , n9049 );
xor ( n9051 , n8883 , n8887 );
xor ( n9052 , n9051 , n8892 );
and ( n9053 , n9049 , n9052 );
and ( n9054 , n9045 , n9052 );
or ( n9055 , n9050 , n9053 , n9054 );
and ( n9056 , n7748 , n7683 );
and ( n9057 , n7767 , n7680 );
nor ( n9058 , n9056 , n9057 );
xnor ( n9059 , n9058 , n7676 );
and ( n9060 , n9055 , n9059 );
xor ( n9061 , n8447 , n8451 );
xor ( n9062 , n9061 , n8456 );
and ( n9063 , n9059 , n9062 );
and ( n9064 , n9055 , n9062 );
or ( n9065 , n9060 , n9063 , n9064 );
xor ( n9066 , n8459 , n8475 );
xor ( n9067 , n9066 , n8480 );
and ( n9068 , n9065 , n9067 );
xor ( n9069 , n8907 , n8909 );
xor ( n9070 , n8574 , n8578 );
xor ( n9071 , n9070 , n8583 );
xor ( n9072 , n8591 , n8599 );
xor ( n9073 , n9072 , n8612 );
and ( n9074 , n9071 , n9073 );
xor ( n9075 , n8895 , n8899 );
xor ( n9076 , n9075 , n8904 );
and ( n9077 , n9073 , n9076 );
and ( n9078 , n9071 , n9076 );
or ( n9079 , n9074 , n9077 , n9078 );
and ( n9080 , n9069 , n9079 );
xor ( n9081 , n5619 , n6562 );
buf ( n536342 , n9081 );
buf ( n536343 , n536342 );
buf ( n9084 , n536343 );
and ( n9085 , n9084 , n8106 );
and ( n9086 , n8604 , n8104 );
nor ( n9087 , n9085 , n9086 );
not ( n9088 , n9087 );
xor ( n9089 , n8924 , n8928 );
xor ( n9090 , n9089 , n8933 );
and ( n9091 , n9088 , n9090 );
and ( n9092 , n8039 , n6852 );
and ( n9093 , n6868 , n6850 );
nor ( n9094 , n9092 , n9093 );
xnor ( n9095 , n9094 , n6862 );
and ( n9096 , n7898 , n7874 );
and ( n9097 , n7929 , n7872 );
nor ( n9098 , n9096 , n9097 );
xnor ( n9099 , n9098 , n7884 );
and ( n9100 , n9095 , n9099 );
and ( n9101 , n9090 , n9100 );
and ( n9102 , n9088 , n9100 );
or ( n9103 , n9091 , n9101 , n9102 );
and ( n9104 , n8021 , n7847 );
and ( n9105 , n6826 , n7845 );
nor ( n9106 , n9104 , n9105 );
xnor ( n9107 , n9106 , n7857 );
and ( n9108 , n7149 , n7036 );
and ( n9109 , n7879 , n7034 );
nor ( n9110 , n9108 , n9109 );
xnor ( n9111 , n9110 , n7125 );
and ( n9112 , n9107 , n9111 );
and ( n9113 , n7783 , n7683 );
and ( n9114 , n7802 , n7680 );
nor ( n9115 , n9113 , n9114 );
xnor ( n9116 , n9115 , n7676 );
and ( n9117 , n7120 , n7762 );
and ( n9118 , n7852 , n7760 );
nor ( n9119 , n9117 , n9118 );
xnor ( n9120 , n9119 , n7772 );
and ( n9121 , n9116 , n9120 );
and ( n9122 , n6816 , n7797 );
and ( n9123 , n7022 , n7795 );
nor ( n9124 , n9122 , n9123 );
xnor ( n9125 , n9124 , n7807 );
and ( n9126 , n9120 , n9125 );
and ( n9127 , n9116 , n9125 );
or ( n9128 , n9121 , n9126 , n9127 );
and ( n9129 , n9112 , n9128 );
and ( n9130 , n6857 , n7826 );
and ( n9131 , n6614 , n7824 );
nor ( n9132 , n9130 , n9131 );
xnor ( n9133 , n9132 , n7836 );
and ( n9134 , n6928 , n6722 );
and ( n9135 , n7130 , n6720 );
nor ( n9136 , n9134 , n9135 );
xnor ( n9137 , n9136 , n6821 );
and ( n9138 , n9133 , n9137 );
and ( n9139 , n7939 , n7144 );
and ( n9140 , n7968 , n7142 );
nor ( n9141 , n9139 , n9140 );
xnor ( n9142 , n9141 , n7154 );
and ( n9143 , n9137 , n9142 );
and ( n9144 , n9133 , n9142 );
or ( n9145 , n9138 , n9143 , n9144 );
and ( n9146 , n9128 , n9145 );
and ( n9147 , n9112 , n9145 );
or ( n9148 , n9129 , n9146 , n9147 );
and ( n9149 , n9103 , n9148 );
and ( n9150 , n8111 , n7963 );
and ( n9151 , n8245 , n7961 );
nor ( n9152 , n9150 , n9151 );
xnor ( n9153 , n9152 , n7973 );
and ( n9154 , n8604 , n8253 );
and ( n9155 , n8609 , n8251 );
nor ( n9156 , n9154 , n9155 );
xnor ( n9157 , n9156 , n8259 );
and ( n9158 , n9153 , n9157 );
xor ( n9159 , n5702 , n6560 );
buf ( n536420 , n9159 );
buf ( n536421 , n536420 );
buf ( n9162 , n536421 );
and ( n9163 , n9162 , n8106 );
and ( n9164 , n9084 , n8104 );
nor ( n9165 , n9163 , n9164 );
not ( n9166 , n9165 );
and ( n9167 , n9157 , n9166 );
and ( n9168 , n9153 , n9166 );
or ( n9169 , n9158 , n9167 , n9168 );
xor ( n9170 , n8949 , n8953 );
xor ( n9171 , n9170 , n8958 );
and ( n9172 , n9169 , n9171 );
xor ( n9173 , n8965 , n8969 );
xor ( n9174 , n9173 , n8974 );
and ( n9175 , n9171 , n9174 );
and ( n9176 , n9169 , n9174 );
or ( n9177 , n9172 , n9175 , n9176 );
and ( n9178 , n9148 , n9177 );
and ( n9179 , n9103 , n9177 );
or ( n9180 , n9149 , n9178 , n9179 );
and ( n9181 , n9079 , n9180 );
and ( n9182 , n9069 , n9180 );
or ( n9183 , n9080 , n9181 , n9182 );
and ( n9184 , n9068 , n9183 );
xor ( n9185 , n8879 , n8910 );
xor ( n9186 , n9185 , n8942 );
and ( n9187 , n9183 , n9186 );
and ( n9188 , n9068 , n9186 );
or ( n9189 , n9184 , n9187 , n9188 );
and ( n9190 , n9029 , n9189 );
xor ( n9191 , n8945 , n9013 );
xor ( n9192 , n9191 , n9016 );
and ( n9193 , n9189 , n9192 );
and ( n9194 , n9029 , n9192 );
or ( n9195 , n9190 , n9193 , n9194 );
and ( n9196 , n9027 , n9195 );
xor ( n9197 , n8874 , n8876 );
xor ( n9198 , n9197 , n9019 );
and ( n9199 , n9195 , n9198 );
and ( n9200 , n9027 , n9198 );
or ( n9201 , n9196 , n9199 , n9200 );
and ( n9202 , n9024 , n9201 );
and ( n9203 , n9022 , n9201 );
or ( n9204 , n9025 , n9202 , n9203 );
xor ( n9205 , n8872 , n9204 );
xor ( n9206 , n9022 , n9024 );
xor ( n9207 , n9206 , n9201 );
xor ( n9208 , n9027 , n9195 );
xor ( n9209 , n9208 , n9198 );
xor ( n9210 , n9005 , n9007 );
xor ( n9211 , n9210 , n9010 );
xor ( n9212 , n8913 , n8915 );
xor ( n9213 , n9212 , n8939 );
xor ( n9214 , n8997 , n8999 );
xor ( n9215 , n9214 , n9002 );
and ( n9216 , n9213 , n9215 );
xor ( n9217 , n9065 , n9067 );
and ( n9218 , n9215 , n9217 );
and ( n9219 , n9213 , n9217 );
or ( n9220 , n9216 , n9218 , n9219 );
and ( n9221 , n9211 , n9220 );
xor ( n9222 , n8918 , n8919 );
xor ( n9223 , n9222 , n8936 );
xor ( n9224 , n8961 , n8977 );
xor ( n9225 , n9224 , n8994 );
and ( n9226 , n9223 , n9225 );
xor ( n9227 , n9055 , n9059 );
xor ( n9228 , n9227 , n9062 );
and ( n9229 , n9225 , n9228 );
and ( n9230 , n9223 , n9228 );
or ( n9231 , n9226 , n9229 , n9230 );
xor ( n9232 , n8982 , n8986 );
xor ( n9233 , n9232 , n8991 );
xor ( n9234 , n9045 , n9049 );
xor ( n9235 , n9234 , n9052 );
and ( n9236 , n9233 , n9235 );
and ( n9237 , n7812 , n7732 );
and ( n9238 , n7831 , n7730 );
nor ( n9239 , n9237 , n9238 );
xnor ( n9240 , n9239 , n7742 );
xor ( n9241 , n9033 , n9037 );
xor ( n9242 , n9241 , n9042 );
and ( n9243 , n9240 , n9242 );
and ( n9244 , n9235 , n9243 );
and ( n9245 , n9233 , n9243 );
or ( n9246 , n9236 , n9244 , n9245 );
xor ( n9247 , n9095 , n9099 );
xor ( n9248 , n9107 , n9111 );
and ( n9249 , n9247 , n9248 );
and ( n9250 , n8076 , n6923 );
and ( n9251 , n7979 , n6921 );
nor ( n9252 , n9250 , n9251 );
xnor ( n9253 , n9252 , n6933 );
and ( n9254 , n8245 , n7924 );
and ( n9255 , n8071 , n7922 );
nor ( n9256 , n9254 , n9255 );
xnor ( n9257 , n9256 , n7934 );
and ( n9258 , n9253 , n9257 );
and ( n9259 , n8091 , n7963 );
and ( n9260 , n8111 , n7961 );
nor ( n9261 , n9259 , n9260 );
xnor ( n9262 , n9261 , n7973 );
and ( n9263 , n9257 , n9262 );
and ( n9264 , n9253 , n9262 );
or ( n9265 , n9258 , n9263 , n9264 );
and ( n9266 , n9248 , n9265 );
and ( n9267 , n9247 , n9265 );
or ( n9268 , n9249 , n9266 , n9267 );
and ( n9269 , n7968 , n7874 );
and ( n9270 , n7898 , n7872 );
nor ( n9271 , n9269 , n9270 );
xnor ( n9272 , n9271 , n7884 );
and ( n9273 , n8000 , n7144 );
and ( n9274 , n7939 , n7142 );
nor ( n9275 , n9273 , n9274 );
xnor ( n9276 , n9275 , n7154 );
and ( n9277 , n9272 , n9276 );
and ( n9278 , n7022 , n7762 );
and ( n9279 , n7120 , n7760 );
nor ( n9280 , n9278 , n9279 );
xnor ( n9281 , n9280 , n7772 );
and ( n9282 , n6826 , n7826 );
and ( n9283 , n6857 , n7824 );
nor ( n9284 , n9282 , n9283 );
xnor ( n9285 , n9284 , n7836 );
and ( n9286 , n9281 , n9285 );
and ( n9287 , n9277 , n9286 );
and ( n9288 , n7831 , n7683 );
and ( n9289 , n7783 , n7680 );
nor ( n9290 , n9288 , n9289 );
xnor ( n9291 , n9290 , n7676 );
and ( n9292 , n6614 , n7797 );
and ( n9293 , n6816 , n7795 );
nor ( n9294 , n9292 , n9293 );
xnor ( n9295 , n9294 , n7807 );
and ( n9296 , n9291 , n9295 );
and ( n9297 , n7879 , n7847 );
and ( n9298 , n8021 , n7845 );
nor ( n9299 , n9297 , n9298 );
xnor ( n9300 , n9299 , n7857 );
and ( n9301 , n9295 , n9300 );
and ( n9302 , n9291 , n9300 );
or ( n9303 , n9296 , n9301 , n9302 );
and ( n9304 , n9286 , n9303 );
and ( n9305 , n9277 , n9303 );
or ( n9306 , n9287 , n9304 , n9305 );
and ( n9307 , n9268 , n9306 );
and ( n9308 , n6868 , n6722 );
and ( n9309 , n6928 , n6720 );
nor ( n9310 , n9308 , n9309 );
xnor ( n9311 , n9310 , n6821 );
and ( n9312 , n7929 , n6852 );
and ( n9313 , n8039 , n6850 );
nor ( n9314 , n9312 , n9313 );
xnor ( n9315 , n9314 , n6862 );
and ( n9316 , n9311 , n9315 );
and ( n9317 , n8609 , n7995 );
and ( n9318 , n8595 , n7993 );
nor ( n9319 , n9317 , n9318 );
xnor ( n9320 , n9319 , n8005 );
and ( n9321 , n9315 , n9320 );
and ( n9322 , n9311 , n9320 );
or ( n9323 , n9316 , n9321 , n9322 );
xor ( n9324 , n9116 , n9120 );
xor ( n9325 , n9324 , n9125 );
and ( n9326 , n9323 , n9325 );
xor ( n9327 , n9133 , n9137 );
xor ( n9328 , n9327 , n9142 );
and ( n9329 , n9325 , n9328 );
and ( n9330 , n9323 , n9328 );
or ( n9331 , n9326 , n9329 , n9330 );
and ( n9332 , n9306 , n9331 );
and ( n9333 , n9268 , n9331 );
or ( n9334 , n9307 , n9332 , n9333 );
and ( n9335 , n9246 , n9334 );
xor ( n9336 , n9088 , n9090 );
xor ( n9337 , n9336 , n9100 );
xor ( n9338 , n9112 , n9128 );
xor ( n9339 , n9338 , n9145 );
and ( n9340 , n9337 , n9339 );
xor ( n9341 , n9169 , n9171 );
xor ( n9342 , n9341 , n9174 );
and ( n9343 , n9339 , n9342 );
and ( n9344 , n9337 , n9342 );
or ( n9345 , n9340 , n9343 , n9344 );
and ( n9346 , n9334 , n9345 );
and ( n9347 , n9246 , n9345 );
or ( n9348 , n9335 , n9346 , n9347 );
and ( n9349 , n9231 , n9348 );
xor ( n9350 , n9069 , n9079 );
xor ( n9351 , n9350 , n9180 );
and ( n9352 , n9348 , n9351 );
and ( n9353 , n9231 , n9351 );
or ( n9354 , n9349 , n9352 , n9353 );
and ( n9355 , n9220 , n9354 );
and ( n9356 , n9211 , n9354 );
or ( n9357 , n9221 , n9355 , n9356 );
xor ( n9358 , n9029 , n9189 );
xor ( n9359 , n9358 , n9192 );
and ( n9360 , n9357 , n9359 );
xor ( n9361 , n9068 , n9183 );
xor ( n9362 , n9361 , n9186 );
xor ( n9363 , n9071 , n9073 );
xor ( n9364 , n9363 , n9076 );
xor ( n9365 , n9103 , n9148 );
xor ( n9366 , n9365 , n9177 );
and ( n9367 , n9364 , n9366 );
xor ( n9368 , n9153 , n9157 );
xor ( n9369 , n9368 , n9166 );
xor ( n9370 , n9240 , n9242 );
and ( n9371 , n9369 , n9370 );
and ( n9372 , n7939 , n7874 );
and ( n9373 , n7968 , n7872 );
nor ( n9374 , n9372 , n9373 );
xnor ( n9375 , n9374 , n7884 );
and ( n9376 , n7979 , n7144 );
and ( n9377 , n8000 , n7142 );
nor ( n9378 , n9376 , n9377 );
xnor ( n9379 , n9378 , n7154 );
and ( n9380 , n9375 , n9379 );
and ( n9381 , n8071 , n6923 );
and ( n9382 , n8076 , n6921 );
nor ( n9383 , n9381 , n9382 );
xnor ( n9384 , n9383 , n6933 );
and ( n9385 , n9379 , n9384 );
and ( n9386 , n9375 , n9384 );
or ( n9387 , n9380 , n9385 , n9386 );
and ( n9388 , n7852 , n7732 );
and ( n9389 , n7812 , n7730 );
nor ( n9390 , n9388 , n9389 );
xnor ( n9391 , n9390 , n7742 );
and ( n9392 , n9387 , n9391 );
and ( n9393 , n7130 , n7036 );
and ( n9394 , n7149 , n7034 );
nor ( n9395 , n9393 , n9394 );
xnor ( n9396 , n9395 , n7125 );
and ( n9397 , n9391 , n9396 );
and ( n9398 , n9387 , n9396 );
or ( n9399 , n9392 , n9397 , n9398 );
and ( n9400 , n9370 , n9399 );
and ( n9401 , n9369 , n9399 );
or ( n9402 , n9371 , n9400 , n9401 );
and ( n9403 , n9084 , n8253 );
and ( n9404 , n8604 , n8251 );
nor ( n9405 , n9403 , n9404 );
xnor ( n9406 , n9405 , n8259 );
xor ( n9407 , n5803 , n6558 );
buf ( n536668 , n9407 );
buf ( n536669 , n536668 );
buf ( n9410 , n536669 );
and ( n9411 , n9410 , n8106 );
and ( n9412 , n9162 , n8104 );
nor ( n9413 , n9411 , n9412 );
not ( n9414 , n9413 );
and ( n9415 , n9406 , n9414 );
xor ( n9416 , n9253 , n9257 );
xor ( n9417 , n9416 , n9262 );
and ( n9418 , n9414 , n9417 );
and ( n9419 , n9406 , n9417 );
or ( n9420 , n9415 , n9418 , n9419 );
xor ( n9421 , n9272 , n9276 );
xor ( n9422 , n9281 , n9285 );
and ( n9423 , n9421 , n9422 );
and ( n9424 , n8111 , n7924 );
and ( n9425 , n8245 , n7922 );
nor ( n9426 , n9424 , n9425 );
xnor ( n9427 , n9426 , n7934 );
and ( n9428 , n8595 , n7963 );
and ( n9429 , n8091 , n7961 );
nor ( n9430 , n9428 , n9429 );
xnor ( n9431 , n9430 , n7973 );
and ( n9432 , n9427 , n9431 );
and ( n9433 , n9422 , n9432 );
and ( n9434 , n9421 , n9432 );
or ( n9435 , n9423 , n9433 , n9434 );
and ( n9436 , n9420 , n9435 );
and ( n9437 , n7812 , n7683 );
and ( n9438 , n7831 , n7680 );
nor ( n9439 , n9437 , n9438 );
xnor ( n9440 , n9439 , n7676 );
and ( n9441 , n6857 , n7797 );
and ( n9442 , n6614 , n7795 );
nor ( n9443 , n9441 , n9442 );
xnor ( n9444 , n9443 , n7807 );
and ( n9445 , n9440 , n9444 );
and ( n9446 , n7149 , n7847 );
and ( n9447 , n7879 , n7845 );
nor ( n9448 , n9446 , n9447 );
xnor ( n9449 , n9448 , n7857 );
and ( n9450 , n9444 , n9449 );
and ( n9451 , n9440 , n9449 );
or ( n9452 , n9445 , n9450 , n9451 );
and ( n9453 , n6928 , n7036 );
and ( n9454 , n7130 , n7034 );
nor ( n9455 , n9453 , n9454 );
xnor ( n9456 , n9455 , n7125 );
and ( n9457 , n8039 , n6722 );
and ( n9458 , n6868 , n6720 );
nor ( n9459 , n9457 , n9458 );
xnor ( n9460 , n9459 , n6821 );
and ( n9461 , n9456 , n9460 );
and ( n9462 , n7898 , n6852 );
and ( n9463 , n7929 , n6850 );
nor ( n9464 , n9462 , n9463 );
xnor ( n9465 , n9464 , n6862 );
and ( n9466 , n9460 , n9465 );
and ( n9467 , n9456 , n9465 );
or ( n9468 , n9461 , n9466 , n9467 );
and ( n9469 , n9452 , n9468 );
and ( n9470 , n8604 , n7995 );
and ( n9471 , n8609 , n7993 );
nor ( n9472 , n9470 , n9471 );
xnor ( n9473 , n9472 , n8005 );
and ( n9474 , n9162 , n8253 );
and ( n9475 , n9084 , n8251 );
nor ( n9476 , n9474 , n9475 );
xnor ( n9477 , n9476 , n8259 );
and ( n9478 , n9473 , n9477 );
xor ( n9479 , n5879 , n6556 );
buf ( n536740 , n9479 );
buf ( n536741 , n536740 );
buf ( n9482 , n536741 );
and ( n9483 , n9482 , n8106 );
and ( n9484 , n9410 , n8104 );
nor ( n9485 , n9483 , n9484 );
not ( n9486 , n9485 );
and ( n9487 , n9477 , n9486 );
and ( n9488 , n9473 , n9486 );
or ( n9489 , n9478 , n9487 , n9488 );
and ( n9490 , n9468 , n9489 );
and ( n9491 , n9452 , n9489 );
or ( n9492 , n9469 , n9490 , n9491 );
and ( n9493 , n9435 , n9492 );
and ( n9494 , n9420 , n9492 );
or ( n9495 , n9436 , n9493 , n9494 );
and ( n9496 , n9402 , n9495 );
xor ( n9497 , n9247 , n9248 );
xor ( n9498 , n9497 , n9265 );
xor ( n9499 , n9277 , n9286 );
xor ( n9500 , n9499 , n9303 );
and ( n9501 , n9498 , n9500 );
xor ( n9502 , n9323 , n9325 );
xor ( n9503 , n9502 , n9328 );
and ( n9504 , n9500 , n9503 );
and ( n9505 , n9498 , n9503 );
or ( n9506 , n9501 , n9504 , n9505 );
and ( n9507 , n9495 , n9506 );
and ( n9508 , n9402 , n9506 );
or ( n9509 , n9496 , n9507 , n9508 );
and ( n9510 , n9366 , n9509 );
and ( n9511 , n9364 , n9509 );
or ( n9512 , n9367 , n9510 , n9511 );
xor ( n9513 , n9233 , n9235 );
xor ( n9514 , n9513 , n9243 );
xor ( n9515 , n9268 , n9306 );
xor ( n9516 , n9515 , n9331 );
and ( n9517 , n9514 , n9516 );
xor ( n9518 , n9337 , n9339 );
xor ( n9519 , n9518 , n9342 );
and ( n9520 , n9516 , n9519 );
and ( n9521 , n9514 , n9519 );
or ( n9522 , n9517 , n9520 , n9521 );
xor ( n9523 , n9223 , n9225 );
xor ( n9524 , n9523 , n9228 );
and ( n9525 , n9522 , n9524 );
xor ( n9526 , n9246 , n9334 );
xor ( n9527 , n9526 , n9345 );
and ( n9528 , n9524 , n9527 );
and ( n9529 , n9522 , n9527 );
or ( n9530 , n9525 , n9528 , n9529 );
and ( n9531 , n9512 , n9530 );
xor ( n9532 , n9213 , n9215 );
xor ( n9533 , n9532 , n9217 );
and ( n9534 , n9530 , n9533 );
and ( n9535 , n9512 , n9533 );
or ( n9536 , n9531 , n9534 , n9535 );
and ( n9537 , n9362 , n9536 );
xor ( n9538 , n9211 , n9220 );
xor ( n9539 , n9538 , n9354 );
and ( n9540 , n9536 , n9539 );
and ( n9541 , n9362 , n9539 );
or ( n9542 , n9537 , n9540 , n9541 );
and ( n9543 , n9359 , n9542 );
and ( n9544 , n9357 , n9542 );
or ( n9545 , n9360 , n9543 , n9544 );
and ( n9546 , n9209 , n9545 );
xor ( n9547 , n9209 , n9545 );
xor ( n9548 , n9357 , n9359 );
xor ( n9549 , n9548 , n9542 );
xor ( n9550 , n9231 , n9348 );
xor ( n9551 , n9550 , n9351 );
and ( n9552 , n6614 , n7762 );
and ( n9553 , n6816 , n7760 );
nor ( n9554 , n9552 , n9553 );
xnor ( n9555 , n9554 , n7772 );
and ( n9556 , n7879 , n7826 );
and ( n9557 , n8021 , n7824 );
nor ( n9558 , n9556 , n9557 );
xnor ( n9559 , n9558 , n7836 );
and ( n9560 , n9555 , n9559 );
and ( n9561 , n7929 , n6722 );
and ( n9562 , n8039 , n6720 );
nor ( n9563 , n9561 , n9562 );
xnor ( n9564 , n9563 , n6821 );
and ( n9565 , n9559 , n9564 );
and ( n9566 , n9555 , n9564 );
or ( n9567 , n9560 , n9565 , n9566 );
and ( n9568 , n7120 , n7732 );
and ( n9569 , n7852 , n7730 );
nor ( n9570 , n9568 , n9569 );
xnor ( n9571 , n9570 , n7742 );
and ( n9572 , n9567 , n9571 );
xor ( n9573 , n9375 , n9379 );
xor ( n9574 , n9573 , n9384 );
and ( n9575 , n9571 , n9574 );
and ( n9576 , n9567 , n9574 );
or ( n9577 , n9572 , n9575 , n9576 );
xor ( n9578 , n9387 , n9391 );
xor ( n9579 , n9578 , n9396 );
and ( n9580 , n9577 , n9579 );
xor ( n9581 , n9291 , n9295 );
xor ( n9582 , n9581 , n9300 );
xor ( n9583 , n9311 , n9315 );
xor ( n9584 , n9583 , n9320 );
and ( n9585 , n9582 , n9584 );
and ( n9586 , n8000 , n7874 );
and ( n9587 , n7939 , n7872 );
nor ( n9588 , n9586 , n9587 );
xnor ( n9589 , n9588 , n7884 );
and ( n9590 , n8076 , n7144 );
and ( n9591 , n7979 , n7142 );
nor ( n9592 , n9590 , n9591 );
xnor ( n9593 , n9592 , n7154 );
and ( n9594 , n9589 , n9593 );
and ( n9595 , n8245 , n6923 );
and ( n9596 , n8071 , n6921 );
nor ( n9597 , n9595 , n9596 );
xnor ( n9598 , n9597 , n6933 );
and ( n9599 , n9593 , n9598 );
and ( n9600 , n9589 , n9598 );
or ( n9601 , n9594 , n9599 , n9600 );
and ( n9602 , n6816 , n7762 );
and ( n9603 , n7022 , n7760 );
nor ( n9604 , n9602 , n9603 );
xnor ( n9605 , n9604 , n7772 );
and ( n9606 , n9601 , n9605 );
and ( n9607 , n8021 , n7826 );
and ( n9608 , n6826 , n7824 );
nor ( n9609 , n9607 , n9608 );
xnor ( n9610 , n9609 , n7836 );
and ( n9611 , n9605 , n9610 );
and ( n9612 , n9601 , n9610 );
or ( n9613 , n9606 , n9611 , n9612 );
and ( n9614 , n9584 , n9613 );
and ( n9615 , n9582 , n9613 );
or ( n9616 , n9585 , n9614 , n9615 );
and ( n9617 , n9580 , n9616 );
xor ( n9618 , n9427 , n9431 );
and ( n9619 , n8609 , n7963 );
and ( n9620 , n8595 , n7961 );
nor ( n9621 , n9619 , n9620 );
xnor ( n9622 , n9621 , n7973 );
and ( n9623 , n9084 , n7995 );
and ( n9624 , n8604 , n7993 );
nor ( n9625 , n9623 , n9624 );
xnor ( n9626 , n9625 , n8005 );
and ( n9627 , n9622 , n9626 );
and ( n9628 , n9618 , n9627 );
and ( n9629 , n7852 , n7683 );
and ( n9630 , n7812 , n7680 );
nor ( n9631 , n9629 , n9630 );
xnor ( n9632 , n9631 , n7676 );
and ( n9633 , n7022 , n7732 );
and ( n9634 , n7120 , n7730 );
nor ( n9635 , n9633 , n9634 );
xnor ( n9636 , n9635 , n7742 );
and ( n9637 , n9632 , n9636 );
and ( n9638 , n6826 , n7797 );
and ( n9639 , n6857 , n7795 );
nor ( n9640 , n9638 , n9639 );
xnor ( n9641 , n9640 , n7807 );
and ( n9642 , n9636 , n9641 );
and ( n9643 , n9632 , n9641 );
or ( n9644 , n9637 , n9642 , n9643 );
and ( n9645 , n9627 , n9644 );
and ( n9646 , n9618 , n9644 );
or ( n9647 , n9628 , n9645 , n9646 );
and ( n9648 , n7130 , n7847 );
and ( n9649 , n7149 , n7845 );
nor ( n9650 , n9648 , n9649 );
xnor ( n9651 , n9650 , n7857 );
and ( n9652 , n6868 , n7036 );
and ( n9653 , n6928 , n7034 );
nor ( n9654 , n9652 , n9653 );
xnor ( n9655 , n9654 , n7125 );
and ( n9656 , n9651 , n9655 );
and ( n9657 , n7968 , n6852 );
and ( n9658 , n7898 , n6850 );
nor ( n9659 , n9657 , n9658 );
xnor ( n9660 , n9659 , n6862 );
and ( n9661 , n9655 , n9660 );
and ( n9662 , n9651 , n9660 );
or ( n9663 , n9656 , n9661 , n9662 );
and ( n9664 , n8091 , n7924 );
and ( n9665 , n8111 , n7922 );
nor ( n9666 , n9664 , n9665 );
xnor ( n9667 , n9666 , n7934 );
and ( n9668 , n9410 , n8253 );
and ( n9669 , n9162 , n8251 );
nor ( n9670 , n9668 , n9669 );
xnor ( n9671 , n9670 , n8259 );
and ( n9672 , n9667 , n9671 );
xor ( n9673 , n5951 , n6554 );
buf ( n536934 , n9673 );
buf ( n536935 , n536934 );
buf ( n9676 , n536935 );
and ( n9677 , n9676 , n8106 );
and ( n9678 , n9482 , n8104 );
nor ( n9679 , n9677 , n9678 );
not ( n9680 , n9679 );
and ( n9681 , n9671 , n9680 );
and ( n9682 , n9667 , n9680 );
or ( n9683 , n9672 , n9681 , n9682 );
and ( n9684 , n9663 , n9683 );
xor ( n9685 , n9440 , n9444 );
xor ( n9686 , n9685 , n9449 );
and ( n9687 , n9683 , n9686 );
and ( n9688 , n9663 , n9686 );
or ( n9689 , n9684 , n9687 , n9688 );
and ( n9690 , n9647 , n9689 );
xor ( n9691 , n9406 , n9414 );
xor ( n9692 , n9691 , n9417 );
and ( n9693 , n9689 , n9692 );
and ( n9694 , n9647 , n9692 );
or ( n9695 , n9690 , n9693 , n9694 );
and ( n9696 , n9616 , n9695 );
and ( n9697 , n9580 , n9695 );
or ( n9698 , n9617 , n9696 , n9697 );
xor ( n9699 , n9369 , n9370 );
xor ( n9700 , n9699 , n9399 );
xor ( n9701 , n9420 , n9435 );
xor ( n9702 , n9701 , n9492 );
and ( n9703 , n9700 , n9702 );
xor ( n9704 , n9498 , n9500 );
xor ( n9705 , n9704 , n9503 );
and ( n9706 , n9702 , n9705 );
and ( n9707 , n9700 , n9705 );
or ( n9708 , n9703 , n9706 , n9707 );
and ( n9709 , n9698 , n9708 );
xor ( n9710 , n9402 , n9495 );
xor ( n9711 , n9710 , n9506 );
and ( n9712 , n9708 , n9711 );
and ( n9713 , n9698 , n9711 );
or ( n9714 , n9709 , n9712 , n9713 );
xor ( n9715 , n9364 , n9366 );
xor ( n9716 , n9715 , n9509 );
and ( n9717 , n9714 , n9716 );
xor ( n9718 , n9522 , n9524 );
xor ( n9719 , n9718 , n9527 );
and ( n9720 , n9716 , n9719 );
and ( n9721 , n9714 , n9719 );
or ( n9722 , n9717 , n9720 , n9721 );
and ( n9723 , n9551 , n9722 );
xor ( n9724 , n9512 , n9530 );
xor ( n9725 , n9724 , n9533 );
and ( n9726 , n9722 , n9725 );
and ( n9727 , n9551 , n9725 );
or ( n9728 , n9723 , n9726 , n9727 );
xor ( n9729 , n9362 , n9536 );
xor ( n9730 , n9729 , n9539 );
and ( n9731 , n9728 , n9730 );
xor ( n9732 , n9728 , n9730 );
xor ( n9733 , n9551 , n9722 );
xor ( n9734 , n9733 , n9725 );
xor ( n9735 , n9514 , n9516 );
xor ( n9736 , n9735 , n9519 );
xor ( n9737 , n9421 , n9422 );
xor ( n9738 , n9737 , n9432 );
xor ( n9739 , n9452 , n9468 );
xor ( n9740 , n9739 , n9489 );
and ( n9741 , n9738 , n9740 );
xor ( n9742 , n9577 , n9579 );
and ( n9743 , n9740 , n9742 );
and ( n9744 , n9738 , n9742 );
or ( n9745 , n9741 , n9743 , n9744 );
xor ( n9746 , n9456 , n9460 );
xor ( n9747 , n9746 , n9465 );
xor ( n9748 , n9473 , n9477 );
xor ( n9749 , n9748 , n9486 );
and ( n9750 , n9747 , n9749 );
xor ( n9751 , n9601 , n9605 );
xor ( n9752 , n9751 , n9610 );
and ( n9753 , n9749 , n9752 );
and ( n9754 , n9747 , n9752 );
or ( n9755 , n9750 , n9753 , n9754 );
xor ( n9756 , n9567 , n9571 );
xor ( n9757 , n9756 , n9574 );
xor ( n9758 , n9589 , n9593 );
xor ( n9759 , n9758 , n9598 );
xor ( n9760 , n9555 , n9559 );
xor ( n9761 , n9760 , n9564 );
and ( n9762 , n9759 , n9761 );
xor ( n9763 , n9622 , n9626 );
and ( n9764 , n9761 , n9763 );
and ( n9765 , n9759 , n9763 );
or ( n9766 , n9762 , n9764 , n9765 );
and ( n9767 , n9757 , n9766 );
and ( n9768 , n6928 , n7847 );
and ( n9769 , n7130 , n7845 );
nor ( n9770 , n9768 , n9769 );
xnor ( n9771 , n9770 , n7857 );
and ( n9772 , n8039 , n7036 );
and ( n9773 , n6868 , n7034 );
nor ( n9774 , n9772 , n9773 );
xnor ( n9775 , n9774 , n7125 );
and ( n9776 , n9771 , n9775 );
and ( n9777 , n7898 , n6722 );
and ( n9778 , n7929 , n6720 );
nor ( n9779 , n9777 , n9778 );
xnor ( n9780 , n9779 , n6821 );
and ( n9781 , n9775 , n9780 );
and ( n9782 , n9771 , n9780 );
or ( n9783 , n9776 , n9781 , n9782 );
and ( n9784 , n6816 , n7732 );
and ( n9785 , n7022 , n7730 );
nor ( n9786 , n9784 , n9785 );
xnor ( n9787 , n9786 , n7742 );
and ( n9788 , n6857 , n7762 );
and ( n9789 , n6614 , n7760 );
nor ( n9790 , n9788 , n9789 );
xnor ( n9791 , n9790 , n7772 );
and ( n9792 , n9787 , n9791 );
and ( n9793 , n8021 , n7797 );
and ( n9794 , n6826 , n7795 );
nor ( n9795 , n9793 , n9794 );
xnor ( n9796 , n9795 , n7807 );
and ( n9797 , n9791 , n9796 );
and ( n9798 , n9787 , n9796 );
or ( n9799 , n9792 , n9797 , n9798 );
and ( n9800 , n9783 , n9799 );
and ( n9801 , n7149 , n7826 );
and ( n9802 , n7879 , n7824 );
nor ( n9803 , n9801 , n9802 );
xnor ( n9804 , n9803 , n7836 );
and ( n9805 , n7939 , n6852 );
and ( n9806 , n7968 , n6850 );
nor ( n9807 , n9805 , n9806 );
xnor ( n9808 , n9807 , n6862 );
and ( n9809 , n9804 , n9808 );
and ( n9810 , n7979 , n7874 );
and ( n537071 , n8000 , n7872 );
nor ( n9812 , n9810 , n537071 );
xnor ( n537073 , n9812 , n7884 );
and ( n9814 , n9808 , n537073 );
and ( n9815 , n9804 , n537073 );
or ( n9816 , n9809 , n9814 , n9815 );
and ( n9817 , n9799 , n9816 );
and ( n9818 , n9783 , n9816 );
or ( n9819 , n9800 , n9817 , n9818 );
and ( n9820 , n9766 , n9819 );
and ( n9821 , n9757 , n9819 );
or ( n9822 , n9767 , n9820 , n9821 );
and ( n9823 , n9755 , n9822 );
and ( n9824 , n8071 , n7144 );
and ( n9825 , n8076 , n7142 );
nor ( n9826 , n9824 , n9825 );
xnor ( n9827 , n9826 , n7154 );
and ( n9828 , n8111 , n6923 );
and ( n9829 , n8245 , n6921 );
nor ( n9830 , n9828 , n9829 );
xnor ( n9831 , n9830 , n6933 );
and ( n9832 , n9827 , n9831 );
and ( n9833 , n8595 , n7924 );
and ( n9834 , n8091 , n7922 );
nor ( n9835 , n9833 , n9834 );
xnor ( n9836 , n9835 , n7934 );
and ( n9837 , n9831 , n9836 );
and ( n9838 , n9827 , n9836 );
or ( n9839 , n9832 , n9837 , n9838 );
and ( n9840 , n8604 , n7963 );
and ( n9841 , n8609 , n7961 );
nor ( n9842 , n9840 , n9841 );
xnor ( n9843 , n9842 , n7973 );
and ( n9844 , n9162 , n7995 );
and ( n9845 , n9084 , n7993 );
nor ( n9846 , n9844 , n9845 );
xnor ( n9847 , n9846 , n8005 );
and ( n9848 , n9843 , n9847 );
and ( n9849 , n9482 , n8253 );
and ( n9850 , n9410 , n8251 );
nor ( n9851 , n9849 , n9850 );
xnor ( n9852 , n9851 , n8259 );
and ( n9853 , n9847 , n9852 );
and ( n9854 , n9843 , n9852 );
or ( n9855 , n9848 , n9853 , n9854 );
and ( n9856 , n9839 , n9855 );
xor ( n9857 , n9632 , n9636 );
xor ( n9858 , n9857 , n9641 );
and ( n9859 , n9855 , n9858 );
and ( n9860 , n9839 , n9858 );
or ( n9861 , n9856 , n9859 , n9860 );
xor ( n9862 , n9618 , n9627 );
xor ( n9863 , n9862 , n9644 );
and ( n9864 , n9861 , n9863 );
xor ( n9865 , n9663 , n9683 );
xor ( n9866 , n9865 , n9686 );
and ( n9867 , n9863 , n9866 );
and ( n9868 , n9861 , n9866 );
or ( n9869 , n9864 , n9867 , n9868 );
and ( n9870 , n9822 , n9869 );
and ( n9871 , n9755 , n9869 );
or ( n9872 , n9823 , n9870 , n9871 );
and ( n9873 , n9745 , n9872 );
xor ( n9874 , n9580 , n9616 );
xor ( n9875 , n9874 , n9695 );
and ( n9876 , n9872 , n9875 );
and ( n9877 , n9745 , n9875 );
or ( n9878 , n9873 , n9876 , n9877 );
and ( n9879 , n9736 , n9878 );
xor ( n9880 , n9698 , n9708 );
xor ( n9881 , n9880 , n9711 );
and ( n9882 , n9878 , n9881 );
and ( n9883 , n9736 , n9881 );
or ( n9884 , n9879 , n9882 , n9883 );
xor ( n9885 , n9714 , n9716 );
xor ( n9886 , n9885 , n9719 );
and ( n9887 , n9884 , n9886 );
xor ( n9888 , n9700 , n9702 );
xor ( n9889 , n9888 , n9705 );
xor ( n9890 , n9582 , n9584 );
xor ( n9891 , n9890 , n9613 );
xor ( n9892 , n9647 , n9689 );
xor ( n9893 , n9892 , n9692 );
and ( n9894 , n9891 , n9893 );
xor ( n9895 , n9651 , n9655 );
xor ( n9896 , n9895 , n9660 );
xor ( n9897 , n9667 , n9671 );
xor ( n9898 , n9897 , n9680 );
and ( n9899 , n9896 , n9898 );
and ( n9900 , n7022 , n7683 );
and ( n9901 , n7120 , n7680 );
nor ( n9902 , n9900 , n9901 );
xnor ( n9903 , n9902 , n7676 );
and ( n9904 , n7130 , n7826 );
and ( n9905 , n7149 , n7824 );
nor ( n9906 , n9904 , n9905 );
xnor ( n9907 , n9906 , n7836 );
and ( n9908 , n9903 , n9907 );
and ( n9909 , n7929 , n7036 );
and ( n9910 , n8039 , n7034 );
nor ( n9911 , n9909 , n9910 );
xnor ( n9912 , n9911 , n7125 );
and ( n9913 , n9907 , n9912 );
and ( n9914 , n9903 , n9912 );
or ( n9915 , n9908 , n9913 , n9914 );
xor ( n9916 , n9771 , n9775 );
xor ( n9917 , n9916 , n9780 );
and ( n9918 , n9915 , n9917 );
and ( n9919 , n9898 , n9918 );
and ( n9920 , n9896 , n9918 );
or ( n9921 , n9899 , n9919 , n9920 );
xor ( n9922 , n6014 , n6552 );
buf ( n537183 , n9922 );
buf ( n537184 , n537183 );
buf ( n9925 , n537184 );
and ( n9926 , n9925 , n8106 );
and ( n9927 , n9676 , n8104 );
nor ( n9928 , n9926 , n9927 );
not ( n9929 , n9928 );
and ( n9930 , n8091 , n6923 );
and ( n9931 , n8111 , n6921 );
nor ( n9932 , n9930 , n9931 );
xnor ( n9933 , n9932 , n6933 );
and ( n9934 , n8609 , n7924 );
and ( n9935 , n8595 , n7922 );
nor ( n9936 , n9934 , n9935 );
xnor ( n9937 , n9936 , n7934 );
and ( n9938 , n9933 , n9937 );
and ( n9939 , n9084 , n7963 );
and ( n9940 , n8604 , n7961 );
nor ( n9941 , n9939 , n9940 );
xnor ( n9942 , n9941 , n7973 );
and ( n9943 , n9937 , n9942 );
and ( n9944 , n9933 , n9942 );
or ( n9945 , n9938 , n9943 , n9944 );
and ( n9946 , n9929 , n9945 );
and ( n9947 , n6826 , n7762 );
and ( n9948 , n6857 , n7760 );
nor ( n9949 , n9947 , n9948 );
xnor ( n9950 , n9949 , n7772 );
and ( n9951 , n8000 , n6852 );
and ( n9952 , n7939 , n6850 );
nor ( n9953 , n9951 , n9952 );
xnor ( n9954 , n9953 , n6862 );
and ( n9955 , n9950 , n9954 );
and ( n9956 , n8076 , n7874 );
and ( n9957 , n7979 , n7872 );
nor ( n9958 , n9956 , n9957 );
xnor ( n9959 , n9958 , n7884 );
and ( n9960 , n9954 , n9959 );
and ( n9961 , n9950 , n9959 );
or ( n9962 , n9955 , n9960 , n9961 );
and ( n9963 , n9945 , n9962 );
and ( n9964 , n9929 , n9962 );
or ( n9965 , n9946 , n9963 , n9964 );
and ( n9966 , n8245 , n7144 );
and ( n9967 , n8071 , n7142 );
nor ( n9968 , n9966 , n9967 );
xnor ( n9969 , n9968 , n7154 );
and ( n9970 , n9410 , n7995 );
and ( n9971 , n9162 , n7993 );
nor ( n9972 , n9970 , n9971 );
xnor ( n9973 , n9972 , n8005 );
and ( n9974 , n9969 , n9973 );
and ( n9975 , n9676 , n8253 );
and ( n9976 , n9482 , n8251 );
nor ( n9977 , n9975 , n9976 );
xnor ( n9978 , n9977 , n8259 );
and ( n9979 , n9973 , n9978 );
and ( n9980 , n9969 , n9978 );
or ( n9981 , n9974 , n9979 , n9980 );
xor ( n9982 , n9787 , n9791 );
xor ( n9983 , n9982 , n9796 );
and ( n9984 , n9981 , n9983 );
xor ( n9985 , n9804 , n9808 );
xor ( n9986 , n9985 , n537073 );
and ( n9987 , n9983 , n9986 );
and ( n9988 , n9981 , n9986 );
or ( n9989 , n9984 , n9987 , n9988 );
and ( n9990 , n9965 , n9989 );
xor ( n9991 , n9759 , n9761 );
xor ( n9992 , n9991 , n9763 );
and ( n9993 , n9989 , n9992 );
and ( n9994 , n9965 , n9992 );
or ( n9995 , n9990 , n9993 , n9994 );
and ( n9996 , n9921 , n9995 );
xor ( n9997 , n9747 , n9749 );
xor ( n9998 , n9997 , n9752 );
and ( n9999 , n9995 , n9998 );
and ( n10000 , n9921 , n9998 );
or ( n10001 , n9996 , n9999 , n10000 );
and ( n10002 , n9893 , n10001 );
and ( n10003 , n9891 , n10001 );
or ( n10004 , n9894 , n10002 , n10003 );
and ( n10005 , n9889 , n10004 );
xor ( n10006 , n9745 , n9872 );
xor ( n10007 , n10006 , n9875 );
and ( n10008 , n10004 , n10007 );
and ( n10009 , n9889 , n10007 );
or ( n10010 , n10005 , n10008 , n10009 );
xor ( n10011 , n9736 , n9878 );
xor ( n10012 , n10011 , n9881 );
and ( n10013 , n10010 , n10012 );
xor ( n10014 , n9738 , n9740 );
xor ( n10015 , n10014 , n9742 );
xor ( n10016 , n9755 , n9822 );
xor ( n10017 , n10016 , n9869 );
and ( n10018 , n10015 , n10017 );
xor ( n10019 , n9757 , n9766 );
xor ( n10020 , n10019 , n9819 );
xor ( n10021 , n9861 , n9863 );
xor ( n10022 , n10021 , n9866 );
and ( n10023 , n10020 , n10022 );
xor ( n10024 , n9783 , n9799 );
xor ( n10025 , n10024 , n9816 );
xor ( n10026 , n9839 , n9855 );
xor ( n10027 , n10026 , n9858 );
and ( n10028 , n10025 , n10027 );
xor ( n10029 , n9827 , n9831 );
xor ( n10030 , n10029 , n9836 );
xor ( n10031 , n9843 , n9847 );
xor ( n10032 , n10031 , n9852 );
and ( n10033 , n10030 , n10032 );
xor ( n10034 , n9915 , n9917 );
and ( n10035 , n10032 , n10034 );
and ( n10036 , n10030 , n10034 );
or ( n10037 , n10033 , n10035 , n10036 );
and ( n10038 , n10027 , n10037 );
and ( n10039 , n10025 , n10037 );
or ( n10040 , n10028 , n10038 , n10039 );
and ( n10041 , n10022 , n10040 );
and ( n10042 , n10020 , n10040 );
or ( n10043 , n10023 , n10041 , n10042 );
and ( n10044 , n10017 , n10043 );
and ( n10045 , n10015 , n10043 );
or ( n10046 , n10018 , n10044 , n10045 );
xor ( n10047 , n9889 , n10004 );
xor ( n10048 , n10047 , n10007 );
and ( n10049 , n10046 , n10048 );
xor ( n10050 , n9891 , n9893 );
xor ( n10051 , n10050 , n10001 );
xor ( n10052 , n6090 , n6550 );
buf ( n537313 , n10052 );
buf ( n537314 , n537313 );
buf ( n10055 , n537314 );
and ( n10056 , n10055 , n8106 );
and ( n10057 , n9925 , n8104 );
nor ( n10058 , n10056 , n10057 );
not ( n10059 , n10058 );
xor ( n10060 , n9903 , n9907 );
xor ( n10061 , n10060 , n9912 );
and ( n10062 , n10059 , n10061 );
and ( n10063 , n6816 , n7683 );
and ( n10064 , n7022 , n7680 );
nor ( n10065 , n10063 , n10064 );
xnor ( n10066 , n10065 , n7676 );
and ( n10067 , n7149 , n7797 );
and ( n10068 , n7879 , n7795 );
nor ( n10069 , n10067 , n10068 );
xnor ( n10070 , n10069 , n7807 );
and ( n10071 , n10066 , n10070 );
and ( n10072 , n7898 , n7036 );
and ( n10073 , n7929 , n7034 );
nor ( n10074 , n10072 , n10073 );
xnor ( n10075 , n10074 , n7125 );
and ( n10076 , n10070 , n10075 );
and ( n10077 , n10066 , n10075 );
or ( n10078 , n10071 , n10076 , n10077 );
and ( n10079 , n10061 , n10078 );
and ( n10080 , n10059 , n10078 );
or ( n10081 , n10062 , n10079 , n10080 );
and ( n10082 , n8604 , n7924 );
and ( n10083 , n8609 , n7922 );
nor ( n10084 , n10082 , n10083 );
xnor ( n10085 , n10084 , n7934 );
and ( n10086 , n9162 , n7963 );
and ( n10087 , n9084 , n7961 );
nor ( n10088 , n10086 , n10087 );
xnor ( n10089 , n10088 , n7973 );
and ( n10090 , n10085 , n10089 );
and ( n10091 , n7939 , n6722 );
and ( n10092 , n7968 , n6720 );
nor ( n10093 , n10091 , n10092 );
xnor ( n10094 , n10093 , n6821 );
and ( n10095 , n7979 , n6852 );
and ( n10096 , n8000 , n6850 );
nor ( n10097 , n10095 , n10096 );
xnor ( n10098 , n10097 , n6862 );
and ( n10099 , n10094 , n10098 );
and ( n10100 , n8071 , n7874 );
and ( n10101 , n8076 , n7872 );
nor ( n10102 , n10100 , n10101 );
xnor ( n10103 , n10102 , n7884 );
and ( n10104 , n10098 , n10103 );
and ( n10105 , n10094 , n10103 );
or ( n10106 , n10099 , n10104 , n10105 );
and ( n10107 , n10090 , n10106 );
and ( n10108 , n9482 , n7995 );
and ( n10109 , n9410 , n7993 );
nor ( n10110 , n10108 , n10109 );
xnor ( n10111 , n10110 , n8005 );
and ( n10112 , n9925 , n8253 );
and ( n10113 , n9676 , n8251 );
nor ( n10114 , n10112 , n10113 );
xnor ( n10115 , n10114 , n8259 );
and ( n10116 , n10111 , n10115 );
xor ( n10117 , n6143 , n6548 );
buf ( n537378 , n10117 );
buf ( n537379 , n537378 );
buf ( n10120 , n537379 );
and ( n10121 , n10120 , n8106 );
and ( n10122 , n10055 , n8104 );
nor ( n10123 , n10121 , n10122 );
not ( n10124 , n10123 );
and ( n10125 , n10115 , n10124 );
and ( n10126 , n10111 , n10124 );
or ( n10127 , n10116 , n10125 , n10126 );
and ( n10128 , n10106 , n10127 );
and ( n10129 , n10090 , n10127 );
or ( n10130 , n10107 , n10128 , n10129 );
and ( n10131 , n10081 , n10130 );
xor ( n10132 , n9929 , n9945 );
xor ( n10133 , n10132 , n9962 );
and ( n10134 , n10130 , n10133 );
and ( n10135 , n10081 , n10133 );
or ( n10136 , n10131 , n10134 , n10135 );
xor ( n10137 , n9896 , n9898 );
xor ( n10138 , n10137 , n9918 );
and ( n10139 , n10136 , n10138 );
xor ( n10140 , n9965 , n9989 );
xor ( n10141 , n10140 , n9992 );
and ( n10142 , n10138 , n10141 );
and ( n10143 , n10136 , n10141 );
or ( n10144 , n10139 , n10142 , n10143 );
xor ( n10145 , n9921 , n9995 );
xor ( n10146 , n10145 , n9998 );
and ( n10147 , n10144 , n10146 );
and ( n10148 , n8609 , n6923 );
and ( n10149 , n8595 , n6921 );
nor ( n10150 , n10148 , n10149 );
xnor ( n10151 , n10150 , n6933 );
and ( n10152 , n9084 , n7924 );
and ( n10153 , n8604 , n7922 );
nor ( n10154 , n10152 , n10153 );
xnor ( n10155 , n10154 , n7934 );
and ( n10156 , n10151 , n10155 );
and ( n10157 , n9410 , n7963 );
and ( n10158 , n9162 , n7961 );
nor ( n10159 , n10157 , n10158 );
xnor ( n10160 , n10159 , n7973 );
and ( n10161 , n10155 , n10160 );
and ( n10162 , n10151 , n10160 );
or ( n10163 , n10156 , n10161 , n10162 );
and ( n10164 , n8111 , n7144 );
and ( n10165 , n8245 , n7142 );
nor ( n10166 , n10164 , n10165 );
xnor ( n10167 , n10166 , n7154 );
and ( n10168 , n10163 , n10167 );
and ( n10169 , n8595 , n6923 );
and ( n10170 , n8091 , n6921 );
nor ( n10171 , n10169 , n10170 );
xnor ( n10172 , n10171 , n6933 );
and ( n10173 , n10167 , n10172 );
and ( n10174 , n10163 , n10172 );
or ( n10175 , n10168 , n10173 , n10174 );
and ( n10176 , n7879 , n7797 );
and ( n10177 , n8021 , n7795 );
nor ( n10178 , n10176 , n10177 );
xnor ( n10179 , n10178 , n7807 );
and ( n10180 , n10175 , n10179 );
and ( n10181 , n6868 , n7847 );
and ( n10182 , n6928 , n7845 );
nor ( n10183 , n10181 , n10182 );
xnor ( n10184 , n10183 , n7857 );
and ( n10185 , n10179 , n10184 );
and ( n10186 , n10175 , n10184 );
or ( n10187 , n10180 , n10185 , n10186 );
and ( n10188 , n6614 , n7732 );
and ( n10189 , n6816 , n7730 );
nor ( n10190 , n10188 , n10189 );
xnor ( n10191 , n10190 , n7742 );
and ( n10192 , n7968 , n6722 );
and ( n10193 , n7898 , n6720 );
nor ( n10194 , n10192 , n10193 );
xnor ( n10195 , n10194 , n6821 );
and ( n10196 , n10191 , n10195 );
xor ( n10197 , n9933 , n9937 );
xor ( n10198 , n10197 , n9942 );
and ( n10199 , n10195 , n10198 );
and ( n10200 , n10191 , n10198 );
or ( n10201 , n10196 , n10199 , n10200 );
and ( n10202 , n10187 , n10201 );
and ( n10203 , n7120 , n7683 );
and ( n10204 , n7852 , n7680 );
nor ( n10205 , n10203 , n10204 );
xnor ( n10206 , n10205 , n7676 );
and ( n10207 , n10201 , n10206 );
and ( n10208 , n10187 , n10206 );
or ( n10209 , n10202 , n10207 , n10208 );
xor ( n10210 , n9981 , n9983 );
xor ( n10211 , n10210 , n9986 );
xor ( n10212 , n9950 , n9954 );
xor ( n10213 , n10212 , n9959 );
xor ( n10214 , n9969 , n9973 );
xor ( n10215 , n10214 , n9978 );
and ( n10216 , n10213 , n10215 );
xor ( n10217 , n10191 , n10195 );
xor ( n10218 , n10217 , n10198 );
and ( n10219 , n10215 , n10218 );
and ( n10220 , n10213 , n10218 );
or ( n10221 , n10216 , n10219 , n10220 );
and ( n10222 , n10211 , n10221 );
xor ( n10223 , n10066 , n10070 );
xor ( n10224 , n10223 , n10075 );
xor ( n10225 , n10085 , n10089 );
and ( n10226 , n10224 , n10225 );
and ( n10227 , n6614 , n7683 );
and ( n10228 , n6816 , n7680 );
nor ( n10229 , n10227 , n10228 );
xnor ( n10230 , n10229 , n7676 );
and ( n10231 , n7879 , n7762 );
and ( n10232 , n8021 , n7760 );
nor ( n10233 , n10231 , n10232 );
xnor ( n10234 , n10233 , n7772 );
and ( n10235 , n10230 , n10234 );
and ( n10236 , n7929 , n7847 );
and ( n10237 , n8039 , n7845 );
nor ( n10238 , n10236 , n10237 );
xnor ( n10239 , n10238 , n7857 );
and ( n10240 , n10234 , n10239 );
and ( n10241 , n10230 , n10239 );
or ( n10242 , n10235 , n10240 , n10241 );
and ( n10243 , n10225 , n10242 );
and ( n10244 , n10224 , n10242 );
or ( n10245 , n10226 , n10243 , n10244 );
and ( n10246 , n6826 , n7732 );
and ( n10247 , n6857 , n7730 );
nor ( n10248 , n10246 , n10247 );
xnor ( n10249 , n10248 , n7742 );
and ( n10250 , n7130 , n7797 );
and ( n10251 , n7149 , n7795 );
nor ( n10252 , n10250 , n10251 );
xnor ( n10253 , n10252 , n7807 );
and ( n10254 , n10249 , n10253 );
and ( n10255 , n6868 , n7826 );
and ( n10256 , n6928 , n7824 );
nor ( n10257 , n10255 , n10256 );
xnor ( n10258 , n10257 , n7836 );
and ( n10259 , n8091 , n7144 );
and ( n10260 , n8111 , n7142 );
nor ( n10261 , n10259 , n10260 );
xnor ( n10262 , n10261 , n7154 );
and ( n10263 , n10258 , n10262 );
and ( n10264 , n9676 , n7995 );
and ( n10265 , n9482 , n7993 );
nor ( n10266 , n10264 , n10265 );
xnor ( n10267 , n10266 , n8005 );
and ( n10268 , n10262 , n10267 );
and ( n10269 , n10258 , n10267 );
or ( n10270 , n10263 , n10268 , n10269 );
and ( n10271 , n10254 , n10270 );
xor ( n10272 , n10094 , n10098 );
xor ( n10273 , n10272 , n10103 );
and ( n10274 , n10270 , n10273 );
and ( n10275 , n10254 , n10273 );
or ( n10276 , n10271 , n10274 , n10275 );
and ( n10277 , n10245 , n10276 );
xor ( n10278 , n10059 , n10061 );
xor ( n10279 , n10278 , n10078 );
and ( n10280 , n10276 , n10279 );
and ( n10281 , n10245 , n10279 );
or ( n10282 , n10277 , n10280 , n10281 );
and ( n10283 , n10221 , n10282 );
and ( n10284 , n10211 , n10282 );
or ( n10285 , n10222 , n10283 , n10284 );
and ( n10286 , n10209 , n10285 );
xor ( n10287 , n10025 , n10027 );
xor ( n10288 , n10287 , n10037 );
and ( n10289 , n10285 , n10288 );
and ( n10290 , n10209 , n10288 );
or ( n10291 , n10286 , n10289 , n10290 );
and ( n10292 , n10146 , n10291 );
and ( n10293 , n10144 , n10291 );
or ( n10294 , n10147 , n10292 , n10293 );
and ( n10295 , n10051 , n10294 );
xor ( n10296 , n10015 , n10017 );
xor ( n10297 , n10296 , n10043 );
and ( n10298 , n10294 , n10297 );
and ( n10299 , n10051 , n10297 );
or ( n10300 , n10295 , n10298 , n10299 );
and ( n10301 , n10048 , n10300 );
and ( n10302 , n10046 , n10300 );
or ( n10303 , n10049 , n10301 , n10302 );
and ( n10304 , n10012 , n10303 );
and ( n10305 , n10010 , n10303 );
or ( n10306 , n10013 , n10304 , n10305 );
and ( n10307 , n9886 , n10306 );
and ( n10308 , n9884 , n10306 );
or ( n10309 , n9887 , n10307 , n10308 );
and ( n10310 , n9734 , n10309 );
xor ( n10311 , n9734 , n10309 );
xor ( n10312 , n9884 , n9886 );
xor ( n10313 , n10312 , n10306 );
xor ( n10314 , n10010 , n10012 );
xor ( n10315 , n10314 , n10303 );
xor ( n10316 , n10046 , n10048 );
xor ( n10317 , n10316 , n10300 );
xor ( n10318 , n10020 , n10022 );
xor ( n10319 , n10318 , n10040 );
xor ( n10320 , n10136 , n10138 );
xor ( n10321 , n10320 , n10141 );
xor ( n10322 , n10030 , n10032 );
xor ( n10323 , n10322 , n10034 );
xor ( n10324 , n10081 , n10130 );
xor ( n10325 , n10324 , n10133 );
and ( n10326 , n10323 , n10325 );
xor ( n10327 , n10187 , n10201 );
xor ( n10328 , n10327 , n10206 );
and ( n10329 , n10325 , n10328 );
and ( n10330 , n10323 , n10328 );
or ( n10331 , n10326 , n10329 , n10330 );
and ( n10332 , n10321 , n10331 );
and ( n10333 , n8604 , n6923 );
and ( n10334 , n8609 , n6921 );
nor ( n10335 , n10333 , n10334 );
xnor ( n10336 , n10335 , n6933 );
and ( n10337 , n9162 , n7924 );
and ( n10338 , n9084 , n7922 );
nor ( n10339 , n10337 , n10338 );
xnor ( n10340 , n10339 , n7934 );
and ( n10341 , n10336 , n10340 );
and ( n10342 , n9482 , n7963 );
and ( n10343 , n9410 , n7961 );
nor ( n10344 , n10342 , n10343 );
xnor ( n10345 , n10344 , n7973 );
and ( n10346 , n10340 , n10345 );
and ( n10347 , n10336 , n10345 );
or ( n10348 , n10341 , n10346 , n10347 );
and ( n10349 , n8000 , n6722 );
and ( n10350 , n7939 , n6720 );
nor ( n10351 , n10349 , n10350 );
xnor ( n10352 , n10351 , n6821 );
and ( n10353 , n10348 , n10352 );
and ( n10354 , n8245 , n7874 );
and ( n10355 , n8071 , n7872 );
nor ( n10356 , n10354 , n10355 );
xnor ( n10357 , n10356 , n7884 );
and ( n10358 , n10352 , n10357 );
and ( n10359 , n10348 , n10357 );
or ( n10360 , n10353 , n10358 , n10359 );
and ( n10361 , n6857 , n7732 );
and ( n10362 , n6614 , n7730 );
nor ( n10363 , n10361 , n10362 );
xnor ( n10364 , n10363 , n7742 );
and ( n10365 , n10360 , n10364 );
and ( n10366 , n8021 , n7762 );
and ( n10367 , n6826 , n7760 );
nor ( n10368 , n10366 , n10367 );
xnor ( n10369 , n10368 , n7772 );
and ( n10370 , n10364 , n10369 );
and ( n10371 , n10360 , n10369 );
or ( n10372 , n10365 , n10370 , n10371 );
and ( n10373 , n6928 , n7826 );
and ( n10374 , n7130 , n7824 );
nor ( n10375 , n10373 , n10374 );
xnor ( n10376 , n10375 , n7836 );
and ( n10377 , n8039 , n7847 );
and ( n10378 , n6868 , n7845 );
nor ( n10379 , n10377 , n10378 );
xnor ( n10380 , n10379 , n7857 );
and ( n10381 , n10376 , n10380 );
xor ( n10382 , n10163 , n10167 );
xor ( n10383 , n10382 , n10172 );
and ( n10384 , n10380 , n10383 );
and ( n10385 , n10376 , n10383 );
or ( n10386 , n10381 , n10384 , n10385 );
and ( n10387 , n10372 , n10386 );
xor ( n10388 , n10175 , n10179 );
xor ( n10389 , n10388 , n10184 );
and ( n10390 , n10386 , n10389 );
and ( n10391 , n10372 , n10389 );
or ( n10392 , n10387 , n10390 , n10391 );
xor ( n10393 , n10090 , n10106 );
xor ( n10394 , n10393 , n10127 );
xor ( n10395 , n10111 , n10115 );
xor ( n10396 , n10395 , n10124 );
and ( n10397 , n7968 , n7036 );
and ( n10398 , n7898 , n7034 );
nor ( n10399 , n10397 , n10398 );
xnor ( n10400 , n10399 , n7125 );
and ( n10401 , n8076 , n6852 );
and ( n10402 , n7979 , n6850 );
nor ( n10403 , n10401 , n10402 );
xnor ( n10404 , n10403 , n6862 );
and ( n10405 , n10400 , n10404 );
xor ( n10406 , n10151 , n10155 );
xor ( n10407 , n10406 , n10160 );
and ( n10408 , n10404 , n10407 );
and ( n10409 , n10400 , n10407 );
or ( n10410 , n10405 , n10408 , n10409 );
and ( n10411 , n10396 , n10410 );
and ( n10412 , n10055 , n8253 );
and ( n10413 , n9925 , n8251 );
nor ( n10414 , n10412 , n10413 );
xnor ( n10415 , n10414 , n8259 );
xor ( n10416 , n6195 , n6546 );
buf ( n537677 , n10416 );
buf ( n537678 , n537677 );
buf ( n10419 , n537678 );
and ( n10420 , n10419 , n8106 );
and ( n10421 , n10120 , n8104 );
nor ( n10422 , n10420 , n10421 );
not ( n10423 , n10422 );
and ( n10424 , n10415 , n10423 );
xor ( n10425 , n10230 , n10234 );
xor ( n10426 , n10425 , n10239 );
and ( n10427 , n10423 , n10426 );
and ( n10428 , n10415 , n10426 );
or ( n10429 , n10424 , n10427 , n10428 );
and ( n10430 , n10410 , n10429 );
and ( n10431 , n10396 , n10429 );
or ( n10432 , n10411 , n10430 , n10431 );
and ( n10433 , n10394 , n10432 );
xor ( n10434 , n10249 , n10253 );
and ( n10435 , n6857 , n7683 );
and ( n10436 , n6614 , n7680 );
nor ( n10437 , n10435 , n10436 );
xnor ( n10438 , n10437 , n7676 );
and ( n10439 , n8021 , n7732 );
and ( n10440 , n6826 , n7730 );
nor ( n10441 , n10439 , n10440 );
xnor ( n10442 , n10441 , n7742 );
and ( n10443 , n10438 , n10442 );
and ( n10444 , n7149 , n7762 );
and ( n10445 , n7879 , n7760 );
nor ( n10446 , n10444 , n10445 );
xnor ( n10447 , n10446 , n7772 );
and ( n10448 , n10442 , n10447 );
and ( n10449 , n10438 , n10447 );
or ( n10450 , n10443 , n10448 , n10449 );
and ( n10451 , n10434 , n10450 );
and ( n10452 , n6928 , n7797 );
and ( n10453 , n7130 , n7795 );
nor ( n10454 , n10452 , n10453 );
xnor ( n10455 , n10454 , n7807 );
and ( n10456 , n8039 , n7826 );
and ( n10457 , n6868 , n7824 );
nor ( n10458 , n10456 , n10457 );
xnor ( n10459 , n10458 , n7836 );
and ( n10460 , n10455 , n10459 );
and ( n10461 , n7898 , n7847 );
and ( n10462 , n7929 , n7845 );
nor ( n10463 , n10461 , n10462 );
xnor ( n10464 , n10463 , n7857 );
and ( n10465 , n10459 , n10464 );
and ( n10466 , n10455 , n10464 );
or ( n10467 , n10460 , n10465 , n10466 );
and ( n10468 , n10450 , n10467 );
and ( n10469 , n10434 , n10467 );
or ( n10470 , n10451 , n10468 , n10469 );
and ( n10471 , n7979 , n6722 );
and ( n10472 , n8000 , n6720 );
nor ( n10473 , n10471 , n10472 );
xnor ( n10474 , n10473 , n6821 );
and ( n10475 , n8111 , n7874 );
and ( n10476 , n8245 , n7872 );
nor ( n10477 , n10475 , n10476 );
xnor ( n10478 , n10477 , n7884 );
and ( n10479 , n10474 , n10478 );
and ( n10480 , n8595 , n7144 );
and ( n10481 , n8091 , n7142 );
nor ( n10482 , n10480 , n10481 );
xnor ( n10483 , n10482 , n7154 );
and ( n10484 , n10478 , n10483 );
and ( n10485 , n10474 , n10483 );
or ( n10486 , n10479 , n10484 , n10485 );
and ( n10487 , n9925 , n7995 );
and ( n10488 , n9676 , n7993 );
nor ( n10489 , n10487 , n10488 );
xnor ( n10490 , n10489 , n8005 );
and ( n10491 , n10120 , n8253 );
and ( n10492 , n10055 , n8251 );
nor ( n10493 , n10491 , n10492 );
xnor ( n10494 , n10493 , n8259 );
and ( n10495 , n10490 , n10494 );
xor ( n10496 , n6228 , n6544 );
buf ( n537757 , n10496 );
buf ( n537758 , n537757 );
buf ( n10499 , n537758 );
and ( n10500 , n10499 , n8106 );
and ( n10501 , n10419 , n8104 );
nor ( n10502 , n10500 , n10501 );
not ( n10503 , n10502 );
and ( n10504 , n10494 , n10503 );
and ( n10505 , n10490 , n10503 );
or ( n10506 , n10495 , n10504 , n10505 );
and ( n10507 , n10486 , n10506 );
xor ( n10508 , n10258 , n10262 );
xor ( n10509 , n10508 , n10267 );
and ( n10510 , n10506 , n10509 );
and ( n10511 , n10486 , n10509 );
or ( n10512 , n10507 , n10510 , n10511 );
and ( n10513 , n10470 , n10512 );
xor ( n10514 , n10224 , n10225 );
xor ( n10515 , n10514 , n10242 );
and ( n10516 , n10512 , n10515 );
and ( n10517 , n10470 , n10515 );
or ( n10518 , n10513 , n10516 , n10517 );
and ( n10519 , n10432 , n10518 );
and ( n10520 , n10394 , n10518 );
or ( n10521 , n10433 , n10519 , n10520 );
and ( n10522 , n10392 , n10521 );
xor ( n10523 , n10211 , n10221 );
xor ( n10524 , n10523 , n10282 );
and ( n10525 , n10521 , n10524 );
and ( n10526 , n10392 , n10524 );
or ( n10527 , n10522 , n10525 , n10526 );
and ( n10528 , n10331 , n10527 );
and ( n10529 , n10321 , n10527 );
or ( n10530 , n10332 , n10528 , n10529 );
and ( n10531 , n10319 , n10530 );
xor ( n10532 , n10144 , n10146 );
xor ( n10533 , n10532 , n10291 );
and ( n10534 , n10530 , n10533 );
and ( n10535 , n10319 , n10533 );
or ( n10536 , n10531 , n10534 , n10535 );
xor ( n10537 , n10051 , n10294 );
xor ( n10538 , n10537 , n10297 );
and ( n10539 , n10536 , n10538 );
xor ( n10540 , n10536 , n10538 );
xor ( n10541 , n10209 , n10285 );
xor ( n10542 , n10541 , n10288 );
xor ( n10543 , n10213 , n10215 );
xor ( n10544 , n10543 , n10218 );
xor ( n10545 , n10245 , n10276 );
xor ( n10546 , n10545 , n10279 );
and ( n10547 , n10544 , n10546 );
xor ( n10548 , n10372 , n10386 );
xor ( n10549 , n10548 , n10389 );
and ( n10550 , n10546 , n10549 );
and ( n10551 , n10544 , n10549 );
or ( n10552 , n10547 , n10550 , n10551 );
xor ( n10553 , n10254 , n10270 );
xor ( n10554 , n10553 , n10273 );
xor ( n10555 , n10360 , n10364 );
xor ( n10556 , n10555 , n10369 );
and ( n10557 , n10554 , n10556 );
xor ( n10558 , n10376 , n10380 );
xor ( n10559 , n10558 , n10383 );
and ( n10560 , n10556 , n10559 );
and ( n10561 , n10554 , n10559 );
or ( n10562 , n10557 , n10560 , n10561 );
and ( n10563 , n7939 , n7036 );
and ( n10564 , n7968 , n7034 );
nor ( n10565 , n10563 , n10564 );
xnor ( n10566 , n10565 , n7125 );
and ( n10567 , n8071 , n6852 );
and ( n10568 , n8076 , n6850 );
nor ( n10569 , n10567 , n10568 );
xnor ( n10570 , n10569 , n6862 );
and ( n10571 , n10566 , n10570 );
xor ( n10572 , n10336 , n10340 );
xor ( n10573 , n10572 , n10345 );
and ( n10574 , n10570 , n10573 );
and ( n10575 , n10566 , n10573 );
or ( n10576 , n10571 , n10574 , n10575 );
xor ( n10577 , n10348 , n10352 );
xor ( n10578 , n10577 , n10357 );
and ( n10579 , n10576 , n10578 );
xor ( n10580 , n10400 , n10404 );
xor ( n10581 , n10580 , n10407 );
and ( n10582 , n10578 , n10581 );
and ( n10583 , n10576 , n10581 );
or ( n10584 , n10579 , n10582 , n10583 );
and ( n10585 , n9084 , n6923 );
and ( n10586 , n8604 , n6921 );
nor ( n10587 , n10585 , n10586 );
xnor ( n10588 , n10587 , n6933 );
and ( n10589 , n9410 , n7924 );
and ( n10590 , n9162 , n7922 );
nor ( n10591 , n10589 , n10590 );
xnor ( n10592 , n10591 , n7934 );
and ( n10593 , n10588 , n10592 );
and ( n10594 , n9676 , n7963 );
and ( n10595 , n9482 , n7961 );
nor ( n10596 , n10594 , n10595 );
xnor ( n10597 , n10596 , n7973 );
and ( n10598 , n10592 , n10597 );
and ( n10599 , n10588 , n10597 );
or ( n10600 , n10593 , n10598 , n10599 );
and ( n10601 , n6826 , n7683 );
and ( n10602 , n6857 , n7680 );
nor ( n10603 , n10601 , n10602 );
xnor ( n10604 , n10603 , n7676 );
and ( n10605 , n7879 , n7732 );
and ( n10606 , n8021 , n7730 );
nor ( n10607 , n10605 , n10606 );
xnor ( n10608 , n10607 , n7742 );
and ( n10609 , n10604 , n10608 );
and ( n10610 , n7130 , n7762 );
and ( n10611 , n7149 , n7760 );
nor ( n10612 , n10610 , n10611 );
xnor ( n10613 , n10612 , n7772 );
and ( n10614 , n10608 , n10613 );
and ( n10615 , n10604 , n10613 );
or ( n10616 , n10609 , n10614 , n10615 );
and ( n10617 , n10600 , n10616 );
and ( n10618 , n6868 , n7797 );
and ( n10619 , n6928 , n7795 );
nor ( n10620 , n10618 , n10619 );
xnor ( n10621 , n10620 , n7807 );
and ( n10622 , n7929 , n7826 );
and ( n10623 , n8039 , n7824 );
nor ( n10624 , n10622 , n10623 );
xnor ( n10625 , n10624 , n7836 );
and ( n10626 , n10621 , n10625 );
and ( n10627 , n7968 , n7847 );
and ( n10628 , n7898 , n7845 );
nor ( n10629 , n10627 , n10628 );
xnor ( n10630 , n10629 , n7857 );
and ( n10631 , n10625 , n10630 );
and ( n10632 , n10621 , n10630 );
or ( n10633 , n10626 , n10631 , n10632 );
and ( n10634 , n10616 , n10633 );
and ( n10635 , n10600 , n10633 );
or ( n10636 , n10617 , n10634 , n10635 );
and ( n10637 , n8000 , n7036 );
and ( n10638 , n7939 , n7034 );
nor ( n10639 , n10637 , n10638 );
xnor ( n10640 , n10639 , n7125 );
and ( n10641 , n8245 , n6852 );
and ( n10642 , n8071 , n6850 );
nor ( n10643 , n10641 , n10642 );
xnor ( n10644 , n10643 , n6862 );
and ( n10645 , n10640 , n10644 );
and ( n10646 , n8091 , n7874 );
and ( n10647 , n8111 , n7872 );
nor ( n10648 , n10646 , n10647 );
xnor ( n10649 , n10648 , n7884 );
and ( n10650 , n10644 , n10649 );
and ( n10651 , n10640 , n10649 );
or ( n10652 , n10645 , n10650 , n10651 );
and ( n10653 , n8609 , n7144 );
and ( n10654 , n8595 , n7142 );
nor ( n10655 , n10653 , n10654 );
xnor ( n10656 , n10655 , n7154 );
and ( n10657 , n10055 , n7995 );
and ( n10658 , n9925 , n7993 );
nor ( n10659 , n10657 , n10658 );
xnor ( n10660 , n10659 , n8005 );
and ( n10661 , n10656 , n10660 );
and ( n10662 , n10419 , n8253 );
and ( n10663 , n10120 , n8251 );
nor ( n10664 , n10662 , n10663 );
xnor ( n10665 , n10664 , n8259 );
and ( n10666 , n10660 , n10665 );
and ( n10667 , n10656 , n10665 );
or ( n10668 , n10661 , n10666 , n10667 );
and ( n10669 , n10652 , n10668 );
xor ( n10670 , n10438 , n10442 );
xor ( n10671 , n10670 , n10447 );
and ( n10672 , n10668 , n10671 );
and ( n10673 , n10652 , n10671 );
or ( n10674 , n10669 , n10672 , n10673 );
and ( n10675 , n10636 , n10674 );
xor ( n10676 , n10455 , n10459 );
xor ( n10677 , n10676 , n10464 );
xor ( n10678 , n10474 , n10478 );
xor ( n10679 , n10678 , n10483 );
and ( n10680 , n10677 , n10679 );
xor ( n10681 , n10490 , n10494 );
xor ( n10682 , n10681 , n10503 );
and ( n10683 , n10679 , n10682 );
and ( n10684 , n10677 , n10682 );
or ( n10685 , n10680 , n10683 , n10684 );
and ( n10686 , n10674 , n10685 );
and ( n10687 , n10636 , n10685 );
or ( n10688 , n10675 , n10686 , n10687 );
and ( n10689 , n10584 , n10688 );
xor ( n10690 , n10415 , n10423 );
xor ( n10691 , n10690 , n10426 );
xor ( n10692 , n10434 , n10450 );
xor ( n10693 , n10692 , n10467 );
and ( n10694 , n10691 , n10693 );
xor ( n10695 , n10486 , n10506 );
xor ( n10696 , n10695 , n10509 );
and ( n10697 , n10693 , n10696 );
and ( n10698 , n10691 , n10696 );
or ( n10699 , n10694 , n10697 , n10698 );
and ( n10700 , n10688 , n10699 );
and ( n10701 , n10584 , n10699 );
or ( n10702 , n10689 , n10700 , n10701 );
and ( n10703 , n10562 , n10702 );
xor ( n10704 , n10394 , n10432 );
xor ( n10705 , n10704 , n10518 );
and ( n10706 , n10702 , n10705 );
and ( n10707 , n10562 , n10705 );
or ( n10708 , n10703 , n10706 , n10707 );
and ( n10709 , n10552 , n10708 );
xor ( n10710 , n10323 , n10325 );
xor ( n10711 , n10710 , n10328 );
and ( n10712 , n10708 , n10711 );
and ( n10713 , n10552 , n10711 );
or ( n10714 , n10709 , n10712 , n10713 );
and ( n10715 , n10542 , n10714 );
xor ( n10716 , n10321 , n10331 );
xor ( n10717 , n10716 , n10527 );
and ( n10718 , n10714 , n10717 );
and ( n10719 , n10542 , n10717 );
or ( n10720 , n10715 , n10718 , n10719 );
xor ( n10721 , n10319 , n10530 );
xor ( n10722 , n10721 , n10533 );
and ( n10723 , n10720 , n10722 );
xor ( n10724 , n10720 , n10722 );
xor ( n10725 , n10392 , n10521 );
xor ( n10726 , n10725 , n10524 );
xor ( n10727 , n10396 , n10410 );
xor ( n10728 , n10727 , n10429 );
xor ( n10729 , n10470 , n10512 );
xor ( n10730 , n10729 , n10515 );
and ( n10731 , n10728 , n10730 );
xor ( n10732 , n10576 , n10578 );
xor ( n10733 , n10732 , n10581 );
xor ( n10734 , n10566 , n10570 );
xor ( n10735 , n10734 , n10573 );
and ( n10736 , n8076 , n6722 );
and ( n10737 , n7979 , n6720 );
nor ( n10738 , n10736 , n10737 );
xnor ( n10739 , n10738 , n6821 );
xor ( n10740 , n10588 , n10592 );
xor ( n10741 , n10740 , n10597 );
and ( n10742 , n10739 , n10741 );
and ( n10743 , n10735 , n10742 );
xor ( n10744 , n6274 , n6542 );
buf ( n538005 , n10744 );
buf ( n538006 , n538005 );
buf ( n10747 , n538006 );
and ( n10748 , n10747 , n8106 );
and ( n10749 , n10499 , n8104 );
nor ( n10750 , n10748 , n10749 );
not ( n10751 , n10750 );
and ( n10752 , n8039 , n7797 );
and ( n10753 , n6868 , n7795 );
nor ( n10754 , n10752 , n10753 );
xnor ( n10755 , n10754 , n7807 );
and ( n10756 , n7898 , n7826 );
and ( n10757 , n7929 , n7824 );
nor ( n10758 , n10756 , n10757 );
xnor ( n10759 , n10758 , n7836 );
and ( n10760 , n10755 , n10759 );
and ( n10761 , n7939 , n7847 );
and ( n10762 , n7968 , n7845 );
nor ( n10763 , n10761 , n10762 );
xnor ( n10764 , n10763 , n7857 );
and ( n10765 , n10759 , n10764 );
and ( n10766 , n10755 , n10764 );
or ( n10767 , n10760 , n10765 , n10766 );
and ( n10768 , n10751 , n10767 );
and ( n10769 , n8604 , n7144 );
and ( n10770 , n8609 , n7142 );
nor ( n10771 , n10769 , n10770 );
xnor ( n10772 , n10771 , n7154 );
and ( n10773 , n9162 , n6923 );
and ( n10774 , n9084 , n6921 );
nor ( n10775 , n10773 , n10774 );
xnor ( n10776 , n10775 , n6933 );
and ( n10777 , n10772 , n10776 );
and ( n10778 , n10767 , n10777 );
and ( n10779 , n10751 , n10777 );
or ( n10780 , n10768 , n10778 , n10779 );
and ( n10781 , n10742 , n10780 );
and ( n10782 , n10735 , n10780 );
or ( n10783 , n10743 , n10781 , n10782 );
and ( n10784 , n10733 , n10783 );
and ( n10785 , n8111 , n6852 );
and ( n10786 , n8245 , n6850 );
nor ( n10787 , n10785 , n10786 );
xnor ( n10788 , n10787 , n6862 );
and ( n10789 , n8595 , n7874 );
and ( n10790 , n8091 , n7872 );
nor ( n10791 , n10789 , n10790 );
xnor ( n10792 , n10791 , n7884 );
and ( n10793 , n10788 , n10792 );
and ( n10794 , n8021 , n7683 );
and ( n10795 , n6826 , n7680 );
nor ( n10796 , n10794 , n10795 );
xnor ( n10797 , n10796 , n7676 );
and ( n10798 , n6928 , n7762 );
and ( n10799 , n7130 , n7760 );
nor ( n10800 , n10798 , n10799 );
xnor ( n10801 , n10800 , n7772 );
and ( n10802 , n10797 , n10801 );
and ( n10803 , n7979 , n7036 );
and ( n10804 , n8000 , n7034 );
nor ( n10805 , n10803 , n10804 );
xnor ( n10806 , n10805 , n7125 );
and ( n10807 , n10801 , n10806 );
and ( n10808 , n10797 , n10806 );
or ( n10809 , n10802 , n10807 , n10808 );
and ( n10810 , n10793 , n10809 );
and ( n10811 , n8071 , n6722 );
and ( n10812 , n8076 , n6720 );
nor ( n10813 , n10811 , n10812 );
xnor ( n10814 , n10813 , n6821 );
and ( n10815 , n9482 , n7924 );
and ( n10816 , n9410 , n7922 );
nor ( n10817 , n10815 , n10816 );
xnor ( n10818 , n10817 , n7934 );
and ( n10819 , n10814 , n10818 );
and ( n10820 , n9925 , n7963 );
and ( n10821 , n9676 , n7961 );
nor ( n10822 , n10820 , n10821 );
xnor ( n10823 , n10822 , n7973 );
and ( n10824 , n10818 , n10823 );
and ( n10825 , n10814 , n10823 );
or ( n10826 , n10819 , n10824 , n10825 );
and ( n10827 , n10809 , n10826 );
and ( n10828 , n10793 , n10826 );
or ( n10829 , n10810 , n10827 , n10828 );
and ( n10830 , n10120 , n7995 );
and ( n10831 , n10055 , n7993 );
nor ( n10832 , n10830 , n10831 );
xnor ( n10833 , n10832 , n8005 );
and ( n10834 , n10499 , n8253 );
and ( n10835 , n10419 , n8251 );
nor ( n10836 , n10834 , n10835 );
xnor ( n10837 , n10836 , n8259 );
and ( n10838 , n10833 , n10837 );
xor ( n10839 , n6316 , n6540 );
buf ( n538100 , n10839 );
buf ( n538101 , n538100 );
buf ( n10842 , n538101 );
and ( n10843 , n10842 , n8106 );
and ( n10844 , n10747 , n8104 );
nor ( n10845 , n10843 , n10844 );
not ( n10846 , n10845 );
and ( n10847 , n10837 , n10846 );
and ( n10848 , n10833 , n10846 );
or ( n10849 , n10838 , n10847 , n10848 );
xor ( n10850 , n10604 , n10608 );
xor ( n10851 , n10850 , n10613 );
and ( n10852 , n10849 , n10851 );
xor ( n10853 , n10621 , n10625 );
xor ( n10854 , n10853 , n10630 );
and ( n10855 , n10851 , n10854 );
and ( n10856 , n10849 , n10854 );
or ( n10857 , n10852 , n10855 , n10856 );
and ( n10858 , n10829 , n10857 );
xor ( n10859 , n10600 , n10616 );
xor ( n10860 , n10859 , n10633 );
and ( n10861 , n10857 , n10860 );
and ( n10862 , n10829 , n10860 );
or ( n10863 , n10858 , n10861 , n10862 );
and ( n10864 , n10783 , n10863 );
and ( n10865 , n10733 , n10863 );
or ( n10866 , n10784 , n10864 , n10865 );
and ( n10867 , n10730 , n10866 );
and ( n10868 , n10728 , n10866 );
or ( n10869 , n10731 , n10867 , n10868 );
xor ( n10870 , n10544 , n10546 );
xor ( n10871 , n10870 , n10549 );
and ( n10872 , n10869 , n10871 );
xor ( n10873 , n10562 , n10702 );
xor ( n10874 , n10873 , n10705 );
and ( n10875 , n10871 , n10874 );
and ( n10876 , n10869 , n10874 );
or ( n10877 , n10872 , n10875 , n10876 );
and ( n10878 , n10726 , n10877 );
xor ( n10879 , n10552 , n10708 );
xor ( n10880 , n10879 , n10711 );
and ( n10881 , n10877 , n10880 );
and ( n10882 , n10726 , n10880 );
or ( n10883 , n10878 , n10881 , n10882 );
xor ( n10884 , n10542 , n10714 );
xor ( n10885 , n10884 , n10717 );
and ( n10886 , n10883 , n10885 );
xor ( n10887 , n10883 , n10885 );
xor ( n10888 , n10726 , n10877 );
xor ( n10889 , n10888 , n10880 );
xor ( n10890 , n10554 , n10556 );
xor ( n10891 , n10890 , n10559 );
xor ( n10892 , n10584 , n10688 );
xor ( n10893 , n10892 , n10699 );
and ( n10894 , n10891 , n10893 );
xor ( n10895 , n10636 , n10674 );
xor ( n10896 , n10895 , n10685 );
xor ( n10897 , n10691 , n10693 );
xor ( n10898 , n10897 , n10696 );
and ( n10899 , n10896 , n10898 );
xor ( n10900 , n10652 , n10668 );
xor ( n10901 , n10900 , n10671 );
xor ( n10902 , n10677 , n10679 );
xor ( n10903 , n10902 , n10682 );
and ( n10904 , n10901 , n10903 );
xor ( n10905 , n10640 , n10644 );
xor ( n10906 , n10905 , n10649 );
xor ( n10907 , n10656 , n10660 );
xor ( n10908 , n10907 , n10665 );
and ( n10909 , n10906 , n10908 );
xor ( n10910 , n10739 , n10741 );
and ( n10911 , n10908 , n10910 );
and ( n10912 , n10906 , n10910 );
or ( n10913 , n10909 , n10911 , n10912 );
and ( n10914 , n10903 , n10913 );
and ( n10915 , n10901 , n10913 );
or ( n10916 , n10904 , n10914 , n10915 );
and ( n10917 , n10898 , n10916 );
and ( n10918 , n10896 , n10916 );
or ( n10919 , n10899 , n10917 , n10918 );
and ( n10920 , n10893 , n10919 );
and ( n10921 , n10891 , n10919 );
or ( n10922 , n10894 , n10920 , n10921 );
xor ( n10923 , n10869 , n10871 );
xor ( n10924 , n10923 , n10874 );
and ( n10925 , n10922 , n10924 );
xor ( n10926 , n10728 , n10730 );
xor ( n10927 , n10926 , n10866 );
xor ( n10928 , n10755 , n10759 );
xor ( n10929 , n10928 , n10764 );
xor ( n10930 , n10772 , n10776 );
and ( n10931 , n10929 , n10930 );
xor ( n10932 , n10788 , n10792 );
and ( n10933 , n10930 , n10932 );
and ( n10934 , n10929 , n10932 );
or ( n10935 , n10931 , n10933 , n10934 );
and ( n10936 , n8609 , n7874 );
and ( n10937 , n8595 , n7872 );
nor ( n10938 , n10936 , n10937 );
xnor ( n10939 , n10938 , n7884 );
and ( n10940 , n9084 , n7144 );
and ( n10941 , n8604 , n7142 );
nor ( n10942 , n10940 , n10941 );
xnor ( n10943 , n10942 , n7154 );
and ( n10944 , n10939 , n10943 );
and ( n10945 , n9410 , n6923 );
and ( n10946 , n9162 , n6921 );
nor ( n10947 , n10945 , n10946 );
xnor ( n10948 , n10947 , n6933 );
and ( n10949 , n10943 , n10948 );
and ( n10950 , n10939 , n10948 );
or ( n10951 , n10944 , n10949 , n10950 );
and ( n10952 , n9676 , n7924 );
and ( n10953 , n9482 , n7922 );
nor ( n10954 , n10952 , n10953 );
xnor ( n10955 , n10954 , n7934 );
and ( n10956 , n10419 , n7995 );
and ( n10957 , n10120 , n7993 );
nor ( n10958 , n10956 , n10957 );
xnor ( n10959 , n10958 , n8005 );
and ( n10960 , n10955 , n10959 );
and ( n10961 , n10951 , n10960 );
and ( n10962 , n7130 , n7732 );
and ( n10963 , n7149 , n7730 );
nor ( n10964 , n10962 , n10963 );
xnor ( n10965 , n10964 , n7742 );
and ( n10966 , n7929 , n7797 );
and ( n10967 , n8039 , n7795 );
nor ( n10968 , n10966 , n10967 );
xnor ( n10969 , n10968 , n7807 );
and ( n10970 , n10965 , n10969 );
and ( n10971 , n10960 , n10970 );
and ( n10972 , n10951 , n10970 );
or ( n10973 , n10961 , n10971 , n10972 );
and ( n10974 , n10935 , n10973 );
and ( n10975 , n7879 , n7683 );
and ( n10976 , n8021 , n7680 );
nor ( n10977 , n10975 , n10976 );
xnor ( n10978 , n10977 , n7676 );
and ( n10979 , n6868 , n7762 );
and ( n10980 , n6928 , n7760 );
nor ( n10981 , n10979 , n10980 );
xnor ( n10982 , n10981 , n7772 );
and ( n10983 , n10978 , n10982 );
and ( n10984 , n7968 , n7826 );
and ( n10985 , n7898 , n7824 );
nor ( n10986 , n10984 , n10985 );
xnor ( n10987 , n10986 , n7836 );
and ( n10988 , n10982 , n10987 );
and ( n10989 , n10978 , n10987 );
or ( n10990 , n10983 , n10988 , n10989 );
and ( n10991 , n8245 , n6722 );
and ( n10992 , n8071 , n6720 );
nor ( n10993 , n10991 , n10992 );
xnor ( n10994 , n10993 , n6821 );
and ( n10995 , n8091 , n6852 );
and ( n10996 , n8111 , n6850 );
nor ( n10997 , n10995 , n10996 );
xnor ( n10998 , n10997 , n6862 );
and ( n10999 , n10994 , n10998 );
and ( n11000 , n10055 , n7963 );
and ( n11001 , n9925 , n7961 );
nor ( n11002 , n11000 , n11001 );
xnor ( n11003 , n11002 , n7973 );
and ( n11004 , n10998 , n11003 );
and ( n11005 , n10994 , n11003 );
or ( n11006 , n10999 , n11004 , n11005 );
and ( n11007 , n10990 , n11006 );
xor ( n11008 , n10797 , n10801 );
xor ( n11009 , n11008 , n10806 );
and ( n11010 , n11006 , n11009 );
and ( n11011 , n10990 , n11009 );
or ( n11012 , n11007 , n11010 , n11011 );
and ( n11013 , n10973 , n11012 );
and ( n11014 , n10935 , n11012 );
or ( n11015 , n10974 , n11013 , n11014 );
xor ( n11016 , n10751 , n10767 );
xor ( n11017 , n11016 , n10777 );
xor ( n11018 , n10793 , n10809 );
xor ( n11019 , n11018 , n10826 );
and ( n11020 , n11017 , n11019 );
xor ( n11021 , n10849 , n10851 );
xor ( n11022 , n11021 , n10854 );
and ( n11023 , n11019 , n11022 );
and ( n11024 , n11017 , n11022 );
or ( n11025 , n11020 , n11023 , n11024 );
and ( n11026 , n11015 , n11025 );
xor ( n11027 , n10735 , n10742 );
xor ( n11028 , n11027 , n10780 );
and ( n11029 , n11025 , n11028 );
and ( n11030 , n11015 , n11028 );
or ( n11031 , n11026 , n11029 , n11030 );
xor ( n11032 , n10733 , n10783 );
xor ( n11033 , n11032 , n10863 );
and ( n11034 , n11031 , n11033 );
xor ( n11035 , n10829 , n10857 );
xor ( n11036 , n11035 , n10860 );
and ( n11037 , n8000 , n7847 );
and ( n11038 , n7939 , n7845 );
nor ( n11039 , n11037 , n11038 );
xnor ( n11040 , n11039 , n7857 );
and ( n11041 , n8076 , n7036 );
and ( n11042 , n7979 , n7034 );
nor ( n11043 , n11041 , n11042 );
xnor ( n11044 , n11043 , n7125 );
and ( n11045 , n11040 , n11044 );
xor ( n11046 , n10939 , n10943 );
xor ( n11047 , n11046 , n10948 );
and ( n11048 , n11044 , n11047 );
and ( n11049 , n11040 , n11047 );
or ( n11050 , n11045 , n11048 , n11049 );
and ( n11051 , n7149 , n7732 );
and ( n11052 , n7879 , n7730 );
nor ( n11053 , n11051 , n11052 );
xnor ( n11054 , n11053 , n7742 );
and ( n11055 , n11050 , n11054 );
xor ( n11056 , n10814 , n10818 );
xor ( n11057 , n11056 , n10823 );
xor ( n11058 , n10833 , n10837 );
xor ( n11059 , n11058 , n10846 );
and ( n11060 , n11057 , n11059 );
and ( n11061 , n10747 , n8253 );
and ( n11062 , n10499 , n8251 );
nor ( n11063 , n11061 , n11062 );
xnor ( n11064 , n11063 , n8259 );
xor ( n11065 , n6349 , n6538 );
buf ( n538326 , n11065 );
buf ( n538327 , n538326 );
buf ( n11068 , n538327 );
and ( n11069 , n11068 , n8106 );
and ( n11070 , n10842 , n8104 );
nor ( n11071 , n11069 , n11070 );
not ( n11072 , n11071 );
and ( n11073 , n11064 , n11072 );
xor ( n11074 , n10955 , n10959 );
and ( n11075 , n11072 , n11074 );
and ( n11076 , n11064 , n11074 );
or ( n11077 , n11073 , n11075 , n11076 );
and ( n11078 , n11059 , n11077 );
and ( n11079 , n11057 , n11077 );
or ( n11080 , n11060 , n11078 , n11079 );
and ( n11081 , n11055 , n11080 );
xor ( n11082 , n10965 , n10969 );
and ( n11083 , n9162 , n7144 );
and ( n11084 , n9084 , n7142 );
nor ( n11085 , n11083 , n11084 );
xnor ( n11086 , n11085 , n7154 );
and ( n11087 , n9482 , n6923 );
and ( n11088 , n9410 , n6921 );
nor ( n11089 , n11087 , n11088 );
xnor ( n11090 , n11089 , n6933 );
and ( n11091 , n11086 , n11090 );
and ( n11092 , n11082 , n11091 );
and ( n11093 , n7149 , n7683 );
and ( n11094 , n7879 , n7680 );
nor ( n11095 , n11093 , n11094 );
xnor ( n11096 , n11095 , n7676 );
and ( n11097 , n6928 , n7732 );
and ( n11098 , n7130 , n7730 );
nor ( n11099 , n11097 , n11098 );
xnor ( n11100 , n11099 , n7742 );
and ( n11101 , n11096 , n11100 );
and ( n11102 , n8039 , n7762 );
and ( n11103 , n6868 , n7760 );
nor ( n11104 , n11102 , n11103 );
xnor ( n11105 , n11104 , n7772 );
and ( n11106 , n11100 , n11105 );
and ( n11107 , n11096 , n11105 );
or ( n11108 , n11101 , n11106 , n11107 );
and ( n11109 , n11091 , n11108 );
and ( n11110 , n11082 , n11108 );
or ( n11111 , n11092 , n11109 , n11110 );
and ( n11112 , n7898 , n7797 );
and ( n11113 , n7929 , n7795 );
nor ( n11114 , n11112 , n11113 );
xnor ( n11115 , n11114 , n7807 );
and ( n11116 , n7939 , n7826 );
and ( n11117 , n7968 , n7824 );
nor ( n11118 , n11116 , n11117 );
xnor ( n11119 , n11118 , n7836 );
and ( n11120 , n11115 , n11119 );
and ( n11121 , n8111 , n6722 );
and ( n11122 , n8245 , n6720 );
nor ( n11123 , n11121 , n11122 );
xnor ( n11124 , n11123 , n6821 );
and ( n11125 , n11119 , n11124 );
and ( n11126 , n11115 , n11124 );
or ( n11127 , n11120 , n11125 , n11126 );
and ( n11128 , n8595 , n6852 );
and ( n11129 , n8091 , n6850 );
nor ( n11130 , n11128 , n11129 );
xnor ( n11131 , n11130 , n6862 );
and ( n11132 , n8604 , n7874 );
and ( n11133 , n8609 , n7872 );
nor ( n11134 , n11132 , n11133 );
xnor ( n11135 , n11134 , n7884 );
and ( n11136 , n11131 , n11135 );
and ( n11137 , n9925 , n7924 );
and ( n11138 , n9676 , n7922 );
nor ( n11139 , n11137 , n11138 );
xnor ( n11140 , n11139 , n7934 );
and ( n11141 , n11135 , n11140 );
and ( n11142 , n11131 , n11140 );
or ( n11143 , n11136 , n11141 , n11142 );
and ( n11144 , n11127 , n11143 );
and ( n11145 , n10120 , n7963 );
and ( n11146 , n10055 , n7961 );
nor ( n11147 , n11145 , n11146 );
xnor ( n11148 , n11147 , n7973 );
and ( n11149 , n10499 , n7995 );
and ( n11150 , n10419 , n7993 );
nor ( n11151 , n11149 , n11150 );
xnor ( n11152 , n11151 , n8005 );
and ( n11153 , n11148 , n11152 );
and ( n11154 , n10842 , n8253 );
and ( n11155 , n10747 , n8251 );
nor ( n11156 , n11154 , n11155 );
xnor ( n11157 , n11156 , n8259 );
and ( n11158 , n11152 , n11157 );
and ( n11159 , n11148 , n11157 );
or ( n11160 , n11153 , n11158 , n11159 );
and ( n11161 , n11143 , n11160 );
and ( n11162 , n11127 , n11160 );
or ( n11163 , n11144 , n11161 , n11162 );
and ( n11164 , n11111 , n11163 );
xor ( n11165 , n10929 , n10930 );
xor ( n11166 , n11165 , n10932 );
and ( n11167 , n11163 , n11166 );
and ( n11168 , n11111 , n11166 );
or ( n11169 , n11164 , n11167 , n11168 );
and ( n11170 , n11080 , n11169 );
and ( n11171 , n11055 , n11169 );
or ( n11172 , n11081 , n11170 , n11171 );
and ( n11173 , n11036 , n11172 );
xor ( n11174 , n10906 , n10908 );
xor ( n11175 , n11174 , n10910 );
xor ( n11176 , n10935 , n10973 );
xor ( n11177 , n11176 , n11012 );
and ( n11178 , n11175 , n11177 );
xor ( n11179 , n11017 , n11019 );
xor ( n11180 , n11179 , n11022 );
and ( n11181 , n11177 , n11180 );
and ( n11182 , n11175 , n11180 );
or ( n11183 , n11178 , n11181 , n11182 );
and ( n11184 , n11172 , n11183 );
and ( n11185 , n11036 , n11183 );
or ( n11186 , n11173 , n11184 , n11185 );
and ( n11187 , n11033 , n11186 );
and ( n11188 , n11031 , n11186 );
or ( n11189 , n11034 , n11187 , n11188 );
and ( n11190 , n10927 , n11189 );
xor ( n11191 , n10891 , n10893 );
xor ( n11192 , n11191 , n10919 );
and ( n11193 , n11189 , n11192 );
and ( n11194 , n10927 , n11192 );
or ( n11195 , n11190 , n11193 , n11194 );
and ( n11196 , n10924 , n11195 );
and ( n11197 , n10922 , n11195 );
or ( n11198 , n10925 , n11196 , n11197 );
and ( n11199 , n10889 , n11198 );
xor ( n11200 , n10889 , n11198 );
xor ( n11201 , n10922 , n10924 );
xor ( n11202 , n11201 , n11195 );
xor ( n11203 , n10896 , n10898 );
xor ( n11204 , n11203 , n10916 );
xor ( n11205 , n10901 , n10903 );
xor ( n11206 , n11205 , n10913 );
xor ( n11207 , n11015 , n11025 );
xor ( n11208 , n11207 , n11028 );
and ( n11209 , n11206 , n11208 );
xor ( n11210 , n10951 , n10960 );
xor ( n11211 , n11210 , n10970 );
xor ( n11212 , n10990 , n11006 );
xor ( n11213 , n11212 , n11009 );
and ( n11214 , n11211 , n11213 );
xor ( n11215 , n11050 , n11054 );
and ( n11216 , n11213 , n11215 );
and ( n11217 , n11211 , n11215 );
or ( n11218 , n11214 , n11216 , n11217 );
xor ( n11219 , n10978 , n10982 );
xor ( n11220 , n11219 , n10987 );
xor ( n11221 , n10994 , n10998 );
xor ( n11222 , n11221 , n11003 );
and ( n11223 , n11220 , n11222 );
xor ( n11224 , n11040 , n11044 );
xor ( n11225 , n11224 , n11047 );
and ( n11226 , n11222 , n11225 );
and ( n11227 , n11220 , n11225 );
or ( n11228 , n11223 , n11226 , n11227 );
and ( n11229 , n8609 , n6852 );
and ( n11230 , n8595 , n6850 );
nor ( n11231 , n11229 , n11230 );
xnor ( n11232 , n11231 , n6862 );
and ( n11233 , n9084 , n7874 );
and ( n11234 , n8604 , n7872 );
nor ( n11235 , n11233 , n11234 );
xnor ( n11236 , n11235 , n7884 );
and ( n11237 , n11232 , n11236 );
and ( n11238 , n9410 , n7144 );
and ( n11239 , n9162 , n7142 );
nor ( n11240 , n11238 , n11239 );
xnor ( n11241 , n11240 , n7154 );
and ( n11242 , n11236 , n11241 );
and ( n11243 , n11232 , n11241 );
or ( n11244 , n11237 , n11242 , n11243 );
and ( n11245 , n7979 , n7847 );
and ( n11246 , n8000 , n7845 );
nor ( n11247 , n11245 , n11246 );
xnor ( n11248 , n11247 , n7857 );
and ( n11249 , n11244 , n11248 );
and ( n11250 , n8071 , n7036 );
and ( n11251 , n8076 , n7034 );
nor ( n11252 , n11250 , n11251 );
xnor ( n11253 , n11252 , n7125 );
and ( n11254 , n11248 , n11253 );
and ( n11255 , n11244 , n11253 );
or ( n11256 , n11249 , n11254 , n11255 );
xor ( n11257 , n6381 , n6536 );
buf ( n538518 , n11257 );
buf ( n538519 , n538518 );
buf ( n11260 , n538519 );
and ( n11261 , n11260 , n8106 );
and ( n11262 , n11068 , n8104 );
nor ( n11263 , n11261 , n11262 );
not ( n11264 , n11263 );
xor ( n11265 , n11086 , n11090 );
and ( n11266 , n11264 , n11265 );
and ( n11267 , n10055 , n7924 );
and ( n11268 , n9925 , n7922 );
nor ( n11269 , n11267 , n11268 );
xnor ( n11270 , n11269 , n7934 );
and ( n11271 , n10419 , n7963 );
and ( n11272 , n10120 , n7961 );
nor ( n11273 , n11271 , n11272 );
xnor ( n11274 , n11273 , n7973 );
and ( n11275 , n11270 , n11274 );
and ( n11276 , n11265 , n11275 );
and ( n11277 , n11264 , n11275 );
or ( n11278 , n11266 , n11276 , n11277 );
and ( n11279 , n11256 , n11278 );
and ( n11280 , n7130 , n7683 );
and ( n11281 , n7149 , n7680 );
nor ( n11282 , n11280 , n11281 );
xnor ( n11283 , n11282 , n7676 );
and ( n11284 , n6868 , n7732 );
and ( n11285 , n6928 , n7730 );
nor ( n11286 , n11284 , n11285 );
xnor ( n11287 , n11286 , n7742 );
and ( n11288 , n11283 , n11287 );
and ( n11289 , n7929 , n7762 );
and ( n11290 , n8039 , n7760 );
nor ( n11291 , n11289 , n11290 );
xnor ( n11292 , n11291 , n7772 );
and ( n11293 , n11287 , n11292 );
and ( n11294 , n11283 , n11292 );
or ( n11295 , n11288 , n11293 , n11294 );
and ( n11296 , n7968 , n7797 );
and ( n11297 , n7898 , n7795 );
nor ( n11298 , n11296 , n11297 );
xnor ( n11299 , n11298 , n7807 );
and ( n11300 , n8245 , n7036 );
and ( n11301 , n8071 , n7034 );
nor ( n11302 , n11300 , n11301 );
xnor ( n11303 , n11302 , n7125 );
and ( n11304 , n11299 , n11303 );
and ( n11305 , n8091 , n6722 );
and ( n11306 , n8111 , n6720 );
nor ( n11307 , n11305 , n11306 );
xnor ( n11308 , n11307 , n6821 );
and ( n11309 , n11303 , n11308 );
and ( n11310 , n11299 , n11308 );
or ( n11311 , n11304 , n11309 , n11310 );
and ( n11312 , n11295 , n11311 );
and ( n11313 , n9676 , n6923 );
and ( n11314 , n9482 , n6921 );
nor ( n11315 , n11313 , n11314 );
xnor ( n11316 , n11315 , n6933 );
and ( n11317 , n10747 , n7995 );
and ( n11318 , n10499 , n7993 );
nor ( n11319 , n11317 , n11318 );
xnor ( n11320 , n11319 , n8005 );
and ( n11321 , n11316 , n11320 );
and ( n11322 , n11068 , n8253 );
and ( n11323 , n10842 , n8251 );
nor ( n11324 , n11322 , n11323 );
xnor ( n11325 , n11324 , n8259 );
and ( n11326 , n11320 , n11325 );
and ( n11327 , n11316 , n11325 );
or ( n11328 , n11321 , n11326 , n11327 );
and ( n11329 , n11311 , n11328 );
and ( n11330 , n11295 , n11328 );
or ( n11331 , n11312 , n11329 , n11330 );
and ( n11332 , n11278 , n11331 );
and ( n11333 , n11256 , n11331 );
or ( n11334 , n11279 , n11332 , n11333 );
and ( n11335 , n11228 , n11334 );
xor ( n11336 , n11096 , n11100 );
xor ( n11337 , n11336 , n11105 );
xor ( n11338 , n11115 , n11119 );
xor ( n11339 , n11338 , n11124 );
and ( n11340 , n11337 , n11339 );
xor ( n11341 , n11131 , n11135 );
xor ( n11342 , n11341 , n11140 );
and ( n11343 , n11339 , n11342 );
and ( n11344 , n11337 , n11342 );
or ( n11345 , n11340 , n11343 , n11344 );
xor ( n11346 , n11064 , n11072 );
xor ( n11347 , n11346 , n11074 );
and ( n11348 , n11345 , n11347 );
xor ( n11349 , n11082 , n11091 );
xor ( n11350 , n11349 , n11108 );
and ( n11351 , n11347 , n11350 );
and ( n11352 , n11345 , n11350 );
or ( n11353 , n11348 , n11351 , n11352 );
and ( n11354 , n11334 , n11353 );
and ( n11355 , n11228 , n11353 );
or ( n11356 , n11335 , n11354 , n11355 );
and ( n11357 , n11218 , n11356 );
xor ( n11358 , n11055 , n11080 );
xor ( n11359 , n11358 , n11169 );
and ( n11360 , n11356 , n11359 );
and ( n11361 , n11218 , n11359 );
or ( n11362 , n11357 , n11360 , n11361 );
and ( n11363 , n11208 , n11362 );
and ( n11364 , n11206 , n11362 );
or ( n11365 , n11209 , n11363 , n11364 );
and ( n11366 , n11204 , n11365 );
xor ( n11367 , n11031 , n11033 );
xor ( n11368 , n11367 , n11186 );
and ( n11369 , n11365 , n11368 );
and ( n11370 , n11204 , n11368 );
or ( n11371 , n11366 , n11369 , n11370 );
xor ( n11372 , n10927 , n11189 );
xor ( n11373 , n11372 , n11192 );
and ( n11374 , n11371 , n11373 );
xor ( n11375 , n11371 , n11373 );
xor ( n11376 , n11036 , n11172 );
xor ( n11377 , n11376 , n11183 );
xor ( n11378 , n11175 , n11177 );
xor ( n11379 , n11378 , n11180 );
xor ( n11380 , n11057 , n11059 );
xor ( n11381 , n11380 , n11077 );
xor ( n11382 , n11111 , n11163 );
xor ( n11383 , n11382 , n11166 );
and ( n11384 , n11381 , n11383 );
xor ( n11385 , n11127 , n11143 );
xor ( n11386 , n11385 , n11160 );
xor ( n11387 , n11148 , n11152 );
xor ( n11388 , n11387 , n11157 );
xor ( n11389 , n11244 , n11248 );
xor ( n11390 , n11389 , n11253 );
and ( n11391 , n11388 , n11390 );
and ( n11392 , n8000 , n7826 );
and ( n11393 , n7939 , n7824 );
nor ( n11394 , n11392 , n11393 );
xnor ( n11395 , n11394 , n7836 );
and ( n11396 , n8076 , n7847 );
and ( n11397 , n7979 , n7845 );
nor ( n11398 , n11396 , n11397 );
xnor ( n11399 , n11398 , n7857 );
and ( n11400 , n11395 , n11399 );
xor ( n11401 , n11232 , n11236 );
xor ( n11402 , n11401 , n11241 );
and ( n11403 , n11399 , n11402 );
and ( n11404 , n11395 , n11402 );
or ( n11405 , n11400 , n11403 , n11404 );
and ( n11406 , n11390 , n11405 );
and ( n11407 , n11388 , n11405 );
or ( n11408 , n11391 , n11406 , n11407 );
and ( n11409 , n11386 , n11408 );
xor ( n11410 , n6409 , n6534 );
buf ( n538671 , n11410 );
buf ( n538672 , n538671 );
buf ( n11413 , n538672 );
and ( n11414 , n11413 , n8106 );
and ( n11415 , n11260 , n8104 );
nor ( n11416 , n11414 , n11415 );
not ( n11417 , n11416 );
xor ( n11418 , n11270 , n11274 );
and ( n11419 , n11417 , n11418 );
and ( n11420 , n8604 , n6852 );
and ( n11421 , n8609 , n6850 );
nor ( n11422 , n11420 , n11421 );
xnor ( n11423 , n11422 , n6862 );
and ( n11424 , n9162 , n7874 );
and ( n11425 , n9084 , n7872 );
nor ( n11426 , n11424 , n11425 );
xnor ( n11427 , n11426 , n7884 );
and ( n11428 , n11423 , n11427 );
and ( n11429 , n9482 , n7144 );
and ( n11430 , n9410 , n7142 );
nor ( n11431 , n11429 , n11430 );
xnor ( n11432 , n11431 , n7154 );
and ( n11433 , n11427 , n11432 );
and ( n11434 , n11423 , n11432 );
or ( n11435 , n11428 , n11433 , n11434 );
and ( n11436 , n11418 , n11435 );
and ( n11437 , n11417 , n11435 );
or ( n11438 , n11419 , n11436 , n11437 );
and ( n11439 , n6928 , n7683 );
and ( n11440 , n7130 , n7680 );
nor ( n11441 , n11439 , n11440 );
xnor ( n11442 , n11441 , n7676 );
and ( n11443 , n8039 , n7732 );
and ( n11444 , n6868 , n7730 );
nor ( n11445 , n11443 , n11444 );
xnor ( n11446 , n11445 , n7742 );
and ( n11447 , n11442 , n11446 );
and ( n11448 , n7898 , n7762 );
and ( n11449 , n7929 , n7760 );
nor ( n11450 , n11448 , n11449 );
xnor ( n11451 , n11450 , n7772 );
and ( n11452 , n11446 , n11451 );
and ( n11453 , n11442 , n11451 );
or ( n11454 , n11447 , n11452 , n11453 );
and ( n11455 , n7939 , n7797 );
and ( n11456 , n7968 , n7795 );
nor ( n11457 , n11455 , n11456 );
xnor ( n11458 , n11457 , n7807 );
and ( n11459 , n7979 , n7826 );
and ( n11460 , n8000 , n7824 );
nor ( n11461 , n11459 , n11460 );
xnor ( n11462 , n11461 , n7836 );
and ( n11463 , n11458 , n11462 );
and ( n11464 , n8071 , n7847 );
and ( n11465 , n8076 , n7845 );
nor ( n11466 , n11464 , n11465 );
xnor ( n11467 , n11466 , n7857 );
and ( n11468 , n11462 , n11467 );
and ( n11469 , n11458 , n11467 );
or ( n11470 , n11463 , n11468 , n11469 );
and ( n11471 , n11454 , n11470 );
and ( n11472 , n8111 , n7036 );
and ( n11473 , n8245 , n7034 );
nor ( n11474 , n11472 , n11473 );
xnor ( n11475 , n11474 , n7125 );
and ( n11476 , n8595 , n6722 );
and ( n11477 , n8091 , n6720 );
nor ( n11478 , n11476 , n11477 );
xnor ( n11479 , n11478 , n6821 );
and ( n11480 , n11475 , n11479 );
and ( n11481 , n9925 , n6923 );
and ( n11482 , n9676 , n6921 );
nor ( n11483 , n11481 , n11482 );
xnor ( n11484 , n11483 , n6933 );
and ( n11485 , n11479 , n11484 );
and ( n11486 , n11475 , n11484 );
or ( n11487 , n11480 , n11485 , n11486 );
and ( n11488 , n11470 , n11487 );
and ( n11489 , n11454 , n11487 );
or ( n11490 , n11471 , n11488 , n11489 );
and ( n11491 , n11438 , n11490 );
and ( n11492 , n10120 , n7924 );
and ( n11493 , n10055 , n7922 );
nor ( n11494 , n11492 , n11493 );
xnor ( n11495 , n11494 , n7934 );
and ( n11496 , n10499 , n7963 );
and ( n11497 , n10419 , n7961 );
nor ( n11498 , n11496 , n11497 );
xnor ( n11499 , n11498 , n7973 );
and ( n11500 , n11495 , n11499 );
and ( n11501 , n10842 , n7995 );
and ( n11502 , n10747 , n7993 );
nor ( n11503 , n11501 , n11502 );
xnor ( n11504 , n11503 , n8005 );
and ( n11505 , n11499 , n11504 );
and ( n11506 , n11495 , n11504 );
or ( n11507 , n11500 , n11505 , n11506 );
xor ( n11508 , n11283 , n11287 );
xor ( n11509 , n11508 , n11292 );
and ( n11510 , n11507 , n11509 );
xor ( n11511 , n11299 , n11303 );
xor ( n11512 , n11511 , n11308 );
and ( n11513 , n11509 , n11512 );
and ( n11514 , n11507 , n11512 );
or ( n11515 , n11510 , n11513 , n11514 );
and ( n11516 , n11490 , n11515 );
and ( n11517 , n11438 , n11515 );
or ( n11518 , n11491 , n11516 , n11517 );
and ( n11519 , n11408 , n11518 );
and ( n11520 , n11386 , n11518 );
or ( n11521 , n11409 , n11519 , n11520 );
and ( n11522 , n11383 , n11521 );
and ( n11523 , n11381 , n11521 );
or ( n11524 , n11384 , n11522 , n11523 );
and ( n11525 , n11379 , n11524 );
xor ( n11526 , n11264 , n11265 );
xor ( n11527 , n11526 , n11275 );
xor ( n11528 , n11295 , n11311 );
xor ( n11529 , n11528 , n11328 );
and ( n11530 , n11527 , n11529 );
xor ( n11531 , n11337 , n11339 );
xor ( n11532 , n11531 , n11342 );
and ( n11533 , n11529 , n11532 );
and ( n11534 , n11527 , n11532 );
or ( n11535 , n11530 , n11533 , n11534 );
xor ( n11536 , n11220 , n11222 );
xor ( n11537 , n11536 , n11225 );
and ( n11538 , n11535 , n11537 );
xor ( n11539 , n11256 , n11278 );
xor ( n11540 , n11539 , n11331 );
and ( n11541 , n11537 , n11540 );
and ( n11542 , n11535 , n11540 );
or ( n11543 , n11538 , n11541 , n11542 );
xor ( n11544 , n11211 , n11213 );
xor ( n11545 , n11544 , n11215 );
and ( n11546 , n11543 , n11545 );
xor ( n11547 , n11228 , n11334 );
xor ( n11548 , n11547 , n11353 );
and ( n11549 , n11545 , n11548 );
and ( n11550 , n11543 , n11548 );
or ( n11551 , n11546 , n11549 , n11550 );
and ( n11552 , n11524 , n11551 );
and ( n11553 , n11379 , n11551 );
or ( n11554 , n11525 , n11552 , n11553 );
and ( n11555 , n11377 , n11554 );
xor ( n11556 , n11206 , n11208 );
xor ( n11557 , n11556 , n11362 );
and ( n11558 , n11554 , n11557 );
and ( n11559 , n11377 , n11557 );
or ( n11560 , n11555 , n11558 , n11559 );
xor ( n11561 , n11204 , n11365 );
xor ( n11562 , n11561 , n11368 );
and ( n11563 , n11560 , n11562 );
xor ( n11564 , n11560 , n11562 );
xor ( n11565 , n11218 , n11356 );
xor ( n11566 , n11565 , n11359 );
xor ( n11567 , n11345 , n11347 );
xor ( n11568 , n11567 , n11350 );
xor ( n11569 , n11316 , n11320 );
xor ( n11570 , n11569 , n11325 );
xor ( n11571 , n11395 , n11399 );
xor ( n11572 , n11571 , n11402 );
and ( n11573 , n11570 , n11572 );
and ( n11574 , n11260 , n8253 );
and ( n11575 , n11068 , n8251 );
nor ( n11576 , n11574 , n11575 );
xnor ( n11577 , n11576 , n8259 );
xor ( n11578 , n6432 , n6532 );
buf ( n538839 , n11578 );
buf ( n538840 , n538839 );
buf ( n11581 , n538840 );
and ( n11582 , n11581 , n8106 );
and ( n11583 , n11413 , n8104 );
nor ( n11584 , n11582 , n11583 );
not ( n11585 , n11584 );
and ( n11586 , n11577 , n11585 );
xor ( n11587 , n11423 , n11427 );
xor ( n11588 , n11587 , n11432 );
and ( n11589 , n11585 , n11588 );
and ( n11590 , n11577 , n11588 );
or ( n11591 , n11586 , n11589 , n11590 );
and ( n11592 , n11572 , n11591 );
and ( n11593 , n11570 , n11591 );
or ( n11594 , n11573 , n11592 , n11593 );
and ( n11595 , n10055 , n6923 );
and ( n11596 , n9925 , n6921 );
nor ( n11597 , n11595 , n11596 );
xnor ( n11598 , n11597 , n6933 );
and ( n11599 , n10419 , n7924 );
and ( n11600 , n10120 , n7922 );
nor ( n11601 , n11599 , n11600 );
xnor ( n11602 , n11601 , n7934 );
and ( n11603 , n11598 , n11602 );
and ( n11604 , n9410 , n7874 );
and ( n11605 , n9162 , n7872 );
nor ( n11606 , n11604 , n11605 );
xnor ( n11607 , n11606 , n7884 );
and ( n11608 , n9676 , n7144 );
and ( n11609 , n9482 , n7142 );
nor ( n11610 , n11608 , n11609 );
xnor ( n11611 , n11610 , n7154 );
and ( n11612 , n11607 , n11611 );
and ( n11613 , n11603 , n11612 );
and ( n11614 , n6868 , n7683 );
and ( n11615 , n6928 , n7680 );
nor ( n11616 , n11614 , n11615 );
xnor ( n11617 , n11616 , n7676 );
and ( n11618 , n7929 , n7732 );
and ( n11619 , n8039 , n7730 );
nor ( n11620 , n11618 , n11619 );
xnor ( n11621 , n11620 , n7742 );
and ( n11622 , n11617 , n11621 );
and ( n11623 , n7968 , n7762 );
and ( n11624 , n7898 , n7760 );
nor ( n11625 , n11623 , n11624 );
xnor ( n11626 , n11625 , n7772 );
and ( n11627 , n11621 , n11626 );
and ( n11628 , n11617 , n11626 );
or ( n11629 , n11622 , n11627 , n11628 );
and ( n11630 , n11612 , n11629 );
and ( n11631 , n11603 , n11629 );
or ( n11632 , n11613 , n11630 , n11631 );
and ( n11633 , n8000 , n7797 );
and ( n11634 , n7939 , n7795 );
nor ( n11635 , n11633 , n11634 );
xnor ( n11636 , n11635 , n7807 );
and ( n11637 , n8076 , n7826 );
and ( n11638 , n7979 , n7824 );
nor ( n11639 , n11637 , n11638 );
xnor ( n11640 , n11639 , n7836 );
and ( n11641 , n11636 , n11640 );
and ( n11642 , n8245 , n7847 );
and ( n11643 , n8071 , n7845 );
nor ( n11644 , n11642 , n11643 );
xnor ( n11645 , n11644 , n7857 );
and ( n11646 , n11640 , n11645 );
and ( n11647 , n11636 , n11645 );
or ( n11648 , n11641 , n11646 , n11647 );
and ( n11649 , n8091 , n7036 );
and ( n11650 , n8111 , n7034 );
nor ( n11651 , n11649 , n11650 );
xnor ( n11652 , n11651 , n7125 );
and ( n11653 , n8609 , n6722 );
and ( n11654 , n8595 , n6720 );
nor ( n11655 , n11653 , n11654 );
xnor ( n11656 , n11655 , n6821 );
and ( n11657 , n11652 , n11656 );
and ( n11658 , n9084 , n6852 );
and ( n11659 , n8604 , n6850 );
nor ( n11660 , n11658 , n11659 );
xnor ( n11661 , n11660 , n6862 );
and ( n11662 , n11656 , n11661 );
and ( n11663 , n11652 , n11661 );
or ( n11664 , n11657 , n11662 , n11663 );
and ( n11665 , n11648 , n11664 );
and ( n11666 , n10747 , n7963 );
and ( n11667 , n10499 , n7961 );
nor ( n11668 , n11666 , n11667 );
xnor ( n11669 , n11668 , n7973 );
and ( n11670 , n11068 , n7995 );
and ( n11671 , n10842 , n7993 );
nor ( n11672 , n11670 , n11671 );
xnor ( n11673 , n11672 , n8005 );
and ( n11674 , n11669 , n11673 );
and ( n11675 , n11413 , n8253 );
and ( n11676 , n11260 , n8251 );
nor ( n11677 , n11675 , n11676 );
xnor ( n11678 , n11677 , n8259 );
and ( n11679 , n11673 , n11678 );
and ( n11680 , n11669 , n11678 );
or ( n11681 , n11674 , n11679 , n11680 );
and ( n11682 , n11664 , n11681 );
and ( n11683 , n11648 , n11681 );
or ( n11684 , n11665 , n11682 , n11683 );
and ( n11685 , n11632 , n11684 );
xor ( n11686 , n11442 , n11446 );
xor ( n11687 , n11686 , n11451 );
xor ( n11688 , n11458 , n11462 );
xor ( n11689 , n11688 , n11467 );
and ( n11690 , n11687 , n11689 );
xor ( n11691 , n11475 , n11479 );
xor ( n11692 , n11691 , n11484 );
and ( n11693 , n11689 , n11692 );
and ( n11694 , n11687 , n11692 );
or ( n11695 , n11690 , n11693 , n11694 );
and ( n11696 , n11684 , n11695 );
and ( n11697 , n11632 , n11695 );
or ( n11698 , n11685 , n11696 , n11697 );
and ( n11699 , n11594 , n11698 );
xor ( n11700 , n11417 , n11418 );
xor ( n11701 , n11700 , n11435 );
xor ( n11702 , n11454 , n11470 );
xor ( n11703 , n11702 , n11487 );
and ( n11704 , n11701 , n11703 );
xor ( n11705 , n11507 , n11509 );
xor ( n11706 , n11705 , n11512 );
and ( n11707 , n11703 , n11706 );
and ( n11708 , n11701 , n11706 );
or ( n11709 , n11704 , n11707 , n11708 );
and ( n11710 , n11698 , n11709 );
and ( n11711 , n11594 , n11709 );
or ( n11712 , n11699 , n11710 , n11711 );
and ( n11713 , n11568 , n11712 );
xor ( n11714 , n11388 , n11390 );
xor ( n11715 , n11714 , n11405 );
xor ( n11716 , n11438 , n11490 );
xor ( n11717 , n11716 , n11515 );
and ( n11718 , n11715 , n11717 );
xor ( n11719 , n11527 , n11529 );
xor ( n11720 , n11719 , n11532 );
and ( n11721 , n11717 , n11720 );
and ( n11722 , n11715 , n11720 );
or ( n11723 , n11718 , n11721 , n11722 );
and ( n11724 , n11712 , n11723 );
and ( n11725 , n11568 , n11723 );
or ( n11726 , n11713 , n11724 , n11725 );
xor ( n11727 , n11381 , n11383 );
xor ( n11728 , n11727 , n11521 );
and ( n11729 , n11726 , n11728 );
xor ( n11730 , n11543 , n11545 );
xor ( n11731 , n11730 , n11548 );
and ( n11732 , n11728 , n11731 );
and ( n11733 , n11726 , n11731 );
or ( n11734 , n11729 , n11732 , n11733 );
and ( n11735 , n11566 , n11734 );
xor ( n11736 , n11379 , n11524 );
xor ( n11737 , n11736 , n11551 );
and ( n11738 , n11734 , n11737 );
and ( n11739 , n11566 , n11737 );
or ( n11740 , n11735 , n11738 , n11739 );
xor ( n11741 , n11377 , n11554 );
xor ( n11742 , n11741 , n11557 );
and ( n11743 , n11740 , n11742 );
xor ( n11744 , n11740 , n11742 );
xor ( n11745 , n11566 , n11734 );
xor ( n11746 , n11745 , n11737 );
xor ( n11747 , n11386 , n11408 );
xor ( n11748 , n11747 , n11518 );
xor ( n11749 , n11535 , n11537 );
xor ( n11750 , n11749 , n11540 );
and ( n11751 , n11748 , n11750 );
xor ( n11752 , n11495 , n11499 );
xor ( n11753 , n11752 , n11504 );
xor ( n11754 , n6454 , n6530 );
buf ( n539015 , n11754 );
buf ( n539016 , n539015 );
buf ( n11757 , n539016 );
and ( n11758 , n11757 , n8106 );
and ( n11759 , n11581 , n8104 );
nor ( n11760 , n11758 , n11759 );
not ( n11761 , n11760 );
xor ( n11762 , n11598 , n11602 );
and ( n11763 , n11761 , n11762 );
xor ( n11764 , n11607 , n11611 );
and ( n11765 , n11762 , n11764 );
and ( n11766 , n11761 , n11764 );
or ( n11767 , n11763 , n11765 , n11766 );
and ( n11768 , n11753 , n11767 );
and ( n11769 , n7939 , n7762 );
and ( n11770 , n7968 , n7760 );
nor ( n11771 , n11769 , n11770 );
xnor ( n11772 , n11771 , n7772 );
and ( n11773 , n7979 , n7797 );
and ( n11774 , n8000 , n7795 );
nor ( n11775 , n11773 , n11774 );
xnor ( n11776 , n11775 , n7807 );
and ( n11777 , n11772 , n11776 );
and ( n11778 , n8039 , n7683 );
and ( n11779 , n6868 , n7680 );
nor ( n11780 , n11778 , n11779 );
xnor ( n11781 , n11780 , n7676 );
and ( n11782 , n7898 , n7732 );
and ( n11783 , n7929 , n7730 );
nor ( n11784 , n11782 , n11783 );
xnor ( n11785 , n11784 , n7742 );
and ( n11786 , n11781 , n11785 );
and ( n11787 , n8071 , n7826 );
and ( n11788 , n8076 , n7824 );
nor ( n11789 , n11787 , n11788 );
xnor ( n11790 , n11789 , n7836 );
and ( n11791 , n11785 , n11790 );
and ( n11792 , n11781 , n11790 );
or ( n11793 , n11786 , n11791 , n11792 );
and ( n11794 , n11777 , n11793 );
and ( n11795 , n8111 , n7847 );
and ( n11796 , n8245 , n7845 );
nor ( n11797 , n11795 , n11796 );
xnor ( n11798 , n11797 , n7857 );
and ( n11799 , n8595 , n7036 );
and ( n11800 , n8091 , n7034 );
nor ( n11801 , n11799 , n11800 );
xnor ( n11802 , n11801 , n7125 );
and ( n11803 , n11798 , n11802 );
and ( n11804 , n8604 , n6722 );
and ( n11805 , n8609 , n6720 );
nor ( n11806 , n11804 , n11805 );
xnor ( n11807 , n11806 , n6821 );
and ( n11808 , n11802 , n11807 );
and ( n11809 , n11798 , n11807 );
or ( n11810 , n11803 , n11808 , n11809 );
and ( n11811 , n11793 , n11810 );
and ( n11812 , n11777 , n11810 );
or ( n11813 , n11794 , n11811 , n11812 );
and ( n11814 , n11767 , n11813 );
and ( n11815 , n11753 , n11813 );
or ( n11816 , n11768 , n11814 , n11815 );
and ( n11817 , n9162 , n6852 );
and ( n11818 , n9084 , n6850 );
nor ( n11819 , n11817 , n11818 );
xnor ( n11820 , n11819 , n6862 );
and ( n11821 , n9482 , n7874 );
and ( n11822 , n9410 , n7872 );
nor ( n11823 , n11821 , n11822 );
xnor ( n11824 , n11823 , n7884 );
and ( n11825 , n11820 , n11824 );
and ( n11826 , n9925 , n7144 );
and ( n11827 , n9676 , n7142 );
nor ( n11828 , n11826 , n11827 );
xnor ( n11829 , n11828 , n7154 );
and ( n11830 , n11824 , n11829 );
and ( n11831 , n11820 , n11829 );
or ( n11832 , n11825 , n11830 , n11831 );
and ( n11833 , n10120 , n6923 );
and ( n11834 , n10055 , n6921 );
nor ( n11835 , n11833 , n11834 );
xnor ( n11836 , n11835 , n6933 );
and ( n11837 , n10499 , n7924 );
and ( n11838 , n10419 , n7922 );
nor ( n11839 , n11837 , n11838 );
xnor ( n11840 , n11839 , n7934 );
and ( n11841 , n11836 , n11840 );
and ( n11842 , n10842 , n7963 );
and ( n11843 , n10747 , n7961 );
nor ( n11844 , n11842 , n11843 );
xnor ( n11845 , n11844 , n7973 );
and ( n11846 , n11840 , n11845 );
and ( n11847 , n11836 , n11845 );
or ( n11848 , n11841 , n11846 , n11847 );
and ( n11849 , n11832 , n11848 );
and ( n11850 , n11260 , n7995 );
and ( n11851 , n11068 , n7993 );
nor ( n11852 , n11850 , n11851 );
xnor ( n11853 , n11852 , n8005 );
and ( n11854 , n11581 , n8253 );
and ( n11855 , n11413 , n8251 );
nor ( n11856 , n11854 , n11855 );
xnor ( n11857 , n11856 , n8259 );
and ( n11858 , n11853 , n11857 );
xor ( n11859 , n6471 , n6528 );
buf ( n539120 , n11859 );
buf ( n539121 , n539120 );
buf ( n11862 , n539121 );
and ( n11863 , n11862 , n8106 );
and ( n11864 , n11757 , n8104 );
nor ( n11865 , n11863 , n11864 );
not ( n11866 , n11865 );
and ( n11867 , n11857 , n11866 );
and ( n11868 , n11853 , n11866 );
or ( n11869 , n11858 , n11867 , n11868 );
and ( n11870 , n11848 , n11869 );
and ( n11871 , n11832 , n11869 );
or ( n11872 , n11849 , n11870 , n11871 );
xor ( n11873 , n11617 , n11621 );
xor ( n11874 , n11873 , n11626 );
xor ( n11875 , n11636 , n11640 );
xor ( n11876 , n11875 , n11645 );
and ( n11877 , n11874 , n11876 );
xor ( n11878 , n11652 , n11656 );
xor ( n11879 , n11878 , n11661 );
and ( n11880 , n11876 , n11879 );
and ( n11881 , n11874 , n11879 );
or ( n11882 , n11877 , n11880 , n11881 );
and ( n11883 , n11872 , n11882 );
xor ( n11884 , n11577 , n11585 );
xor ( n11885 , n11884 , n11588 );
and ( n11886 , n11882 , n11885 );
and ( n11887 , n11872 , n11885 );
or ( n11888 , n11883 , n11886 , n11887 );
and ( n11889 , n11816 , n11888 );
xor ( n11890 , n11603 , n11612 );
xor ( n11891 , n11890 , n11629 );
xor ( n11892 , n11648 , n11664 );
xor ( n11893 , n11892 , n11681 );
and ( n11894 , n11891 , n11893 );
xor ( n11895 , n11687 , n11689 );
xor ( n11896 , n11895 , n11692 );
and ( n11897 , n11893 , n11896 );
and ( n11898 , n11891 , n11896 );
or ( n11899 , n11894 , n11897 , n11898 );
and ( n11900 , n11888 , n11899 );
and ( n11901 , n11816 , n11899 );
or ( n11902 , n11889 , n11900 , n11901 );
xor ( n11903 , n11570 , n11572 );
xor ( n11904 , n11903 , n11591 );
xor ( n11905 , n11632 , n11684 );
xor ( n11906 , n11905 , n11695 );
and ( n11907 , n11904 , n11906 );
xor ( n11908 , n11701 , n11703 );
xor ( n11909 , n11908 , n11706 );
and ( n11910 , n11906 , n11909 );
and ( n11911 , n11904 , n11909 );
or ( n11912 , n11907 , n11910 , n11911 );
and ( n11913 , n11902 , n11912 );
xor ( n11914 , n11594 , n11698 );
xor ( n11915 , n11914 , n11709 );
and ( n11916 , n11912 , n11915 );
and ( n11917 , n11902 , n11915 );
or ( n11918 , n11913 , n11916 , n11917 );
and ( n11919 , n11750 , n11918 );
and ( n11920 , n11748 , n11918 );
or ( n11921 , n11751 , n11919 , n11920 );
xor ( n11922 , n11726 , n11728 );
xor ( n11923 , n11922 , n11731 );
and ( n11924 , n11921 , n11923 );
xor ( n11925 , n11568 , n11712 );
xor ( n11926 , n11925 , n11723 );
xor ( n11927 , n11715 , n11717 );
xor ( n11928 , n11927 , n11720 );
xor ( n11929 , n11669 , n11673 );
xor ( n11930 , n11929 , n11678 );
xor ( n11931 , n11772 , n11776 );
and ( n11932 , n7929 , n7683 );
and ( n11933 , n8039 , n7680 );
nor ( n11934 , n11932 , n11933 );
xnor ( n11935 , n11934 , n7676 );
and ( n11936 , n7968 , n7732 );
and ( n11937 , n7898 , n7730 );
nor ( n11938 , n11936 , n11937 );
xnor ( n11939 , n11938 , n7742 );
and ( n11940 , n11935 , n11939 );
and ( n11941 , n8000 , n7762 );
and ( n11942 , n7939 , n7760 );
nor ( n11943 , n11941 , n11942 );
xnor ( n11944 , n11943 , n7772 );
and ( n11945 , n11939 , n11944 );
and ( n11946 , n11935 , n11944 );
or ( n11947 , n11940 , n11945 , n11946 );
and ( n11948 , n11931 , n11947 );
and ( n11949 , n8076 , n7797 );
and ( n11950 , n7979 , n7795 );
nor ( n11951 , n11949 , n11950 );
xnor ( n11952 , n11951 , n7807 );
and ( n11953 , n8245 , n7826 );
and ( n11954 , n8071 , n7824 );
nor ( n11955 , n11953 , n11954 );
xnor ( n11956 , n11955 , n7836 );
and ( n11957 , n11952 , n11956 );
and ( n11958 , n8091 , n7847 );
and ( n11959 , n8111 , n7845 );
nor ( n11960 , n11958 , n11959 );
xnor ( n11961 , n11960 , n7857 );
and ( n11962 , n11956 , n11961 );
and ( n11963 , n11952 , n11961 );
or ( n11964 , n11957 , n11962 , n11963 );
and ( n11965 , n11947 , n11964 );
and ( n11966 , n11931 , n11964 );
or ( n11967 , n11948 , n11965 , n11966 );
and ( n11968 , n11930 , n11967 );
and ( n11969 , n8609 , n7036 );
and ( n11970 , n8595 , n7034 );
nor ( n11971 , n11969 , n11970 );
xnor ( n11972 , n11971 , n7125 );
and ( n11973 , n9084 , n6722 );
and ( n11974 , n8604 , n6720 );
nor ( n11975 , n11973 , n11974 );
xnor ( n11976 , n11975 , n6821 );
and ( n11977 , n11972 , n11976 );
and ( n11978 , n9410 , n6852 );
and ( n11979 , n9162 , n6850 );
nor ( n11980 , n11978 , n11979 );
xnor ( n11981 , n11980 , n6862 );
and ( n11982 , n11976 , n11981 );
and ( n11983 , n11972 , n11981 );
or ( n11984 , n11977 , n11982 , n11983 );
and ( n11985 , n9676 , n7874 );
and ( n11986 , n9482 , n7872 );
nor ( n11987 , n11985 , n11986 );
xnor ( n11988 , n11987 , n7884 );
and ( n11989 , n10055 , n7144 );
and ( n11990 , n9925 , n7142 );
nor ( n11991 , n11989 , n11990 );
xnor ( n11992 , n11991 , n7154 );
and ( n11993 , n11988 , n11992 );
and ( n11994 , n10419 , n6923 );
and ( n11995 , n10120 , n6921 );
nor ( n11996 , n11994 , n11995 );
xnor ( n11997 , n11996 , n6933 );
and ( n11998 , n11992 , n11997 );
and ( n11999 , n11988 , n11997 );
or ( n12000 , n11993 , n11998 , n11999 );
and ( n12001 , n11984 , n12000 );
and ( n12002 , n10747 , n7924 );
and ( n12003 , n10499 , n7922 );
nor ( n12004 , n12002 , n12003 );
xnor ( n12005 , n12004 , n7934 );
and ( n12006 , n11068 , n7963 );
and ( n12007 , n10842 , n7961 );
nor ( n12008 , n12006 , n12007 );
xnor ( n12009 , n12008 , n7973 );
and ( n12010 , n12005 , n12009 );
and ( n12011 , n11413 , n7995 );
and ( n12012 , n11260 , n7993 );
nor ( n12013 , n12011 , n12012 );
xnor ( n12014 , n12013 , n8005 );
and ( n12015 , n12009 , n12014 );
and ( n12016 , n12005 , n12014 );
or ( n12017 , n12010 , n12015 , n12016 );
and ( n12018 , n12000 , n12017 );
and ( n12019 , n11984 , n12017 );
or ( n12020 , n12001 , n12018 , n12019 );
and ( n12021 , n11967 , n12020 );
and ( n12022 , n11930 , n12020 );
or ( n12023 , n11968 , n12021 , n12022 );
xor ( n12024 , n11781 , n11785 );
xor ( n12025 , n12024 , n11790 );
xor ( n12026 , n11798 , n11802 );
xor ( n12027 , n12026 , n11807 );
and ( n12028 , n12025 , n12027 );
xor ( n12029 , n11820 , n11824 );
xor ( n12030 , n12029 , n11829 );
and ( n12031 , n12027 , n12030 );
and ( n12032 , n12025 , n12030 );
or ( n12033 , n12028 , n12031 , n12032 );
xor ( n12034 , n11761 , n11762 );
xor ( n12035 , n12034 , n11764 );
and ( n12036 , n12033 , n12035 );
xor ( n12037 , n11777 , n11793 );
xor ( n12038 , n12037 , n11810 );
and ( n12039 , n12035 , n12038 );
and ( n12040 , n12033 , n12038 );
or ( n12041 , n12036 , n12039 , n12040 );
and ( n12042 , n12023 , n12041 );
xor ( n12043 , n11753 , n11767 );
xor ( n12044 , n12043 , n11813 );
and ( n12045 , n12041 , n12044 );
and ( n12046 , n12023 , n12044 );
or ( n12047 , n12042 , n12045 , n12046 );
xor ( n12048 , n11816 , n11888 );
xor ( n12049 , n12048 , n11899 );
and ( n12050 , n12047 , n12049 );
xor ( n12051 , n11904 , n11906 );
xor ( n12052 , n12051 , n11909 );
and ( n12053 , n12049 , n12052 );
and ( n12054 , n12047 , n12052 );
or ( n12055 , n12050 , n12053 , n12054 );
and ( n12056 , n11928 , n12055 );
xor ( n12057 , n11902 , n11912 );
xor ( n12058 , n12057 , n11915 );
and ( n12059 , n12055 , n12058 );
and ( n12060 , n11928 , n12058 );
or ( n12061 , n12056 , n12059 , n12060 );
and ( n12062 , n11926 , n12061 );
xor ( n12063 , n11748 , n11750 );
xor ( n12064 , n12063 , n11918 );
and ( n12065 , n12061 , n12064 );
and ( n12066 , n11926 , n12064 );
or ( n12067 , n12062 , n12065 , n12066 );
and ( n12068 , n11923 , n12067 );
and ( n12069 , n11921 , n12067 );
or ( n12070 , n11924 , n12068 , n12069 );
and ( n12071 , n11746 , n12070 );
xor ( n12072 , n11746 , n12070 );
xor ( n12073 , n11921 , n11923 );
xor ( n12074 , n12073 , n12067 );
xor ( n12075 , n11926 , n12061 );
xor ( n12076 , n12075 , n12064 );
xor ( n12077 , n11928 , n12055 );
xor ( n12078 , n12077 , n12058 );
xor ( n12079 , n11872 , n11882 );
xor ( n12080 , n12079 , n11885 );
xor ( n12081 , n11891 , n11893 );
xor ( n12082 , n12081 , n11896 );
and ( n12083 , n12080 , n12082 );
xor ( n12084 , n11832 , n11848 );
xor ( n12085 , n12084 , n11869 );
xor ( n12086 , n11874 , n11876 );
xor ( n12087 , n12086 , n11879 );
and ( n12088 , n12085 , n12087 );
xor ( n12089 , n11836 , n11840 );
xor ( n12090 , n12089 , n11845 );
xor ( n12091 , n11853 , n11857 );
xor ( n12092 , n12091 , n11866 );
and ( n12093 , n12090 , n12092 );
and ( n12094 , n11757 , n8253 );
and ( n12095 , n11581 , n8251 );
nor ( n12096 , n12094 , n12095 );
xnor ( n12097 , n12096 , n8259 );
xor ( n12098 , n6487 , n6526 );
buf ( n539359 , n12098 );
buf ( n539360 , n539359 );
buf ( n12101 , n539360 );
and ( n12102 , n12101 , n8106 );
and ( n12103 , n11862 , n8104 );
nor ( n12104 , n12102 , n12103 );
not ( n12105 , n12104 );
and ( n12106 , n12097 , n12105 );
and ( n12107 , n8111 , n7826 );
and ( n12108 , n8245 , n7824 );
nor ( n12109 , n12107 , n12108 );
xnor ( n12110 , n12109 , n7836 );
and ( n12111 , n8595 , n7847 );
and ( n12112 , n8091 , n7845 );
nor ( n12113 , n12111 , n12112 );
xnor ( n12114 , n12113 , n7857 );
and ( n12115 , n12110 , n12114 );
and ( n12116 , n12105 , n12115 );
and ( n12117 , n12097 , n12115 );
or ( n12118 , n12106 , n12116 , n12117 );
and ( n12119 , n12092 , n12118 );
and ( n12120 , n12090 , n12118 );
or ( n12121 , n12093 , n12119 , n12120 );
and ( n12122 , n12087 , n12121 );
and ( n12123 , n12085 , n12121 );
or ( n12124 , n12088 , n12122 , n12123 );
and ( n12125 , n12082 , n12124 );
and ( n12126 , n12080 , n12124 );
or ( n12127 , n12083 , n12125 , n12126 );
xor ( n12128 , n12047 , n12049 );
xor ( n12129 , n12128 , n12052 );
and ( n12130 , n12127 , n12129 );
and ( n12131 , n7939 , n7732 );
and ( n12132 , n7968 , n7730 );
nor ( n12133 , n12131 , n12132 );
xnor ( n12134 , n12133 , n7742 );
and ( n12135 , n8071 , n7797 );
and ( n12136 , n8076 , n7795 );
nor ( n12137 , n12135 , n12136 );
xnor ( n12138 , n12137 , n7807 );
and ( n12139 , n12134 , n12138 );
and ( n12140 , n7898 , n7683 );
and ( n12141 , n7929 , n7680 );
nor ( n12142 , n12140 , n12141 );
xnor ( n12143 , n12142 , n7676 );
and ( n12144 , n7979 , n7762 );
and ( n12145 , n8000 , n7760 );
nor ( n12146 , n12144 , n12145 );
xnor ( n12147 , n12146 , n7772 );
and ( n12148 , n12143 , n12147 );
and ( n12149 , n8604 , n7036 );
and ( n12150 , n8609 , n7034 );
nor ( n12151 , n12149 , n12150 );
xnor ( n12152 , n12151 , n7125 );
and ( n12153 , n12147 , n12152 );
and ( n12154 , n12143 , n12152 );
or ( n12155 , n12148 , n12153 , n12154 );
and ( n12156 , n12139 , n12155 );
and ( n12157 , n9162 , n6722 );
and ( n12158 , n9084 , n6720 );
nor ( n12159 , n12157 , n12158 );
xnor ( n12160 , n12159 , n6821 );
and ( n12161 , n9482 , n6852 );
and ( n12162 , n9410 , n6850 );
nor ( n12163 , n12161 , n12162 );
xnor ( n12164 , n12163 , n6862 );
and ( n12165 , n12160 , n12164 );
and ( n12166 , n9925 , n7874 );
and ( n12167 , n9676 , n7872 );
nor ( n12168 , n12166 , n12167 );
xnor ( n12169 , n12168 , n7884 );
and ( n12170 , n12164 , n12169 );
and ( n12171 , n12160 , n12169 );
or ( n12172 , n12165 , n12170 , n12171 );
and ( n12173 , n12155 , n12172 );
and ( n12174 , n12139 , n12172 );
or ( n12175 , n12156 , n12173 , n12174 );
and ( n12176 , n10120 , n7144 );
and ( n12177 , n10055 , n7142 );
nor ( n12178 , n12176 , n12177 );
xnor ( n12179 , n12178 , n7154 );
and ( n12180 , n10499 , n6923 );
and ( n12181 , n10419 , n6921 );
nor ( n12182 , n12180 , n12181 );
xnor ( n12183 , n12182 , n6933 );
and ( n12184 , n12179 , n12183 );
and ( n12185 , n10842 , n7924 );
and ( n12186 , n10747 , n7922 );
nor ( n12187 , n12185 , n12186 );
xnor ( n12188 , n12187 , n7934 );
and ( n12189 , n12183 , n12188 );
and ( n12190 , n12179 , n12188 );
or ( n12191 , n12184 , n12189 , n12190 );
and ( n12192 , n11260 , n7963 );
and ( n12193 , n11068 , n7961 );
nor ( n12194 , n12192 , n12193 );
xnor ( n12195 , n12194 , n7973 );
and ( n12196 , n11581 , n7995 );
and ( n12197 , n11413 , n7993 );
nor ( n12198 , n12196 , n12197 );
xnor ( n12199 , n12198 , n8005 );
and ( n12200 , n12195 , n12199 );
and ( n12201 , n11862 , n8253 );
and ( n12202 , n11757 , n8251 );
nor ( n12203 , n12201 , n12202 );
xnor ( n12204 , n12203 , n8259 );
and ( n12205 , n12199 , n12204 );
and ( n12206 , n12195 , n12204 );
or ( n12207 , n12200 , n12205 , n12206 );
and ( n12208 , n12191 , n12207 );
xor ( n12209 , n11935 , n11939 );
xor ( n12210 , n12209 , n11944 );
and ( n12211 , n12207 , n12210 );
and ( n12212 , n12191 , n12210 );
or ( n12213 , n12208 , n12211 , n12212 );
and ( n12214 , n12175 , n12213 );
xor ( n12215 , n11952 , n11956 );
xor ( n12216 , n12215 , n11961 );
xor ( n12217 , n11972 , n11976 );
xor ( n12218 , n12217 , n11981 );
and ( n12219 , n12216 , n12218 );
xor ( n12220 , n11988 , n11992 );
xor ( n12221 , n12220 , n11997 );
and ( n12222 , n12218 , n12221 );
and ( n12223 , n12216 , n12221 );
or ( n12224 , n12219 , n12222 , n12223 );
and ( n12225 , n12213 , n12224 );
and ( n12226 , n12175 , n12224 );
or ( n12227 , n12214 , n12225 , n12226 );
xor ( n12228 , n11931 , n11947 );
xor ( n12229 , n12228 , n11964 );
xor ( n12230 , n11984 , n12000 );
xor ( n12231 , n12230 , n12017 );
and ( n12232 , n12229 , n12231 );
xor ( n12233 , n12025 , n12027 );
xor ( n12234 , n12233 , n12030 );
and ( n12235 , n12231 , n12234 );
and ( n12236 , n12229 , n12234 );
or ( n12237 , n12232 , n12235 , n12236 );
and ( n12238 , n12227 , n12237 );
xor ( n12239 , n11930 , n11967 );
xor ( n12240 , n12239 , n12020 );
and ( n12241 , n12237 , n12240 );
and ( n12242 , n12227 , n12240 );
or ( n12243 , n12238 , n12241 , n12242 );
xor ( n12244 , n12023 , n12041 );
xor ( n12245 , n12244 , n12044 );
and ( n12246 , n12243 , n12245 );
xor ( n12247 , n12033 , n12035 );
xor ( n12248 , n12247 , n12038 );
xor ( n12249 , n12005 , n12009 );
xor ( n12250 , n12249 , n12014 );
xor ( n12251 , n6499 , n6524 );
buf ( n539512 , n12251 );
buf ( n539513 , n539512 );
buf ( n12254 , n539513 );
and ( n12255 , n12254 , n8106 );
and ( n12256 , n12101 , n8104 );
nor ( n12257 , n12255 , n12256 );
not ( n12258 , n12257 );
xor ( n12259 , n12110 , n12114 );
and ( n12260 , n12258 , n12259 );
xor ( n12261 , n12134 , n12138 );
and ( n12262 , n12259 , n12261 );
and ( n12263 , n12258 , n12261 );
or ( n12264 , n12260 , n12262 , n12263 );
and ( n12265 , n12250 , n12264 );
and ( n12266 , n10419 , n7144 );
and ( n12267 , n10120 , n7142 );
nor ( n12268 , n12266 , n12267 );
xnor ( n12269 , n12268 , n7154 );
and ( n12270 , n10747 , n6923 );
and ( n12271 , n10499 , n6921 );
nor ( n12272 , n12270 , n12271 );
xnor ( n12273 , n12272 , n6933 );
and ( n12274 , n12269 , n12273 );
and ( n12275 , n7968 , n7683 );
and ( n12276 , n7898 , n7680 );
nor ( n12277 , n12275 , n12276 );
xnor ( n12278 , n12277 , n7676 );
and ( n12279 , n8000 , n7732 );
and ( n12280 , n7939 , n7730 );
nor ( n12281 , n12279 , n12280 );
xnor ( n12282 , n12281 , n7742 );
and ( n12283 , n12278 , n12282 );
and ( n12284 , n8076 , n7762 );
and ( n12285 , n7979 , n7760 );
nor ( n12286 , n12284 , n12285 );
xnor ( n12287 , n12286 , n7772 );
and ( n12288 , n12282 , n12287 );
and ( n12289 , n12278 , n12287 );
or ( n12290 , n12283 , n12288 , n12289 );
and ( n12291 , n12274 , n12290 );
and ( n12292 , n8245 , n7797 );
and ( n12293 , n8071 , n7795 );
nor ( n12294 , n12292 , n12293 );
xnor ( n12295 , n12294 , n7807 );
and ( n12296 , n8091 , n7826 );
and ( n12297 , n8111 , n7824 );
nor ( n12298 , n12296 , n12297 );
xnor ( n12299 , n12298 , n7836 );
and ( n12300 , n12295 , n12299 );
and ( n12301 , n8609 , n7847 );
and ( n12302 , n8595 , n7845 );
nor ( n12303 , n12301 , n12302 );
xnor ( n12304 , n12303 , n7857 );
and ( n12305 , n12299 , n12304 );
and ( n12306 , n12295 , n12304 );
or ( n12307 , n12300 , n12305 , n12306 );
and ( n12308 , n12290 , n12307 );
and ( n12309 , n12274 , n12307 );
or ( n12310 , n12291 , n12308 , n12309 );
and ( n12311 , n12264 , n12310 );
and ( n12312 , n12250 , n12310 );
or ( n12313 , n12265 , n12311 , n12312 );
and ( n12314 , n9084 , n7036 );
and ( n12315 , n8604 , n7034 );
nor ( n12316 , n12314 , n12315 );
xnor ( n12317 , n12316 , n7125 );
and ( n12318 , n9410 , n6722 );
and ( n12319 , n9162 , n6720 );
nor ( n12320 , n12318 , n12319 );
xnor ( n12321 , n12320 , n6821 );
and ( n12322 , n12317 , n12321 );
and ( n12323 , n9676 , n6852 );
and ( n12324 , n9482 , n6850 );
nor ( n12325 , n12323 , n12324 );
xnor ( n12326 , n12325 , n6862 );
and ( n12327 , n12321 , n12326 );
and ( n12328 , n12317 , n12326 );
or ( n12329 , n12322 , n12327 , n12328 );
and ( n12330 , n10055 , n7874 );
and ( n12331 , n9925 , n7872 );
nor ( n12332 , n12330 , n12331 );
xnor ( n12333 , n12332 , n7884 );
and ( n12334 , n11068 , n7924 );
and ( n12335 , n10842 , n7922 );
nor ( n12336 , n12334 , n12335 );
xnor ( n12337 , n12336 , n7934 );
and ( n12338 , n12333 , n12337 );
and ( n12339 , n11413 , n7963 );
and ( n12340 , n11260 , n7961 );
nor ( n12341 , n12339 , n12340 );
xnor ( n12342 , n12341 , n7973 );
and ( n12343 , n12337 , n12342 );
and ( n12344 , n12333 , n12342 );
or ( n12345 , n12338 , n12343 , n12344 );
and ( n12346 , n12329 , n12345 );
and ( n12347 , n11757 , n7995 );
and ( n12348 , n11581 , n7993 );
nor ( n12349 , n12347 , n12348 );
xnor ( n12350 , n12349 , n8005 );
and ( n12351 , n12101 , n8253 );
and ( n12352 , n11862 , n8251 );
nor ( n12353 , n12351 , n12352 );
xnor ( n12354 , n12353 , n8259 );
and ( n12355 , n12350 , n12354 );
xor ( n12356 , n6506 , n6522 );
buf ( n539617 , n12356 );
buf ( n539618 , n539617 );
buf ( n12359 , n539618 );
and ( n12360 , n12359 , n8106 );
and ( n12361 , n12254 , n8104 );
nor ( n12362 , n12360 , n12361 );
not ( n12363 , n12362 );
and ( n12364 , n12354 , n12363 );
and ( n12365 , n12350 , n12363 );
or ( n12366 , n12355 , n12364 , n12365 );
and ( n12367 , n12345 , n12366 );
and ( n12368 , n12329 , n12366 );
or ( n12369 , n12346 , n12367 , n12368 );
xor ( n12370 , n12143 , n12147 );
xor ( n12371 , n12370 , n12152 );
xor ( n12372 , n12160 , n12164 );
xor ( n12373 , n12372 , n12169 );
and ( n12374 , n12371 , n12373 );
xor ( n12375 , n12179 , n12183 );
xor ( n12376 , n12375 , n12188 );
and ( n12377 , n12373 , n12376 );
and ( n12378 , n12371 , n12376 );
or ( n12379 , n12374 , n12377 , n12378 );
and ( n12380 , n12369 , n12379 );
xor ( n12381 , n12097 , n12105 );
xor ( n12382 , n12381 , n12115 );
and ( n12383 , n12379 , n12382 );
and ( n12384 , n12369 , n12382 );
or ( n12385 , n12380 , n12383 , n12384 );
and ( n12386 , n12313 , n12385 );
xor ( n12387 , n12139 , n12155 );
xor ( n12388 , n12387 , n12172 );
xor ( n12389 , n12191 , n12207 );
xor ( n12390 , n12389 , n12210 );
and ( n12391 , n12388 , n12390 );
xor ( n12392 , n12216 , n12218 );
xor ( n12393 , n12392 , n12221 );
and ( n12394 , n12390 , n12393 );
and ( n12395 , n12388 , n12393 );
or ( n12396 , n12391 , n12394 , n12395 );
and ( n12397 , n12385 , n12396 );
and ( n12398 , n12313 , n12396 );
or ( n12399 , n12386 , n12397 , n12398 );
and ( n12400 , n12248 , n12399 );
xor ( n12401 , n12090 , n12092 );
xor ( n12402 , n12401 , n12118 );
xor ( n12403 , n12175 , n12213 );
xor ( n12404 , n12403 , n12224 );
and ( n12405 , n12402 , n12404 );
xor ( n12406 , n12229 , n12231 );
xor ( n12407 , n12406 , n12234 );
and ( n12408 , n12404 , n12407 );
and ( n12409 , n12402 , n12407 );
or ( n12410 , n12405 , n12408 , n12409 );
and ( n12411 , n12399 , n12410 );
and ( n12412 , n12248 , n12410 );
or ( n12413 , n12400 , n12411 , n12412 );
and ( n12414 , n12245 , n12413 );
and ( n12415 , n12243 , n12413 );
or ( n12416 , n12246 , n12414 , n12415 );
and ( n12417 , n12129 , n12416 );
and ( n12418 , n12127 , n12416 );
or ( n12419 , n12130 , n12417 , n12418 );
and ( n12420 , n12078 , n12419 );
xor ( n12421 , n12078 , n12419 );
xor ( n12422 , n12080 , n12082 );
xor ( n12423 , n12422 , n12124 );
xor ( n12424 , n12085 , n12087 );
xor ( n12425 , n12424 , n12121 );
xor ( n12426 , n12227 , n12237 );
xor ( n12427 , n12426 , n12240 );
and ( n12428 , n12425 , n12427 );
xor ( n12429 , n12195 , n12199 );
xor ( n12430 , n12429 , n12204 );
xor ( n12431 , n12269 , n12273 );
and ( n12432 , n10499 , n7144 );
and ( n12433 , n10419 , n7142 );
nor ( n12434 , n12432 , n12433 );
xnor ( n12435 , n12434 , n7154 );
and ( n12436 , n10842 , n6923 );
and ( n12437 , n10747 , n6921 );
nor ( n12438 , n12436 , n12437 );
xnor ( n12439 , n12438 , n6933 );
and ( n12440 , n12435 , n12439 );
and ( n12441 , n12431 , n12440 );
and ( n12442 , n7939 , n7683 );
and ( n12443 , n7968 , n7680 );
nor ( n12444 , n12442 , n12443 );
xnor ( n12445 , n12444 , n7676 );
and ( n12446 , n8071 , n7762 );
and ( n12447 , n8076 , n7760 );
nor ( n12448 , n12446 , n12447 );
xnor ( n12449 , n12448 , n7772 );
and ( n12450 , n12445 , n12449 );
and ( n12451 , n12440 , n12450 );
and ( n12452 , n12431 , n12450 );
or ( n12453 , n12441 , n12451 , n12452 );
and ( n12454 , n12430 , n12453 );
and ( n12455 , n7979 , n7732 );
and ( n12456 , n8000 , n7730 );
nor ( n12457 , n12455 , n12456 );
xnor ( n12458 , n12457 , n7742 );
and ( n12459 , n8111 , n7797 );
and ( n12460 , n8245 , n7795 );
nor ( n12461 , n12459 , n12460 );
xnor ( n12462 , n12461 , n7807 );
and ( n12463 , n12458 , n12462 );
and ( n12464 , n8595 , n7826 );
and ( n12465 , n8091 , n7824 );
nor ( n12466 , n12464 , n12465 );
xnor ( n12467 , n12466 , n7836 );
and ( n12468 , n12462 , n12467 );
and ( n12469 , n12458 , n12467 );
or ( n12470 , n12463 , n12468 , n12469 );
and ( n12471 , n8604 , n7847 );
and ( n12472 , n8609 , n7845 );
nor ( n12473 , n12471 , n12472 );
xnor ( n12474 , n12473 , n7857 );
and ( n12475 , n9162 , n7036 );
and ( n12476 , n9084 , n7034 );
nor ( n12477 , n12475 , n12476 );
xnor ( n12478 , n12477 , n7125 );
and ( n12479 , n12474 , n12478 );
and ( n12480 , n9482 , n6722 );
and ( n12481 , n9410 , n6720 );
nor ( n12482 , n12480 , n12481 );
xnor ( n12483 , n12482 , n6821 );
and ( n12484 , n12478 , n12483 );
and ( n12485 , n12474 , n12483 );
or ( n12486 , n12479 , n12484 , n12485 );
and ( n12487 , n12470 , n12486 );
and ( n12488 , n9925 , n6852 );
and ( n12489 , n9676 , n6850 );
nor ( n12490 , n12488 , n12489 );
xnor ( n12491 , n12490 , n6862 );
and ( n12492 , n10120 , n7874 );
and ( n12493 , n10055 , n7872 );
nor ( n12494 , n12492 , n12493 );
xnor ( n12495 , n12494 , n7884 );
and ( n12496 , n12491 , n12495 );
and ( n12497 , n11260 , n7924 );
and ( n12498 , n11068 , n7922 );
nor ( n12499 , n12497 , n12498 );
xnor ( n12500 , n12499 , n7934 );
and ( n12501 , n12495 , n12500 );
and ( n12502 , n12491 , n12500 );
or ( n12503 , n12496 , n12501 , n12502 );
and ( n12504 , n12486 , n12503 );
and ( n12505 , n12470 , n12503 );
or ( n12506 , n12487 , n12504 , n12505 );
and ( n12507 , n12453 , n12506 );
and ( n12508 , n12430 , n12506 );
or ( n12509 , n12454 , n12507 , n12508 );
and ( n12510 , n11581 , n7963 );
and ( n12511 , n11413 , n7961 );
nor ( n12512 , n12510 , n12511 );
xnor ( n12513 , n12512 , n7973 );
and ( n12514 , n12254 , n8253 );
and ( n12515 , n12101 , n8251 );
nor ( n12516 , n12514 , n12515 );
xnor ( n12517 , n12516 , n8259 );
and ( n12518 , n12513 , n12517 );
xor ( n12519 , n6512 , n6520 );
buf ( n539780 , n12519 );
buf ( n539781 , n539780 );
buf ( n12522 , n539781 );
and ( n12523 , n12522 , n8106 );
and ( n12524 , n12359 , n8104 );
nor ( n12525 , n12523 , n12524 );
not ( n12526 , n12525 );
and ( n12527 , n12517 , n12526 );
and ( n12528 , n12513 , n12526 );
or ( n12529 , n12518 , n12527 , n12528 );
xor ( n12530 , n12278 , n12282 );
xor ( n12531 , n12530 , n12287 );
and ( n12532 , n12529 , n12531 );
xor ( n12533 , n12295 , n12299 );
xor ( n12534 , n12533 , n12304 );
and ( n12535 , n12531 , n12534 );
and ( n12536 , n12529 , n12534 );
or ( n12537 , n12532 , n12535 , n12536 );
xor ( n12538 , n12317 , n12321 );
xor ( n12539 , n12538 , n12326 );
xor ( n12540 , n12333 , n12337 );
xor ( n12541 , n12540 , n12342 );
and ( n12542 , n12539 , n12541 );
xor ( n12543 , n12350 , n12354 );
xor ( n12544 , n12543 , n12363 );
and ( n12545 , n12541 , n12544 );
and ( n12546 , n12539 , n12544 );
or ( n12547 , n12542 , n12545 , n12546 );
and ( n12548 , n12537 , n12547 );
xor ( n12549 , n12258 , n12259 );
xor ( n12550 , n12549 , n12261 );
and ( n12551 , n12547 , n12550 );
and ( n12552 , n12537 , n12550 );
or ( n12553 , n12548 , n12551 , n12552 );
and ( n12554 , n12509 , n12553 );
xor ( n12555 , n12274 , n12290 );
xor ( n12556 , n12555 , n12307 );
xor ( n12557 , n12329 , n12345 );
xor ( n12558 , n12557 , n12366 );
and ( n12559 , n12556 , n12558 );
xor ( n12560 , n12371 , n12373 );
xor ( n12561 , n12560 , n12376 );
and ( n12562 , n12558 , n12561 );
and ( n12563 , n12556 , n12561 );
or ( n12564 , n12559 , n12562 , n12563 );
and ( n12565 , n12553 , n12564 );
and ( n12566 , n12509 , n12564 );
or ( n12567 , n12554 , n12565 , n12566 );
xor ( n12568 , n12250 , n12264 );
xor ( n12569 , n12568 , n12310 );
xor ( n12570 , n12369 , n12379 );
xor ( n12571 , n12570 , n12382 );
and ( n12572 , n12569 , n12571 );
xor ( n12573 , n12388 , n12390 );
xor ( n12574 , n12573 , n12393 );
and ( n12575 , n12571 , n12574 );
and ( n12576 , n12569 , n12574 );
or ( n12577 , n12572 , n12575 , n12576 );
and ( n12578 , n12567 , n12577 );
xor ( n12579 , n12313 , n12385 );
xor ( n12580 , n12579 , n12396 );
and ( n12581 , n12577 , n12580 );
and ( n12582 , n12567 , n12580 );
or ( n12583 , n12578 , n12581 , n12582 );
and ( n12584 , n12427 , n12583 );
and ( n12585 , n12425 , n12583 );
or ( n12586 , n12428 , n12584 , n12585 );
and ( n12587 , n12423 , n12586 );
xor ( n12588 , n12243 , n12245 );
xor ( n12589 , n12588 , n12413 );
and ( n12590 , n12586 , n12589 );
and ( n12591 , n12423 , n12589 );
or ( n12592 , n12587 , n12590 , n12591 );
xor ( n12593 , n12127 , n12129 );
xor ( n12594 , n12593 , n12416 );
and ( n12595 , n12592 , n12594 );
xor ( n12596 , n12592 , n12594 );
xor ( n12597 , n12248 , n12399 );
xor ( n12598 , n12597 , n12410 );
xor ( n12599 , n12402 , n12404 );
xor ( n12600 , n12599 , n12407 );
and ( n12601 , n12101 , n7995 );
and ( n12602 , n11862 , n7993 );
nor ( n12603 , n12601 , n12602 );
xnor ( n12604 , n12603 , n8005 );
and ( n12605 , n12359 , n8253 );
and ( n12606 , n12254 , n8251 );
nor ( n12607 , n12605 , n12606 );
xnor ( n12608 , n12607 , n8259 );
and ( n12609 , n12604 , n12608 );
and ( n12610 , n11862 , n7995 );
and ( n12611 , n11757 , n7993 );
nor ( n12612 , n12610 , n12611 );
xnor ( n12613 , n12612 , n8005 );
and ( n12614 , n12609 , n12613 );
xor ( n12615 , n12435 , n12439 );
xor ( n12616 , n12445 , n12449 );
and ( n12617 , n12615 , n12616 );
and ( n12618 , n10055 , n6852 );
and ( n12619 , n9925 , n6850 );
nor ( n12620 , n12618 , n12619 );
xnor ( n12621 , n12620 , n6862 );
and ( n12622 , n10419 , n7874 );
and ( n12623 , n10120 , n7872 );
nor ( n12624 , n12622 , n12623 );
xnor ( n12625 , n12624 , n7884 );
and ( n12626 , n12621 , n12625 );
and ( n12627 , n12616 , n12626 );
and ( n12628 , n12615 , n12626 );
or ( n12629 , n12617 , n12627 , n12628 );
and ( n12630 , n12614 , n12629 );
and ( n12631 , n8000 , n7683 );
and ( n12632 , n7939 , n7680 );
nor ( n12633 , n12631 , n12632 );
xnor ( n12634 , n12633 , n7676 );
and ( n12635 , n8076 , n7732 );
and ( n12636 , n7979 , n7730 );
nor ( n12637 , n12635 , n12636 );
xnor ( n12638 , n12637 , n7742 );
and ( n12639 , n12634 , n12638 );
and ( n12640 , n8245 , n7762 );
and ( n12641 , n8071 , n7760 );
nor ( n12642 , n12640 , n12641 );
xnor ( n12643 , n12642 , n7772 );
and ( n12644 , n12638 , n12643 );
and ( n12645 , n12634 , n12643 );
or ( n12646 , n12639 , n12644 , n12645 );
and ( n12647 , n8091 , n7797 );
and ( n12648 , n8111 , n7795 );
nor ( n12649 , n12647 , n12648 );
xnor ( n12650 , n12649 , n7807 );
and ( n12651 , n8609 , n7826 );
and ( n12652 , n8595 , n7824 );
nor ( n12653 , n12651 , n12652 );
xnor ( n12654 , n12653 , n7836 );
and ( n12655 , n12650 , n12654 );
and ( n12656 , n9084 , n7847 );
and ( n12657 , n8604 , n7845 );
nor ( n12658 , n12656 , n12657 );
xnor ( n12659 , n12658 , n7857 );
and ( n12660 , n12654 , n12659 );
and ( n12661 , n12650 , n12659 );
or ( n12662 , n12655 , n12660 , n12661 );
and ( n12663 , n12646 , n12662 );
and ( n12664 , n9410 , n7036 );
and ( n12665 , n9162 , n7034 );
nor ( n12666 , n12664 , n12665 );
xnor ( n12667 , n12666 , n7125 );
and ( n12668 , n9676 , n6722 );
and ( n12669 , n9482 , n6720 );
nor ( n12670 , n12668 , n12669 );
xnor ( n12671 , n12670 , n6821 );
and ( n12672 , n12667 , n12671 );
and ( n12673 , n10747 , n7144 );
and ( n12674 , n10499 , n7142 );
nor ( n12675 , n12673 , n12674 );
xnor ( n12676 , n12675 , n7154 );
and ( n12677 , n12671 , n12676 );
and ( n12678 , n12667 , n12676 );
or ( n12679 , n12672 , n12677 , n12678 );
and ( n12680 , n12662 , n12679 );
and ( n12681 , n12646 , n12679 );
or ( n12682 , n12663 , n12680 , n12681 );
and ( n12683 , n12629 , n12682 );
and ( n12684 , n12614 , n12682 );
or ( n12685 , n12630 , n12683 , n12684 );
and ( n12686 , n11068 , n6923 );
and ( n12687 , n10842 , n6921 );
nor ( n12688 , n12686 , n12687 );
xnor ( n12689 , n12688 , n6933 );
and ( n12690 , n11413 , n7924 );
and ( n12691 , n11260 , n7922 );
nor ( n12692 , n12690 , n12691 );
xnor ( n12693 , n12692 , n7934 );
and ( n12694 , n12689 , n12693 );
and ( n12695 , n11757 , n7963 );
and ( n12696 , n11581 , n7961 );
nor ( n12697 , n12695 , n12696 );
xnor ( n12698 , n12697 , n7973 );
and ( n12699 , n12693 , n12698 );
and ( n12700 , n12689 , n12698 );
or ( n12701 , n12694 , n12699 , n12700 );
xor ( n12702 , n12458 , n12462 );
xor ( n12703 , n12702 , n12467 );
and ( n12704 , n12701 , n12703 );
xor ( n12705 , n12474 , n12478 );
xor ( n12706 , n12705 , n12483 );
and ( n12707 , n12703 , n12706 );
and ( n12708 , n12701 , n12706 );
or ( n12709 , n12704 , n12707 , n12708 );
xor ( n12710 , n12431 , n12440 );
xor ( n12711 , n12710 , n12450 );
and ( n12712 , n12709 , n12711 );
xor ( n12713 , n12470 , n12486 );
xor ( n12714 , n12713 , n12503 );
and ( n12715 , n12711 , n12714 );
and ( n12716 , n12709 , n12714 );
or ( n12717 , n12712 , n12715 , n12716 );
and ( n12718 , n12685 , n12717 );
xor ( n12719 , n12430 , n12453 );
xor ( n12720 , n12719 , n12506 );
and ( n12721 , n12717 , n12720 );
and ( n12722 , n12685 , n12720 );
or ( n12723 , n12718 , n12721 , n12722 );
xor ( n12724 , n12509 , n12553 );
xor ( n12725 , n12724 , n12564 );
and ( n12726 , n12723 , n12725 );
xor ( n12727 , n12569 , n12571 );
xor ( n12728 , n12727 , n12574 );
and ( n12729 , n12725 , n12728 );
and ( n12730 , n12723 , n12728 );
or ( n12731 , n12726 , n12729 , n12730 );
and ( n12732 , n12600 , n12731 );
xor ( n12733 , n12567 , n12577 );
xor ( n12734 , n12733 , n12580 );
and ( n12735 , n12731 , n12734 );
and ( n12736 , n12600 , n12734 );
or ( n12737 , n12732 , n12735 , n12736 );
and ( n12738 , n12598 , n12737 );
xor ( n12739 , n12425 , n12427 );
xor ( n12740 , n12739 , n12583 );
and ( n12741 , n12737 , n12740 );
and ( n12742 , n12598 , n12740 );
or ( n12743 , n12738 , n12741 , n12742 );
xor ( n12744 , n12423 , n12586 );
xor ( n12745 , n12744 , n12589 );
and ( n12746 , n12743 , n12745 );
xor ( n12747 , n12743 , n12745 );
xor ( n12748 , n12598 , n12737 );
xor ( n12749 , n12748 , n12740 );
xor ( n12750 , n12600 , n12731 );
xor ( n12751 , n12750 , n12734 );
xor ( n12752 , n12537 , n12547 );
xor ( n12753 , n12752 , n12550 );
xor ( n12754 , n12556 , n12558 );
xor ( n12755 , n12754 , n12561 );
and ( n12756 , n12753 , n12755 );
xor ( n12757 , n12529 , n12531 );
xor ( n12758 , n12757 , n12534 );
xor ( n12759 , n12539 , n12541 );
xor ( n12760 , n12759 , n12544 );
and ( n12761 , n12758 , n12760 );
xor ( n12762 , n12491 , n12495 );
xor ( n12763 , n12762 , n12500 );
xor ( n12764 , n12513 , n12517 );
xor ( n12765 , n12764 , n12526 );
and ( n12766 , n12763 , n12765 );
xor ( n12767 , n12609 , n12613 );
and ( n12768 , n12765 , n12767 );
and ( n12769 , n12763 , n12767 );
or ( n12770 , n12766 , n12768 , n12769 );
and ( n12771 , n12760 , n12770 );
and ( n12772 , n12758 , n12770 );
or ( n12773 , n12761 , n12771 , n12772 );
and ( n12774 , n12755 , n12773 );
and ( n12775 , n12753 , n12773 );
or ( n12776 , n12756 , n12774 , n12775 );
xor ( n12777 , n12723 , n12725 );
xor ( n12778 , n12777 , n12728 );
and ( n12779 , n12776 , n12778 );
xor ( n12780 , n6516 , n6519 );
buf ( n540041 , n12780 );
buf ( n540042 , n540041 );
buf ( n12783 , n540042 );
and ( n12784 , n12783 , n8106 );
and ( n12785 , n12522 , n8104 );
nor ( n12786 , n12784 , n12785 );
not ( n12787 , n12786 );
xor ( n12788 , n12604 , n12608 );
and ( n12789 , n12787 , n12788 );
xor ( n12790 , n12621 , n12625 );
and ( n12791 , n12788 , n12790 );
and ( n12792 , n12787 , n12790 );
or ( n12793 , n12789 , n12791 , n12792 );
and ( n12794 , n7979 , n7683 );
and ( n12795 , n8000 , n7680 );
nor ( n12796 , n12794 , n12795 );
xnor ( n12797 , n12796 , n7676 );
and ( n12798 , n8071 , n7732 );
and ( n12799 , n8076 , n7730 );
nor ( n12800 , n12798 , n12799 );
xnor ( n12801 , n12800 , n7742 );
and ( n12802 , n12797 , n12801 );
and ( n12803 , n8111 , n7762 );
and ( n12804 , n8245 , n7760 );
nor ( n12805 , n12803 , n12804 );
xnor ( n12806 , n12805 , n7772 );
and ( n12807 , n12801 , n12806 );
and ( n12808 , n12797 , n12806 );
or ( n12809 , n12802 , n12807 , n12808 );
and ( n12810 , n8604 , n7826 );
and ( n12811 , n8609 , n7824 );
nor ( n12812 , n12810 , n12811 );
xnor ( n12813 , n12812 , n7836 );
and ( n12814 , n9162 , n7847 );
and ( n12815 , n9084 , n7845 );
nor ( n12816 , n12814 , n12815 );
xnor ( n12817 , n12816 , n7857 );
and ( n12818 , n12813 , n12817 );
and ( n12819 , n10120 , n6852 );
and ( n12820 , n10055 , n6850 );
nor ( n12821 , n12819 , n12820 );
xnor ( n12822 , n12821 , n6862 );
and ( n12823 , n12817 , n12822 );
and ( n12824 , n12813 , n12822 );
or ( n12825 , n12818 , n12823 , n12824 );
and ( n12826 , n12809 , n12825 );
and ( n12827 , n10499 , n7874 );
and ( n12828 , n10419 , n7872 );
nor ( n12829 , n12827 , n12828 );
xnor ( n12830 , n12829 , n7884 );
and ( n12831 , n10842 , n7144 );
and ( n12832 , n10747 , n7142 );
nor ( n12833 , n12831 , n12832 );
xnor ( n12834 , n12833 , n7154 );
and ( n12835 , n12830 , n12834 );
and ( n12836 , n11260 , n6923 );
and ( n12837 , n11068 , n6921 );
nor ( n12838 , n12836 , n12837 );
xnor ( n12839 , n12838 , n6933 );
and ( n12840 , n12834 , n12839 );
and ( n12841 , n12830 , n12839 );
or ( n12842 , n12835 , n12840 , n12841 );
and ( n12843 , n12825 , n12842 );
and ( n12844 , n12809 , n12842 );
or ( n12845 , n12826 , n12843 , n12844 );
and ( n12846 , n12793 , n12845 );
and ( n12847 , n11581 , n7924 );
and ( n12848 , n11413 , n7922 );
nor ( n12849 , n12847 , n12848 );
xnor ( n12850 , n12849 , n7934 );
and ( n12851 , n11862 , n7963 );
and ( n12852 , n11757 , n7961 );
nor ( n12853 , n12851 , n12852 );
xnor ( n12854 , n12853 , n7973 );
and ( n12855 , n12850 , n12854 );
and ( n12856 , n12254 , n7995 );
and ( n12857 , n12101 , n7993 );
nor ( n12858 , n12856 , n12857 );
xnor ( n12859 , n12858 , n8005 );
and ( n12860 , n12854 , n12859 );
and ( n12861 , n12850 , n12859 );
or ( n12862 , n12855 , n12860 , n12861 );
xor ( n12863 , n12634 , n12638 );
xor ( n12864 , n12863 , n12643 );
and ( n12865 , n12862 , n12864 );
xor ( n12866 , n12650 , n12654 );
xor ( n12867 , n12866 , n12659 );
and ( n12868 , n12864 , n12867 );
and ( n12869 , n12862 , n12867 );
or ( n12870 , n12865 , n12868 , n12869 );
and ( n12871 , n12845 , n12870 );
and ( n12872 , n12793 , n12870 );
or ( n12873 , n12846 , n12871 , n12872 );
xor ( n12874 , n12615 , n12616 );
xor ( n12875 , n12874 , n12626 );
xor ( n12876 , n12646 , n12662 );
xor ( n12877 , n12876 , n12679 );
and ( n12878 , n12875 , n12877 );
xor ( n12879 , n12701 , n12703 );
xor ( n12880 , n12879 , n12706 );
and ( n12881 , n12877 , n12880 );
and ( n12882 , n12875 , n12880 );
or ( n12883 , n12878 , n12881 , n12882 );
and ( n12884 , n12873 , n12883 );
xor ( n12885 , n12614 , n12629 );
xor ( n12886 , n12885 , n12682 );
and ( n12887 , n12883 , n12886 );
and ( n12888 , n12873 , n12886 );
or ( n12889 , n12884 , n12887 , n12888 );
xor ( n12890 , n12685 , n12717 );
xor ( n12891 , n12890 , n12720 );
and ( n12892 , n12889 , n12891 );
xor ( n12893 , n12709 , n12711 );
xor ( n12894 , n12893 , n12714 );
xor ( n12895 , n12667 , n12671 );
xor ( n12896 , n12895 , n12676 );
xor ( n12897 , n12689 , n12693 );
xor ( n12898 , n12897 , n12698 );
and ( n12899 , n12896 , n12898 );
and ( n12900 , n12522 , n8253 );
and ( n12901 , n12359 , n8251 );
nor ( n12902 , n12900 , n12901 );
xnor ( n12903 , n12902 , n8259 );
buf ( n12904 , n6517 );
buf ( n540165 , n12904 );
buf ( n540166 , n540165 );
buf ( n12907 , n540166 );
and ( n12908 , n12907 , n8106 );
and ( n12909 , n12783 , n8104 );
nor ( n12910 , n12908 , n12909 );
not ( n12911 , n12910 );
and ( n12912 , n12903 , n12911 );
and ( n12913 , n8091 , n7762 );
and ( n12914 , n8111 , n7760 );
nor ( n12915 , n12913 , n12914 );
xnor ( n12916 , n12915 , n7772 );
and ( n12917 , n10747 , n7874 );
and ( n12918 , n10499 , n7872 );
nor ( n12919 , n12917 , n12918 );
xnor ( n12920 , n12919 , n7884 );
and ( n12921 , n12916 , n12920 );
and ( n12922 , n11413 , n6923 );
and ( n12923 , n11260 , n6921 );
nor ( n12924 , n12922 , n12923 );
xnor ( n12925 , n12924 , n6933 );
and ( n12926 , n12920 , n12925 );
and ( n12927 , n12916 , n12925 );
or ( n12928 , n12921 , n12926 , n12927 );
and ( n12929 , n12911 , n12928 );
and ( n12930 , n12903 , n12928 );
or ( n12931 , n12912 , n12929 , n12930 );
and ( n12932 , n12898 , n12931 );
and ( n12933 , n12896 , n12931 );
or ( n12934 , n12899 , n12932 , n12933 );
and ( n12935 , n12101 , n7963 );
and ( n12936 , n11862 , n7961 );
nor ( n12937 , n12935 , n12936 );
xnor ( n12938 , n12937 , n7973 );
and ( n12939 , n12783 , n8253 );
and ( n12940 , n12522 , n8251 );
nor ( n12941 , n12939 , n12940 );
xnor ( n12942 , n12941 , n8259 );
and ( n12943 , n12938 , n12942 );
and ( n12944 , n12907 , n8104 );
and ( n12945 , n12942 , n12944 );
and ( n12946 , n12938 , n12944 );
or ( n12947 , n12943 , n12945 , n12946 );
xor ( n12948 , n12797 , n12801 );
xor ( n12949 , n12948 , n12806 );
and ( n12950 , n12947 , n12949 );
xor ( n12951 , n12813 , n12817 );
xor ( n12952 , n12951 , n12822 );
and ( n12953 , n12949 , n12952 );
and ( n12954 , n12947 , n12952 );
or ( n12955 , n12950 , n12953 , n12954 );
xor ( n12956 , n12787 , n12788 );
xor ( n12957 , n12956 , n12790 );
and ( n12958 , n12955 , n12957 );
xor ( n12959 , n12809 , n12825 );
xor ( n12960 , n12959 , n12842 );
and ( n12961 , n12957 , n12960 );
and ( n12962 , n12955 , n12960 );
or ( n12963 , n12958 , n12961 , n12962 );
and ( n12964 , n12934 , n12963 );
xor ( n12965 , n12763 , n12765 );
xor ( n12966 , n12965 , n12767 );
and ( n12967 , n12963 , n12966 );
and ( n12968 , n12934 , n12966 );
or ( n12969 , n12964 , n12967 , n12968 );
and ( n12970 , n12894 , n12969 );
xor ( n12971 , n12758 , n12760 );
xor ( n12972 , n12971 , n12770 );
and ( n12973 , n12969 , n12972 );
and ( n12974 , n12894 , n12972 );
or ( n12975 , n12970 , n12973 , n12974 );
and ( n12976 , n12891 , n12975 );
and ( n12977 , n12889 , n12975 );
or ( n12978 , n12892 , n12976 , n12977 );
and ( n12979 , n12778 , n12978 );
and ( n12980 , n12776 , n12978 );
or ( n12981 , n12779 , n12979 , n12980 );
and ( n12982 , n12751 , n12981 );
xor ( n12983 , n12751 , n12981 );
xor ( n12984 , n12753 , n12755 );
xor ( n12985 , n12984 , n12773 );
xor ( n12986 , n12873 , n12883 );
xor ( n12987 , n12986 , n12886 );
xor ( n12988 , n12793 , n12845 );
xor ( n12989 , n12988 , n12870 );
xor ( n12990 , n12875 , n12877 );
xor ( n12991 , n12990 , n12880 );
and ( n12992 , n12989 , n12991 );
xor ( n12993 , n12862 , n12864 );
xor ( n12994 , n12993 , n12867 );
xor ( n12995 , n12830 , n12834 );
xor ( n12996 , n12995 , n12839 );
xor ( n12997 , n12850 , n12854 );
xor ( n12998 , n12997 , n12859 );
and ( n12999 , n12996 , n12998 );
and ( n13000 , n12254 , n7963 );
and ( n13001 , n12101 , n7961 );
nor ( n13002 , n13000 , n13001 );
xnor ( n13003 , n13002 , n7973 );
and ( n13004 , n12907 , n8251 );
not ( n13005 , n13004 );
and ( n13006 , n13005 , n8259 );
and ( n13007 , n13003 , n13006 );
and ( n13008 , n11757 , n7924 );
and ( n13009 , n11581 , n7922 );
nor ( n13010 , n13008 , n13009 );
xnor ( n13011 , n13010 , n7934 );
and ( n13012 , n13007 , n13011 );
and ( n13013 , n12359 , n7995 );
and ( n13014 , n12254 , n7993 );
nor ( n13015 , n13013 , n13014 );
xnor ( n13016 , n13015 , n8005 );
and ( n13017 , n13011 , n13016 );
and ( n13018 , n13007 , n13016 );
or ( n13019 , n13012 , n13017 , n13018 );
and ( n13020 , n12998 , n13019 );
and ( n13021 , n12996 , n13019 );
or ( n13022 , n12999 , n13020 , n13021 );
and ( n13023 , n12994 , n13022 );
and ( n13024 , n11862 , n7924 );
and ( n13025 , n11757 , n7922 );
nor ( n13026 , n13024 , n13025 );
xnor ( n13027 , n13026 , n7934 );
and ( n13028 , n12522 , n7995 );
and ( n13029 , n12359 , n7993 );
nor ( n13030 , n13028 , n13029 );
xnor ( n13031 , n13030 , n8005 );
and ( n13032 , n13027 , n13031 );
and ( n13033 , n12907 , n8253 );
and ( n13034 , n12783 , n8251 );
nor ( n13035 , n13033 , n13034 );
xnor ( n13036 , n13035 , n8259 );
and ( n13037 , n13031 , n13036 );
and ( n13038 , n13027 , n13036 );
or ( n13039 , n13032 , n13037 , n13038 );
xor ( n13040 , n12916 , n12920 );
xor ( n13041 , n13040 , n12925 );
and ( n13042 , n13039 , n13041 );
xor ( n13043 , n12938 , n12942 );
xor ( n13044 , n13043 , n12944 );
and ( n13045 , n13041 , n13044 );
and ( n13046 , n13039 , n13044 );
or ( n13047 , n13042 , n13045 , n13046 );
xor ( n13048 , n12903 , n12911 );
xor ( n13049 , n13048 , n12928 );
and ( n13050 , n13047 , n13049 );
xor ( n13051 , n12947 , n12949 );
xor ( n13052 , n13051 , n12952 );
and ( n13053 , n13049 , n13052 );
and ( n13054 , n13047 , n13052 );
or ( n13055 , n13050 , n13053 , n13054 );
and ( n13056 , n13022 , n13055 );
and ( n13057 , n12994 , n13055 );
or ( n13058 , n13023 , n13056 , n13057 );
and ( n13059 , n12991 , n13058 );
and ( n13060 , n12989 , n13058 );
or ( n13061 , n12992 , n13059 , n13060 );
and ( n13062 , n12987 , n13061 );
xor ( n13063 , n12894 , n12969 );
xor ( n13064 , n13063 , n12972 );
and ( n13065 , n13061 , n13064 );
and ( n13066 , n12987 , n13064 );
or ( n13067 , n13062 , n13065 , n13066 );
and ( n13068 , n12985 , n13067 );
xor ( n13069 , n12889 , n12891 );
xor ( n13070 , n13069 , n12975 );
and ( n13071 , n13067 , n13070 );
and ( n13072 , n12985 , n13070 );
or ( n13073 , n13068 , n13071 , n13072 );
xor ( n13074 , n12776 , n12778 );
xor ( n13075 , n13074 , n12978 );
and ( n13076 , n13073 , n13075 );
xor ( n13077 , n13073 , n13075 );
xor ( n13078 , n12985 , n13067 );
xor ( n13079 , n13078 , n13070 );
xor ( n13080 , n12934 , n12963 );
xor ( n13081 , n13080 , n12966 );
xor ( n13082 , n12896 , n12898 );
xor ( n13083 , n13082 , n12931 );
xor ( n13084 , n12955 , n12957 );
xor ( n13085 , n13084 , n12960 );
and ( n13086 , n13083 , n13085 );
xor ( n13087 , n13003 , n13006 );
and ( n13088 , n12101 , n7924 );
and ( n13089 , n11862 , n7922 );
nor ( n13090 , n13088 , n13089 );
xnor ( n13091 , n13090 , n7934 );
and ( n13092 , n12359 , n7963 );
and ( n13093 , n12254 , n7961 );
nor ( n13094 , n13092 , n13093 );
xnor ( n13095 , n13094 , n7973 );
and ( n13096 , n13091 , n13095 );
and ( n13097 , n13095 , n13004 );
and ( n13098 , n13091 , n13004 );
or ( n13099 , n13096 , n13097 , n13098 );
and ( n13100 , n13087 , n13099 );
and ( n13101 , n11581 , n6923 );
and ( n13102 , n11413 , n6921 );
nor ( n13103 , n13101 , n13102 );
xnor ( n13104 , n13103 , n6933 );
and ( n13105 , n13099 , n13104 );
and ( n13106 , n13087 , n13104 );
or ( n13107 , n13100 , n13105 , n13106 );
and ( n13108 , n11068 , n7144 );
and ( n13109 , n10842 , n7142 );
nor ( n13110 , n13108 , n13109 );
xnor ( n13111 , n13110 , n7154 );
and ( n13112 , n13107 , n13111 );
xor ( n13113 , n13007 , n13011 );
xor ( n13114 , n13113 , n13016 );
and ( n13115 , n13111 , n13114 );
and ( n13116 , n13107 , n13114 );
or ( n13117 , n13112 , n13115 , n13116 );
xor ( n13118 , n12996 , n12998 );
xor ( n13119 , n13118 , n13019 );
and ( n13120 , n13117 , n13119 );
xor ( n13121 , n13047 , n13049 );
xor ( n13122 , n13121 , n13052 );
and ( n13123 , n13119 , n13122 );
and ( n13124 , n13117 , n13122 );
or ( n13125 , n13120 , n13123 , n13124 );
and ( n13126 , n13085 , n13125 );
and ( n13127 , n13083 , n13125 );
or ( n13128 , n13086 , n13126 , n13127 );
and ( n13129 , n13081 , n13128 );
xor ( n13130 , n12989 , n12991 );
xor ( n13131 , n13130 , n13058 );
and ( n13132 , n13128 , n13131 );
and ( n13133 , n13081 , n13131 );
or ( n13134 , n13129 , n13132 , n13133 );
xor ( n13135 , n12987 , n13061 );
xor ( n13136 , n13135 , n13064 );
and ( n13137 , n13134 , n13136 );
xor ( n13138 , n12994 , n13022 );
xor ( n13139 , n13138 , n13055 );
and ( n13140 , n10055 , n6722 );
and ( n13141 , n9925 , n6720 );
nor ( n13142 , n13140 , n13141 );
xnor ( n13143 , n13142 , n6821 );
and ( n13144 , n10419 , n6852 );
and ( n13145 , n10120 , n6850 );
nor ( n13146 , n13144 , n13145 );
xnor ( n13147 , n13146 , n6862 );
and ( n13148 , n13143 , n13147 );
xor ( n13149 , n13107 , n13111 );
xor ( n13150 , n13149 , n13114 );
and ( n13151 , n13147 , n13150 );
and ( n13152 , n13143 , n13150 );
or ( n13153 , n13148 , n13151 , n13152 );
and ( n13154 , n9482 , n7036 );
and ( n13155 , n9410 , n7034 );
nor ( n13156 , n13154 , n13155 );
xnor ( n13157 , n13156 , n7125 );
and ( n13158 , n13153 , n13157 );
and ( n13159 , n9925 , n6722 );
and ( n13160 , n9676 , n6720 );
nor ( n13161 , n13159 , n13160 );
xnor ( n13162 , n13161 , n6821 );
and ( n13163 , n13157 , n13162 );
and ( n13164 , n13153 , n13162 );
or ( n13165 , n13158 , n13163 , n13164 );
and ( n13166 , n13139 , n13165 );
xor ( n13167 , n13083 , n13085 );
xor ( n13168 , n13167 , n13125 );
and ( n13169 , n13165 , n13168 );
and ( n13170 , n13139 , n13168 );
or ( n13171 , n13166 , n13169 , n13170 );
xor ( n13172 , n13081 , n13128 );
xor ( n13173 , n13172 , n13131 );
and ( n13174 , n13171 , n13173 );
and ( n13175 , n12254 , n7924 );
and ( n13176 , n12101 , n7922 );
nor ( n13177 , n13175 , n13176 );
xnor ( n13178 , n13177 , n7934 );
and ( n13179 , n12907 , n7993 );
not ( n13180 , n13179 );
and ( n13181 , n13180 , n8005 );
xor ( n13182 , n13178 , n13181 );
and ( n13183 , n12101 , n6923 );
and ( n13184 , n11862 , n6921 );
nor ( n13185 , n13183 , n13184 );
xnor ( n13186 , n13185 , n6933 );
and ( n13187 , n12359 , n7924 );
and ( n13188 , n12254 , n7922 );
nor ( n13189 , n13187 , n13188 );
xnor ( n13190 , n13189 , n7934 );
and ( n13191 , n13186 , n13190 );
and ( n13192 , n13190 , n13179 );
and ( n13193 , n13186 , n13179 );
or ( n13194 , n13191 , n13192 , n13193 );
and ( n13195 , n13182 , n13194 );
and ( n13196 , n11581 , n7144 );
and ( n13197 , n11413 , n7142 );
nor ( n13198 , n13196 , n13197 );
xnor ( n13199 , n13198 , n7154 );
and ( n13200 , n13194 , n13199 );
and ( n13201 , n13182 , n13199 );
or ( n13202 , n13195 , n13200 , n13201 );
and ( n13203 , n11068 , n7874 );
and ( n13204 , n10842 , n7872 );
nor ( n13205 , n13203 , n13204 );
xnor ( n13206 , n13205 , n7884 );
and ( n13207 , n13202 , n13206 );
and ( n13208 , n13178 , n13181 );
and ( n13209 , n11757 , n6923 );
and ( n13210 , n11581 , n6921 );
nor ( n13211 , n13209 , n13210 );
xnor ( n13212 , n13211 , n6933 );
xor ( n13213 , n13208 , n13212 );
and ( n13214 , n12783 , n7995 );
and ( n13215 , n12522 , n7993 );
nor ( n13216 , n13214 , n13215 );
xnor ( n13217 , n13216 , n8005 );
xor ( n13218 , n13213 , n13217 );
and ( n13219 , n13206 , n13218 );
and ( n13220 , n13202 , n13218 );
or ( n13221 , n13207 , n13219 , n13220 );
and ( n13222 , n10120 , n6722 );
and ( n13223 , n10055 , n6720 );
nor ( n13224 , n13222 , n13223 );
xnor ( n13225 , n13224 , n6821 );
and ( n13226 , n13221 , n13225 );
and ( n13227 , n13208 , n13212 );
and ( n13228 , n13212 , n13217 );
and ( n13229 , n13208 , n13217 );
or ( n13230 , n13227 , n13228 , n13229 );
and ( n13231 , n11260 , n7144 );
and ( n13232 , n11068 , n7142 );
nor ( n13233 , n13231 , n13232 );
xnor ( n13234 , n13233 , n7154 );
xor ( n13235 , n13230 , n13234 );
xor ( n13236 , n13027 , n13031 );
xor ( n13237 , n13236 , n13036 );
xor ( n13238 , n13235 , n13237 );
and ( n13239 , n13225 , n13238 );
and ( n13240 , n13221 , n13238 );
or ( n13241 , n13226 , n13239 , n13240 );
and ( n13242 , n9084 , n7826 );
and ( n13243 , n8604 , n7824 );
nor ( n13244 , n13242 , n13243 );
xnor ( n13245 , n13244 , n7836 );
and ( n13246 , n13241 , n13245 );
and ( n13247 , n9410 , n7847 );
and ( n13248 , n9162 , n7845 );
nor ( n13249 , n13247 , n13248 );
xnor ( n13250 , n13249 , n7857 );
and ( n13251 , n13245 , n13250 );
and ( n13252 , n13241 , n13250 );
or ( n13253 , n13246 , n13251 , n13252 );
and ( n13254 , n8595 , n7797 );
and ( n13255 , n8091 , n7795 );
nor ( n13256 , n13254 , n13255 );
xnor ( n13257 , n13256 , n7807 );
and ( n13258 , n13253 , n13257 );
xor ( n13259 , n13153 , n13157 );
xor ( n13260 , n13259 , n13162 );
and ( n13261 , n13257 , n13260 );
and ( n13262 , n13253 , n13260 );
or ( n13263 , n13258 , n13261 , n13262 );
and ( n13264 , n11862 , n6923 );
and ( n13265 , n11757 , n6921 );
nor ( n13266 , n13264 , n13265 );
xnor ( n13267 , n13266 , n6933 );
and ( n13268 , n12522 , n7963 );
and ( n13269 , n12359 , n7961 );
nor ( n13270 , n13268 , n13269 );
xnor ( n13271 , n13270 , n7973 );
and ( n13272 , n13267 , n13271 );
and ( n13273 , n12907 , n7995 );
and ( n13274 , n12783 , n7993 );
nor ( n13275 , n13273 , n13274 );
xnor ( n13276 , n13275 , n8005 );
and ( n13277 , n13271 , n13276 );
and ( n13278 , n13267 , n13276 );
or ( n13279 , n13272 , n13277 , n13278 );
and ( n13280 , n11413 , n7144 );
and ( n13281 , n11260 , n7142 );
nor ( n13282 , n13280 , n13281 );
xnor ( n13283 , n13282 , n7154 );
and ( n13284 , n13279 , n13283 );
xor ( n13285 , n13091 , n13095 );
xor ( n13286 , n13285 , n13004 );
and ( n13287 , n13283 , n13286 );
and ( n13288 , n13279 , n13286 );
or ( n13289 , n13284 , n13287 , n13288 );
and ( n13290 , n10842 , n7874 );
and ( n13291 , n10747 , n7872 );
nor ( n13292 , n13290 , n13291 );
xnor ( n13293 , n13292 , n7884 );
and ( n13294 , n13289 , n13293 );
xor ( n13295 , n13087 , n13099 );
xor ( n13296 , n13295 , n13104 );
and ( n13297 , n13293 , n13296 );
and ( n13298 , n13289 , n13296 );
or ( n13299 , n13294 , n13297 , n13298 );
and ( n13300 , n9676 , n7036 );
and ( n13301 , n9482 , n7034 );
nor ( n13302 , n13300 , n13301 );
xnor ( n13303 , n13302 , n7125 );
and ( n13304 , n13299 , n13303 );
xor ( n13305 , n13117 , n13119 );
xor ( n13306 , n13305 , n13122 );
and ( n13307 , n13304 , n13306 );
xor ( n13308 , n13039 , n13041 );
xor ( n13309 , n13308 , n13044 );
and ( n13310 , n13230 , n13234 );
and ( n13311 , n13234 , n13237 );
and ( n13312 , n13230 , n13237 );
or ( n13313 , n13310 , n13311 , n13312 );
and ( n13314 , n13309 , n13313 );
xor ( n13315 , n13299 , n13303 );
and ( n13316 , n13313 , n13315 );
and ( n13317 , n13309 , n13315 );
or ( n13318 , n13314 , n13316 , n13317 );
and ( n13319 , n13306 , n13318 );
and ( n13320 , n13304 , n13318 );
or ( n13321 , n13307 , n13319 , n13320 );
and ( n13322 , n13263 , n13321 );
xor ( n13323 , n13139 , n13165 );
xor ( n13324 , n13323 , n13168 );
and ( n13325 , n13321 , n13324 );
and ( n13326 , n13263 , n13324 );
or ( n13327 , n13322 , n13325 , n13326 );
and ( n13328 , n13173 , n13327 );
and ( n13329 , n13171 , n13327 );
or ( n13330 , n13174 , n13328 , n13329 );
and ( n13331 , n13136 , n13330 );
and ( n13332 , n13134 , n13330 );
or ( n13333 , n13137 , n13331 , n13332 );
and ( n13334 , n13079 , n13333 );
xor ( n13335 , n13079 , n13333 );
xor ( n13336 , n13134 , n13136 );
xor ( n13337 , n13336 , n13330 );
xor ( n13338 , n13171 , n13173 );
xor ( n13339 , n13338 , n13327 );
and ( n13340 , n8604 , n7797 );
and ( n13341 , n8609 , n7795 );
nor ( n13342 , n13340 , n13341 );
xnor ( n13343 , n13342 , n7807 );
and ( n13344 , n9162 , n7826 );
and ( n13345 , n9084 , n7824 );
nor ( n13346 , n13344 , n13345 );
xnor ( n13347 , n13346 , n7836 );
and ( n13348 , n13343 , n13347 );
xor ( n13349 , n13221 , n13225 );
xor ( n13350 , n13349 , n13238 );
and ( n13351 , n13347 , n13350 );
and ( n13352 , n13343 , n13350 );
or ( n13353 , n13348 , n13351 , n13352 );
and ( n13354 , n8245 , n7732 );
and ( n13355 , n8071 , n7730 );
nor ( n13356 , n13354 , n13355 );
xnor ( n13357 , n13356 , n7742 );
and ( n13358 , n13353 , n13357 );
xor ( n13359 , n13241 , n13245 );
xor ( n13360 , n13359 , n13250 );
and ( n13361 , n13357 , n13360 );
and ( n13362 , n13353 , n13360 );
or ( n13363 , n13358 , n13361 , n13362 );
xor ( n13364 , n13253 , n13257 );
xor ( n13365 , n13364 , n13260 );
and ( n13366 , n13363 , n13365 );
xor ( n13367 , n13263 , n13321 );
xor ( n13368 , n13367 , n13324 );
and ( n13369 , n13366 , n13368 );
and ( n13370 , n12254 , n6923 );
and ( n13371 , n12101 , n6921 );
nor ( n13372 , n13370 , n13371 );
xnor ( n13373 , n13372 , n6933 );
and ( n13374 , n12907 , n7961 );
not ( n13375 , n13374 );
and ( n13376 , n13375 , n7973 );
and ( n13377 , n13373 , n13376 );
and ( n13378 , n11757 , n7144 );
and ( n13379 , n11581 , n7142 );
nor ( n13380 , n13378 , n13379 );
xnor ( n13381 , n13380 , n7154 );
and ( n13382 , n13377 , n13381 );
and ( n13383 , n12783 , n7963 );
and ( n13384 , n12522 , n7961 );
nor ( n13385 , n13383 , n13384 );
xnor ( n13386 , n13385 , n7973 );
and ( n13387 , n13381 , n13386 );
and ( n13388 , n13377 , n13386 );
or ( n13389 , n13382 , n13387 , n13388 );
and ( n13390 , n11260 , n7874 );
and ( n13391 , n11068 , n7872 );
nor ( n13392 , n13390 , n13391 );
xnor ( n13393 , n13392 , n7884 );
and ( n13394 , n13389 , n13393 );
xor ( n13395 , n13267 , n13271 );
xor ( n13396 , n13395 , n13276 );
and ( n13397 , n13393 , n13396 );
and ( n13398 , n13389 , n13396 );
or ( n13399 , n13394 , n13397 , n13398 );
and ( n13400 , n10747 , n6852 );
and ( n13401 , n10499 , n6850 );
nor ( n13402 , n13400 , n13401 );
xnor ( n13403 , n13402 , n6862 );
and ( n13404 , n13399 , n13403 );
xor ( n13405 , n13279 , n13283 );
xor ( n13406 , n13405 , n13286 );
and ( n13407 , n13403 , n13406 );
and ( n13408 , n13399 , n13406 );
or ( n13409 , n13404 , n13407 , n13408 );
and ( n13410 , n10499 , n6852 );
and ( n13411 , n10419 , n6850 );
nor ( n13412 , n13410 , n13411 );
xnor ( n13413 , n13412 , n6862 );
and ( n13414 , n13409 , n13413 );
xor ( n13415 , n13289 , n13293 );
xor ( n13416 , n13415 , n13296 );
and ( n13417 , n13413 , n13416 );
and ( n13418 , n13409 , n13416 );
or ( n13419 , n13414 , n13417 , n13418 );
and ( n13420 , n8609 , n7797 );
and ( n13421 , n8595 , n7795 );
nor ( n13422 , n13420 , n13421 );
xnor ( n13423 , n13422 , n7807 );
and ( n13424 , n13419 , n13423 );
xor ( n13425 , n13143 , n13147 );
xor ( n13426 , n13425 , n13150 );
and ( n13427 , n13423 , n13426 );
and ( n13428 , n13419 , n13426 );
or ( n13429 , n13424 , n13427 , n13428 );
xor ( n13430 , n13304 , n13306 );
xor ( n13431 , n13430 , n13318 );
and ( n13432 , n13429 , n13431 );
xor ( n13433 , n13363 , n13365 );
and ( n13434 , n13431 , n13433 );
and ( n13435 , n13429 , n13433 );
or ( n13436 , n13432 , n13434 , n13435 );
and ( n13437 , n13368 , n13436 );
and ( n13438 , n13366 , n13436 );
or ( n13439 , n13369 , n13437 , n13438 );
and ( n13440 , n13339 , n13439 );
and ( n13441 , n11862 , n7144 );
and ( n13442 , n11757 , n7142 );
nor ( n13443 , n13441 , n13442 );
xnor ( n13444 , n13443 , n7154 );
and ( n13445 , n12522 , n7924 );
and ( n13446 , n12359 , n7922 );
nor ( n13447 , n13445 , n13446 );
xnor ( n13448 , n13447 , n7934 );
and ( n13449 , n13444 , n13448 );
and ( n13450 , n12907 , n7963 );
and ( n13451 , n12783 , n7961 );
nor ( n13452 , n13450 , n13451 );
xnor ( n13453 , n13452 , n7973 );
and ( n13454 , n13448 , n13453 );
and ( n13455 , n13444 , n13453 );
or ( n13456 , n13449 , n13454 , n13455 );
and ( n13457 , n11413 , n7874 );
and ( n13458 , n11260 , n7872 );
nor ( n13459 , n13457 , n13458 );
xnor ( n13460 , n13459 , n7884 );
and ( n13461 , n13456 , n13460 );
xor ( n13462 , n13186 , n13190 );
xor ( n13463 , n13462 , n13179 );
and ( n13464 , n13460 , n13463 );
and ( n13465 , n13456 , n13463 );
or ( n13466 , n13461 , n13464 , n13465 );
and ( n13467 , n10842 , n6852 );
and ( n13468 , n10747 , n6850 );
nor ( n13469 , n13467 , n13468 );
xnor ( n13470 , n13469 , n6862 );
and ( n13471 , n13466 , n13470 );
xor ( n13472 , n13182 , n13194 );
xor ( n13473 , n13472 , n13199 );
and ( n13474 , n13470 , n13473 );
and ( n13475 , n13466 , n13473 );
or ( n13476 , n13471 , n13474 , n13475 );
and ( n13477 , n9676 , n7847 );
and ( n13478 , n9482 , n7845 );
nor ( n13479 , n13477 , n13478 );
xnor ( n13480 , n13479 , n7857 );
and ( n13481 , n13476 , n13480 );
xor ( n13482 , n13399 , n13403 );
xor ( n13483 , n13482 , n13406 );
and ( n13484 , n13480 , n13483 );
and ( n13485 , n13476 , n13483 );
or ( n13486 , n13481 , n13484 , n13485 );
and ( n13487 , n8595 , n7762 );
and ( n13488 , n8091 , n7760 );
nor ( n13489 , n13487 , n13488 );
xnor ( n13490 , n13489 , n7772 );
and ( n13491 , n13486 , n13490 );
xor ( n13492 , n13409 , n13413 );
xor ( n13493 , n13492 , n13416 );
and ( n13494 , n13490 , n13493 );
and ( n13495 , n13486 , n13493 );
or ( n13496 , n13491 , n13494 , n13495 );
and ( n13497 , n8076 , n7683 );
and ( n13498 , n7979 , n7680 );
nor ( n13499 , n13497 , n13498 );
xnor ( n13500 , n13499 , n7676 );
and ( n13501 , n13496 , n13500 );
xor ( n13502 , n13419 , n13423 );
xor ( n13503 , n13502 , n13426 );
and ( n13504 , n13500 , n13503 );
and ( n13505 , n13496 , n13503 );
or ( n13506 , n13501 , n13504 , n13505 );
and ( n13507 , n10055 , n7036 );
and ( n13508 , n9925 , n7034 );
nor ( n13509 , n13507 , n13508 );
xnor ( n13510 , n13509 , n7125 );
and ( n13511 , n10419 , n6722 );
and ( n13512 , n10120 , n6720 );
nor ( n13513 , n13511 , n13512 );
xnor ( n13514 , n13513 , n6821 );
and ( n13515 , n13510 , n13514 );
xor ( n13516 , n13202 , n13206 );
xor ( n13517 , n13516 , n13218 );
and ( n13518 , n13514 , n13517 );
and ( n13519 , n13510 , n13517 );
or ( n13520 , n13515 , n13518 , n13519 );
and ( n13521 , n9482 , n7847 );
and ( n13522 , n9410 , n7845 );
nor ( n13523 , n13521 , n13522 );
xnor ( n13524 , n13523 , n7857 );
and ( n13525 , n13520 , n13524 );
and ( n13526 , n9925 , n7036 );
and ( n13527 , n9676 , n7034 );
nor ( n13528 , n13526 , n13527 );
xnor ( n13529 , n13528 , n7125 );
and ( n13530 , n13524 , n13529 );
and ( n13531 , n13520 , n13529 );
or ( n13532 , n13525 , n13530 , n13531 );
xor ( n13533 , n13309 , n13313 );
xor ( n13534 , n13533 , n13315 );
and ( n13535 , n13532 , n13534 );
xor ( n13536 , n13373 , n13376 );
and ( n13537 , n12101 , n7144 );
and ( n13538 , n11862 , n7142 );
nor ( n13539 , n13537 , n13538 );
xnor ( n13540 , n13539 , n7154 );
and ( n13541 , n12783 , n7924 );
and ( n13542 , n12522 , n7922 );
nor ( n13543 , n13541 , n13542 );
xnor ( n13544 , n13543 , n7934 );
and ( n13545 , n13540 , n13544 );
and ( n13546 , n13544 , n13374 );
and ( n13547 , n13540 , n13374 );
or ( n13548 , n13545 , n13546 , n13547 );
and ( n13549 , n13536 , n13548 );
and ( n13550 , n11581 , n7874 );
and ( n13551 , n11413 , n7872 );
nor ( n13552 , n13550 , n13551 );
xnor ( n13553 , n13552 , n7884 );
and ( n13554 , n13548 , n13553 );
and ( n13555 , n13536 , n13553 );
or ( n13556 , n13549 , n13554 , n13555 );
and ( n13557 , n11068 , n6852 );
and ( n13558 , n10842 , n6850 );
nor ( n13559 , n13557 , n13558 );
xnor ( n13560 , n13559 , n6862 );
and ( n13561 , n13556 , n13560 );
xor ( n13562 , n13377 , n13381 );
xor ( n13563 , n13562 , n13386 );
and ( n13564 , n13560 , n13563 );
and ( n13565 , n13556 , n13563 );
or ( n13566 , n13561 , n13564 , n13565 );
and ( n13567 , n10499 , n6722 );
and ( n13568 , n10419 , n6720 );
nor ( n13569 , n13567 , n13568 );
xnor ( n13570 , n13569 , n6821 );
and ( n13571 , n13566 , n13570 );
xor ( n13572 , n13389 , n13393 );
xor ( n13573 , n13572 , n13396 );
and ( n13574 , n13570 , n13573 );
and ( n13575 , n13566 , n13573 );
or ( n13576 , n13571 , n13574 , n13575 );
and ( n13577 , n9410 , n7826 );
and ( n13578 , n9162 , n7824 );
nor ( n13579 , n13577 , n13578 );
xnor ( n13580 , n13579 , n7836 );
and ( n13581 , n13576 , n13580 );
xor ( n13582 , n13510 , n13514 );
xor ( n13583 , n13582 , n13517 );
and ( n13584 , n13580 , n13583 );
and ( n13585 , n13576 , n13583 );
or ( n13586 , n13581 , n13584 , n13585 );
and ( n13587 , n8071 , n7683 );
and ( n13588 , n8076 , n7680 );
nor ( n13589 , n13587 , n13588 );
xnor ( n13590 , n13589 , n7676 );
and ( n13591 , n13586 , n13590 );
xor ( n13592 , n13343 , n13347 );
xor ( n13593 , n13592 , n13350 );
and ( n13594 , n13590 , n13593 );
and ( n13595 , n13586 , n13593 );
or ( n13596 , n13591 , n13594 , n13595 );
and ( n13597 , n13534 , n13596 );
and ( n13598 , n13532 , n13596 );
or ( n13599 , n13535 , n13597 , n13598 );
and ( n13600 , n13506 , n13599 );
and ( n13601 , n10055 , n7847 );
and ( n13602 , n9925 , n7845 );
nor ( n13603 , n13601 , n13602 );
xnor ( n13604 , n13603 , n7857 );
and ( n13605 , n10419 , n7036 );
and ( n13606 , n10120 , n7034 );
nor ( n13607 , n13605 , n13606 );
xnor ( n13608 , n13607 , n7125 );
and ( n13609 , n13604 , n13608 );
xor ( n13610 , n13556 , n13560 );
xor ( n13611 , n13610 , n13563 );
and ( n13612 , n13608 , n13611 );
and ( n13613 , n13604 , n13611 );
or ( n13614 , n13609 , n13612 , n13613 );
and ( n13615 , n9482 , n7826 );
and ( n13616 , n9410 , n7824 );
nor ( n13617 , n13615 , n13616 );
xnor ( n13618 , n13617 , n7836 );
and ( n13619 , n13614 , n13618 );
and ( n13620 , n9925 , n7847 );
and ( n13621 , n9676 , n7845 );
nor ( n13622 , n13620 , n13621 );
xnor ( n13623 , n13622 , n7857 );
and ( n13624 , n13618 , n13623 );
and ( n13625 , n13614 , n13623 );
or ( n13626 , n13619 , n13624 , n13625 );
and ( n13627 , n8091 , n7732 );
and ( n13628 , n8111 , n7730 );
nor ( n13629 , n13627 , n13628 );
xnor ( n13630 , n13629 , n7742 );
and ( n13631 , n13626 , n13630 );
xor ( n13632 , n13476 , n13480 );
xor ( n13633 , n13632 , n13483 );
and ( n13634 , n13630 , n13633 );
and ( n13635 , n13626 , n13633 );
or ( n13636 , n13631 , n13634 , n13635 );
and ( n13637 , n8604 , n7762 );
and ( n13638 , n8609 , n7760 );
nor ( n13639 , n13637 , n13638 );
xnor ( n13640 , n13639 , n7772 );
and ( n13641 , n9162 , n7797 );
and ( n13642 , n9084 , n7795 );
nor ( n13643 , n13641 , n13642 );
xnor ( n13644 , n13643 , n7807 );
and ( n13645 , n13640 , n13644 );
xor ( n13646 , n13566 , n13570 );
xor ( n13647 , n13646 , n13573 );
and ( n13648 , n13644 , n13647 );
and ( n13649 , n13640 , n13647 );
or ( n13650 , n13645 , n13648 , n13649 );
and ( n13651 , n8245 , n7683 );
and ( n13652 , n8071 , n7680 );
nor ( n13653 , n13651 , n13652 );
xnor ( n13654 , n13653 , n7676 );
and ( n13655 , n13650 , n13654 );
xor ( n13656 , n13576 , n13580 );
xor ( n13657 , n13656 , n13583 );
and ( n13658 , n13654 , n13657 );
and ( n13659 , n13650 , n13657 );
or ( n13660 , n13655 , n13658 , n13659 );
and ( n13661 , n13636 , n13660 );
xor ( n13662 , n13486 , n13490 );
xor ( n13663 , n13662 , n13493 );
and ( n13664 , n13660 , n13663 );
and ( n13665 , n13636 , n13663 );
or ( n13666 , n13661 , n13664 , n13665 );
xor ( n13667 , n13353 , n13357 );
xor ( n13668 , n13667 , n13360 );
and ( n13669 , n13666 , n13668 );
xor ( n13670 , n13496 , n13500 );
xor ( n13671 , n13670 , n13503 );
and ( n13672 , n13668 , n13671 );
and ( n13673 , n13666 , n13671 );
or ( n13674 , n13669 , n13672 , n13673 );
and ( n13675 , n13599 , n13674 );
and ( n13676 , n13506 , n13674 );
or ( n13677 , n13600 , n13675 , n13676 );
xor ( n13678 , n13366 , n13368 );
xor ( n13679 , n13678 , n13436 );
and ( n13680 , n13677 , n13679 );
xor ( n13681 , n13429 , n13431 );
xor ( n13682 , n13681 , n13433 );
and ( n13683 , n12254 , n7144 );
and ( n13684 , n12101 , n7142 );
nor ( n13685 , n13683 , n13684 );
xnor ( n13686 , n13685 , n7154 );
and ( n13687 , n12907 , n7922 );
not ( n13688 , n13687 );
and ( n13689 , n13688 , n7934 );
and ( n13690 , n13686 , n13689 );
and ( n13691 , n11757 , n7874 );
and ( n13692 , n11581 , n7872 );
nor ( n13693 , n13691 , n13692 );
xnor ( n13694 , n13693 , n7884 );
and ( n13695 , n13690 , n13694 );
and ( n13696 , n12359 , n6923 );
and ( n13697 , n12254 , n6921 );
nor ( n13698 , n13696 , n13697 );
xnor ( n13699 , n13698 , n6933 );
and ( n13700 , n13694 , n13699 );
and ( n13701 , n13690 , n13699 );
or ( n13702 , n13695 , n13700 , n13701 );
and ( n13703 , n11260 , n6852 );
and ( n13704 , n11068 , n6850 );
nor ( n13705 , n13703 , n13704 );
xnor ( n13706 , n13705 , n6862 );
and ( n13707 , n13702 , n13706 );
xor ( n13708 , n13444 , n13448 );
xor ( n13709 , n13708 , n13453 );
and ( n13710 , n13706 , n13709 );
and ( n13711 , n13702 , n13709 );
or ( n13712 , n13707 , n13710 , n13711 );
and ( n13713 , n10747 , n6722 );
and ( n13714 , n10499 , n6720 );
nor ( n13715 , n13713 , n13714 );
xnor ( n13716 , n13715 , n6821 );
and ( n13717 , n13712 , n13716 );
xor ( n13718 , n13456 , n13460 );
xor ( n13719 , n13718 , n13463 );
and ( n13720 , n13716 , n13719 );
and ( n13721 , n13712 , n13719 );
or ( n13722 , n13717 , n13720 , n13721 );
and ( n13723 , n10120 , n7036 );
and ( n13724 , n10055 , n7034 );
nor ( n13725 , n13723 , n13724 );
xnor ( n13726 , n13725 , n7125 );
and ( n13727 , n13722 , n13726 );
xor ( n13728 , n13466 , n13470 );
xor ( n13729 , n13728 , n13473 );
and ( n13730 , n13726 , n13729 );
and ( n13731 , n13722 , n13729 );
or ( n13732 , n13727 , n13730 , n13731 );
and ( n13733 , n8609 , n7762 );
and ( n13734 , n8595 , n7760 );
nor ( n13735 , n13733 , n13734 );
xnor ( n13736 , n13735 , n7772 );
and ( n13737 , n13732 , n13736 );
and ( n13738 , n9084 , n7797 );
and ( n13739 , n8604 , n7795 );
nor ( n13740 , n13738 , n13739 );
xnor ( n13741 , n13740 , n7807 );
and ( n13742 , n13736 , n13741 );
and ( n13743 , n13732 , n13741 );
or ( n13744 , n13737 , n13742 , n13743 );
and ( n13745 , n8111 , n7732 );
and ( n13746 , n8245 , n7730 );
nor ( n13747 , n13745 , n13746 );
xnor ( n13748 , n13747 , n7742 );
and ( n13749 , n13744 , n13748 );
xor ( n13750 , n13520 , n13524 );
xor ( n13751 , n13750 , n13529 );
and ( n13752 , n13748 , n13751 );
and ( n13753 , n13744 , n13751 );
or ( n13754 , n13749 , n13752 , n13753 );
xor ( n13755 , n13532 , n13534 );
xor ( n13756 , n13755 , n13596 );
and ( n13757 , n13754 , n13756 );
xor ( n13758 , n13666 , n13668 );
xor ( n13759 , n13758 , n13671 );
and ( n13760 , n13756 , n13759 );
and ( n13761 , n13754 , n13759 );
or ( n13762 , n13757 , n13760 , n13761 );
and ( n13763 , n13682 , n13762 );
xor ( n13764 , n13506 , n13599 );
xor ( n13765 , n13764 , n13674 );
and ( n13766 , n13762 , n13765 );
and ( n13767 , n13682 , n13765 );
or ( n13768 , n13763 , n13766 , n13767 );
and ( n13769 , n13679 , n13768 );
and ( n13770 , n13677 , n13768 );
or ( n13771 , n13680 , n13769 , n13770 );
and ( n13772 , n13439 , n13771 );
and ( n13773 , n13339 , n13771 );
or ( n13774 , n13440 , n13772 , n13773 );
and ( n13775 , n13337 , n13774 );
xor ( n13776 , n13337 , n13774 );
xor ( n13777 , n13339 , n13439 );
xor ( n13778 , n13777 , n13771 );
xor ( n13779 , n13677 , n13679 );
xor ( n13780 , n13779 , n13768 );
xor ( n13781 , n13744 , n13748 );
xor ( n13782 , n13781 , n13751 );
xor ( n13783 , n13586 , n13590 );
xor ( n13784 , n13783 , n13593 );
and ( n13785 , n13782 , n13784 );
xor ( n13786 , n13636 , n13660 );
xor ( n13787 , n13786 , n13663 );
and ( n13788 , n13784 , n13787 );
and ( n13789 , n13782 , n13787 );
or ( n13790 , n13785 , n13788 , n13789 );
and ( n13791 , n12522 , n7144 );
and ( n13792 , n12359 , n7142 );
nor ( n13793 , n13791 , n13792 );
xnor ( n13794 , n13793 , n7154 );
and ( n13795 , n12907 , n6921 );
not ( n13796 , n13795 );
and ( n13797 , n13796 , n6933 );
and ( n13798 , n13794 , n13797 );
and ( n13799 , n11757 , n6852 );
and ( n13800 , n11581 , n6850 );
nor ( n13801 , n13799 , n13800 );
xnor ( n13802 , n13801 , n6862 );
and ( n13803 , n13798 , n13802 );
and ( n13804 , n12783 , n6923 );
and ( n13805 , n12522 , n6921 );
nor ( n13806 , n13804 , n13805 );
xnor ( n13807 , n13806 , n6933 );
and ( n13808 , n13802 , n13807 );
and ( n13809 , n13798 , n13807 );
or ( n13810 , n13803 , n13808 , n13809 );
and ( n13811 , n11260 , n6722 );
and ( n13812 , n11068 , n6720 );
nor ( n13813 , n13811 , n13812 );
xnor ( n13814 , n13813 , n6821 );
and ( n13815 , n13810 , n13814 );
and ( n13816 , n11862 , n7874 );
and ( n13817 , n11757 , n7872 );
nor ( n13818 , n13816 , n13817 );
xnor ( n13819 , n13818 , n7884 );
and ( n13820 , n12522 , n6923 );
and ( n13821 , n12359 , n6921 );
nor ( n13822 , n13820 , n13821 );
xnor ( n13823 , n13822 , n6933 );
xor ( n13824 , n13819 , n13823 );
and ( n13825 , n12907 , n7924 );
and ( n13826 , n12783 , n7922 );
nor ( n13827 , n13825 , n13826 );
xnor ( n13828 , n13827 , n7934 );
xor ( n13829 , n13824 , n13828 );
and ( n13830 , n13814 , n13829 );
and ( n13831 , n13810 , n13829 );
or ( n13832 , n13815 , n13830 , n13831 );
and ( n13833 , n10747 , n7036 );
and ( n13834 , n10499 , n7034 );
nor ( n13835 , n13833 , n13834 );
xnor ( n13836 , n13835 , n7125 );
and ( n13837 , n13832 , n13836 );
and ( n13838 , n13819 , n13823 );
and ( n13839 , n13823 , n13828 );
and ( n13840 , n13819 , n13828 );
or ( n13841 , n13838 , n13839 , n13840 );
and ( n13842 , n11413 , n6852 );
and ( n13843 , n11260 , n6850 );
nor ( n13844 , n13842 , n13843 );
xnor ( n13845 , n13844 , n6862 );
xor ( n13846 , n13841 , n13845 );
xor ( n13847 , n13540 , n13544 );
xor ( n13848 , n13847 , n13374 );
xor ( n13849 , n13846 , n13848 );
and ( n13850 , n13836 , n13849 );
and ( n13851 , n13832 , n13849 );
or ( n13852 , n13837 , n13850 , n13851 );
and ( n13853 , n10499 , n7036 );
and ( n13854 , n10419 , n7034 );
nor ( n13855 , n13853 , n13854 );
xnor ( n13856 , n13855 , n7125 );
and ( n13857 , n13852 , n13856 );
and ( n13858 , n13841 , n13845 );
and ( n13859 , n13845 , n13848 );
and ( n13860 , n13841 , n13848 );
or ( n13861 , n13858 , n13859 , n13860 );
and ( n13862 , n10842 , n6722 );
and ( n13863 , n10747 , n6720 );
nor ( n13864 , n13862 , n13863 );
xnor ( n13865 , n13864 , n6821 );
xor ( n13866 , n13861 , n13865 );
xor ( n13867 , n13536 , n13548 );
xor ( n13868 , n13867 , n13553 );
xor ( n13869 , n13866 , n13868 );
and ( n13870 , n13856 , n13869 );
and ( n13871 , n13852 , n13869 );
or ( n13872 , n13857 , n13870 , n13871 );
and ( n13873 , n8609 , n7732 );
and ( n13874 , n8595 , n7730 );
nor ( n13875 , n13873 , n13874 );
xnor ( n13876 , n13875 , n7742 );
and ( n13877 , n13872 , n13876 );
and ( n13878 , n9084 , n7762 );
and ( n13879 , n8604 , n7760 );
nor ( n13880 , n13878 , n13879 );
xnor ( n13881 , n13880 , n7772 );
and ( n13882 , n13876 , n13881 );
and ( n13883 , n13872 , n13881 );
or ( n13884 , n13877 , n13882 , n13883 );
and ( n13885 , n8595 , n7732 );
and ( n13886 , n8091 , n7730 );
nor ( n13887 , n13885 , n13886 );
xnor ( n13888 , n13887 , n7742 );
and ( n13889 , n13884 , n13888 );
xor ( n13890 , n13614 , n13618 );
xor ( n13891 , n13890 , n13623 );
and ( n13892 , n13888 , n13891 );
and ( n13893 , n13884 , n13891 );
or ( n13894 , n13889 , n13892 , n13893 );
and ( n13895 , n13861 , n13865 );
and ( n13896 , n13865 , n13868 );
and ( n13897 , n13861 , n13868 );
or ( n13898 , n13895 , n13896 , n13897 );
and ( n13899 , n9676 , n7826 );
and ( n13900 , n9482 , n7824 );
nor ( n13901 , n13899 , n13900 );
xnor ( n13902 , n13901 , n7836 );
and ( n13903 , n13898 , n13902 );
xor ( n13904 , n13712 , n13716 );
xor ( n13905 , n13904 , n13719 );
and ( n13906 , n13902 , n13905 );
and ( n13907 , n13898 , n13905 );
or ( n13908 , n13903 , n13906 , n13907 );
and ( n13909 , n8111 , n7683 );
and ( n13910 , n8245 , n7680 );
nor ( n13911 , n13909 , n13910 );
xnor ( n13912 , n13911 , n7676 );
and ( n13913 , n13908 , n13912 );
xor ( n13914 , n13722 , n13726 );
xor ( n13915 , n13914 , n13729 );
and ( n13916 , n13912 , n13915 );
and ( n13917 , n13908 , n13915 );
or ( n13918 , n13913 , n13916 , n13917 );
and ( n13919 , n13894 , n13918 );
xor ( n13920 , n13732 , n13736 );
xor ( n13921 , n13920 , n13741 );
and ( n13922 , n13918 , n13921 );
and ( n13923 , n13894 , n13921 );
or ( n13924 , n13919 , n13922 , n13923 );
xor ( n13925 , n13686 , n13689 );
and ( n13926 , n12101 , n7874 );
and ( n13927 , n11862 , n7872 );
nor ( n13928 , n13926 , n13927 );
xnor ( n13929 , n13928 , n7884 );
and ( n13930 , n12359 , n7144 );
and ( n13931 , n12254 , n7142 );
nor ( n13932 , n13930 , n13931 );
xnor ( n13933 , n13932 , n7154 );
and ( n13934 , n13929 , n13933 );
and ( n13935 , n13933 , n13687 );
and ( n13936 , n13929 , n13687 );
or ( n13937 , n13934 , n13935 , n13936 );
and ( n13938 , n13925 , n13937 );
and ( n13939 , n11581 , n6852 );
and ( n13940 , n11413 , n6850 );
nor ( n13941 , n13939 , n13940 );
xnor ( n13942 , n13941 , n6862 );
and ( n13943 , n13937 , n13942 );
and ( n13944 , n13925 , n13942 );
or ( n13945 , n13938 , n13943 , n13944 );
and ( n13946 , n11068 , n6722 );
and ( n13947 , n10842 , n6720 );
nor ( n13948 , n13946 , n13947 );
xnor ( n13949 , n13948 , n6821 );
and ( n13950 , n13945 , n13949 );
xor ( n13951 , n13690 , n13694 );
xor ( n13952 , n13951 , n13699 );
and ( n13953 , n13949 , n13952 );
and ( n13954 , n13945 , n13952 );
or ( n13955 , n13950 , n13953 , n13954 );
and ( n13956 , n10120 , n7847 );
and ( n13957 , n10055 , n7845 );
nor ( n13958 , n13956 , n13957 );
xnor ( n13959 , n13958 , n7857 );
and ( n13960 , n13955 , n13959 );
xor ( n13961 , n13702 , n13706 );
xor ( n13962 , n13961 , n13709 );
and ( n13963 , n13959 , n13962 );
and ( n13964 , n13955 , n13962 );
or ( n13965 , n13960 , n13963 , n13964 );
and ( n13966 , n9410 , n7797 );
and ( n13967 , n9162 , n7795 );
nor ( n13968 , n13966 , n13967 );
xnor ( n13969 , n13968 , n7807 );
and ( n13970 , n13965 , n13969 );
xor ( n13971 , n13604 , n13608 );
xor ( n13972 , n13971 , n13611 );
and ( n13973 , n13969 , n13972 );
and ( n13974 , n13965 , n13972 );
or ( n13975 , n13970 , n13973 , n13974 );
xor ( n13976 , n13640 , n13644 );
xor ( n13977 , n13976 , n13647 );
and ( n13978 , n13975 , n13977 );
xor ( n13979 , n13908 , n13912 );
xor ( n13980 , n13979 , n13915 );
and ( n13981 , n13977 , n13980 );
and ( n13982 , n13975 , n13980 );
or ( n13983 , n13978 , n13981 , n13982 );
xor ( n13984 , n13626 , n13630 );
xor ( n13985 , n13984 , n13633 );
and ( n13986 , n13983 , n13985 );
xor ( n13987 , n13650 , n13654 );
xor ( n13988 , n13987 , n13657 );
and ( n13989 , n13985 , n13988 );
and ( n13990 , n13983 , n13988 );
or ( n13991 , n13986 , n13989 , n13990 );
and ( n13992 , n13924 , n13991 );
xor ( n13993 , n13782 , n13784 );
xor ( n13994 , n13993 , n13787 );
and ( n13995 , n13991 , n13994 );
and ( n13996 , n13924 , n13994 );
or ( n13997 , n13992 , n13995 , n13996 );
and ( n13998 , n13790 , n13997 );
xor ( n13999 , n13754 , n13756 );
xor ( n14000 , n13999 , n13759 );
and ( n14001 , n13997 , n14000 );
and ( n14002 , n13790 , n14000 );
or ( n14003 , n13998 , n14001 , n14002 );
xor ( n14004 , n13682 , n13762 );
xor ( n14005 , n14004 , n13765 );
and ( n14006 , n14003 , n14005 );
xor ( n14007 , n14003 , n14005 );
xor ( n14008 , n13790 , n13997 );
xor ( n14009 , n14008 , n14000 );
xor ( n14010 , n13924 , n13991 );
xor ( n14011 , n14010 , n13994 );
and ( n14012 , n10055 , n7826 );
and ( n14013 , n9925 , n7824 );
nor ( n14014 , n14012 , n14013 );
xnor ( n14015 , n14014 , n7836 );
and ( n14016 , n10419 , n7847 );
and ( n14017 , n10120 , n7845 );
nor ( n14018 , n14016 , n14017 );
xnor ( n14019 , n14018 , n7857 );
and ( n14020 , n14015 , n14019 );
xor ( n14021 , n13945 , n13949 );
xor ( n14022 , n14021 , n13952 );
and ( n14023 , n14019 , n14022 );
and ( n14024 , n14015 , n14022 );
or ( n14025 , n14020 , n14023 , n14024 );
and ( n14026 , n9482 , n7797 );
and ( n14027 , n9410 , n7795 );
nor ( n14028 , n14026 , n14027 );
xnor ( n14029 , n14028 , n7807 );
and ( n14030 , n14025 , n14029 );
and ( n14031 , n9925 , n7826 );
and ( n14032 , n9676 , n7824 );
nor ( n14033 , n14031 , n14032 );
xnor ( n14034 , n14033 , n7836 );
and ( n14035 , n14029 , n14034 );
and ( n14036 , n14025 , n14034 );
or ( n14037 , n14030 , n14035 , n14036 );
and ( n14038 , n8091 , n7683 );
and ( n14039 , n8111 , n7680 );
nor ( n14040 , n14038 , n14039 );
xnor ( n14041 , n14040 , n7676 );
and ( n14042 , n14037 , n14041 );
xor ( n14043 , n13898 , n13902 );
xor ( n14044 , n14043 , n13905 );
and ( n14045 , n14041 , n14044 );
and ( n14046 , n14037 , n14044 );
or ( n14047 , n14042 , n14045 , n14046 );
and ( n14048 , n8604 , n7732 );
and ( n14049 , n8609 , n7730 );
nor ( n14050 , n14048 , n14049 );
xnor ( n14051 , n14050 , n7742 );
and ( n14052 , n9162 , n7762 );
and ( n14053 , n9084 , n7760 );
nor ( n14054 , n14052 , n14053 );
xnor ( n14055 , n14054 , n7772 );
and ( n14056 , n14051 , n14055 );
xor ( n14057 , n13955 , n13959 );
xor ( n14058 , n14057 , n13962 );
and ( n14059 , n14055 , n14058 );
and ( n14060 , n14051 , n14058 );
or ( n14061 , n14056 , n14059 , n14060 );
xor ( n14062 , n13872 , n13876 );
xor ( n14063 , n14062 , n13881 );
and ( n14064 , n14061 , n14063 );
xor ( n14065 , n13965 , n13969 );
xor ( n14066 , n14065 , n13972 );
and ( n14067 , n14063 , n14066 );
and ( n14068 , n14061 , n14066 );
or ( n14069 , n14064 , n14067 , n14068 );
and ( n14070 , n14047 , n14069 );
xor ( n14071 , n13884 , n13888 );
xor ( n14072 , n14071 , n13891 );
and ( n14073 , n14069 , n14072 );
and ( n14074 , n14047 , n14072 );
or ( n14075 , n14070 , n14073 , n14074 );
xor ( n14076 , n13894 , n13918 );
xor ( n14077 , n14076 , n13921 );
and ( n14078 , n14075 , n14077 );
xor ( n14079 , n13983 , n13985 );
xor ( n14080 , n14079 , n13988 );
and ( n14081 , n14077 , n14080 );
and ( n14082 , n14075 , n14080 );
or ( n14083 , n14078 , n14081 , n14082 );
and ( n14084 , n14011 , n14083 );
xor ( n14085 , n14075 , n14077 );
xor ( n14086 , n14085 , n14080 );
xor ( n14087 , n13975 , n13977 );
xor ( n14088 , n14087 , n13980 );
and ( n14089 , n8595 , n7683 );
and ( n14090 , n8091 , n7680 );
nor ( n14091 , n14089 , n14090 );
xnor ( n14092 , n14091 , n7676 );
and ( n14093 , n8609 , n7683 );
and ( n14094 , n8595 , n7680 );
nor ( n14095 , n14093 , n14094 );
xnor ( n14096 , n14095 , n7676 );
and ( n14097 , n9084 , n7732 );
and ( n14098 , n8604 , n7730 );
nor ( n14099 , n14097 , n14098 );
xnor ( n14100 , n14099 , n7742 );
and ( n14101 , n14096 , n14100 );
and ( n14102 , n9410 , n7762 );
and ( n14103 , n9162 , n7760 );
nor ( n14104 , n14102 , n14103 );
xnor ( n14105 , n14104 , n7772 );
and ( n14106 , n14100 , n14105 );
and ( n14107 , n14096 , n14105 );
or ( n14108 , n14101 , n14106 , n14107 );
and ( n14109 , n14092 , n14108 );
and ( n14110 , n9676 , n7797 );
and ( n14111 , n9482 , n7795 );
nor ( n14112 , n14110 , n14111 );
xnor ( n14113 , n14112 , n7807 );
and ( n14114 , n8604 , n7683 );
and ( n14115 , n8609 , n7680 );
nor ( n14116 , n14114 , n14115 );
xnor ( n14117 , n14116 , n7676 );
and ( n14118 , n9162 , n7732 );
and ( n14119 , n9084 , n7730 );
nor ( n14120 , n14118 , n14119 );
xnor ( n14121 , n14120 , n7742 );
and ( n14122 , n14117 , n14121 );
and ( n14123 , n14113 , n14122 );
and ( n14124 , n9482 , n7762 );
and ( n14125 , n9410 , n7760 );
nor ( n14126 , n14124 , n14125 );
xnor ( n14127 , n14126 , n7772 );
and ( n14128 , n9925 , n7797 );
and ( n14129 , n9676 , n7795 );
nor ( n14130 , n14128 , n14129 );
xnor ( n14131 , n14130 , n7807 );
and ( n14132 , n14127 , n14131 );
and ( n14133 , n10120 , n7826 );
and ( n14134 , n10055 , n7824 );
nor ( n14135 , n14133 , n14134 );
xnor ( n14136 , n14135 , n7836 );
and ( n14137 , n14131 , n14136 );
and ( n14138 , n14127 , n14136 );
or ( n14139 , n14132 , n14137 , n14138 );
and ( n14140 , n14122 , n14139 );
and ( n14141 , n14113 , n14139 );
or ( n14142 , n14123 , n14140 , n14141 );
and ( n14143 , n14108 , n14142 );
and ( n14144 , n14092 , n14142 );
or ( n14145 , n14109 , n14143 , n14144 );
xor ( n14146 , n14096 , n14100 );
xor ( n14147 , n14146 , n14105 );
and ( n14148 , n10499 , n7847 );
and ( n14149 , n10419 , n7845 );
nor ( n14150 , n14148 , n14149 );
xnor ( n14151 , n14150 , n7857 );
and ( n14152 , n10842 , n7036 );
and ( n14153 , n10747 , n7034 );
nor ( n14154 , n14152 , n14153 );
xnor ( n14155 , n14154 , n7125 );
and ( n14156 , n14151 , n14155 );
xor ( n14157 , n14117 , n14121 );
and ( n14158 , n14155 , n14157 );
and ( n14159 , n14151 , n14157 );
or ( n14160 , n14156 , n14158 , n14159 );
and ( n14161 , n14147 , n14160 );
and ( n14162 , n9084 , n7683 );
and ( n14163 , n8604 , n7680 );
nor ( n14164 , n14162 , n14163 );
xnor ( n14165 , n14164 , n7676 );
and ( n14166 , n9676 , n7762 );
and ( n14167 , n9482 , n7760 );
nor ( n14168 , n14166 , n14167 );
xnor ( n14169 , n14168 , n7772 );
and ( n14170 , n14165 , n14169 );
and ( n14171 , n10055 , n7797 );
and ( n14172 , n9925 , n7795 );
nor ( n14173 , n14171 , n14172 );
xnor ( n14174 , n14173 , n7807 );
and ( n14175 , n14169 , n14174 );
and ( n14176 , n14165 , n14174 );
or ( n14177 , n14170 , n14175 , n14176 );
and ( n14178 , n10419 , n7826 );
and ( n14179 , n10120 , n7824 );
nor ( n14180 , n14178 , n14179 );
xnor ( n14181 , n14180 , n7836 );
and ( n14182 , n10747 , n7847 );
and ( n14183 , n10499 , n7845 );
nor ( n14184 , n14182 , n14183 );
xnor ( n14185 , n14184 , n7857 );
and ( n14186 , n14181 , n14185 );
and ( n14187 , n11068 , n7036 );
and ( n14188 , n10842 , n7034 );
nor ( n14189 , n14187 , n14188 );
xnor ( n14190 , n14189 , n7125 );
and ( n14191 , n14185 , n14190 );
and ( n14192 , n14181 , n14190 );
or ( n14193 , n14186 , n14191 , n14192 );
and ( n14194 , n14177 , n14193 );
xor ( n14195 , n14127 , n14131 );
xor ( n14196 , n14195 , n14136 );
and ( n14197 , n14193 , n14196 );
and ( n14198 , n14177 , n14196 );
or ( n14199 , n14194 , n14197 , n14198 );
and ( n14200 , n14160 , n14199 );
and ( n14201 , n14147 , n14199 );
or ( n14202 , n14161 , n14200 , n14201 );
xor ( n14203 , n14092 , n14108 );
xor ( n14204 , n14203 , n14142 );
and ( n14205 , n14202 , n14204 );
xor ( n14206 , n14113 , n14122 );
xor ( n14207 , n14206 , n14139 );
xor ( n14208 , n13925 , n13937 );
xor ( n14209 , n14208 , n13942 );
and ( n14210 , n11413 , n6722 );
and ( n14211 , n11260 , n6720 );
nor ( n14212 , n14210 , n14211 );
xnor ( n14213 , n14212 , n6821 );
xor ( n14214 , n13929 , n13933 );
xor ( n14215 , n14214 , n13687 );
and ( n14216 , n14213 , n14215 );
and ( n14217 , n11862 , n6852 );
and ( n14218 , n11757 , n6850 );
nor ( n14219 , n14217 , n14218 );
xnor ( n14220 , n14219 , n6862 );
and ( n14221 , n12254 , n7874 );
and ( n14222 , n12101 , n7872 );
nor ( n14223 , n14221 , n14222 );
xnor ( n14224 , n14223 , n7884 );
and ( n14225 , n14220 , n14224 );
and ( n14226 , n12907 , n6923 );
and ( n14227 , n12783 , n6921 );
nor ( n14228 , n14226 , n14227 );
xnor ( n14229 , n14228 , n6933 );
and ( n14230 , n14224 , n14229 );
and ( n14231 , n14220 , n14229 );
or ( n14232 , n14225 , n14230 , n14231 );
and ( n14233 , n14215 , n14232 );
and ( n14234 , n14213 , n14232 );
or ( n14235 , n14216 , n14233 , n14234 );
and ( n14236 , n14209 , n14235 );
xor ( n14237 , n14151 , n14155 );
xor ( n14238 , n14237 , n14157 );
and ( n14239 , n14235 , n14238 );
and ( n14240 , n14209 , n14238 );
or ( n14241 , n14236 , n14239 , n14240 );
and ( n14242 , n14207 , n14241 );
xor ( n14243 , n14147 , n14160 );
xor ( n14244 , n14243 , n14199 );
and ( n14245 , n14241 , n14244 );
and ( n14246 , n14207 , n14244 );
or ( n14247 , n14242 , n14245 , n14246 );
and ( n14248 , n14204 , n14247 );
and ( n14249 , n14202 , n14247 );
or ( n14250 , n14205 , n14248 , n14249 );
and ( n14251 , n14145 , n14250 );
xor ( n14252 , n14037 , n14041 );
xor ( n14253 , n14252 , n14044 );
and ( n14254 , n14250 , n14253 );
and ( n14255 , n14145 , n14253 );
or ( n14256 , n14251 , n14254 , n14255 );
and ( n14257 , n14088 , n14256 );
xor ( n14258 , n14047 , n14069 );
xor ( n14259 , n14258 , n14072 );
and ( n14260 , n14256 , n14259 );
and ( n14261 , n14088 , n14259 );
or ( n14262 , n14257 , n14260 , n14261 );
and ( n14263 , n14086 , n14262 );
xor ( n14264 , n14025 , n14029 );
xor ( n14265 , n14264 , n14034 );
xor ( n14266 , n13852 , n13856 );
xor ( n14267 , n14266 , n13869 );
and ( n14268 , n14265 , n14267 );
xor ( n14269 , n14051 , n14055 );
xor ( n14270 , n14269 , n14058 );
and ( n14271 , n14267 , n14270 );
and ( n14272 , n14265 , n14270 );
or ( n14273 , n14268 , n14271 , n14272 );
xor ( n14274 , n14061 , n14063 );
xor ( n14275 , n14274 , n14066 );
and ( n14276 , n14273 , n14275 );
xor ( n14277 , n14015 , n14019 );
xor ( n14278 , n14277 , n14022 );
xor ( n14279 , n13832 , n13836 );
xor ( n14280 , n14279 , n13849 );
and ( n14281 , n14278 , n14280 );
xor ( n14282 , n14177 , n14193 );
xor ( n14283 , n14282 , n14196 );
xor ( n14284 , n13810 , n13814 );
xor ( n14285 , n14284 , n13829 );
and ( n14286 , n14283 , n14285 );
xor ( n14287 , n14165 , n14169 );
xor ( n14288 , n14287 , n14174 );
xor ( n14289 , n14181 , n14185 );
xor ( n14290 , n14289 , n14190 );
and ( n14291 , n14288 , n14290 );
xor ( n14292 , n13798 , n13802 );
xor ( n14293 , n14292 , n13807 );
and ( n14294 , n14290 , n14293 );
and ( n14295 , n14288 , n14293 );
or ( n14296 , n14291 , n14294 , n14295 );
and ( n14297 , n14285 , n14296 );
and ( n14298 , n14283 , n14296 );
or ( n14299 , n14286 , n14297 , n14298 );
and ( n14300 , n14280 , n14299 );
and ( n14301 , n14278 , n14299 );
or ( n14302 , n14281 , n14300 , n14301 );
xor ( n14303 , n14202 , n14204 );
xor ( n14304 , n14303 , n14247 );
and ( n14305 , n14302 , n14304 );
xor ( n14306 , n14207 , n14241 );
xor ( n14307 , n14306 , n14244 );
xor ( n14308 , n14209 , n14235 );
xor ( n14309 , n14308 , n14238 );
and ( n14310 , n12359 , n7874 );
and ( n14311 , n12254 , n7872 );
nor ( n14312 , n14310 , n14311 );
xnor ( n14313 , n14312 , n7884 );
and ( n14314 , n12783 , n7144 );
and ( n14315 , n12522 , n7142 );
nor ( n14316 , n14314 , n14315 );
xnor ( n14317 , n14316 , n7154 );
and ( n14318 , n14313 , n14317 );
and ( n14319 , n14317 , n13795 );
and ( n14320 , n14313 , n13795 );
or ( n14321 , n14318 , n14319 , n14320 );
xor ( n14322 , n13794 , n13797 );
and ( n14323 , n14321 , n14322 );
xor ( n14324 , n14213 , n14215 );
xor ( n14325 , n14324 , n14232 );
and ( n14326 , n14323 , n14325 );
and ( n14327 , n12254 , n6852 );
and ( n14328 , n12101 , n6850 );
nor ( n14329 , n14327 , n14328 );
xnor ( n14330 , n14329 , n6862 );
and ( n14331 , n12907 , n7142 );
not ( n14332 , n14331 );
and ( n14333 , n14332 , n7154 );
and ( n14334 , n14330 , n14333 );
and ( n14335 , n11757 , n6722 );
and ( n14336 , n11581 , n6720 );
nor ( n14337 , n14335 , n14336 );
xnor ( n14338 , n14337 , n6821 );
and ( n14339 , n14334 , n14338 );
and ( n14340 , n12101 , n6852 );
and ( n14341 , n11862 , n6850 );
nor ( n14342 , n14340 , n14341 );
xnor ( n14343 , n14342 , n6862 );
and ( n14344 , n14338 , n14343 );
and ( n14345 , n14334 , n14343 );
or ( n14346 , n14339 , n14344 , n14345 );
and ( n14347 , n11260 , n7036 );
and ( n14348 , n11068 , n7034 );
nor ( n14349 , n14347 , n14348 );
xnor ( n14350 , n14349 , n7125 );
and ( n14351 , n14346 , n14350 );
xor ( n14352 , n14220 , n14224 );
xor ( n14353 , n14352 , n14229 );
and ( n14354 , n14350 , n14353 );
and ( n14355 , n14346 , n14353 );
or ( n14356 , n14351 , n14354 , n14355 );
and ( n14357 , n14325 , n14356 );
and ( n14358 , n14323 , n14356 );
or ( n14359 , n14326 , n14357 , n14358 );
and ( n14360 , n14309 , n14359 );
xor ( n14361 , n14283 , n14285 );
xor ( n14362 , n14361 , n14296 );
and ( n14363 , n14359 , n14362 );
and ( n14364 , n14309 , n14362 );
or ( n14365 , n14360 , n14363 , n14364 );
and ( n14366 , n14307 , n14365 );
xor ( n14367 , n14278 , n14280 );
xor ( n14368 , n14367 , n14299 );
and ( n14369 , n14365 , n14368 );
and ( n14370 , n14307 , n14368 );
or ( n14371 , n14366 , n14369 , n14370 );
and ( n14372 , n14304 , n14371 );
and ( n14373 , n14302 , n14371 );
or ( n14374 , n14305 , n14372 , n14373 );
and ( n14375 , n14275 , n14374 );
and ( n14376 , n14273 , n14374 );
or ( n14377 , n14276 , n14375 , n14376 );
xor ( n14378 , n14088 , n14256 );
xor ( n14379 , n14378 , n14259 );
and ( n14380 , n14377 , n14379 );
xor ( n14381 , n14145 , n14250 );
xor ( n14382 , n14381 , n14253 );
xor ( n14383 , n14273 , n14275 );
xor ( n14384 , n14383 , n14374 );
and ( n14385 , n14382 , n14384 );
xor ( n14386 , n14265 , n14267 );
xor ( n14387 , n14386 , n14270 );
xor ( n14388 , n14302 , n14304 );
xor ( n14389 , n14388 , n14371 );
and ( n14390 , n14387 , n14389 );
xor ( n14391 , n14307 , n14365 );
xor ( n14392 , n14391 , n14368 );
and ( n14393 , n10120 , n7797 );
and ( n14394 , n10055 , n7795 );
nor ( n14395 , n14393 , n14394 );
xnor ( n14396 , n14395 , n7807 );
and ( n14397 , n11581 , n6722 );
and ( n14398 , n11413 , n6720 );
nor ( n14399 , n14397 , n14398 );
xnor ( n14400 , n14399 , n6821 );
and ( n14401 , n14396 , n14400 );
xor ( n14402 , n14321 , n14322 );
and ( n14403 , n14400 , n14402 );
and ( n14404 , n14396 , n14402 );
or ( n14405 , n14401 , n14403 , n14404 );
xor ( n14406 , n14288 , n14290 );
xor ( n14407 , n14406 , n14293 );
and ( n14408 , n14405 , n14407 );
xor ( n14409 , n14346 , n14350 );
xor ( n14410 , n14409 , n14353 );
xor ( n14411 , n14330 , n14333 );
and ( n14412 , n12522 , n7874 );
and ( n14413 , n12359 , n7872 );
nor ( n14414 , n14412 , n14413 );
xnor ( n14415 , n14414 , n7884 );
and ( n14416 , n14411 , n14415 );
and ( n14417 , n12907 , n7144 );
and ( n14418 , n12783 , n7142 );
nor ( n14419 , n14417 , n14418 );
xnor ( n14420 , n14419 , n7154 );
and ( n14421 , n14415 , n14420 );
and ( n14422 , n14411 , n14420 );
or ( n14423 , n14416 , n14421 , n14422 );
and ( n14424 , n11413 , n7036 );
and ( n14425 , n11260 , n7034 );
nor ( n14426 , n14424 , n14425 );
xnor ( n14427 , n14426 , n7125 );
and ( n14428 , n14423 , n14427 );
xor ( n14429 , n14313 , n14317 );
xor ( n14430 , n14429 , n13795 );
and ( n14431 , n14427 , n14430 );
and ( n14432 , n14423 , n14430 );
or ( n14433 , n14428 , n14431 , n14432 );
and ( n14434 , n14410 , n14433 );
xor ( n14435 , n14396 , n14400 );
xor ( n14436 , n14435 , n14402 );
and ( n14437 , n14433 , n14436 );
and ( n14438 , n14410 , n14436 );
or ( n14439 , n14434 , n14437 , n14438 );
and ( n14440 , n14407 , n14439 );
and ( n14441 , n14405 , n14439 );
or ( n14442 , n14408 , n14440 , n14441 );
xor ( n14443 , n14309 , n14359 );
xor ( n14444 , n14443 , n14362 );
and ( n14445 , n14442 , n14444 );
and ( n14446 , n12101 , n6722 );
and ( n14447 , n11862 , n6720 );
nor ( n14448 , n14446 , n14447 );
xnor ( n14449 , n14448 , n6821 );
and ( n14450 , n12359 , n6852 );
and ( n14451 , n12254 , n6850 );
nor ( n14452 , n14450 , n14451 );
xnor ( n14453 , n14452 , n6862 );
and ( n14454 , n14449 , n14453 );
and ( n14455 , n14453 , n14331 );
and ( n14456 , n14449 , n14331 );
or ( n14457 , n14454 , n14455 , n14456 );
and ( n14458 , n11862 , n6722 );
and ( n14459 , n11757 , n6720 );
nor ( n14460 , n14458 , n14459 );
xnor ( n14461 , n14460 , n6821 );
and ( n14462 , n14457 , n14461 );
xor ( n14463 , n14411 , n14415 );
xor ( n14464 , n14463 , n14420 );
and ( n14465 , n14461 , n14464 );
and ( n14466 , n14457 , n14464 );
or ( n14467 , n14462 , n14465 , n14466 );
xor ( n14468 , n14334 , n14338 );
xor ( n14469 , n14468 , n14343 );
and ( n14470 , n14467 , n14469 );
xor ( n14471 , n14423 , n14427 );
xor ( n14472 , n14471 , n14430 );
and ( n14473 , n14469 , n14472 );
and ( n14474 , n14467 , n14472 );
or ( n14475 , n14470 , n14473 , n14474 );
and ( n14476 , n10499 , n7826 );
and ( n14477 , n10419 , n7824 );
nor ( n14478 , n14476 , n14477 );
xnor ( n14479 , n14478 , n7836 );
and ( n14480 , n14475 , n14479 );
and ( n14481 , n10842 , n7847 );
and ( n14482 , n10747 , n7845 );
nor ( n14483 , n14481 , n14482 );
xnor ( n14484 , n14483 , n7857 );
and ( n14485 , n14479 , n14484 );
and ( n14486 , n14475 , n14484 );
or ( n14487 , n14480 , n14485 , n14486 );
and ( n14488 , n9410 , n7732 );
and ( n14489 , n9162 , n7730 );
nor ( n14490 , n14488 , n14489 );
xnor ( n14491 , n14490 , n7742 );
and ( n14492 , n14487 , n14491 );
and ( n14493 , n14444 , n14492 );
and ( n14494 , n14442 , n14492 );
or ( n14495 , n14445 , n14493 , n14494 );
and ( n14496 , n14392 , n14495 );
xor ( n14497 , n14323 , n14325 );
xor ( n14498 , n14497 , n14356 );
xor ( n14499 , n14405 , n14407 );
xor ( n14500 , n14499 , n14439 );
and ( n14501 , n14498 , n14500 );
xor ( n14502 , n14487 , n14491 );
and ( n14503 , n14500 , n14502 );
and ( n14504 , n14498 , n14502 );
or ( n14505 , n14501 , n14503 , n14504 );
xor ( n14506 , n14442 , n14444 );
xor ( n14507 , n14506 , n14492 );
and ( n14508 , n14505 , n14507 );
and ( n14509 , n10055 , n7762 );
and ( n14510 , n9925 , n7760 );
nor ( n14511 , n14509 , n14510 );
xnor ( n14512 , n14511 , n7772 );
and ( n14513 , n10419 , n7797 );
and ( n14514 , n10120 , n7795 );
nor ( n14515 , n14513 , n14514 );
xnor ( n14516 , n14515 , n7807 );
and ( n14517 , n14512 , n14516 );
xor ( n14518 , n14467 , n14469 );
xor ( n14519 , n14518 , n14472 );
and ( n14520 , n14516 , n14519 );
and ( n14521 , n14512 , n14519 );
or ( n14522 , n14517 , n14520 , n14521 );
and ( n14523 , n9482 , n7732 );
and ( n14524 , n9410 , n7730 );
nor ( n14525 , n14523 , n14524 );
xnor ( n14526 , n14525 , n7742 );
and ( n14527 , n14522 , n14526 );
and ( n14528 , n9925 , n7762 );
and ( n14529 , n9676 , n7760 );
nor ( n14530 , n14528 , n14529 );
xnor ( n14531 , n14530 , n7772 );
and ( n14532 , n14526 , n14531 );
and ( n14533 , n14522 , n14531 );
or ( n14534 , n14527 , n14532 , n14533 );
and ( n14535 , n12254 , n6722 );
and ( n14536 , n12101 , n6720 );
nor ( n14537 , n14535 , n14536 );
xnor ( n14538 , n14537 , n6821 );
and ( n14539 , n12907 , n7872 );
not ( n14540 , n14539 );
and ( n14541 , n14540 , n7884 );
xor ( n14542 , n14538 , n14541 );
and ( n14543 , n12522 , n6852 );
and ( n14544 , n12359 , n6850 );
nor ( n14545 , n14543 , n14544 );
xnor ( n14546 , n14545 , n6862 );
and ( n14547 , n14542 , n14546 );
and ( n14548 , n12907 , n7874 );
and ( n14549 , n12783 , n7872 );
nor ( n14550 , n14548 , n14549 );
xnor ( n14551 , n14550 , n7884 );
and ( n14552 , n14546 , n14551 );
and ( n14553 , n14542 , n14551 );
or ( n14554 , n14547 , n14552 , n14553 );
and ( n14555 , n11413 , n7847 );
and ( n14556 , n11260 , n7845 );
nor ( n14557 , n14555 , n14556 );
xnor ( n14558 , n14557 , n7857 );
and ( n14559 , n14554 , n14558 );
xor ( n14560 , n14449 , n14453 );
xor ( n14561 , n14560 , n14331 );
and ( n14562 , n14558 , n14561 );
and ( n14563 , n14554 , n14561 );
or ( n14564 , n14559 , n14562 , n14563 );
and ( n14565 , n11260 , n7847 );
and ( n14566 , n11068 , n7845 );
nor ( n14567 , n14565 , n14566 );
xnor ( n14568 , n14567 , n7857 );
and ( n14569 , n14564 , n14568 );
and ( n14570 , n14538 , n14541 );
and ( n14571 , n11757 , n7036 );
and ( n14572 , n11581 , n7034 );
nor ( n14573 , n14571 , n14572 );
xnor ( n14574 , n14573 , n7125 );
and ( n14575 , n14570 , n14574 );
and ( n14576 , n12783 , n7874 );
and ( n14577 , n12522 , n7872 );
nor ( n14578 , n14576 , n14577 );
xnor ( n14579 , n14578 , n7884 );
and ( n14580 , n14574 , n14579 );
and ( n14581 , n14570 , n14579 );
or ( n14582 , n14575 , n14580 , n14581 );
and ( n14583 , n11581 , n7036 );
and ( n14584 , n11413 , n7034 );
nor ( n14585 , n14583 , n14584 );
xnor ( n14586 , n14585 , n7125 );
xor ( n14587 , n14582 , n14586 );
xor ( n14588 , n14457 , n14461 );
xor ( n14589 , n14588 , n14464 );
xor ( n14590 , n14587 , n14589 );
and ( n14591 , n14568 , n14590 );
and ( n14592 , n14564 , n14590 );
or ( n14593 , n14569 , n14591 , n14592 );
and ( n14594 , n9676 , n7732 );
and ( n14595 , n9482 , n7730 );
nor ( n14596 , n14594 , n14595 );
xnor ( n14597 , n14596 , n7742 );
and ( n14598 , n14593 , n14597 );
and ( n14599 , n14582 , n14586 );
and ( n14600 , n14586 , n14589 );
and ( n14601 , n14582 , n14589 );
or ( n14602 , n14599 , n14600 , n14601 );
and ( n14603 , n10747 , n7826 );
and ( n14604 , n10499 , n7824 );
nor ( n14605 , n14603 , n14604 );
xnor ( n14606 , n14605 , n7836 );
xor ( n14607 , n14602 , n14606 );
and ( n14608 , n11068 , n7847 );
and ( n14609 , n10842 , n7845 );
nor ( n14610 , n14608 , n14609 );
xnor ( n14611 , n14610 , n7857 );
xor ( n14612 , n14607 , n14611 );
and ( n14613 , n14597 , n14612 );
and ( n14614 , n14593 , n14612 );
or ( n14615 , n14598 , n14613 , n14614 );
and ( n14616 , n9162 , n7683 );
and ( n14617 , n9084 , n7680 );
nor ( n14618 , n14616 , n14617 );
xnor ( n14619 , n14618 , n7676 );
and ( n14620 , n14615 , n14619 );
xor ( n14621 , n14475 , n14479 );
xor ( n14622 , n14621 , n14484 );
and ( n14623 , n14619 , n14622 );
and ( n14624 , n14615 , n14622 );
or ( n14625 , n14620 , n14623 , n14624 );
and ( n14626 , n14534 , n14625 );
xor ( n14627 , n14410 , n14433 );
xor ( n14628 , n14627 , n14436 );
and ( n14629 , n14602 , n14606 );
and ( n14630 , n14606 , n14611 );
and ( n14631 , n14602 , n14611 );
or ( n14632 , n14629 , n14630 , n14631 );
and ( n14633 , n14628 , n14632 );
xor ( n14634 , n14522 , n14526 );
xor ( n14635 , n14634 , n14531 );
and ( n14636 , n14632 , n14635 );
and ( n14637 , n14628 , n14635 );
or ( n14638 , n14633 , n14636 , n14637 );
and ( n14639 , n14625 , n14638 );
and ( n14640 , n14534 , n14638 );
or ( n14641 , n14626 , n14639 , n14640 );
and ( n14642 , n14507 , n14641 );
and ( n14643 , n14505 , n14641 );
or ( n14644 , n14508 , n14642 , n14643 );
and ( n14645 , n14495 , n14644 );
and ( n14646 , n14392 , n14644 );
or ( n14647 , n14496 , n14645 , n14646 );
and ( n14648 , n14389 , n14647 );
and ( n14649 , n14387 , n14647 );
or ( n14650 , n14390 , n14648 , n14649 );
and ( n14651 , n14384 , n14650 );
and ( n14652 , n14382 , n14650 );
or ( n14653 , n14385 , n14651 , n14652 );
and ( n14654 , n14379 , n14653 );
and ( n14655 , n14377 , n14653 );
or ( n14656 , n14380 , n14654 , n14655 );
and ( n14657 , n14262 , n14656 );
and ( n14658 , n14086 , n14656 );
or ( n14659 , n14263 , n14657 , n14658 );
and ( n14660 , n14083 , n14659 );
and ( n14661 , n14011 , n14659 );
or ( n14662 , n14084 , n14660 , n14661 );
and ( n14663 , n14009 , n14662 );
xor ( n14664 , n14009 , n14662 );
xor ( n14665 , n14011 , n14083 );
xor ( n14666 , n14665 , n14659 );
xor ( n14667 , n14086 , n14262 );
xor ( n14668 , n14667 , n14656 );
xor ( n14669 , n14377 , n14379 );
xor ( n14670 , n14669 , n14653 );
xor ( n14671 , n14382 , n14384 );
xor ( n14672 , n14671 , n14650 );
xor ( n14673 , n14387 , n14389 );
xor ( n14674 , n14673 , n14647 );
xor ( n14675 , n14392 , n14495 );
xor ( n14676 , n14675 , n14644 );
xor ( n14677 , n14498 , n14500 );
xor ( n14678 , n14677 , n14502 );
and ( n14679 , n10055 , n7732 );
and ( n14680 , n9925 , n7730 );
nor ( n14681 , n14679 , n14680 );
xnor ( n14682 , n14681 , n7742 );
and ( n14683 , n10419 , n7762 );
and ( n14684 , n10120 , n7760 );
nor ( n14685 , n14683 , n14684 );
xnor ( n14686 , n14685 , n7772 );
and ( n14687 , n14682 , n14686 );
and ( n14688 , n12359 , n6722 );
and ( n14689 , n12254 , n6720 );
nor ( n14690 , n14688 , n14689 );
xnor ( n14691 , n14690 , n6821 );
and ( n14692 , n12783 , n6852 );
and ( n14693 , n12522 , n6850 );
nor ( n14694 , n14692 , n14693 );
xnor ( n14695 , n14694 , n6862 );
and ( n14696 , n14691 , n14695 );
and ( n14697 , n14695 , n14539 );
and ( n14698 , n14691 , n14539 );
or ( n14699 , n14696 , n14697 , n14698 );
and ( n14700 , n11862 , n7036 );
and ( n14701 , n11757 , n7034 );
nor ( n14702 , n14700 , n14701 );
xnor ( n14703 , n14702 , n7125 );
and ( n14704 , n14699 , n14703 );
xor ( n14705 , n14542 , n14546 );
xor ( n14706 , n14705 , n14551 );
and ( n14707 , n14703 , n14706 );
and ( n14708 , n14699 , n14706 );
or ( n14709 , n14704 , n14707 , n14708 );
xor ( n14710 , n14570 , n14574 );
xor ( n14711 , n14710 , n14579 );
xor ( n14712 , n14709 , n14711 );
xor ( n14713 , n14554 , n14558 );
xor ( n14714 , n14713 , n14561 );
xor ( n14715 , n14712 , n14714 );
and ( n14716 , n14686 , n14715 );
and ( n14717 , n14682 , n14715 );
or ( n14718 , n14687 , n14716 , n14717 );
and ( n14719 , n9482 , n7683 );
and ( n14720 , n9410 , n7680 );
nor ( n14721 , n14719 , n14720 );
xnor ( n14722 , n14721 , n7676 );
and ( n14723 , n14718 , n14722 );
and ( n14724 , n9925 , n7732 );
and ( n14725 , n9676 , n7730 );
nor ( n14726 , n14724 , n14725 );
xnor ( n14727 , n14726 , n7742 );
and ( n14728 , n14722 , n14727 );
and ( n14729 , n14718 , n14727 );
or ( n14730 , n14723 , n14728 , n14729 );
xor ( n14731 , n14593 , n14597 );
xor ( n14732 , n14731 , n14612 );
and ( n14733 , n14730 , n14732 );
xor ( n14734 , n14512 , n14516 );
xor ( n14735 , n14734 , n14519 );
and ( n14736 , n14732 , n14735 );
and ( n14737 , n14730 , n14735 );
or ( n14738 , n14733 , n14736 , n14737 );
xor ( n14739 , n14615 , n14619 );
xor ( n14740 , n14739 , n14622 );
and ( n14741 , n14738 , n14740 );
and ( n14742 , n14678 , n14741 );
xor ( n14743 , n14534 , n14625 );
xor ( n14744 , n14743 , n14638 );
and ( n14745 , n14741 , n14744 );
and ( n14746 , n14678 , n14744 );
or ( n14747 , n14742 , n14745 , n14746 );
xor ( n14748 , n14505 , n14507 );
xor ( n14749 , n14748 , n14641 );
and ( n14750 , n14747 , n14749 );
and ( n14751 , n14709 , n14711 );
and ( n14752 , n14711 , n14714 );
and ( n14753 , n14709 , n14714 );
or ( n14754 , n14751 , n14752 , n14753 );
and ( n14755 , n10120 , n7762 );
and ( n14756 , n10055 , n7760 );
nor ( n14757 , n14755 , n14756 );
xnor ( n14758 , n14757 , n7772 );
and ( n14759 , n14754 , n14758 );
and ( n14760 , n10842 , n7826 );
and ( n14761 , n10747 , n7824 );
nor ( n14762 , n14760 , n14761 );
xnor ( n14763 , n14762 , n7836 );
and ( n14764 , n14758 , n14763 );
and ( n14765 , n14754 , n14763 );
or ( n14766 , n14759 , n14764 , n14765 );
and ( n14767 , n12522 , n6722 );
and ( n14768 , n12359 , n6720 );
nor ( n14769 , n14767 , n14768 );
xnor ( n14770 , n14769 , n6821 );
and ( n14771 , n12907 , n6850 );
not ( n14772 , n14771 );
and ( n14773 , n14772 , n6862 );
and ( n14774 , n14770 , n14773 );
and ( n14775 , n12101 , n7036 );
and ( n14776 , n11862 , n7034 );
nor ( n14777 , n14775 , n14776 );
xnor ( n14778 , n14777 , n7125 );
and ( n14779 , n14774 , n14778 );
xor ( n14780 , n14691 , n14695 );
xor ( n14781 , n14780 , n14539 );
and ( n14782 , n14778 , n14781 );
and ( n14783 , n14774 , n14781 );
or ( n14784 , n14779 , n14782 , n14783 );
and ( n14785 , n11581 , n7847 );
and ( n14786 , n11413 , n7845 );
nor ( n14787 , n14785 , n14786 );
xnor ( n14788 , n14787 , n7857 );
and ( n14789 , n14784 , n14788 );
xor ( n14790 , n14699 , n14703 );
xor ( n14791 , n14790 , n14706 );
and ( n14792 , n14788 , n14791 );
and ( n14793 , n14784 , n14791 );
or ( n14794 , n14789 , n14792 , n14793 );
and ( n14795 , n10747 , n7797 );
and ( n14796 , n10499 , n7795 );
nor ( n14797 , n14795 , n14796 );
xnor ( n14798 , n14797 , n7807 );
and ( n14799 , n14794 , n14798 );
and ( n14800 , n11068 , n7826 );
and ( n14801 , n10842 , n7824 );
nor ( n14802 , n14800 , n14801 );
xnor ( n14803 , n14802 , n7836 );
and ( n14804 , n14798 , n14803 );
and ( n14805 , n14794 , n14803 );
or ( n14806 , n14799 , n14804 , n14805 );
and ( n14807 , n10499 , n7797 );
and ( n14808 , n10419 , n7795 );
nor ( n14809 , n14807 , n14808 );
xnor ( n14810 , n14809 , n7807 );
and ( n14811 , n14806 , n14810 );
xor ( n14812 , n14564 , n14568 );
xor ( n14813 , n14812 , n14590 );
and ( n14814 , n14810 , n14813 );
and ( n14815 , n14806 , n14813 );
or ( n14816 , n14811 , n14814 , n14815 );
and ( n14817 , n14766 , n14816 );
and ( n14818 , n9410 , n7683 );
and ( n14819 , n9162 , n7680 );
nor ( n14820 , n14818 , n14819 );
xnor ( n14821 , n14820 , n7676 );
and ( n14822 , n14816 , n14821 );
and ( n14823 , n14766 , n14821 );
or ( n14824 , n14817 , n14822 , n14823 );
xor ( n14825 , n14628 , n14632 );
xor ( n14826 , n14825 , n14635 );
and ( n14827 , n14824 , n14826 );
xor ( n14828 , n14738 , n14740 );
and ( n14829 , n14826 , n14828 );
and ( n14830 , n14824 , n14828 );
or ( n14831 , n14827 , n14829 , n14830 );
xor ( n14832 , n14678 , n14741 );
xor ( n14833 , n14832 , n14744 );
and ( n14834 , n14831 , n14833 );
xor ( n14835 , n14770 , n14773 );
and ( n14836 , n12254 , n7036 );
and ( n14837 , n12101 , n7034 );
nor ( n14838 , n14836 , n14837 );
xnor ( n14839 , n14838 , n7125 );
and ( n14840 , n14835 , n14839 );
and ( n14841 , n12907 , n6852 );
and ( n14842 , n12783 , n6850 );
nor ( n14843 , n14841 , n14842 );
xnor ( n14844 , n14843 , n6862 );
and ( n14845 , n14839 , n14844 );
and ( n14846 , n14835 , n14844 );
or ( n14847 , n14840 , n14845 , n14846 );
and ( n14848 , n11757 , n7847 );
and ( n14849 , n11581 , n7845 );
nor ( n14850 , n14848 , n14849 );
xnor ( n14851 , n14850 , n7857 );
and ( n14852 , n14847 , n14851 );
xor ( n14853 , n14774 , n14778 );
xor ( n14854 , n14853 , n14781 );
and ( n14855 , n14851 , n14854 );
and ( n14856 , n14847 , n14854 );
or ( n14857 , n14852 , n14855 , n14856 );
and ( n14858 , n10842 , n7797 );
and ( n14859 , n10747 , n7795 );
nor ( n14860 , n14858 , n14859 );
xnor ( n14861 , n14860 , n7807 );
and ( n14862 , n14857 , n14861 );
and ( n14863 , n11260 , n7826 );
and ( n14864 , n11068 , n7824 );
nor ( n14865 , n14863 , n14864 );
xnor ( n14866 , n14865 , n7836 );
and ( n14867 , n14861 , n14866 );
and ( n14868 , n14857 , n14866 );
or ( n14869 , n14862 , n14867 , n14868 );
and ( n14870 , n9676 , n7683 );
and ( n14871 , n9482 , n7680 );
nor ( n14872 , n14870 , n14871 );
xnor ( n14873 , n14872 , n7676 );
and ( n14874 , n14869 , n14873 );
xor ( n14875 , n14794 , n14798 );
xor ( n14876 , n14875 , n14803 );
and ( n14877 , n14873 , n14876 );
and ( n14878 , n14869 , n14876 );
or ( n14879 , n14874 , n14877 , n14878 );
xor ( n14880 , n14754 , n14758 );
xor ( n14881 , n14880 , n14763 );
and ( n14882 , n14879 , n14881 );
xor ( n14883 , n14806 , n14810 );
xor ( n14884 , n14883 , n14813 );
and ( n14885 , n14881 , n14884 );
and ( n14886 , n14879 , n14884 );
or ( n14887 , n14882 , n14885 , n14886 );
xor ( n14888 , n14766 , n14816 );
xor ( n14889 , n14888 , n14821 );
and ( n14890 , n14887 , n14889 );
xor ( n14891 , n14730 , n14732 );
xor ( n14892 , n14891 , n14735 );
and ( n14893 , n14889 , n14892 );
and ( n14894 , n14887 , n14892 );
or ( n14895 , n14890 , n14893 , n14894 );
xor ( n14896 , n14824 , n14826 );
xor ( n14897 , n14896 , n14828 );
and ( n14898 , n14895 , n14897 );
xor ( n14899 , n14887 , n14889 );
xor ( n14900 , n14899 , n14892 );
xor ( n14901 , n14718 , n14722 );
xor ( n14902 , n14901 , n14727 );
xor ( n14903 , n14879 , n14881 );
xor ( n14904 , n14903 , n14884 );
and ( n14905 , n14902 , n14904 );
xor ( n14906 , n14682 , n14686 );
xor ( n14907 , n14906 , n14715 );
and ( n14908 , n12359 , n7036 );
and ( n14909 , n12254 , n7034 );
nor ( n14910 , n14908 , n14909 );
xnor ( n14911 , n14910 , n7125 );
and ( n14912 , n12783 , n6722 );
and ( n14913 , n12522 , n6720 );
nor ( n14914 , n14912 , n14913 );
xnor ( n14915 , n14914 , n6821 );
and ( n14916 , n14911 , n14915 );
and ( n14917 , n14915 , n14771 );
and ( n14918 , n14911 , n14771 );
or ( n14919 , n14916 , n14917 , n14918 );
and ( n14920 , n11862 , n7847 );
and ( n14921 , n11757 , n7845 );
nor ( n14922 , n14920 , n14921 );
xnor ( n14923 , n14922 , n7857 );
and ( n14924 , n14919 , n14923 );
xor ( n14925 , n14835 , n14839 );
xor ( n14926 , n14925 , n14844 );
and ( n14927 , n14923 , n14926 );
and ( n14928 , n14919 , n14926 );
or ( n14929 , n14924 , n14927 , n14928 );
and ( n14930 , n11413 , n7826 );
and ( n14931 , n11260 , n7824 );
nor ( n14932 , n14930 , n14931 );
xnor ( n14933 , n14932 , n7836 );
and ( n14934 , n14929 , n14933 );
xor ( n14935 , n14847 , n14851 );
xor ( n14936 , n14935 , n14854 );
and ( n14937 , n14933 , n14936 );
and ( n14938 , n14929 , n14936 );
or ( n14939 , n14934 , n14937 , n14938 );
and ( n14940 , n10120 , n7732 );
and ( n14941 , n10055 , n7730 );
nor ( n14942 , n14940 , n14941 );
xnor ( n14943 , n14942 , n7742 );
and ( n14944 , n14939 , n14943 );
xor ( n14945 , n14784 , n14788 );
xor ( n14946 , n14945 , n14791 );
and ( n14947 , n14943 , n14946 );
and ( n14948 , n14939 , n14946 );
or ( n14949 , n14944 , n14947 , n14948 );
and ( n14950 , n14907 , n14949 );
and ( n14951 , n10499 , n7762 );
and ( n14952 , n10419 , n7760 );
nor ( n14953 , n14951 , n14952 );
xnor ( n14954 , n14953 , n7772 );
xor ( n14955 , n14857 , n14861 );
xor ( n14956 , n14955 , n14866 );
and ( n14957 , n14954 , n14956 );
and ( n14958 , n12522 , n7036 );
and ( n14959 , n12359 , n7034 );
nor ( n14960 , n14958 , n14959 );
xnor ( n14961 , n14960 , n7125 );
and ( n14962 , n12907 , n6720 );
not ( n14963 , n14962 );
and ( n14964 , n14963 , n6821 );
and ( n14965 , n14961 , n14964 );
and ( n14966 , n12101 , n7847 );
and ( n14967 , n11862 , n7845 );
nor ( n14968 , n14966 , n14967 );
xnor ( n14969 , n14968 , n7857 );
and ( n14970 , n14965 , n14969 );
xor ( n14971 , n14911 , n14915 );
xor ( n14972 , n14971 , n14771 );
and ( n14973 , n14969 , n14972 );
and ( n14974 , n14965 , n14972 );
or ( n14975 , n14970 , n14973 , n14974 );
and ( n14976 , n11581 , n7826 );
and ( n14977 , n11413 , n7824 );
nor ( n14978 , n14976 , n14977 );
xnor ( n14979 , n14978 , n7836 );
and ( n14980 , n14975 , n14979 );
xor ( n14981 , n14919 , n14923 );
xor ( n14982 , n14981 , n14926 );
and ( n14983 , n14979 , n14982 );
and ( n14984 , n14975 , n14982 );
or ( n14985 , n14980 , n14983 , n14984 );
and ( n14986 , n11068 , n7797 );
and ( n14987 , n10842 , n7795 );
nor ( n14988 , n14986 , n14987 );
xnor ( n14989 , n14988 , n7807 );
and ( n14990 , n14985 , n14989 );
and ( n14991 , n14956 , n14990 );
and ( n14992 , n14954 , n14990 );
or ( n14993 , n14957 , n14991 , n14992 );
and ( n14994 , n14949 , n14993 );
and ( n14995 , n14907 , n14993 );
or ( n14996 , n14950 , n14994 , n14995 );
and ( n14997 , n14904 , n14996 );
and ( n14998 , n14902 , n14996 );
or ( n14999 , n14905 , n14997 , n14998 );
and ( n15000 , n14900 , n14999 );
xor ( n15001 , n14961 , n14964 );
and ( n15002 , n12254 , n7847 );
and ( n15003 , n12101 , n7845 );
nor ( n15004 , n15002 , n15003 );
xnor ( n15005 , n15004 , n7857 );
and ( n15006 , n15001 , n15005 );
and ( n15007 , n12907 , n6722 );
and ( n15008 , n12783 , n6720 );
nor ( n15009 , n15007 , n15008 );
xnor ( n15010 , n15009 , n6821 );
and ( n15011 , n15005 , n15010 );
and ( n15012 , n15001 , n15010 );
or ( n15013 , n15006 , n15011 , n15012 );
and ( n15014 , n11413 , n7797 );
and ( n15015 , n11260 , n7795 );
nor ( n15016 , n15014 , n15015 );
xnor ( n15017 , n15016 , n7807 );
and ( n15018 , n15013 , n15017 );
and ( n15019 , n11757 , n7826 );
and ( n15020 , n11581 , n7824 );
nor ( n15021 , n15019 , n15020 );
xnor ( n15022 , n15021 , n7836 );
and ( n15023 , n15017 , n15022 );
and ( n15024 , n15013 , n15022 );
or ( n15025 , n15018 , n15023 , n15024 );
and ( n15026 , n11260 , n7797 );
and ( n15027 , n11068 , n7795 );
nor ( n15028 , n15026 , n15027 );
xnor ( n15029 , n15028 , n7807 );
and ( n15030 , n15025 , n15029 );
xor ( n15031 , n14975 , n14979 );
xor ( n15032 , n15031 , n14982 );
and ( n15033 , n15029 , n15032 );
and ( n15034 , n15025 , n15032 );
or ( n15035 , n15030 , n15033 , n15034 );
and ( n15036 , n10419 , n7732 );
and ( n15037 , n10120 , n7730 );
nor ( n15038 , n15036 , n15037 );
xnor ( n15039 , n15038 , n7742 );
and ( n15040 , n15035 , n15039 );
xor ( n15041 , n14929 , n14933 );
xor ( n15042 , n15041 , n14936 );
and ( n15043 , n15039 , n15042 );
and ( n15044 , n15035 , n15042 );
or ( n15045 , n15040 , n15043 , n15044 );
and ( n15046 , n9925 , n7683 );
and ( n15047 , n9676 , n7680 );
nor ( n15048 , n15046 , n15047 );
xnor ( n15049 , n15048 , n7676 );
and ( n15050 , n15045 , n15049 );
xor ( n15051 , n14939 , n14943 );
xor ( n15052 , n15051 , n14946 );
and ( n15053 , n15049 , n15052 );
and ( n15054 , n15045 , n15052 );
or ( n15055 , n15050 , n15053 , n15054 );
xor ( n15056 , n14869 , n14873 );
xor ( n15057 , n15056 , n14876 );
and ( n15058 , n15055 , n15057 );
xor ( n15059 , n14902 , n14904 );
xor ( n15060 , n15059 , n14996 );
and ( n15061 , n15058 , n15060 );
xor ( n15062 , n14907 , n14949 );
xor ( n15063 , n15062 , n14993 );
xor ( n15064 , n15055 , n15057 );
and ( n15065 , n15063 , n15064 );
and ( n15066 , n10055 , n7683 );
and ( n15067 , n9925 , n7680 );
nor ( n15068 , n15066 , n15067 );
xnor ( n15069 , n15068 , n7676 );
and ( n15070 , n10747 , n7762 );
and ( n15071 , n10499 , n7760 );
nor ( n15072 , n15070 , n15071 );
xnor ( n15073 , n15072 , n7772 );
and ( n15074 , n15069 , n15073 );
xor ( n15075 , n14985 , n14989 );
and ( n15076 , n15073 , n15075 );
and ( n15077 , n15069 , n15075 );
or ( n15078 , n15074 , n15076 , n15077 );
xor ( n15079 , n14954 , n14956 );
xor ( n15080 , n15079 , n14990 );
and ( n15081 , n15078 , n15080 );
xor ( n15082 , n15045 , n15049 );
xor ( n15083 , n15082 , n15052 );
and ( n15084 , n15080 , n15083 );
and ( n15085 , n15078 , n15083 );
or ( n15086 , n15081 , n15084 , n15085 );
and ( n15087 , n15064 , n15086 );
and ( n15088 , n15063 , n15086 );
or ( n15089 , n15065 , n15087 , n15088 );
and ( n15090 , n15060 , n15089 );
and ( n15091 , n15058 , n15089 );
or ( n15092 , n15061 , n15090 , n15091 );
and ( n15093 , n14999 , n15092 );
and ( n15094 , n14900 , n15092 );
or ( n15095 , n15000 , n15093 , n15094 );
and ( n15096 , n14897 , n15095 );
and ( n15097 , n14895 , n15095 );
or ( n15098 , n14898 , n15096 , n15097 );
and ( n15099 , n14833 , n15098 );
and ( n15100 , n14831 , n15098 );
or ( n15101 , n14834 , n15099 , n15100 );
and ( n15102 , n14749 , n15101 );
and ( n15103 , n14747 , n15101 );
or ( n15104 , n14750 , n15102 , n15103 );
and ( n15105 , n14676 , n15104 );
xor ( n15106 , n14676 , n15104 );
xor ( n15107 , n14747 , n14749 );
xor ( n15108 , n15107 , n15101 );
xor ( n15109 , n14831 , n14833 );
xor ( n15110 , n15109 , n15098 );
xor ( n15111 , n14895 , n14897 );
xor ( n15112 , n15111 , n15095 );
xor ( n15113 , n14900 , n14999 );
xor ( n15114 , n15113 , n15092 );
xor ( n15115 , n15058 , n15060 );
xor ( n15116 , n15115 , n15089 );
and ( n15117 , n12522 , n7847 );
and ( n15118 , n12359 , n7845 );
nor ( n15119 , n15117 , n15118 );
xnor ( n15120 , n15119 , n7857 );
and ( n15121 , n12907 , n7034 );
not ( n15122 , n15121 );
and ( n15123 , n15122 , n7125 );
and ( n15124 , n15120 , n15123 );
and ( n15125 , n12101 , n7826 );
and ( n15126 , n11862 , n7824 );
nor ( n15127 , n15125 , n15126 );
xnor ( n15128 , n15127 , n7836 );
and ( n15129 , n15124 , n15128 );
and ( n15130 , n12359 , n7847 );
and ( n15131 , n12254 , n7845 );
nor ( n15132 , n15130 , n15131 );
xnor ( n15133 , n15132 , n7857 );
and ( n15134 , n12783 , n7036 );
and ( n15135 , n12522 , n7034 );
nor ( n15136 , n15134 , n15135 );
xnor ( n15137 , n15136 , n7125 );
xor ( n15138 , n15133 , n15137 );
xor ( n15139 , n15138 , n14962 );
and ( n15140 , n15128 , n15139 );
and ( n15141 , n15124 , n15139 );
or ( n15142 , n15129 , n15140 , n15141 );
and ( n15143 , n11581 , n7797 );
and ( n15144 , n11413 , n7795 );
nor ( n15145 , n15143 , n15144 );
xnor ( n15146 , n15145 , n7807 );
and ( n15147 , n15142 , n15146 );
and ( n15148 , n15133 , n15137 );
and ( n15149 , n15137 , n14962 );
and ( n15150 , n15133 , n14962 );
or ( n15151 , n15148 , n15149 , n15150 );
and ( n15152 , n11862 , n7826 );
and ( n15153 , n11757 , n7824 );
nor ( n15154 , n15152 , n15153 );
xnor ( n15155 , n15154 , n7836 );
xor ( n15156 , n15151 , n15155 );
xor ( n15157 , n15001 , n15005 );
xor ( n15158 , n15157 , n15010 );
xor ( n15159 , n15156 , n15158 );
and ( n15160 , n15146 , n15159 );
and ( n15161 , n15142 , n15159 );
or ( n15162 , n15147 , n15160 , n15161 );
and ( n15163 , n10747 , n7732 );
and ( n15164 , n10499 , n7730 );
nor ( n15165 , n15163 , n15164 );
xnor ( n15166 , n15165 , n7742 );
and ( n15167 , n15162 , n15166 );
and ( n15168 , n11068 , n7762 );
and ( n15169 , n10842 , n7760 );
nor ( n15170 , n15168 , n15169 );
xnor ( n15171 , n15170 , n7772 );
and ( n15172 , n15166 , n15171 );
and ( n15173 , n15162 , n15171 );
or ( n15174 , n15167 , n15172 , n15173 );
and ( n15175 , n10120 , n7683 );
and ( n15176 , n10055 , n7680 );
nor ( n15177 , n15175 , n15176 );
xnor ( n15178 , n15177 , n7676 );
and ( n15179 , n15174 , n15178 );
and ( n15180 , n10499 , n7732 );
and ( n15181 , n10419 , n7730 );
nor ( n15182 , n15180 , n15181 );
xnor ( n15183 , n15182 , n7742 );
and ( n15184 , n15178 , n15183 );
and ( n15185 , n15174 , n15183 );
or ( n15186 , n15179 , n15184 , n15185 );
xor ( n15187 , n15035 , n15039 );
xor ( n15188 , n15187 , n15042 );
and ( n15189 , n15186 , n15188 );
and ( n15190 , n10842 , n7762 );
and ( n15191 , n10747 , n7760 );
nor ( n15192 , n15190 , n15191 );
xnor ( n15193 , n15192 , n7772 );
and ( n15194 , n15151 , n15155 );
and ( n15195 , n15155 , n15158 );
and ( n15196 , n15151 , n15158 );
or ( n15197 , n15194 , n15195 , n15196 );
xor ( n15198 , n15013 , n15017 );
xor ( n15199 , n15198 , n15022 );
and ( n15200 , n15197 , n15199 );
xor ( n15201 , n14965 , n14969 );
xor ( n15202 , n15201 , n14972 );
and ( n15203 , n15199 , n15202 );
and ( n15204 , n15197 , n15202 );
or ( n15205 , n15200 , n15203 , n15204 );
and ( n15206 , n15193 , n15205 );
xor ( n15207 , n15025 , n15029 );
xor ( n15208 , n15207 , n15032 );
and ( n15209 , n15205 , n15208 );
and ( n15210 , n15193 , n15208 );
or ( n15211 , n15206 , n15209 , n15210 );
xor ( n15212 , n15069 , n15073 );
xor ( n15213 , n15212 , n15075 );
and ( n15214 , n15211 , n15213 );
xor ( n15215 , n15186 , n15188 );
and ( n15216 , n15213 , n15215 );
and ( n15217 , n15211 , n15215 );
or ( n15218 , n15214 , n15216 , n15217 );
and ( n15219 , n15189 , n15218 );
xor ( n15220 , n15078 , n15080 );
xor ( n15221 , n15220 , n15083 );
and ( n15222 , n15218 , n15221 );
and ( n15223 , n15189 , n15221 );
or ( n15224 , n15219 , n15222 , n15223 );
xor ( n15225 , n15063 , n15064 );
xor ( n15226 , n15225 , n15086 );
and ( n15227 , n15224 , n15226 );
xor ( n15228 , n15224 , n15226 );
xor ( n15229 , n15189 , n15218 );
xor ( n15230 , n15229 , n15221 );
xor ( n15231 , n15174 , n15178 );
xor ( n15232 , n15231 , n15183 );
xor ( n15233 , n15120 , n15123 );
and ( n15234 , n12254 , n7826 );
and ( n15235 , n12101 , n7824 );
nor ( n15236 , n15234 , n15235 );
xnor ( n15237 , n15236 , n7836 );
and ( n15238 , n15233 , n15237 );
and ( n15239 , n12907 , n7036 );
and ( n15240 , n12783 , n7034 );
nor ( n15241 , n15239 , n15240 );
xnor ( n15242 , n15241 , n7125 );
and ( n15243 , n15237 , n15242 );
and ( n15244 , n15233 , n15242 );
or ( n15245 , n15238 , n15243 , n15244 );
and ( n15246 , n11757 , n7797 );
and ( n15247 , n11581 , n7795 );
nor ( n15248 , n15246 , n15247 );
xnor ( n15249 , n15248 , n7807 );
and ( n15250 , n15245 , n15249 );
xor ( n15251 , n15124 , n15128 );
xor ( n15252 , n15251 , n15139 );
and ( n15253 , n15249 , n15252 );
and ( n15254 , n15245 , n15252 );
or ( n15255 , n15250 , n15253 , n15254 );
and ( n15256 , n11260 , n7762 );
and ( n15257 , n11068 , n7760 );
nor ( n15258 , n15256 , n15257 );
xnor ( n15259 , n15258 , n7772 );
and ( n15260 , n15255 , n15259 );
xor ( n15261 , n15142 , n15146 );
xor ( n15262 , n15261 , n15159 );
and ( n15263 , n15259 , n15262 );
and ( n15264 , n15255 , n15262 );
or ( n15265 , n15260 , n15263 , n15264 );
and ( n15266 , n10419 , n7683 );
and ( n15267 , n10120 , n7680 );
nor ( n15268 , n15266 , n15267 );
xnor ( n15269 , n15268 , n7676 );
and ( n15270 , n15265 , n15269 );
xor ( n15271 , n15197 , n15199 );
xor ( n15272 , n15271 , n15202 );
and ( n15273 , n15269 , n15272 );
and ( n15274 , n15265 , n15272 );
or ( n15275 , n15270 , n15273 , n15274 );
and ( n15276 , n15232 , n15275 );
xor ( n15277 , n15193 , n15205 );
xor ( n15278 , n15277 , n15208 );
and ( n15279 , n15275 , n15278 );
and ( n15280 , n15232 , n15278 );
or ( n15281 , n15276 , n15279 , n15280 );
xor ( n15282 , n15211 , n15213 );
xor ( n15283 , n15282 , n15215 );
and ( n15284 , n15281 , n15283 );
xor ( n15285 , n15281 , n15283 );
and ( n15286 , n12359 , n7826 );
and ( n15287 , n12254 , n7824 );
nor ( n15288 , n15286 , n15287 );
xnor ( n15289 , n15288 , n7836 );
and ( n15290 , n12783 , n7847 );
and ( n15291 , n12522 , n7845 );
nor ( n15292 , n15290 , n15291 );
xnor ( n15293 , n15292 , n7857 );
and ( n15294 , n15289 , n15293 );
and ( n15295 , n15293 , n15121 );
and ( n15296 , n15289 , n15121 );
or ( n15297 , n15294 , n15295 , n15296 );
and ( n15298 , n11862 , n7797 );
and ( n15299 , n11757 , n7795 );
nor ( n15300 , n15298 , n15299 );
xnor ( n15301 , n15300 , n7807 );
and ( n15302 , n15297 , n15301 );
xor ( n15303 , n15233 , n15237 );
xor ( n15304 , n15303 , n15242 );
and ( n15305 , n15301 , n15304 );
and ( n15306 , n15297 , n15304 );
or ( n15307 , n15302 , n15305 , n15306 );
and ( n15308 , n11413 , n7762 );
and ( n15309 , n11260 , n7760 );
nor ( n15310 , n15308 , n15309 );
xnor ( n15311 , n15310 , n7772 );
and ( n15312 , n15307 , n15311 );
xor ( n15313 , n15245 , n15249 );
xor ( n15314 , n15313 , n15252 );
and ( n15315 , n15311 , n15314 );
and ( n15316 , n15307 , n15314 );
or ( n15317 , n15312 , n15315 , n15316 );
and ( n15318 , n10499 , n7683 );
and ( n15319 , n10419 , n7680 );
nor ( n15320 , n15318 , n15319 );
xnor ( n15321 , n15320 , n7676 );
and ( n15322 , n15317 , n15321 );
and ( n15323 , n10842 , n7732 );
and ( n15324 , n10747 , n7730 );
nor ( n15325 , n15323 , n15324 );
xnor ( n15326 , n15325 , n7742 );
and ( n15327 , n15321 , n15326 );
and ( n15328 , n15317 , n15326 );
or ( n15329 , n15322 , n15327 , n15328 );
xor ( n15330 , n15162 , n15166 );
xor ( n15331 , n15330 , n15171 );
and ( n15332 , n15329 , n15331 );
xor ( n15333 , n15265 , n15269 );
xor ( n15334 , n15333 , n15272 );
and ( n15335 , n15331 , n15334 );
and ( n15336 , n15329 , n15334 );
or ( n15337 , n15332 , n15335 , n15336 );
xor ( n15338 , n15232 , n15275 );
xor ( n15339 , n15338 , n15278 );
and ( n15340 , n15337 , n15339 );
xor ( n15341 , n15337 , n15339 );
and ( n15342 , n12522 , n7826 );
and ( n15343 , n12359 , n7824 );
nor ( n15344 , n15342 , n15343 );
xnor ( n15345 , n15344 , n7836 );
and ( n15346 , n12907 , n7845 );
not ( n15347 , n15346 );
and ( n15348 , n15347 , n7857 );
and ( n15349 , n15345 , n15348 );
and ( n15350 , n12101 , n7797 );
and ( n15351 , n11862 , n7795 );
nor ( n15352 , n15350 , n15351 );
xnor ( n15353 , n15352 , n7807 );
and ( n15354 , n15349 , n15353 );
xor ( n15355 , n15289 , n15293 );
xor ( n15356 , n15355 , n15121 );
and ( n15357 , n15353 , n15356 );
and ( n15358 , n15349 , n15356 );
or ( n15359 , n15354 , n15357 , n15358 );
and ( n15360 , n11581 , n7762 );
and ( n15361 , n11413 , n7760 );
nor ( n15362 , n15360 , n15361 );
xnor ( n15363 , n15362 , n7772 );
and ( n15364 , n15359 , n15363 );
xor ( n15365 , n15297 , n15301 );
xor ( n15366 , n15365 , n15304 );
and ( n15367 , n15363 , n15366 );
and ( n15368 , n15359 , n15366 );
or ( n15369 , n15364 , n15367 , n15368 );
and ( n15370 , n10747 , n7683 );
and ( n15371 , n10499 , n7680 );
nor ( n15372 , n15370 , n15371 );
xnor ( n15373 , n15372 , n7676 );
and ( n15374 , n15369 , n15373 );
and ( n15375 , n11068 , n7732 );
and ( n15376 , n10842 , n7730 );
nor ( n15377 , n15375 , n15376 );
xnor ( n15378 , n15377 , n7742 );
and ( n15379 , n15373 , n15378 );
and ( n15380 , n15369 , n15378 );
or ( n15381 , n15374 , n15379 , n15380 );
xor ( n15382 , n15317 , n15321 );
xor ( n15383 , n15382 , n15326 );
and ( n15384 , n15381 , n15383 );
xor ( n15385 , n15255 , n15259 );
xor ( n15386 , n15385 , n15262 );
and ( n15387 , n15383 , n15386 );
and ( n15388 , n15381 , n15386 );
or ( n15389 , n15384 , n15387 , n15388 );
xor ( n15390 , n15329 , n15331 );
xor ( n15391 , n15390 , n15334 );
and ( n15392 , n15389 , n15391 );
xor ( n15393 , n15389 , n15391 );
xor ( n15394 , n15381 , n15383 );
xor ( n15395 , n15394 , n15386 );
xor ( n15396 , n15345 , n15348 );
and ( n15397 , n12254 , n7797 );
and ( n15398 , n12101 , n7795 );
nor ( n15399 , n15397 , n15398 );
xnor ( n15400 , n15399 , n7807 );
and ( n15401 , n15396 , n15400 );
and ( n15402 , n12907 , n7847 );
and ( n15403 , n12783 , n7845 );
nor ( n15404 , n15402 , n15403 );
xnor ( n15405 , n15404 , n7857 );
and ( n15406 , n15400 , n15405 );
and ( n15407 , n15396 , n15405 );
or ( n15408 , n15401 , n15406 , n15407 );
and ( n15409 , n11757 , n7762 );
and ( n15410 , n11581 , n7760 );
nor ( n15411 , n15409 , n15410 );
xnor ( n15412 , n15411 , n7772 );
and ( n15413 , n15408 , n15412 );
xor ( n15414 , n15349 , n15353 );
xor ( n15415 , n15414 , n15356 );
and ( n15416 , n15412 , n15415 );
and ( n15417 , n15408 , n15415 );
or ( n15418 , n15413 , n15416 , n15417 );
and ( n15419 , n11260 , n7732 );
and ( n15420 , n11068 , n7730 );
nor ( n15421 , n15419 , n15420 );
xnor ( n15422 , n15421 , n7742 );
and ( n15423 , n15418 , n15422 );
xor ( n15424 , n15359 , n15363 );
xor ( n15425 , n15424 , n15366 );
and ( n15426 , n15422 , n15425 );
and ( n15427 , n15418 , n15425 );
or ( n15428 , n15423 , n15426 , n15427 );
xor ( n15429 , n15369 , n15373 );
xor ( n15430 , n15429 , n15378 );
and ( n15431 , n15428 , n15430 );
xor ( n15432 , n15307 , n15311 );
xor ( n15433 , n15432 , n15314 );
and ( n15434 , n15430 , n15433 );
and ( n15435 , n15428 , n15433 );
or ( n15436 , n15431 , n15434 , n15435 );
and ( n15437 , n15395 , n15436 );
xor ( n15438 , n15395 , n15436 );
xor ( n15439 , n15428 , n15430 );
xor ( n15440 , n15439 , n15433 );
and ( n15441 , n12359 , n7797 );
and ( n15442 , n12254 , n7795 );
nor ( n15443 , n15441 , n15442 );
xnor ( n15444 , n15443 , n7807 );
and ( n15445 , n12783 , n7826 );
and ( n15446 , n12522 , n7824 );
nor ( n15447 , n15445 , n15446 );
xnor ( n15448 , n15447 , n7836 );
and ( n15449 , n15444 , n15448 );
and ( n15450 , n15448 , n15346 );
and ( n15451 , n15444 , n15346 );
or ( n15452 , n15449 , n15450 , n15451 );
and ( n15453 , n11862 , n7762 );
and ( n15454 , n11757 , n7760 );
nor ( n15455 , n15453 , n15454 );
xnor ( n15456 , n15455 , n7772 );
and ( n15457 , n15452 , n15456 );
xor ( n15458 , n15396 , n15400 );
xor ( n15459 , n15458 , n15405 );
and ( n15460 , n15456 , n15459 );
and ( n15461 , n15452 , n15459 );
or ( n15462 , n15457 , n15460 , n15461 );
and ( n15463 , n11413 , n7732 );
and ( n15464 , n11260 , n7730 );
nor ( n15465 , n15463 , n15464 );
xnor ( n15466 , n15465 , n7742 );
and ( n15467 , n15462 , n15466 );
xor ( n15468 , n15408 , n15412 );
xor ( n15469 , n15468 , n15415 );
and ( n15470 , n15466 , n15469 );
and ( n15471 , n15462 , n15469 );
or ( n15472 , n15467 , n15470 , n15471 );
and ( n15473 , n10842 , n7683 );
and ( n15474 , n10747 , n7680 );
nor ( n15475 , n15473 , n15474 );
xnor ( n15476 , n15475 , n7676 );
and ( n15477 , n15472 , n15476 );
xor ( n15478 , n15418 , n15422 );
xor ( n15479 , n15478 , n15425 );
and ( n15480 , n15476 , n15479 );
and ( n15481 , n15472 , n15479 );
or ( n15482 , n15477 , n15480 , n15481 );
and ( n15483 , n15440 , n15482 );
xor ( n15484 , n15440 , n15482 );
and ( n15485 , n12522 , n7797 );
and ( n15486 , n12359 , n7795 );
nor ( n15487 , n15485 , n15486 );
xnor ( n15488 , n15487 , n7807 );
and ( n15489 , n12907 , n7824 );
not ( n15490 , n15489 );
and ( n15491 , n15490 , n7836 );
and ( n15492 , n15488 , n15491 );
and ( n15493 , n12101 , n7762 );
and ( n15494 , n11862 , n7760 );
nor ( n15495 , n15493 , n15494 );
xnor ( n15496 , n15495 , n7772 );
and ( n15497 , n15492 , n15496 );
xor ( n15498 , n15444 , n15448 );
xor ( n15499 , n15498 , n15346 );
and ( n15500 , n15496 , n15499 );
and ( n15501 , n15492 , n15499 );
or ( n15502 , n15497 , n15500 , n15501 );
and ( n15503 , n11581 , n7732 );
and ( n15504 , n11413 , n7730 );
nor ( n15505 , n15503 , n15504 );
xnor ( n15506 , n15505 , n7742 );
and ( n15507 , n15502 , n15506 );
xor ( n15508 , n15452 , n15456 );
xor ( n15509 , n15508 , n15459 );
and ( n15510 , n15506 , n15509 );
and ( n15511 , n15502 , n15509 );
or ( n15512 , n15507 , n15510 , n15511 );
and ( n15513 , n11068 , n7683 );
and ( n15514 , n10842 , n7680 );
nor ( n15515 , n15513 , n15514 );
xnor ( n15516 , n15515 , n7676 );
and ( n15517 , n15512 , n15516 );
xor ( n15518 , n15462 , n15466 );
xor ( n15519 , n15518 , n15469 );
and ( n15520 , n15516 , n15519 );
and ( n15521 , n15512 , n15519 );
or ( n15522 , n15517 , n15520 , n15521 );
xor ( n15523 , n15472 , n15476 );
xor ( n15524 , n15523 , n15479 );
and ( n15525 , n15522 , n15524 );
xor ( n15526 , n15522 , n15524 );
xor ( n15527 , n15512 , n15516 );
xor ( n15528 , n15527 , n15519 );
xor ( n15529 , n15488 , n15491 );
and ( n15530 , n12254 , n7762 );
and ( n15531 , n12101 , n7760 );
nor ( n15532 , n15530 , n15531 );
xnor ( n15533 , n15532 , n7772 );
and ( n15534 , n15529 , n15533 );
and ( n15535 , n12907 , n7826 );
and ( n15536 , n12783 , n7824 );
nor ( n15537 , n15535 , n15536 );
xnor ( n15538 , n15537 , n7836 );
and ( n15539 , n15533 , n15538 );
and ( n15540 , n15529 , n15538 );
or ( n15541 , n15534 , n15539 , n15540 );
and ( n15542 , n11757 , n7732 );
and ( n15543 , n11581 , n7730 );
nor ( n15544 , n15542 , n15543 );
xnor ( n15545 , n15544 , n7742 );
and ( n15546 , n15541 , n15545 );
xor ( n15547 , n15492 , n15496 );
xor ( n15548 , n15547 , n15499 );
and ( n15549 , n15545 , n15548 );
and ( n15550 , n15541 , n15548 );
or ( n15551 , n15546 , n15549 , n15550 );
and ( n15552 , n11260 , n7683 );
and ( n15553 , n11068 , n7680 );
nor ( n15554 , n15552 , n15553 );
xnor ( n15555 , n15554 , n7676 );
and ( n15556 , n15551 , n15555 );
xor ( n15557 , n15502 , n15506 );
xor ( n15558 , n15557 , n15509 );
and ( n15559 , n15555 , n15558 );
and ( n15560 , n15551 , n15558 );
or ( n15561 , n15556 , n15559 , n15560 );
and ( n15562 , n15528 , n15561 );
xor ( n15563 , n15528 , n15561 );
and ( n15564 , n12359 , n7762 );
and ( n15565 , n12254 , n7760 );
nor ( n15566 , n15564 , n15565 );
xnor ( n15567 , n15566 , n7772 );
and ( n15568 , n12783 , n7797 );
and ( n15569 , n12522 , n7795 );
nor ( n15570 , n15568 , n15569 );
xnor ( n15571 , n15570 , n7807 );
and ( n15572 , n15567 , n15571 );
and ( n15573 , n15571 , n15489 );
and ( n15574 , n15567 , n15489 );
or ( n15575 , n15572 , n15573 , n15574 );
and ( n15576 , n11862 , n7732 );
and ( n15577 , n11757 , n7730 );
nor ( n15578 , n15576 , n15577 );
xnor ( n15579 , n15578 , n7742 );
and ( n15580 , n15575 , n15579 );
xor ( n15581 , n15529 , n15533 );
xor ( n15582 , n15581 , n15538 );
and ( n15583 , n15579 , n15582 );
and ( n15584 , n15575 , n15582 );
or ( n15585 , n15580 , n15583 , n15584 );
and ( n15586 , n11413 , n7683 );
and ( n15587 , n11260 , n7680 );
nor ( n15588 , n15586 , n15587 );
xnor ( n15589 , n15588 , n7676 );
and ( n15590 , n15585 , n15589 );
xor ( n15591 , n15541 , n15545 );
xor ( n15592 , n15591 , n15548 );
and ( n15593 , n15589 , n15592 );
and ( n15594 , n15585 , n15592 );
or ( n15595 , n15590 , n15593 , n15594 );
xor ( n15596 , n15551 , n15555 );
xor ( n15597 , n15596 , n15558 );
and ( n15598 , n15595 , n15597 );
xor ( n15599 , n15595 , n15597 );
xor ( n15600 , n15585 , n15589 );
xor ( n15601 , n15600 , n15592 );
and ( n15602 , n12522 , n7762 );
and ( n15603 , n12359 , n7760 );
nor ( n15604 , n15602 , n15603 );
xnor ( n15605 , n15604 , n7772 );
and ( n15606 , n12907 , n7795 );
not ( n15607 , n15606 );
and ( n15608 , n15607 , n7807 );
and ( n15609 , n15605 , n15608 );
and ( n15610 , n12101 , n7732 );
and ( n15611 , n11862 , n7730 );
nor ( n15612 , n15610 , n15611 );
xnor ( n15613 , n15612 , n7742 );
and ( n15614 , n15609 , n15613 );
xor ( n15615 , n15567 , n15571 );
xor ( n15616 , n15615 , n15489 );
and ( n15617 , n15613 , n15616 );
and ( n15618 , n15609 , n15616 );
or ( n15619 , n15614 , n15617 , n15618 );
and ( n15620 , n11581 , n7683 );
and ( n15621 , n11413 , n7680 );
nor ( n15622 , n15620 , n15621 );
xnor ( n15623 , n15622 , n7676 );
and ( n15624 , n15619 , n15623 );
xor ( n15625 , n15575 , n15579 );
xor ( n15626 , n15625 , n15582 );
and ( n15627 , n15623 , n15626 );
and ( n15628 , n15619 , n15626 );
or ( n15629 , n15624 , n15627 , n15628 );
and ( n15630 , n15601 , n15629 );
xor ( n15631 , n15601 , n15629 );
xor ( n15632 , n15605 , n15608 );
and ( n15633 , n12254 , n7732 );
and ( n15634 , n12101 , n7730 );
nor ( n15635 , n15633 , n15634 );
xnor ( n15636 , n15635 , n7742 );
and ( n15637 , n15632 , n15636 );
and ( n15638 , n12907 , n7797 );
and ( n15639 , n12783 , n7795 );
nor ( n15640 , n15638 , n15639 );
xnor ( n15641 , n15640 , n7807 );
and ( n15642 , n15636 , n15641 );
and ( n15643 , n15632 , n15641 );
or ( n15644 , n15637 , n15642 , n15643 );
and ( n15645 , n11757 , n7683 );
and ( n15646 , n11581 , n7680 );
nor ( n15647 , n15645 , n15646 );
xnor ( n15648 , n15647 , n7676 );
and ( n15649 , n15644 , n15648 );
xor ( n15650 , n15609 , n15613 );
xor ( n15651 , n15650 , n15616 );
and ( n15652 , n15648 , n15651 );
and ( n15653 , n15644 , n15651 );
or ( n15654 , n15649 , n15652 , n15653 );
xor ( n15655 , n15619 , n15623 );
xor ( n15656 , n15655 , n15626 );
and ( n15657 , n15654 , n15656 );
xor ( n15658 , n15654 , n15656 );
xor ( n15659 , n15644 , n15648 );
xor ( n15660 , n15659 , n15651 );
and ( n15661 , n12907 , n7760 );
not ( n15662 , n15661 );
and ( n15663 , n15662 , n7772 );
and ( n15664 , n12907 , n7762 );
and ( n15665 , n12783 , n7760 );
nor ( n15666 , n15664 , n15665 );
xnor ( n15667 , n15666 , n7772 );
and ( n15668 , n15663 , n15667 );
and ( n15669 , n12783 , n7762 );
and ( n15670 , n12522 , n7760 );
nor ( n15671 , n15669 , n15670 );
xnor ( n15672 , n15671 , n7772 );
and ( n15673 , n15668 , n15672 );
and ( n15674 , n15672 , n15606 );
and ( n15675 , n15668 , n15606 );
or ( n15676 , n15673 , n15674 , n15675 );
and ( n15677 , n11862 , n7683 );
and ( n15678 , n11757 , n7680 );
nor ( n15679 , n15677 , n15678 );
xnor ( n15680 , n15679 , n7676 );
and ( n15681 , n15676 , n15680 );
xor ( n15682 , n15632 , n15636 );
xor ( n15683 , n15682 , n15641 );
and ( n15684 , n15680 , n15683 );
and ( n15685 , n15676 , n15683 );
or ( n15686 , n15681 , n15684 , n15685 );
and ( n15687 , n15660 , n15686 );
xor ( n15688 , n15660 , n15686 );
xor ( n15689 , n15676 , n15680 );
xor ( n15690 , n15689 , n15683 );
and ( n15691 , n12101 , n7683 );
and ( n15692 , n11862 , n7680 );
nor ( n15693 , n15691 , n15692 );
xnor ( n15694 , n15693 , n7676 );
and ( n15695 , n12359 , n7732 );
and ( n15696 , n12254 , n7730 );
nor ( n15697 , n15695 , n15696 );
xnor ( n15698 , n15697 , n7742 );
and ( n15699 , n15694 , n15698 );
xor ( n15700 , n15668 , n15672 );
xor ( n15701 , n15700 , n15606 );
and ( n15702 , n15698 , n15701 );
and ( n15703 , n15694 , n15701 );
or ( n15704 , n15699 , n15702 , n15703 );
and ( n15705 , n15690 , n15704 );
xor ( n15706 , n15690 , n15704 );
xor ( n15707 , n15694 , n15698 );
xor ( n15708 , n15707 , n15701 );
xor ( n15709 , n15663 , n15667 );
and ( n15710 , n12907 , n7730 );
not ( n15711 , n15710 );
and ( n15712 , n15711 , n7742 );
and ( n15713 , n12907 , n7732 );
and ( n15714 , n12783 , n7730 );
nor ( n15715 , n15713 , n15714 );
xnor ( n15716 , n15715 , n7742 );
and ( n15717 , n15712 , n15716 );
and ( n15718 , n12783 , n7732 );
and ( n15719 , n12522 , n7730 );
nor ( n15720 , n15718 , n15719 );
xnor ( n15721 , n15720 , n7742 );
and ( n15722 , n15717 , n15721 );
and ( n15723 , n15721 , n15661 );
and ( n15724 , n15717 , n15661 );
or ( n15725 , n15722 , n15723 , n15724 );
and ( n15726 , n15709 , n15725 );
and ( n15727 , n12522 , n7732 );
and ( n15728 , n12359 , n7730 );
nor ( n15729 , n15727 , n15728 );
xnor ( n15730 , n15729 , n7742 );
and ( n15731 , n15725 , n15730 );
and ( n15732 , n15709 , n15730 );
or ( n15733 , n15726 , n15731 , n15732 );
and ( n15734 , n15708 , n15733 );
xor ( n15735 , n15708 , n15733 );
and ( n15736 , n12254 , n7683 );
and ( n15737 , n12101 , n7680 );
nor ( n15738 , n15736 , n15737 );
xnor ( n15739 , n15738 , n7676 );
xor ( n15740 , n15709 , n15725 );
xor ( n15741 , n15740 , n15730 );
and ( n15742 , n15739 , n15741 );
xor ( n15743 , n15739 , n15741 );
and ( n15744 , n12359 , n7683 );
and ( n15745 , n12254 , n7680 );
nor ( n15746 , n15744 , n15745 );
xnor ( n15747 , n15746 , n7676 );
xor ( n15748 , n15717 , n15721 );
xor ( n15749 , n15748 , n15661 );
and ( n15750 , n15747 , n15749 );
xor ( n15751 , n15747 , n15749 );
and ( n15752 , n12522 , n7683 );
and ( n15753 , n12359 , n7680 );
nor ( n15754 , n15752 , n15753 );
xnor ( n15755 , n15754 , n7676 );
xor ( n15756 , n15712 , n15716 );
and ( n15757 , n15755 , n15756 );
xor ( n15758 , n15755 , n15756 );
and ( n15759 , n12783 , n7683 );
and ( n15760 , n12522 , n7680 );
nor ( n15761 , n15759 , n15760 );
xnor ( n15762 , n15761 , n7676 );
and ( n15763 , n15762 , n15710 );
xor ( n15764 , n15762 , n15710 );
and ( n15765 , n12907 , n7683 );
and ( n15766 , n12783 , n7680 );
nor ( n15767 , n15765 , n15766 );
xnor ( n15768 , n15767 , n7676 );
and ( n15769 , n12907 , n7680 );
not ( n15770 , n15769 );
and ( n15771 , n15770 , n7676 );
and ( n15772 , n15768 , n15771 );
and ( n15773 , n15764 , n15772 );
or ( n15774 , n15763 , n15773 );
and ( n15775 , n15758 , n15774 );
or ( n15776 , n15757 , n15775 );
and ( n15777 , n15751 , n15776 );
or ( n15778 , n15750 , n15777 );
and ( n15779 , n15743 , n15778 );
or ( n15780 , n15742 , n15779 );
and ( n15781 , n15735 , n15780 );
or ( n15782 , n15734 , n15781 );
and ( n15783 , n15706 , n15782 );
or ( n15784 , n15705 , n15783 );
and ( n15785 , n15688 , n15784 );
or ( n15786 , n15687 , n15785 );
and ( n15787 , n15658 , n15786 );
or ( n15788 , n15657 , n15787 );
and ( n15789 , n15631 , n15788 );
or ( n15790 , n15630 , n15789 );
and ( n15791 , n15599 , n15790 );
or ( n15792 , n15598 , n15791 );
and ( n15793 , n15563 , n15792 );
or ( n15794 , n15562 , n15793 );
and ( n15795 , n15526 , n15794 );
or ( n15796 , n15525 , n15795 );
and ( n15797 , n15484 , n15796 );
or ( n15798 , n15483 , n15797 );
and ( n15799 , n15438 , n15798 );
or ( n15800 , n15437 , n15799 );
and ( n15801 , n15393 , n15800 );
or ( n15802 , n15392 , n15801 );
and ( n15803 , n15341 , n15802 );
or ( n15804 , n15340 , n15803 );
and ( n15805 , n15285 , n15804 );
or ( n15806 , n15284 , n15805 );
and ( n15807 , n15230 , n15806 );
and ( n15808 , n15228 , n15807 );
or ( n15809 , n15227 , n15808 );
and ( n15810 , n15116 , n15809 );
and ( n15811 , n15114 , n15810 );
and ( n15812 , n15112 , n15811 );
and ( n15813 , n15110 , n15812 );
and ( n15814 , n15108 , n15813 );
and ( n15815 , n15106 , n15814 );
or ( n15816 , n15105 , n15815 );
and ( n15817 , n14674 , n15816 );
and ( n15818 , n14672 , n15817 );
and ( n15819 , n14670 , n15818 );
and ( n15820 , n14668 , n15819 );
and ( n15821 , n14666 , n15820 );
and ( n15822 , n14664 , n15821 );
or ( n15823 , n14663 , n15822 );
and ( n15824 , n14007 , n15823 );
or ( n15825 , n14006 , n15824 );
and ( n15826 , n13780 , n15825 );
and ( n15827 , n13778 , n15826 );
and ( n15828 , n13776 , n15827 );
or ( n15829 , n13775 , n15828 );
and ( n15830 , n13335 , n15829 );
or ( n15831 , n13334 , n15830 );
and ( n15832 , n13077 , n15831 );
or ( n15833 , n13076 , n15832 );
and ( n15834 , n12983 , n15833 );
or ( n15835 , n12982 , n15834 );
and ( n15836 , n12749 , n15835 );
and ( n15837 , n12747 , n15836 );
or ( n15838 , n12746 , n15837 );
and ( n15839 , n12596 , n15838 );
or ( n15840 , n12595 , n15839 );
and ( n15841 , n12421 , n15840 );
or ( n15842 , n12420 , n15841 );
and ( n15843 , n12076 , n15842 );
and ( n15844 , n12074 , n15843 );
and ( n15845 , n12072 , n15844 );
or ( n15846 , n12071 , n15845 );
and ( n15847 , n11744 , n15846 );
or ( n15848 , n11743 , n15847 );
and ( n15849 , n11564 , n15848 );
or ( n15850 , n11563 , n15849 );
and ( n15851 , n11375 , n15850 );
or ( n15852 , n11374 , n15851 );
and ( n15853 , n11202 , n15852 );
and ( n15854 , n11200 , n15853 );
or ( n15855 , n11199 , n15854 );
and ( n15856 , n10887 , n15855 );
or ( n15857 , n10886 , n15856 );
and ( n15858 , n10724 , n15857 );
or ( n15859 , n10723 , n15858 );
and ( n15860 , n10540 , n15859 );
or ( n15861 , n10539 , n15860 );
and ( n15862 , n10317 , n15861 );
and ( n15863 , n10315 , n15862 );
and ( n15864 , n10313 , n15863 );
and ( n15865 , n10311 , n15864 );
or ( n15866 , n10310 , n15865 );
and ( n15867 , n9732 , n15866 );
or ( n15868 , n9731 , n15867 );
and ( n15869 , n9549 , n15868 );
and ( n15870 , n9547 , n15869 );
or ( n15871 , n9546 , n15870 );
and ( n15872 , n9207 , n15871 );
xor ( n15873 , n9205 , n15872 );
buf ( n543134 , n15873 );
buf ( n543135 , n543134 );
xor ( n15876 , n9207 , n15871 );
buf ( n543137 , n15876 );
buf ( n543138 , n543137 );
xor ( n15879 , n9547 , n15869 );
buf ( n543140 , n15879 );
buf ( n543141 , n543140 );
xor ( n15882 , n9549 , n15868 );
buf ( n543143 , n15882 );
buf ( n543144 , n543143 );
xor ( n15885 , n9732 , n15866 );
buf ( n543146 , n15885 );
buf ( n543147 , n543146 );
xor ( n15888 , n10311 , n15864 );
buf ( n543149 , n15888 );
buf ( n543150 , n543149 );
xor ( n15891 , n10313 , n15863 );
buf ( n543152 , n15891 );
buf ( n543153 , n543152 );
xor ( n15894 , n10315 , n15862 );
buf ( n543155 , n15894 );
buf ( n543156 , n543155 );
xor ( n15897 , n10317 , n15861 );
buf ( n543158 , n15897 );
buf ( n543159 , n543158 );
xor ( n15900 , n10540 , n15859 );
buf ( n543161 , n15900 );
buf ( n543162 , n543161 );
xor ( n15903 , n10724 , n15857 );
buf ( n543164 , n15903 );
buf ( n543165 , n543164 );
xor ( n15906 , n10887 , n15855 );
buf ( n543167 , n15906 );
buf ( n543168 , n543167 );
xor ( n15909 , n11200 , n15853 );
buf ( n543170 , n15909 );
buf ( n543171 , n543170 );
xor ( n15912 , n11202 , n15852 );
buf ( n543173 , n15912 );
buf ( n543174 , n543173 );
xor ( n15915 , n11375 , n15850 );
buf ( n543176 , n15915 );
buf ( n543177 , n543176 );
xor ( n15918 , n11564 , n15848 );
buf ( n543179 , n15918 );
buf ( n543180 , n543179 );
xor ( n15921 , n11744 , n15846 );
buf ( n543182 , n15921 );
buf ( n543183 , n543182 );
xor ( n15924 , n12072 , n15844 );
buf ( n543185 , n15924 );
buf ( n543186 , n543185 );
xor ( n15927 , n12074 , n15843 );
buf ( n543188 , n15927 );
buf ( n543189 , n543188 );
xor ( n15930 , n12076 , n15842 );
buf ( n543191 , n15930 );
buf ( n543192 , n543191 );
xor ( n15933 , n12421 , n15840 );
buf ( n543194 , n15933 );
buf ( n543195 , n543194 );
xor ( n15936 , n12596 , n15838 );
buf ( n543197 , n15936 );
buf ( n543198 , n543197 );
xor ( n15939 , n12747 , n15836 );
buf ( n543200 , n15939 );
buf ( n543201 , n543200 );
xor ( n15942 , n12749 , n15835 );
buf ( n543203 , n15942 );
buf ( n543204 , n543203 );
xor ( n15945 , n12983 , n15833 );
buf ( n543206 , n15945 );
buf ( n543207 , n543206 );
xor ( n15948 , n13077 , n15831 );
buf ( n543209 , n15948 );
buf ( n543210 , n543209 );
xor ( n15951 , n13335 , n15829 );
buf ( n543212 , n15951 );
buf ( n543213 , n543212 );
xor ( n15954 , n13776 , n15827 );
buf ( n543215 , n15954 );
buf ( n543216 , n543215 );
xor ( n15957 , n13778 , n15826 );
buf ( n543218 , n15957 );
buf ( n543219 , n543218 );
xor ( n15960 , n13780 , n15825 );
buf ( n543221 , n15960 );
buf ( n543222 , n543221 );
xor ( n15963 , n14007 , n15823 );
buf ( n543224 , n15963 );
buf ( n543225 , n543224 );
xor ( n15966 , n14664 , n15821 );
buf ( n543227 , n15966 );
buf ( n543228 , n543227 );
xor ( n15969 , n14666 , n15820 );
buf ( n543230 , n15969 );
buf ( n543231 , n543230 );
xor ( n15972 , n14668 , n15819 );
buf ( n543233 , n15972 );
buf ( n543234 , n543233 );
xor ( n15975 , n14670 , n15818 );
buf ( n543236 , n15975 );
buf ( n543237 , n543236 );
xor ( n15978 , n14672 , n15817 );
buf ( n543239 , n15978 );
buf ( n543240 , n543239 );
xor ( n15981 , n14674 , n15816 );
buf ( n543242 , n15981 );
buf ( n543243 , n543242 );
xor ( n15984 , n15106 , n15814 );
buf ( n543245 , n15984 );
buf ( n543246 , n543245 );
xor ( n15987 , n15108 , n15813 );
buf ( n543248 , n15987 );
buf ( n543249 , n543248 );
xor ( n15990 , n15110 , n15812 );
buf ( n543251 , n15990 );
buf ( n543252 , n543251 );
xor ( n15993 , n15112 , n15811 );
buf ( n543254 , n15993 );
buf ( n543255 , n543254 );
xor ( n15996 , n15114 , n15810 );
buf ( n543257 , n15996 );
buf ( n543258 , n543257 );
xor ( n15999 , n15116 , n15809 );
buf ( n543260 , n15999 );
buf ( n543261 , n543260 );
xor ( n16002 , n15228 , n15807 );
buf ( n543263 , n16002 );
buf ( n543264 , n543263 );
xor ( n16005 , n15230 , n15806 );
buf ( n543266 , n16005 );
buf ( n543267 , n543266 );
xor ( n16008 , n15285 , n15804 );
buf ( n543269 , n16008 );
buf ( n543270 , n543269 );
xor ( n16011 , n15341 , n15802 );
buf ( n543272 , n16011 );
buf ( n543273 , n543272 );
xor ( n16014 , n15393 , n15800 );
buf ( n543275 , n16014 );
buf ( n543276 , n543275 );
xor ( n16017 , n15438 , n15798 );
buf ( n543278 , n16017 );
buf ( n543279 , n543278 );
xor ( n16020 , n15484 , n15796 );
buf ( n543281 , n16020 );
buf ( n543282 , n543281 );
xor ( n16023 , n15526 , n15794 );
buf ( n543284 , n16023 );
buf ( n543285 , n543284 );
xor ( n16026 , n15563 , n15792 );
buf ( n543287 , n16026 );
buf ( n543288 , n543287 );
xor ( n16029 , n15599 , n15790 );
buf ( n543290 , n16029 );
buf ( n543291 , n543290 );
xor ( n16032 , n15631 , n15788 );
buf ( n543293 , n16032 );
buf ( n543294 , n543293 );
xor ( n16035 , n15658 , n15786 );
buf ( n543296 , n16035 );
buf ( n543297 , n543296 );
xor ( n16038 , n15688 , n15784 );
buf ( n543299 , n16038 );
buf ( n543300 , n543299 );
xor ( n16041 , n15706 , n15782 );
buf ( n543302 , n16041 );
buf ( n543303 , n543302 );
xor ( n16044 , n15735 , n15780 );
buf ( n543305 , n16044 );
buf ( n543306 , n543305 );
xor ( n16047 , n15743 , n15778 );
buf ( n543308 , n16047 );
buf ( n543309 , n543308 );
xor ( n16050 , n15751 , n15776 );
buf ( n543311 , n16050 );
buf ( n543312 , n543311 );
xor ( n16053 , n15758 , n15774 );
buf ( n543314 , n16053 );
buf ( n543315 , n543314 );
xor ( n16056 , n15764 , n15772 );
buf ( n543317 , n16056 );
buf ( n543318 , n543317 );
xor ( n16059 , n15768 , n15771 );
buf ( n543320 , n16059 );
buf ( n543321 , n543320 );
buf ( n16062 , n15769 );
buf ( n543323 , n16062 );
buf ( n543324 , n543323 );
buf ( n543325 , n1090 );
buf ( n16066 , n543325 );
buf ( n543327 , n1156 );
buf ( n16068 , n543327 );
buf ( n543329 , n1157 );
buf ( n16070 , n543329 );
xor ( n16071 , n16068 , n16070 );
buf ( n543332 , n1158 );
buf ( n16073 , n543332 );
xor ( n16074 , n16070 , n16073 );
not ( n16075 , n16074 );
and ( n16076 , n16071 , n16075 );
and ( n16077 , n16066 , n16076 );
not ( n16078 , n16077 );
and ( n16079 , n16070 , n16073 );
not ( n16080 , n16079 );
and ( n16081 , n16068 , n16080 );
xnor ( n16082 , n16078 , n16081 );
not ( n16083 , n16082 );
buf ( n543344 , n1092 );
buf ( n16085 , n543344 );
buf ( n543346 , n1154 );
buf ( n16087 , n543346 );
buf ( n543348 , n1155 );
buf ( n16089 , n543348 );
xor ( n16090 , n16087 , n16089 );
xor ( n16091 , n16089 , n16068 );
not ( n16092 , n16091 );
and ( n16093 , n16090 , n16092 );
and ( n16094 , n16085 , n16093 );
buf ( n543355 , n1091 );
buf ( n16096 , n543355 );
and ( n16097 , n16096 , n16091 );
nor ( n16098 , n16094 , n16097 );
and ( n16099 , n16089 , n16068 );
not ( n16100 , n16099 );
and ( n16101 , n16087 , n16100 );
xnor ( n16102 , n16098 , n16101 );
and ( n16103 , n16083 , n16102 );
buf ( n543364 , n1093 );
buf ( n16105 , n543364 );
and ( n16106 , n16105 , n16087 );
and ( n16107 , n16102 , n16106 );
and ( n16108 , n16083 , n16106 );
or ( n16109 , n16103 , n16107 , n16108 );
buf ( n16110 , n16082 );
xor ( n16111 , n16109 , n16110 );
not ( n16112 , n16081 );
and ( n16113 , n16096 , n16093 );
and ( n16114 , n16066 , n16091 );
nor ( n16115 , n16113 , n16114 );
xnor ( n16116 , n16115 , n16101 );
xor ( n16117 , n16112 , n16116 );
and ( n16118 , n16085 , n16087 );
xor ( n16119 , n16117 , n16118 );
xor ( n16120 , n16111 , n16119 );
buf ( n543381 , n1159 );
buf ( n16122 , n543381 );
buf ( n543383 , n1160 );
buf ( n16124 , n543383 );
and ( n16125 , n16122 , n16124 );
not ( n16126 , n16125 );
and ( n16127 , n16073 , n16126 );
not ( n16128 , n16127 );
and ( n16129 , n16096 , n16076 );
and ( n16130 , n16066 , n16074 );
nor ( n16131 , n16129 , n16130 );
xnor ( n16132 , n16131 , n16081 );
and ( n16133 , n16128 , n16132 );
buf ( n543394 , n1094 );
buf ( n16135 , n543394 );
and ( n16136 , n16135 , n16087 );
and ( n16137 , n16132 , n16136 );
and ( n16138 , n16128 , n16136 );
or ( n16139 , n16133 , n16137 , n16138 );
and ( n16140 , n16085 , n16076 );
and ( n16141 , n16096 , n16074 );
nor ( n16142 , n16140 , n16141 );
xnor ( n16143 , n16142 , n16081 );
and ( n16144 , n16135 , n16093 );
and ( n16145 , n16105 , n16091 );
nor ( n16146 , n16144 , n16145 );
xnor ( n16147 , n16146 , n16101 );
and ( n16148 , n16143 , n16147 );
buf ( n543409 , n1095 );
buf ( n16150 , n543409 );
and ( n16151 , n16150 , n16087 );
and ( n16152 , n16147 , n16151 );
and ( n16153 , n16143 , n16151 );
or ( n16154 , n16148 , n16152 , n16153 );
xor ( n16155 , n16073 , n16122 );
xor ( n16156 , n16122 , n16124 );
not ( n16157 , n16156 );
and ( n16158 , n16155 , n16157 );
and ( n16159 , n16066 , n16158 );
not ( n16160 , n16159 );
xnor ( n16161 , n16160 , n16127 );
buf ( n16162 , n16161 );
and ( n16163 , n16154 , n16162 );
and ( n16164 , n16105 , n16093 );
and ( n16165 , n16085 , n16091 );
nor ( n16166 , n16164 , n16165 );
xnor ( n16167 , n16166 , n16101 );
and ( n16168 , n16162 , n16167 );
and ( n16169 , n16154 , n16167 );
or ( n16170 , n16163 , n16168 , n16169 );
and ( n16171 , n16139 , n16170 );
xor ( n16172 , n16083 , n16102 );
xor ( n16173 , n16172 , n16106 );
and ( n16174 , n16170 , n16173 );
and ( n16175 , n16139 , n16173 );
or ( n16176 , n16171 , n16174 , n16175 );
xor ( n16177 , n16120 , n16176 );
xor ( n16178 , n16139 , n16170 );
xor ( n16179 , n16178 , n16173 );
buf ( n543440 , n1161 );
buf ( n16181 , n543440 );
buf ( n543442 , n1162 );
buf ( n16183 , n543442 );
and ( n16184 , n16181 , n16183 );
not ( n16185 , n16184 );
and ( n16186 , n16124 , n16185 );
not ( n16187 , n16186 );
and ( n16188 , n16096 , n16158 );
and ( n16189 , n16066 , n16156 );
nor ( n16190 , n16188 , n16189 );
xnor ( n16191 , n16190 , n16127 );
and ( n16192 , n16187 , n16191 );
and ( n16193 , n16150 , n16093 );
and ( n16194 , n16135 , n16091 );
nor ( n16195 , n16193 , n16194 );
xnor ( n16196 , n16195 , n16101 );
and ( n16197 , n16191 , n16196 );
and ( n16198 , n16187 , n16196 );
or ( n16199 , n16192 , n16197 , n16198 );
not ( n16200 , n16161 );
and ( n16201 , n16199 , n16200 );
xor ( n16202 , n16143 , n16147 );
xor ( n16203 , n16202 , n16151 );
and ( n16204 , n16200 , n16203 );
and ( n16205 , n16199 , n16203 );
or ( n16206 , n16201 , n16204 , n16205 );
xor ( n16207 , n16128 , n16132 );
xor ( n16208 , n16207 , n16136 );
and ( n16209 , n16206 , n16208 );
xor ( n16210 , n16154 , n16162 );
xor ( n16211 , n16210 , n16167 );
and ( n16212 , n16208 , n16211 );
and ( n16213 , n16206 , n16211 );
or ( n16214 , n16209 , n16212 , n16213 );
and ( n16215 , n16179 , n16214 );
xor ( n16216 , n16206 , n16208 );
xor ( n16217 , n16216 , n16211 );
and ( n16218 , n16085 , n16158 );
and ( n16219 , n16096 , n16156 );
nor ( n16220 , n16218 , n16219 );
xnor ( n16221 , n16220 , n16127 );
buf ( n16222 , n16221 );
and ( n16223 , n16105 , n16076 );
and ( n16224 , n16085 , n16074 );
nor ( n16225 , n16223 , n16224 );
xnor ( n16226 , n16225 , n16081 );
and ( n16227 , n16222 , n16226 );
buf ( n543488 , n1096 );
buf ( n16229 , n543488 );
and ( n16230 , n16229 , n16087 );
and ( n16231 , n16226 , n16230 );
and ( n16232 , n16222 , n16230 );
or ( n16233 , n16227 , n16231 , n16232 );
xor ( n16234 , n16124 , n16181 );
xor ( n16235 , n16181 , n16183 );
not ( n16236 , n16235 );
and ( n16237 , n16234 , n16236 );
and ( n16238 , n16066 , n16237 );
not ( n16239 , n16238 );
xnor ( n16240 , n16239 , n16186 );
and ( n16241 , n16229 , n16093 );
and ( n16242 , n16150 , n16091 );
nor ( n16243 , n16241 , n16242 );
xnor ( n16244 , n16243 , n16101 );
and ( n16245 , n16240 , n16244 );
buf ( n543506 , n1097 );
buf ( n16247 , n543506 );
and ( n16248 , n16247 , n16087 );
and ( n16249 , n16244 , n16248 );
and ( n16250 , n16240 , n16248 );
or ( n16251 , n16245 , n16249 , n16250 );
xor ( n16252 , n16187 , n16191 );
xor ( n16253 , n16252 , n16196 );
and ( n16254 , n16251 , n16253 );
xor ( n16255 , n16222 , n16226 );
xor ( n16256 , n16255 , n16230 );
and ( n16257 , n16253 , n16256 );
and ( n16258 , n16251 , n16256 );
or ( n16259 , n16254 , n16257 , n16258 );
and ( n16260 , n16233 , n16259 );
xor ( n16261 , n16199 , n16200 );
xor ( n16262 , n16261 , n16203 );
and ( n16263 , n16259 , n16262 );
and ( n16264 , n16233 , n16262 );
or ( n16265 , n16260 , n16263 , n16264 );
and ( n16266 , n16217 , n16265 );
xor ( n16267 , n16233 , n16259 );
xor ( n16268 , n16267 , n16262 );
and ( n16269 , n16105 , n16158 );
and ( n16270 , n16085 , n16156 );
nor ( n16271 , n16269 , n16270 );
xnor ( n16272 , n16271 , n16127 );
and ( n16273 , n16247 , n16093 );
and ( n16274 , n16229 , n16091 );
nor ( n16275 , n16273 , n16274 );
xnor ( n16276 , n16275 , n16101 );
and ( n16277 , n16272 , n16276 );
buf ( n543538 , n1098 );
buf ( n16279 , n543538 );
and ( n16280 , n16279 , n16087 );
and ( n16281 , n16276 , n16280 );
and ( n16282 , n16272 , n16280 );
or ( n16283 , n16277 , n16281 , n16282 );
not ( n16284 , n16221 );
and ( n16285 , n16283 , n16284 );
and ( n16286 , n16135 , n16076 );
and ( n16287 , n16105 , n16074 );
nor ( n16288 , n16286 , n16287 );
xnor ( n16289 , n16288 , n16081 );
and ( n16290 , n16284 , n16289 );
and ( n16291 , n16283 , n16289 );
or ( n16292 , n16285 , n16290 , n16291 );
buf ( n543553 , n1163 );
buf ( n16294 , n543553 );
buf ( n543555 , n1164 );
buf ( n16296 , n543555 );
and ( n16297 , n16294 , n16296 );
not ( n16298 , n16297 );
and ( n16299 , n16183 , n16298 );
not ( n16300 , n16299 );
and ( n16301 , n16096 , n16237 );
and ( n16302 , n16066 , n16235 );
nor ( n16303 , n16301 , n16302 );
xnor ( n16304 , n16303 , n16186 );
and ( n16305 , n16300 , n16304 );
and ( n16306 , n16150 , n16076 );
and ( n16307 , n16135 , n16074 );
nor ( n16308 , n16306 , n16307 );
xnor ( n16309 , n16308 , n16081 );
and ( n16310 , n16304 , n16309 );
and ( n16311 , n16300 , n16309 );
or ( n16312 , n16305 , n16310 , n16311 );
xor ( n16313 , n16240 , n16244 );
xor ( n16314 , n16313 , n16248 );
and ( n16315 , n16312 , n16314 );
xor ( n16316 , n16283 , n16284 );
xor ( n16317 , n16316 , n16289 );
and ( n16318 , n16314 , n16317 );
and ( n16319 , n16312 , n16317 );
or ( n16320 , n16315 , n16318 , n16319 );
and ( n16321 , n16292 , n16320 );
xor ( n16322 , n16251 , n16253 );
xor ( n16323 , n16322 , n16256 );
and ( n16324 , n16320 , n16323 );
and ( n16325 , n16292 , n16323 );
or ( n16326 , n16321 , n16324 , n16325 );
and ( n16327 , n16268 , n16326 );
xor ( n16328 , n16183 , n16294 );
xor ( n16329 , n16294 , n16296 );
not ( n16330 , n16329 );
and ( n16331 , n16328 , n16330 );
and ( n16332 , n16066 , n16331 );
not ( n16333 , n16332 );
xnor ( n16334 , n16333 , n16299 );
and ( n16335 , n16229 , n16076 );
and ( n16336 , n16150 , n16074 );
nor ( n16337 , n16335 , n16336 );
xnor ( n16338 , n16337 , n16081 );
and ( n16339 , n16334 , n16338 );
and ( n16340 , n16279 , n16093 );
and ( n16341 , n16247 , n16091 );
nor ( n16342 , n16340 , n16341 );
xnor ( n16343 , n16342 , n16101 );
and ( n16344 , n16338 , n16343 );
and ( n16345 , n16334 , n16343 );
or ( n16346 , n16339 , n16344 , n16345 );
and ( n16347 , n16085 , n16237 );
and ( n16348 , n16096 , n16235 );
nor ( n16349 , n16347 , n16348 );
xnor ( n16350 , n16349 , n16186 );
buf ( n16351 , n16350 );
and ( n16352 , n16346 , n16351 );
xor ( n16353 , n16272 , n16276 );
xor ( n16354 , n16353 , n16280 );
and ( n16355 , n16351 , n16354 );
and ( n16356 , n16346 , n16354 );
or ( n16357 , n16352 , n16355 , n16356 );
not ( n16358 , n16350 );
and ( n16359 , n16135 , n16158 );
and ( n16360 , n16105 , n16156 );
nor ( n16361 , n16359 , n16360 );
xnor ( n16362 , n16361 , n16127 );
and ( n16363 , n16358 , n16362 );
buf ( n543624 , n1099 );
buf ( n16365 , n543624 );
and ( n16366 , n16365 , n16087 );
and ( n16367 , n16362 , n16366 );
and ( n16368 , n16358 , n16366 );
or ( n16369 , n16363 , n16367 , n16368 );
xor ( n16370 , n16300 , n16304 );
xor ( n16371 , n16370 , n16309 );
and ( n16372 , n16369 , n16371 );
xor ( n16373 , n16346 , n16351 );
xor ( n16374 , n16373 , n16354 );
and ( n16375 , n16371 , n16374 );
and ( n16376 , n16369 , n16374 );
or ( n16377 , n16372 , n16375 , n16376 );
and ( n16378 , n16357 , n16377 );
xor ( n16379 , n16312 , n16314 );
xor ( n16380 , n16379 , n16317 );
and ( n16381 , n16377 , n16380 );
and ( n16382 , n16357 , n16380 );
or ( n16383 , n16378 , n16381 , n16382 );
xor ( n16384 , n16292 , n16320 );
xor ( n16385 , n16384 , n16323 );
and ( n16386 , n16383 , n16385 );
xor ( n16387 , n16357 , n16377 );
xor ( n16388 , n16387 , n16380 );
buf ( n543649 , n1165 );
buf ( n16390 , n543649 );
buf ( n543651 , n1166 );
buf ( n16392 , n543651 );
and ( n16393 , n16390 , n16392 );
not ( n16394 , n16393 );
and ( n16395 , n16296 , n16394 );
not ( n16396 , n16395 );
and ( n16397 , n16096 , n16331 );
and ( n16398 , n16066 , n16329 );
nor ( n16399 , n16397 , n16398 );
xnor ( n16400 , n16399 , n16299 );
and ( n16401 , n16396 , n16400 );
and ( n16402 , n16150 , n16158 );
and ( n16403 , n16135 , n16156 );
nor ( n16404 , n16402 , n16403 );
xnor ( n16405 , n16404 , n16127 );
and ( n16406 , n16400 , n16405 );
and ( n16407 , n16396 , n16405 );
or ( n16408 , n16401 , n16406 , n16407 );
and ( n16409 , n16105 , n16237 );
and ( n16410 , n16085 , n16235 );
nor ( n16411 , n16409 , n16410 );
xnor ( n16412 , n16411 , n16186 );
and ( n16413 , n16247 , n16076 );
and ( n16414 , n16229 , n16074 );
nor ( n16415 , n16413 , n16414 );
xnor ( n16416 , n16415 , n16081 );
and ( n16417 , n16412 , n16416 );
and ( n16418 , n16365 , n16093 );
and ( n16419 , n16279 , n16091 );
nor ( n16420 , n16418 , n16419 );
xnor ( n16421 , n16420 , n16101 );
and ( n16422 , n16416 , n16421 );
and ( n16423 , n16412 , n16421 );
or ( n16424 , n16417 , n16422 , n16423 );
and ( n16425 , n16408 , n16424 );
xor ( n16426 , n16334 , n16338 );
xor ( n16427 , n16426 , n16343 );
and ( n16428 , n16424 , n16427 );
and ( n16429 , n16408 , n16427 );
or ( n16430 , n16425 , n16428 , n16429 );
and ( n16431 , n16085 , n16331 );
and ( n16432 , n16096 , n16329 );
nor ( n16433 , n16431 , n16432 );
xnor ( n16434 , n16433 , n16299 );
and ( n16435 , n16229 , n16158 );
and ( n16436 , n16150 , n16156 );
nor ( n16437 , n16435 , n16436 );
xnor ( n16438 , n16437 , n16127 );
and ( n16439 , n16434 , n16438 );
and ( n16440 , n16279 , n16076 );
and ( n16441 , n16247 , n16074 );
nor ( n16442 , n16440 , n16441 );
xnor ( n16443 , n16442 , n16081 );
and ( n16444 , n16438 , n16443 );
and ( n16445 , n16434 , n16443 );
or ( n16446 , n16439 , n16444 , n16445 );
xor ( n16447 , n16296 , n16390 );
xor ( n16448 , n16390 , n16392 );
not ( n16449 , n16448 );
and ( n16450 , n16447 , n16449 );
and ( n16451 , n16066 , n16450 );
not ( n16452 , n16451 );
xnor ( n16453 , n16452 , n16395 );
buf ( n16454 , n16453 );
and ( n16455 , n16446 , n16454 );
buf ( n543716 , n1100 );
buf ( n16457 , n543716 );
and ( n16458 , n16457 , n16087 );
and ( n16459 , n16454 , n16458 );
and ( n16460 , n16446 , n16458 );
or ( n16461 , n16455 , n16459 , n16460 );
and ( n16462 , n16135 , n16237 );
and ( n16463 , n16105 , n16235 );
nor ( n16464 , n16462 , n16463 );
xnor ( n16465 , n16464 , n16186 );
and ( n16466 , n16457 , n16093 );
and ( n16467 , n16365 , n16091 );
nor ( n16468 , n16466 , n16467 );
xnor ( n16469 , n16468 , n16101 );
and ( n16470 , n16465 , n16469 );
buf ( n543731 , n1101 );
buf ( n16472 , n543731 );
and ( n16473 , n16472 , n16087 );
and ( n16474 , n16469 , n16473 );
and ( n16475 , n16465 , n16473 );
or ( n16476 , n16470 , n16474 , n16475 );
xor ( n16477 , n16396 , n16400 );
xor ( n16478 , n16477 , n16405 );
and ( n16479 , n16476 , n16478 );
xor ( n16480 , n16412 , n16416 );
xor ( n16481 , n16480 , n16421 );
and ( n16482 , n16478 , n16481 );
and ( n16483 , n16476 , n16481 );
or ( n16484 , n16479 , n16482 , n16483 );
and ( n16485 , n16461 , n16484 );
xor ( n16486 , n16358 , n16362 );
xor ( n16487 , n16486 , n16366 );
and ( n16488 , n16484 , n16487 );
and ( n16489 , n16461 , n16487 );
or ( n16490 , n16485 , n16488 , n16489 );
and ( n16491 , n16430 , n16490 );
xor ( n16492 , n16369 , n16371 );
xor ( n16493 , n16492 , n16374 );
and ( n16494 , n16490 , n16493 );
and ( n16495 , n16430 , n16493 );
or ( n16496 , n16491 , n16494 , n16495 );
and ( n16497 , n16388 , n16496 );
xor ( n16498 , n16430 , n16490 );
xor ( n16499 , n16498 , n16493 );
and ( n16500 , n16105 , n16331 );
and ( n16501 , n16085 , n16329 );
nor ( n16502 , n16500 , n16501 );
xnor ( n16503 , n16502 , n16299 );
and ( n16504 , n16247 , n16158 );
and ( n16505 , n16229 , n16156 );
nor ( n16506 , n16504 , n16505 );
xnor ( n16507 , n16506 , n16127 );
and ( n16508 , n16503 , n16507 );
buf ( n543769 , n1102 );
buf ( n16510 , n543769 );
and ( n16511 , n16510 , n16087 );
and ( n16512 , n16507 , n16511 );
and ( n16513 , n16503 , n16511 );
or ( n16514 , n16508 , n16512 , n16513 );
buf ( n543775 , n1167 );
buf ( n16516 , n543775 );
buf ( n543777 , n1168 );
buf ( n16518 , n543777 );
and ( n16519 , n16516 , n16518 );
not ( n16520 , n16519 );
and ( n16521 , n16392 , n16520 );
not ( n16522 , n16521 );
and ( n16523 , n16096 , n16450 );
and ( n16524 , n16066 , n16448 );
nor ( n16525 , n16523 , n16524 );
xnor ( n16526 , n16525 , n16395 );
and ( n16527 , n16522 , n16526 );
and ( n16528 , n16150 , n16237 );
and ( n16529 , n16135 , n16235 );
nor ( n16530 , n16528 , n16529 );
xnor ( n16531 , n16530 , n16186 );
and ( n16532 , n16526 , n16531 );
and ( n16533 , n16522 , n16531 );
or ( n16534 , n16527 , n16532 , n16533 );
and ( n16535 , n16514 , n16534 );
not ( n16536 , n16453 );
and ( n16537 , n16534 , n16536 );
and ( n16538 , n16514 , n16536 );
or ( n16539 , n16535 , n16537 , n16538 );
xor ( n16540 , n16392 , n16516 );
xor ( n16541 , n16516 , n16518 );
not ( n16542 , n16541 );
and ( n16543 , n16540 , n16542 );
and ( n16544 , n16066 , n16543 );
not ( n16545 , n16544 );
xnor ( n16546 , n16545 , n16521 );
buf ( n16547 , n16546 );
and ( n16548 , n16365 , n16076 );
and ( n16549 , n16279 , n16074 );
nor ( n16550 , n16548 , n16549 );
xnor ( n16551 , n16550 , n16081 );
and ( n16552 , n16547 , n16551 );
and ( n16553 , n16472 , n16093 );
and ( n16554 , n16457 , n16091 );
nor ( n16555 , n16553 , n16554 );
xnor ( n16556 , n16555 , n16101 );
and ( n16557 , n16551 , n16556 );
and ( n16558 , n16547 , n16556 );
or ( n16559 , n16552 , n16557 , n16558 );
xor ( n16560 , n16465 , n16469 );
xor ( n16561 , n16560 , n16473 );
and ( n16562 , n16559 , n16561 );
xor ( n16563 , n16434 , n16438 );
xor ( n16564 , n16563 , n16443 );
and ( n16565 , n16561 , n16564 );
and ( n16566 , n16559 , n16564 );
or ( n16567 , n16562 , n16565 , n16566 );
and ( n16568 , n16539 , n16567 );
xor ( n16569 , n16446 , n16454 );
xor ( n16570 , n16569 , n16458 );
and ( n16571 , n16567 , n16570 );
and ( n16572 , n16539 , n16570 );
or ( n16573 , n16568 , n16571 , n16572 );
xor ( n16574 , n16408 , n16424 );
xor ( n16575 , n16574 , n16427 );
and ( n16576 , n16573 , n16575 );
xor ( n16577 , n16461 , n16484 );
xor ( n16578 , n16577 , n16487 );
and ( n16579 , n16575 , n16578 );
and ( n16580 , n16573 , n16578 );
or ( n16581 , n16576 , n16579 , n16580 );
and ( n16582 , n16499 , n16581 );
xor ( n16583 , n16573 , n16575 );
xor ( n16584 , n16583 , n16578 );
and ( n16585 , n16135 , n16331 );
and ( n16586 , n16105 , n16329 );
nor ( n16587 , n16585 , n16586 );
xnor ( n16588 , n16587 , n16299 );
and ( n16589 , n16279 , n16158 );
and ( n16590 , n16247 , n16156 );
nor ( n16591 , n16589 , n16590 );
xnor ( n16592 , n16591 , n16127 );
and ( n16593 , n16588 , n16592 );
and ( n16594 , n16457 , n16076 );
and ( n16595 , n16365 , n16074 );
nor ( n16596 , n16594 , n16595 );
xnor ( n16597 , n16596 , n16081 );
and ( n16598 , n16592 , n16597 );
and ( n16599 , n16588 , n16597 );
or ( n16600 , n16593 , n16598 , n16599 );
and ( n16601 , n16085 , n16450 );
and ( n16602 , n16096 , n16448 );
nor ( n16603 , n16601 , n16602 );
xnor ( n16604 , n16603 , n16395 );
and ( n16605 , n16229 , n16237 );
and ( n16606 , n16150 , n16235 );
nor ( n16607 , n16605 , n16606 );
xnor ( n16608 , n16607 , n16186 );
and ( n16609 , n16604 , n16608 );
buf ( n543870 , n1103 );
buf ( n16611 , n543870 );
and ( n16612 , n16611 , n16087 );
and ( n16613 , n16608 , n16612 );
and ( n16614 , n16604 , n16612 );
or ( n16615 , n16609 , n16613 , n16614 );
and ( n16616 , n16600 , n16615 );
xor ( n16617 , n16522 , n16526 );
xor ( n16618 , n16617 , n16531 );
and ( n16619 , n16615 , n16618 );
and ( n16620 , n16600 , n16618 );
or ( n16621 , n16616 , n16619 , n16620 );
xor ( n16622 , n16514 , n16534 );
xor ( n16623 , n16622 , n16536 );
and ( n16624 , n16621 , n16623 );
xor ( n16625 , n16559 , n16561 );
xor ( n16626 , n16625 , n16564 );
and ( n16627 , n16623 , n16626 );
and ( n16628 , n16621 , n16626 );
or ( n16629 , n16624 , n16627 , n16628 );
xor ( n16630 , n16476 , n16478 );
xor ( n16631 , n16630 , n16481 );
and ( n16632 , n16629 , n16631 );
xor ( n16633 , n16539 , n16567 );
xor ( n16634 , n16633 , n16570 );
and ( n16635 , n16631 , n16634 );
and ( n16636 , n16629 , n16634 );
or ( n16637 , n16632 , n16635 , n16636 );
and ( n16638 , n16584 , n16637 );
xor ( n16639 , n16629 , n16631 );
xor ( n16640 , n16639 , n16634 );
buf ( n543901 , n1169 );
buf ( n16642 , n543901 );
buf ( n543903 , n1170 );
buf ( n16644 , n543903 );
and ( n16645 , n16642 , n16644 );
not ( n16646 , n16645 );
and ( n16647 , n16518 , n16646 );
not ( n16648 , n16647 );
and ( n16649 , n16096 , n16543 );
and ( n16650 , n16066 , n16541 );
nor ( n16651 , n16649 , n16650 );
xnor ( n16652 , n16651 , n16521 );
and ( n16653 , n16648 , n16652 );
and ( n16654 , n16150 , n16331 );
and ( n16655 , n16135 , n16329 );
nor ( n16656 , n16654 , n16655 );
xnor ( n16657 , n16656 , n16299 );
and ( n16658 , n16652 , n16657 );
and ( n16659 , n16648 , n16657 );
or ( n16660 , n16653 , n16658 , n16659 );
not ( n16661 , n16546 );
and ( n16662 , n16660 , n16661 );
and ( n16663 , n16510 , n16093 );
and ( n16664 , n16472 , n16091 );
nor ( n16665 , n16663 , n16664 );
xnor ( n16666 , n16665 , n16101 );
and ( n16667 , n16661 , n16666 );
and ( n16668 , n16660 , n16666 );
or ( n16669 , n16662 , n16667 , n16668 );
xor ( n16670 , n16503 , n16507 );
xor ( n16671 , n16670 , n16511 );
and ( n16672 , n16669 , n16671 );
xor ( n16673 , n16547 , n16551 );
xor ( n16674 , n16673 , n16556 );
and ( n16675 , n16671 , n16674 );
and ( n16676 , n16669 , n16674 );
or ( n16677 , n16672 , n16675 , n16676 );
and ( n16678 , n16247 , n16237 );
and ( n16679 , n16229 , n16235 );
nor ( n16680 , n16678 , n16679 );
xnor ( n16681 , n16680 , n16186 );
and ( n16682 , n16611 , n16093 );
and ( n16683 , n16510 , n16091 );
nor ( n16684 , n16682 , n16683 );
xnor ( n16685 , n16684 , n16101 );
and ( n16686 , n16681 , n16685 );
buf ( n543947 , n1104 );
buf ( n16688 , n543947 );
and ( n16689 , n16688 , n16087 );
and ( n16690 , n16685 , n16689 );
and ( n16691 , n16681 , n16689 );
or ( n16692 , n16686 , n16690 , n16691 );
and ( n16693 , n16105 , n16450 );
and ( n16694 , n16085 , n16448 );
nor ( n16695 , n16693 , n16694 );
xnor ( n16696 , n16695 , n16395 );
and ( n16697 , n16365 , n16158 );
and ( n16698 , n16279 , n16156 );
nor ( n16699 , n16697 , n16698 );
xnor ( n16700 , n16699 , n16127 );
and ( n16701 , n16696 , n16700 );
and ( n16702 , n16472 , n16076 );
and ( n16703 , n16457 , n16074 );
nor ( n16704 , n16702 , n16703 );
xnor ( n16705 , n16704 , n16081 );
and ( n16706 , n16700 , n16705 );
and ( n16707 , n16696 , n16705 );
or ( n16708 , n16701 , n16706 , n16707 );
and ( n16709 , n16692 , n16708 );
xor ( n16710 , n16588 , n16592 );
xor ( n16711 , n16710 , n16597 );
and ( n16712 , n16708 , n16711 );
and ( n16713 , n16692 , n16711 );
or ( n16714 , n16709 , n16712 , n16713 );
and ( n16715 , n16229 , n16331 );
and ( n16716 , n16150 , n16329 );
nor ( n16717 , n16715 , n16716 );
xnor ( n16718 , n16717 , n16299 );
and ( n16719 , n16688 , n16093 );
and ( n16720 , n16611 , n16091 );
nor ( n16721 , n16719 , n16720 );
xnor ( n16722 , n16721 , n16101 );
and ( n16723 , n16718 , n16722 );
buf ( n543984 , n1105 );
buf ( n16725 , n543984 );
and ( n16726 , n16725 , n16087 );
and ( n16727 , n16722 , n16726 );
and ( n16728 , n16718 , n16726 );
or ( n16729 , n16723 , n16727 , n16728 );
and ( n16730 , n16085 , n16543 );
and ( n16731 , n16096 , n16541 );
nor ( n16732 , n16730 , n16731 );
xnor ( n16733 , n16732 , n16521 );
and ( n16734 , n16135 , n16450 );
and ( n16735 , n16105 , n16448 );
nor ( n16736 , n16734 , n16735 );
xnor ( n16737 , n16736 , n16395 );
and ( n16738 , n16733 , n16737 );
and ( n16739 , n16279 , n16237 );
and ( n16740 , n16247 , n16235 );
nor ( n16741 , n16739 , n16740 );
xnor ( n16742 , n16741 , n16186 );
and ( n16743 , n16737 , n16742 );
and ( n16744 , n16733 , n16742 );
or ( n16745 , n16738 , n16743 , n16744 );
and ( n16746 , n16729 , n16745 );
xor ( n16747 , n16518 , n16642 );
xor ( n16748 , n16642 , n16644 );
not ( n16749 , n16748 );
and ( n16750 , n16747 , n16749 );
and ( n16751 , n16066 , n16750 );
not ( n16752 , n16751 );
xnor ( n16753 , n16752 , n16647 );
buf ( n16754 , n16753 );
and ( n16755 , n16745 , n16754 );
and ( n16756 , n16729 , n16754 );
or ( n16757 , n16746 , n16755 , n16756 );
xor ( n16758 , n16604 , n16608 );
xor ( n16759 , n16758 , n16612 );
and ( n16760 , n16757 , n16759 );
xor ( n16761 , n16660 , n16661 );
xor ( n16762 , n16761 , n16666 );
and ( n16763 , n16759 , n16762 );
and ( n16764 , n16757 , n16762 );
or ( n16765 , n16760 , n16763 , n16764 );
and ( n16766 , n16714 , n16765 );
xor ( n16767 , n16600 , n16615 );
xor ( n16768 , n16767 , n16618 );
and ( n16769 , n16765 , n16768 );
and ( n16770 , n16714 , n16768 );
or ( n16771 , n16766 , n16769 , n16770 );
and ( n16772 , n16677 , n16771 );
xor ( n16773 , n16621 , n16623 );
xor ( n16774 , n16773 , n16626 );
and ( n16775 , n16771 , n16774 );
and ( n16776 , n16677 , n16774 );
or ( n16777 , n16772 , n16775 , n16776 );
and ( n16778 , n16640 , n16777 );
xor ( n16779 , n16681 , n16685 );
xor ( n16780 , n16779 , n16689 );
xor ( n16781 , n16696 , n16700 );
xor ( n16782 , n16781 , n16705 );
and ( n16783 , n16780 , n16782 );
xor ( n16784 , n16648 , n16652 );
xor ( n16785 , n16784 , n16657 );
and ( n16786 , n16782 , n16785 );
and ( n16787 , n16780 , n16785 );
or ( n16788 , n16783 , n16786 , n16787 );
xor ( n16789 , n16692 , n16708 );
xor ( n16790 , n16789 , n16711 );
and ( n16791 , n16788 , n16790 );
xor ( n16792 , n16757 , n16759 );
xor ( n16793 , n16792 , n16762 );
and ( n16794 , n16790 , n16793 );
and ( n16795 , n16788 , n16793 );
or ( n16796 , n16791 , n16794 , n16795 );
xor ( n16797 , n16669 , n16671 );
xor ( n16798 , n16797 , n16674 );
and ( n16799 , n16796 , n16798 );
xor ( n16800 , n16714 , n16765 );
xor ( n16801 , n16800 , n16768 );
and ( n16802 , n16798 , n16801 );
and ( n16803 , n16796 , n16801 );
or ( n16804 , n16799 , n16802 , n16803 );
xor ( n16805 , n16677 , n16771 );
xor ( n16806 , n16805 , n16774 );
and ( n16807 , n16804 , n16806 );
xor ( n16808 , n16796 , n16798 );
xor ( n16809 , n16808 , n16801 );
and ( n16810 , n16105 , n16543 );
and ( n16811 , n16085 , n16541 );
nor ( n16812 , n16810 , n16811 );
xnor ( n16813 , n16812 , n16521 );
and ( n16814 , n16365 , n16237 );
and ( n16815 , n16279 , n16235 );
nor ( n16816 , n16814 , n16815 );
xnor ( n16817 , n16816 , n16186 );
and ( n16818 , n16813 , n16817 );
buf ( n544079 , n1106 );
buf ( n16820 , n544079 );
and ( n16821 , n16820 , n16087 );
and ( n16822 , n16817 , n16821 );
and ( n16823 , n16813 , n16821 );
or ( n16824 , n16818 , n16822 , n16823 );
and ( n16825 , n16247 , n16331 );
and ( n16826 , n16229 , n16329 );
nor ( n16827 , n16825 , n16826 );
xnor ( n16828 , n16827 , n16299 );
and ( n16829 , n16611 , n16076 );
and ( n16830 , n16510 , n16074 );
nor ( n16831 , n16829 , n16830 );
xnor ( n16832 , n16831 , n16081 );
and ( n16833 , n16828 , n16832 );
and ( n16834 , n16725 , n16093 );
and ( n16835 , n16688 , n16091 );
nor ( n16836 , n16834 , n16835 );
xnor ( n16837 , n16836 , n16101 );
and ( n16838 , n16832 , n16837 );
and ( n16839 , n16828 , n16837 );
or ( n16840 , n16833 , n16838 , n16839 );
and ( n16841 , n16824 , n16840 );
buf ( n544102 , n1171 );
buf ( n16843 , n544102 );
buf ( n544104 , n1172 );
buf ( n16845 , n544104 );
and ( n16846 , n16843 , n16845 );
not ( n16847 , n16846 );
and ( n16848 , n16644 , n16847 );
not ( n16849 , n16848 );
and ( n16850 , n16096 , n16750 );
and ( n16851 , n16066 , n16748 );
nor ( n16852 , n16850 , n16851 );
xnor ( n16853 , n16852 , n16647 );
and ( n16854 , n16849 , n16853 );
and ( n16855 , n16150 , n16450 );
and ( n16856 , n16135 , n16448 );
nor ( n16857 , n16855 , n16856 );
xnor ( n16858 , n16857 , n16395 );
and ( n16859 , n16853 , n16858 );
and ( n16860 , n16849 , n16858 );
or ( n16861 , n16854 , n16859 , n16860 );
and ( n16862 , n16840 , n16861 );
and ( n16863 , n16824 , n16861 );
or ( n16864 , n16841 , n16862 , n16863 );
not ( n16865 , n16753 );
and ( n16866 , n16457 , n16158 );
and ( n16867 , n16365 , n16156 );
nor ( n16868 , n16866 , n16867 );
xnor ( n16869 , n16868 , n16127 );
and ( n16870 , n16865 , n16869 );
and ( n16871 , n16510 , n16076 );
and ( n16872 , n16472 , n16074 );
nor ( n16873 , n16871 , n16872 );
xnor ( n16874 , n16873 , n16081 );
and ( n16875 , n16869 , n16874 );
and ( n16876 , n16865 , n16874 );
or ( n16877 , n16870 , n16875 , n16876 );
and ( n16878 , n16864 , n16877 );
xor ( n16879 , n16729 , n16745 );
xor ( n16880 , n16879 , n16754 );
and ( n16881 , n16877 , n16880 );
and ( n16882 , n16864 , n16880 );
or ( n16883 , n16878 , n16881 , n16882 );
xor ( n16884 , n16718 , n16722 );
xor ( n16885 , n16884 , n16726 );
xor ( n16886 , n16733 , n16737 );
xor ( n16887 , n16886 , n16742 );
and ( n16888 , n16885 , n16887 );
xor ( n16889 , n16865 , n16869 );
xor ( n16890 , n16889 , n16874 );
and ( n16891 , n16887 , n16890 );
and ( n16892 , n16885 , n16890 );
or ( n16893 , n16888 , n16891 , n16892 );
and ( n16894 , n16229 , n16450 );
and ( n16895 , n16150 , n16448 );
nor ( n16896 , n16894 , n16895 );
xnor ( n16897 , n16896 , n16395 );
and ( n16898 , n16688 , n16076 );
and ( n16899 , n16611 , n16074 );
nor ( n16900 , n16898 , n16899 );
xnor ( n16901 , n16900 , n16081 );
and ( n16902 , n16897 , n16901 );
and ( n16903 , n16820 , n16093 );
and ( n16904 , n16725 , n16091 );
nor ( n16905 , n16903 , n16904 );
xnor ( n16906 , n16905 , n16101 );
and ( n16907 , n16901 , n16906 );
and ( n16908 , n16897 , n16906 );
or ( n16909 , n16902 , n16907 , n16908 );
xor ( n16910 , n16644 , n16843 );
xor ( n16911 , n16843 , n16845 );
not ( n16912 , n16911 );
and ( n16913 , n16910 , n16912 );
and ( n16914 , n16066 , n16913 );
not ( n16915 , n16914 );
xnor ( n16916 , n16915 , n16848 );
buf ( n16917 , n16916 );
and ( n16918 , n16909 , n16917 );
and ( n16919 , n16472 , n16158 );
and ( n16920 , n16457 , n16156 );
nor ( n16921 , n16919 , n16920 );
xnor ( n16922 , n16921 , n16127 );
and ( n16923 , n16917 , n16922 );
and ( n16924 , n16909 , n16922 );
or ( n16925 , n16918 , n16923 , n16924 );
and ( n16926 , n16085 , n16750 );
and ( n16927 , n16096 , n16748 );
nor ( n16928 , n16926 , n16927 );
xnor ( n16929 , n16928 , n16647 );
and ( n16930 , n16279 , n16331 );
and ( n16931 , n16247 , n16329 );
nor ( n16932 , n16930 , n16931 );
xnor ( n16933 , n16932 , n16299 );
and ( n16934 , n16929 , n16933 );
buf ( n544195 , n1107 );
buf ( n16936 , n544195 );
and ( n16937 , n16936 , n16087 );
and ( n16938 , n16933 , n16937 );
and ( n16939 , n16929 , n16937 );
or ( n16940 , n16934 , n16938 , n16939 );
and ( n16941 , n16135 , n16543 );
and ( n16942 , n16105 , n16541 );
nor ( n16943 , n16941 , n16942 );
xnor ( n16944 , n16943 , n16521 );
and ( n16945 , n16457 , n16237 );
and ( n16946 , n16365 , n16235 );
nor ( n16947 , n16945 , n16946 );
xnor ( n16948 , n16947 , n16186 );
and ( n16949 , n16944 , n16948 );
and ( n16950 , n16510 , n16158 );
and ( n16951 , n16472 , n16156 );
nor ( n16952 , n16950 , n16951 );
xnor ( n16953 , n16952 , n16127 );
and ( n16954 , n16948 , n16953 );
and ( n16955 , n16944 , n16953 );
or ( n544216 , n16949 , n16954 , n16955 );
and ( n544217 , n16940 , n544216 );
xor ( n16958 , n16813 , n16817 );
xor ( n544219 , n16958 , n16821 );
and ( n16960 , n544216 , n544219 );
and ( n16961 , n16940 , n544219 );
or ( n16962 , n544217 , n16960 , n16961 );
and ( n16963 , n16925 , n16962 );
xor ( n16964 , n16824 , n16840 );
xor ( n16965 , n16964 , n16861 );
and ( n16966 , n16962 , n16965 );
and ( n16967 , n16925 , n16965 );
or ( n16968 , n16963 , n16966 , n16967 );
and ( n16969 , n16893 , n16968 );
xor ( n16970 , n16780 , n16782 );
xor ( n16971 , n16970 , n16785 );
and ( n16972 , n16968 , n16971 );
and ( n16973 , n16893 , n16971 );
or ( n16974 , n16969 , n16972 , n16973 );
and ( n16975 , n16883 , n16974 );
xor ( n16976 , n16788 , n16790 );
xor ( n16977 , n16976 , n16793 );
and ( n16978 , n16974 , n16977 );
and ( n16979 , n16883 , n16977 );
or ( n16980 , n16975 , n16978 , n16979 );
and ( n16981 , n16809 , n16980 );
xor ( n16982 , n16883 , n16974 );
xor ( n16983 , n16982 , n16977 );
xor ( n16984 , n16828 , n16832 );
xor ( n16985 , n16984 , n16837 );
xor ( n16986 , n16849 , n16853 );
xor ( n16987 , n16986 , n16858 );
and ( n16988 , n16985 , n16987 );
xor ( n16989 , n16909 , n16917 );
xor ( n16990 , n16989 , n16922 );
and ( n16991 , n16987 , n16990 );
and ( n16992 , n16985 , n16990 );
or ( n16993 , n16988 , n16991 , n16992 );
buf ( n544254 , n1173 );
buf ( n16995 , n544254 );
buf ( n544256 , n1174 );
buf ( n16997 , n544256 );
and ( n16998 , n16995 , n16997 );
not ( n16999 , n16998 );
and ( n17000 , n16845 , n16999 );
not ( n17001 , n17000 );
and ( n17002 , n16096 , n16913 );
and ( n17003 , n16066 , n16911 );
nor ( n17004 , n17002 , n17003 );
xnor ( n17005 , n17004 , n16848 );
and ( n17006 , n17001 , n17005 );
and ( n17007 , n16150 , n16543 );
and ( n17008 , n16135 , n16541 );
nor ( n17009 , n17007 , n17008 );
xnor ( n17010 , n17009 , n16521 );
and ( n17011 , n17005 , n17010 );
and ( n17012 , n17001 , n17010 );
or ( n17013 , n17006 , n17011 , n17012 );
and ( n17014 , n16247 , n16450 );
and ( n17015 , n16229 , n16448 );
nor ( n17016 , n17014 , n17015 );
xnor ( n17017 , n17016 , n16395 );
and ( n17018 , n16611 , n16158 );
and ( n17019 , n16510 , n16156 );
nor ( n17020 , n17018 , n17019 );
xnor ( n17021 , n17020 , n16127 );
and ( n17022 , n17017 , n17021 );
and ( n17023 , n16725 , n16076 );
and ( n17024 , n16688 , n16074 );
nor ( n17025 , n17023 , n17024 );
xnor ( n17026 , n17025 , n16081 );
and ( n17027 , n17021 , n17026 );
and ( n17028 , n17017 , n17026 );
or ( n17029 , n17022 , n17027 , n17028 );
and ( n17030 , n17013 , n17029 );
not ( n17031 , n16916 );
and ( n17032 , n17029 , n17031 );
and ( n17033 , n17013 , n17031 );
or ( n17034 , n17030 , n17032 , n17033 );
and ( n17035 , n16105 , n16750 );
and ( n17036 , n16085 , n16748 );
nor ( n17037 , n17035 , n17036 );
xnor ( n17038 , n17037 , n16647 );
and ( n17039 , n16936 , n16093 );
and ( n17040 , n16820 , n16091 );
nor ( n17041 , n17039 , n17040 );
xnor ( n17042 , n17041 , n16101 );
and ( n17043 , n17038 , n17042 );
buf ( n544304 , n1108 );
buf ( n17045 , n544304 );
and ( n17046 , n17045 , n16087 );
and ( n17047 , n17042 , n17046 );
and ( n17048 , n17038 , n17046 );
or ( n17049 , n17043 , n17047 , n17048 );
xor ( n17050 , n16897 , n16901 );
xor ( n17051 , n17050 , n16906 );
and ( n17052 , n17049 , n17051 );
xor ( n17053 , n16929 , n16933 );
xor ( n17054 , n17053 , n16937 );
and ( n17055 , n17051 , n17054 );
and ( n17056 , n17049 , n17054 );
or ( n17057 , n17052 , n17055 , n17056 );
and ( n17058 , n17034 , n17057 );
xor ( n17059 , n16940 , n544216 );
xor ( n17060 , n17059 , n544219 );
and ( n17061 , n17057 , n17060 );
and ( n17062 , n17034 , n17060 );
or ( n17063 , n17058 , n17061 , n17062 );
and ( n17064 , n16993 , n17063 );
xor ( n17065 , n16885 , n16887 );
xor ( n17066 , n17065 , n16890 );
and ( n17067 , n17063 , n17066 );
and ( n17068 , n16993 , n17066 );
or ( n17069 , n17064 , n17067 , n17068 );
xor ( n17070 , n16864 , n16877 );
xor ( n17071 , n17070 , n16880 );
and ( n17072 , n17069 , n17071 );
xor ( n17073 , n16893 , n16968 );
xor ( n17074 , n17073 , n16971 );
and ( n17075 , n17071 , n17074 );
and ( n17076 , n17069 , n17074 );
or ( n17077 , n17072 , n17075 , n17076 );
and ( n17078 , n16983 , n17077 );
xor ( n17079 , n17069 , n17071 );
xor ( n17080 , n17079 , n17074 );
and ( n17081 , n16229 , n16543 );
and ( n17082 , n16150 , n16541 );
nor ( n17083 , n17081 , n17082 );
xnor ( n17084 , n17083 , n16521 );
and ( n17085 , n16688 , n16158 );
and ( n17086 , n16611 , n16156 );
nor ( n17087 , n17085 , n17086 );
xnor ( n17088 , n17087 , n16127 );
and ( n17089 , n17084 , n17088 );
and ( n17090 , n16820 , n16076 );
and ( n17091 , n16725 , n16074 );
nor ( n17092 , n17090 , n17091 );
xnor ( n17093 , n17092 , n16081 );
and ( n17094 , n17088 , n17093 );
and ( n17095 , n17084 , n17093 );
or ( n17096 , n17089 , n17094 , n17095 );
and ( n17097 , n16279 , n16450 );
and ( n17098 , n16247 , n16448 );
nor ( n17099 , n17097 , n17098 );
xnor ( n17100 , n17099 , n16395 );
and ( n17101 , n17045 , n16093 );
and ( n17102 , n16936 , n16091 );
nor ( n17103 , n17101 , n17102 );
xnor ( n17104 , n17103 , n16101 );
and ( n17105 , n17100 , n17104 );
buf ( n544366 , n1109 );
buf ( n17107 , n544366 );
and ( n17108 , n17107 , n16087 );
and ( n17109 , n17104 , n17108 );
and ( n17110 , n17100 , n17108 );
or ( n17111 , n17105 , n17109 , n17110 );
and ( n17112 , n17096 , n17111 );
xor ( n17113 , n16845 , n16995 );
xor ( n17114 , n16995 , n16997 );
not ( n17115 , n17114 );
and ( n17116 , n17113 , n17115 );
and ( n17117 , n16066 , n17116 );
not ( n17118 , n17117 );
xnor ( n17119 , n17118 , n17000 );
and ( n17120 , n16135 , n16750 );
and ( n17121 , n16105 , n16748 );
nor ( n17122 , n17120 , n17121 );
xnor ( n17123 , n17122 , n16647 );
and ( n17124 , n17119 , n17123 );
and ( n17125 , n16457 , n16331 );
and ( n17126 , n16365 , n16329 );
nor ( n17127 , n17125 , n17126 );
xnor ( n17128 , n17127 , n16299 );
and ( n17129 , n17123 , n17128 );
and ( n17130 , n17119 , n17128 );
or ( n17131 , n17124 , n17129 , n17130 );
and ( n17132 , n17111 , n17131 );
and ( n17133 , n17096 , n17131 );
or ( n17134 , n17112 , n17132 , n17133 );
and ( n17135 , n16085 , n16913 );
and ( n17136 , n16096 , n16911 );
nor ( n17137 , n17135 , n17136 );
xnor ( n17138 , n17137 , n16848 );
buf ( n17139 , n17138 );
and ( n17140 , n16365 , n16331 );
and ( n17141 , n16279 , n16329 );
nor ( n17142 , n17140 , n17141 );
xnor ( n17143 , n17142 , n16299 );
and ( n17144 , n17139 , n17143 );
and ( n17145 , n16472 , n16237 );
and ( n17146 , n16457 , n16235 );
nor ( n17147 , n17145 , n17146 );
xnor ( n17148 , n17147 , n16186 );
and ( n17149 , n17143 , n17148 );
and ( n17150 , n17139 , n17148 );
or ( n17151 , n17144 , n17149 , n17150 );
and ( n17152 , n17134 , n17151 );
xor ( n17153 , n16944 , n16948 );
xor ( n17154 , n17153 , n16953 );
and ( n17155 , n17151 , n17154 );
and ( n17156 , n17134 , n17154 );
or ( n17157 , n17152 , n17155 , n17156 );
xor ( n17158 , n17038 , n17042 );
xor ( n17159 , n17158 , n17046 );
xor ( n17160 , n17001 , n17005 );
xor ( n17161 , n17160 , n17010 );
and ( n17162 , n17159 , n17161 );
xor ( n17163 , n17017 , n17021 );
xor ( n17164 , n17163 , n17026 );
and ( n17165 , n17161 , n17164 );
and ( n17166 , n17159 , n17164 );
or ( n17167 , n17162 , n17165 , n17166 );
xor ( n17168 , n17013 , n17029 );
xor ( n17169 , n17168 , n17031 );
and ( n17170 , n17167 , n17169 );
xor ( n17171 , n17049 , n17051 );
xor ( n17172 , n17171 , n17054 );
and ( n17173 , n17169 , n17172 );
and ( n17174 , n17167 , n17172 );
or ( n17175 , n17170 , n17173 , n17174 );
and ( n17176 , n17157 , n17175 );
xor ( n17177 , n16985 , n16987 );
xor ( n17178 , n17177 , n16990 );
and ( n17179 , n17175 , n17178 );
and ( n17180 , n17157 , n17178 );
or ( n17181 , n17176 , n17179 , n17180 );
xor ( n17182 , n16925 , n16962 );
xor ( n17183 , n17182 , n16965 );
and ( n17184 , n17181 , n17183 );
xor ( n17185 , n16993 , n17063 );
xor ( n17186 , n17185 , n17066 );
and ( n17187 , n17183 , n17186 );
and ( n17188 , n17181 , n17186 );
or ( n17189 , n17184 , n17187 , n17188 );
and ( n17190 , n17080 , n17189 );
xor ( n17191 , n17181 , n17183 );
xor ( n17192 , n17191 , n17186 );
and ( n17193 , n16247 , n16543 );
and ( n17194 , n16229 , n16541 );
nor ( n17195 , n17193 , n17194 );
xnor ( n17196 , n17195 , n16521 );
and ( n17197 , n16611 , n16237 );
and ( n17198 , n16510 , n16235 );
nor ( n17199 , n17197 , n17198 );
xnor ( n17200 , n17199 , n16186 );
and ( n17201 , n17196 , n17200 );
and ( n17202 , n16725 , n16158 );
and ( n17203 , n16688 , n16156 );
nor ( n17204 , n17202 , n17203 );
xnor ( n17205 , n17204 , n16127 );
and ( n17206 , n17200 , n17205 );
and ( n17207 , n17196 , n17205 );
or ( n17208 , n17201 , n17206 , n17207 );
buf ( n544469 , n1175 );
buf ( n17210 , n544469 );
buf ( n544471 , n1176 );
buf ( n17212 , n544471 );
and ( n17213 , n17210 , n17212 );
not ( n17214 , n17213 );
and ( n17215 , n16997 , n17214 );
not ( n17216 , n17215 );
and ( n17217 , n16096 , n17116 );
and ( n17218 , n16066 , n17114 );
nor ( n17219 , n17217 , n17218 );
xnor ( n17220 , n17219 , n17000 );
and ( n17221 , n17216 , n17220 );
and ( n17222 , n16150 , n16750 );
and ( n17223 , n16135 , n16748 );
nor ( n17224 , n17222 , n17223 );
xnor ( n17225 , n17224 , n16647 );
and ( n17226 , n17220 , n17225 );
and ( n17227 , n17216 , n17225 );
or ( n17228 , n17221 , n17226 , n17227 );
and ( n17229 , n17208 , n17228 );
and ( n17230 , n16365 , n16450 );
and ( n17231 , n16279 , n16448 );
nor ( n17232 , n17230 , n17231 );
xnor ( n17233 , n17232 , n16395 );
and ( n17234 , n16472 , n16331 );
and ( n17235 , n16457 , n16329 );
nor ( n17236 , n17234 , n17235 );
xnor ( n17237 , n17236 , n16299 );
and ( n17238 , n17233 , n17237 );
buf ( n544499 , n1110 );
buf ( n17240 , n544499 );
and ( n17241 , n17240 , n16087 );
and ( n17242 , n17237 , n17241 );
and ( n17243 , n17233 , n17241 );
or ( n17244 , n17238 , n17242 , n17243 );
and ( n17245 , n17228 , n17244 );
and ( n17246 , n17208 , n17244 );
or ( n17247 , n17229 , n17245 , n17246 );
and ( n17248 , n16105 , n16913 );
and ( n17249 , n16085 , n16911 );
nor ( n17250 , n17248 , n17249 );
xnor ( n17251 , n17250 , n16848 );
and ( n17252 , n16936 , n16076 );
and ( n17253 , n16820 , n16074 );
nor ( n17254 , n17252 , n17253 );
xnor ( n17255 , n17254 , n16081 );
and ( n17256 , n17251 , n17255 );
and ( n17257 , n17107 , n16093 );
and ( n17258 , n17045 , n16091 );
nor ( n17259 , n17257 , n17258 );
xnor ( n17260 , n17259 , n16101 );
and ( n17261 , n17255 , n17260 );
and ( n17262 , n17251 , n17260 );
or ( n17263 , n17256 , n17261 , n17262 );
not ( n17264 , n17138 );
and ( n17265 , n17263 , n17264 );
and ( n17266 , n16510 , n16237 );
and ( n17267 , n16472 , n16235 );
nor ( n17268 , n17266 , n17267 );
xnor ( n17269 , n17268 , n16186 );
and ( n17270 , n17264 , n17269 );
and ( n17271 , n17263 , n17269 );
or ( n17272 , n17265 , n17270 , n17271 );
and ( n17273 , n17247 , n17272 );
xor ( n17274 , n17139 , n17143 );
xor ( n17275 , n17274 , n17148 );
and ( n17276 , n17272 , n17275 );
and ( n17277 , n17247 , n17275 );
or ( n17278 , n17273 , n17276 , n17277 );
xor ( n17279 , n17084 , n17088 );
xor ( n17280 , n17279 , n17093 );
xor ( n17281 , n17100 , n17104 );
xor ( n17282 , n17281 , n17108 );
and ( n17283 , n17280 , n17282 );
xor ( n17284 , n17119 , n17123 );
xor ( n17285 , n17284 , n17128 );
and ( n17286 , n17282 , n17285 );
and ( n17287 , n17280 , n17285 );
or ( n17288 , n17283 , n17286 , n17287 );
xor ( n17289 , n17096 , n17111 );
xor ( n17290 , n17289 , n17131 );
and ( n17291 , n17288 , n17290 );
xor ( n17292 , n17159 , n17161 );
xor ( n17293 , n17292 , n17164 );
and ( n17294 , n17290 , n17293 );
and ( n17295 , n17288 , n17293 );
or ( n17296 , n17291 , n17294 , n17295 );
and ( n17297 , n17278 , n17296 );
xor ( n17298 , n17134 , n17151 );
xor ( n17299 , n17298 , n17154 );
and ( n17300 , n17296 , n17299 );
and ( n17301 , n17278 , n17299 );
or ( n17302 , n17297 , n17300 , n17301 );
xor ( n17303 , n17034 , n17057 );
xor ( n17304 , n17303 , n17060 );
and ( n17305 , n17302 , n17304 );
xor ( n17306 , n17157 , n17175 );
xor ( n17307 , n17306 , n17178 );
and ( n17308 , n17304 , n17307 );
and ( n17309 , n17302 , n17307 );
or ( n17310 , n17305 , n17308 , n17309 );
and ( n17311 , n17192 , n17310 );
xor ( n17312 , n17302 , n17304 );
xor ( n17313 , n17312 , n17307 );
xor ( n17314 , n16997 , n17210 );
xor ( n17315 , n17210 , n17212 );
not ( n17316 , n17315 );
and ( n17317 , n17314 , n17316 );
and ( n17318 , n16066 , n17317 );
not ( n17319 , n17318 );
xnor ( n17320 , n17319 , n17215 );
and ( n17321 , n16135 , n16913 );
and ( n17322 , n16105 , n16911 );
nor ( n17323 , n17321 , n17322 );
xnor ( n17324 , n17323 , n16848 );
and ( n17325 , n17320 , n17324 );
buf ( n544586 , n1111 );
buf ( n17327 , n544586 );
and ( n17328 , n17327 , n16087 );
and ( n17329 , n17324 , n17328 );
and ( n17330 , n17320 , n17328 );
or ( n17331 , n17325 , n17329 , n17330 );
and ( n17332 , n16229 , n16750 );
and ( n17333 , n16150 , n16748 );
nor ( n17334 , n17332 , n17333 );
xnor ( n17335 , n17334 , n16647 );
and ( n17336 , n16688 , n16237 );
and ( n17337 , n16611 , n16235 );
nor ( n17338 , n17336 , n17337 );
xnor ( n17339 , n17338 , n16186 );
and ( n17340 , n17335 , n17339 );
and ( n17341 , n16820 , n16158 );
and ( n17342 , n16725 , n16156 );
nor ( n17343 , n17341 , n17342 );
xnor ( n17344 , n17343 , n16127 );
and ( n17345 , n17339 , n17344 );
and ( n17346 , n17335 , n17344 );
or ( n17347 , n17340 , n17345 , n17346 );
and ( n17348 , n17331 , n17347 );
and ( n17349 , n16085 , n17116 );
and ( n17350 , n16096 , n17114 );
nor ( n17351 , n17349 , n17350 );
xnor ( n17352 , n17351 , n17000 );
buf ( n17353 , n17352 );
and ( n17354 , n17347 , n17353 );
and ( n17355 , n17331 , n17353 );
or ( n17356 , n17348 , n17354 , n17355 );
xor ( n17357 , n17208 , n17228 );
xor ( n17358 , n17357 , n17244 );
and ( n17359 , n17356 , n17358 );
xor ( n17360 , n17263 , n17264 );
xor ( n17361 , n17360 , n17269 );
and ( n17362 , n17358 , n17361 );
and ( n17363 , n17356 , n17361 );
or ( n17364 , n17359 , n17362 , n17363 );
xor ( n17365 , n17247 , n17272 );
xor ( n17366 , n17365 , n17275 );
and ( n17367 , n17364 , n17366 );
xor ( n17368 , n17288 , n17290 );
xor ( n17369 , n17368 , n17293 );
and ( n17370 , n17366 , n17369 );
and ( n17371 , n17364 , n17369 );
or ( n17372 , n17367 , n17370 , n17371 );
xor ( n17373 , n17167 , n17169 );
xor ( n17374 , n17373 , n17172 );
and ( n17375 , n17372 , n17374 );
xor ( n17376 , n17278 , n17296 );
xor ( n17377 , n17376 , n17299 );
and ( n17378 , n17374 , n17377 );
and ( n17379 , n17372 , n17377 );
or ( n17380 , n17375 , n17378 , n17379 );
and ( n17381 , n17313 , n17380 );
xor ( n17382 , n17372 , n17374 );
xor ( n17383 , n17382 , n17377 );
not ( n17384 , n17352 );
and ( n17385 , n16457 , n16450 );
and ( n17386 , n16365 , n16448 );
nor ( n17387 , n17385 , n17386 );
xnor ( n17388 , n17387 , n16395 );
and ( n17389 , n17384 , n17388 );
and ( n17390 , n16510 , n16331 );
and ( n17391 , n16472 , n16329 );
nor ( n17392 , n17390 , n17391 );
xnor ( n17393 , n17392 , n16299 );
and ( n17394 , n17388 , n17393 );
and ( n17395 , n17384 , n17393 );
or ( n17396 , n17389 , n17394 , n17395 );
xor ( n17397 , n17196 , n17200 );
xor ( n17398 , n17397 , n17205 );
and ( n17399 , n17396 , n17398 );
xor ( n17400 , n17216 , n17220 );
xor ( n17401 , n17400 , n17225 );
and ( n17402 , n17398 , n17401 );
and ( n17403 , n17396 , n17401 );
or ( n17404 , n17399 , n17402 , n17403 );
and ( n17405 , n16279 , n16543 );
and ( n17406 , n16247 , n16541 );
nor ( n17407 , n17405 , n17406 );
xnor ( n17408 , n17407 , n16521 );
and ( n17409 , n17045 , n16076 );
and ( n17410 , n16936 , n16074 );
nor ( n17411 , n17409 , n17410 );
xnor ( n17412 , n17411 , n16081 );
and ( n17413 , n17408 , n17412 );
and ( n17414 , n17240 , n16093 );
and ( n17415 , n17107 , n16091 );
nor ( n17416 , n17414 , n17415 );
xnor ( n17417 , n17416 , n16101 );
and ( n17418 , n17412 , n17417 );
and ( n17419 , n17408 , n17417 );
or ( n17420 , n17413 , n17418 , n17419 );
xor ( n17421 , n17233 , n17237 );
xor ( n17422 , n17421 , n17241 );
and ( n17423 , n17420 , n17422 );
xor ( n17424 , n17251 , n17255 );
xor ( n17425 , n17424 , n17260 );
and ( n17426 , n17422 , n17425 );
and ( n17427 , n17420 , n17425 );
or ( n17428 , n17423 , n17426 , n17427 );
and ( n17429 , n17404 , n17428 );
xor ( n17430 , n17280 , n17282 );
xor ( n17431 , n17430 , n17285 );
and ( n17432 , n17428 , n17431 );
and ( n17433 , n17404 , n17431 );
or ( n17434 , n17429 , n17432 , n17433 );
and ( n17435 , n16105 , n17116 );
and ( n17436 , n16085 , n17114 );
nor ( n17437 , n17435 , n17436 );
xnor ( n17438 , n17437 , n17000 );
and ( n17439 , n16936 , n16158 );
and ( n17440 , n16820 , n16156 );
nor ( n17441 , n17439 , n17440 );
xnor ( n17442 , n17441 , n16127 );
and ( n17443 , n17438 , n17442 );
and ( n17444 , n17107 , n16076 );
and ( n17445 , n17045 , n16074 );
nor ( n17446 , n17444 , n17445 );
xnor ( n17447 , n17446 , n16081 );
and ( n17448 , n17442 , n17447 );
and ( n17449 , n17438 , n17447 );
or ( n17450 , n17443 , n17448 , n17449 );
buf ( n544711 , n1177 );
buf ( n17452 , n544711 );
buf ( n544713 , n1178 );
buf ( n17454 , n544713 );
and ( n17455 , n17452 , n17454 );
not ( n17456 , n17455 );
and ( n17457 , n17212 , n17456 );
not ( n17458 , n17457 );
and ( n17459 , n16096 , n17317 );
and ( n17460 , n16066 , n17315 );
nor ( n17461 , n17459 , n17460 );
xnor ( n17462 , n17461 , n17215 );
and ( n17463 , n17458 , n17462 );
and ( n17464 , n16150 , n16913 );
and ( n17465 , n16135 , n16911 );
nor ( n17466 , n17464 , n17465 );
xnor ( n17467 , n17466 , n16848 );
and ( n17468 , n17462 , n17467 );
and ( n17469 , n17458 , n17467 );
or ( n17470 , n17463 , n17468 , n17469 );
and ( n17471 , n17450 , n17470 );
and ( n17472 , n16365 , n16543 );
and ( n17473 , n16279 , n16541 );
nor ( n17474 , n17472 , n17473 );
xnor ( n17475 , n17474 , n16521 );
and ( n17476 , n17327 , n16093 );
and ( n17477 , n17240 , n16091 );
nor ( n17478 , n17476 , n17477 );
xnor ( n17479 , n17478 , n16101 );
and ( n17480 , n17475 , n17479 );
buf ( n544741 , n1112 );
buf ( n17482 , n544741 );
and ( n17483 , n17482 , n16087 );
and ( n17484 , n17479 , n17483 );
and ( n17485 , n17475 , n17483 );
or ( n17486 , n17480 , n17484 , n17485 );
and ( n17487 , n17470 , n17486 );
and ( n17488 , n17450 , n17486 );
or ( n17489 , n17471 , n17487 , n17488 );
and ( n17490 , n16247 , n16750 );
and ( n17491 , n16229 , n16748 );
nor ( n17492 , n17490 , n17491 );
xnor ( n17493 , n17492 , n16647 );
and ( n17494 , n16611 , n16331 );
and ( n17495 , n16510 , n16329 );
nor ( n17496 , n17494 , n17495 );
xnor ( n17497 , n17496 , n16299 );
and ( n17498 , n17493 , n17497 );
and ( n17499 , n16725 , n16237 );
and ( n17500 , n16688 , n16235 );
nor ( n17501 , n17499 , n17500 );
xnor ( n17502 , n17501 , n16186 );
and ( n17503 , n17497 , n17502 );
and ( n17504 , n17493 , n17502 );
or ( n17505 , n17498 , n17503 , n17504 );
xor ( n17506 , n17320 , n17324 );
xor ( n17507 , n17506 , n17328 );
and ( n17508 , n17505 , n17507 );
xor ( n17509 , n17335 , n17339 );
xor ( n17510 , n17509 , n17344 );
and ( n17511 , n17507 , n17510 );
and ( n17512 , n17505 , n17510 );
or ( n17513 , n17508 , n17511 , n17512 );
and ( n17514 , n17489 , n17513 );
xor ( n17515 , n17331 , n17347 );
xor ( n17516 , n17515 , n17353 );
and ( n17517 , n17513 , n17516 );
and ( n17518 , n17489 , n17516 );
or ( n17519 , n17514 , n17517 , n17518 );
and ( n17520 , n16135 , n17116 );
and ( n17521 , n16105 , n17114 );
nor ( n17522 , n17520 , n17521 );
xnor ( n17523 , n17522 , n17000 );
and ( n17524 , n16510 , n16450 );
and ( n17525 , n16472 , n16448 );
nor ( n17526 , n17524 , n17525 );
xnor ( n17527 , n17526 , n16395 );
and ( n17528 , n17523 , n17527 );
buf ( n544789 , n1113 );
buf ( n17530 , n544789 );
and ( n17531 , n17530 , n16087 );
and ( n17532 , n17527 , n17531 );
and ( n17533 , n17523 , n17531 );
or ( n17534 , n17528 , n17532 , n17533 );
and ( n17535 , n16229 , n16913 );
and ( n17536 , n16150 , n16911 );
nor ( n17537 , n17535 , n17536 );
xnor ( n17538 , n17537 , n16848 );
and ( n17539 , n16688 , n16331 );
and ( n17540 , n16611 , n16329 );
nor ( n17541 , n17539 , n17540 );
xnor ( n17542 , n17541 , n16299 );
and ( n17543 , n17538 , n17542 );
and ( n17544 , n16820 , n16237 );
and ( n17545 , n16725 , n16235 );
nor ( n17546 , n17544 , n17545 );
xnor ( n17547 , n17546 , n16186 );
and ( n17548 , n17542 , n17547 );
and ( n17549 , n17538 , n17547 );
or ( n17550 , n17543 , n17548 , n17549 );
and ( n17551 , n17534 , n17550 );
xor ( n17552 , n17212 , n17452 );
xor ( n17553 , n17452 , n17454 );
not ( n17554 , n17553 );
and ( n17555 , n17552 , n17554 );
and ( n17556 , n16066 , n17555 );
not ( n17557 , n17556 );
xnor ( n17558 , n17557 , n17457 );
and ( n17559 , n16457 , n16543 );
and ( n17560 , n16365 , n16541 );
nor ( n17561 , n17559 , n17560 );
xnor ( n17562 , n17561 , n16521 );
and ( n17563 , n17558 , n17562 );
and ( n17564 , n17482 , n16093 );
and ( n17565 , n17327 , n16091 );
nor ( n17566 , n17564 , n17565 );
xnor ( n17567 , n17566 , n16101 );
and ( n17568 , n17562 , n17567 );
and ( n17569 , n17558 , n17567 );
or ( n17570 , n17563 , n17568 , n17569 );
and ( n17571 , n17550 , n17570 );
and ( n17572 , n17534 , n17570 );
or ( n17573 , n17551 , n17571 , n17572 );
xor ( n17574 , n17408 , n17412 );
xor ( n17575 , n17574 , n17417 );
and ( n17576 , n17573 , n17575 );
xor ( n17577 , n17384 , n17388 );
xor ( n17578 , n17577 , n17393 );
and ( n17579 , n17575 , n17578 );
and ( n17580 , n17573 , n17578 );
or ( n17581 , n17576 , n17579 , n17580 );
xor ( n17582 , n17396 , n17398 );
xor ( n17583 , n17582 , n17401 );
and ( n17584 , n17581 , n17583 );
xor ( n17585 , n17420 , n17422 );
xor ( n17586 , n17585 , n17425 );
and ( n17587 , n17583 , n17586 );
and ( n17588 , n17581 , n17586 );
or ( n17589 , n17584 , n17587 , n17588 );
and ( n17590 , n17519 , n17589 );
xor ( n17591 , n17356 , n17358 );
xor ( n17592 , n17591 , n17361 );
and ( n17593 , n17589 , n17592 );
and ( n17594 , n17519 , n17592 );
or ( n17595 , n17590 , n17593 , n17594 );
and ( n17596 , n17434 , n17595 );
xor ( n17597 , n17364 , n17366 );
xor ( n17598 , n17597 , n17369 );
and ( n17599 , n17595 , n17598 );
and ( n17600 , n17434 , n17598 );
or ( n17601 , n17596 , n17599 , n17600 );
and ( n17602 , n17383 , n17601 );
xor ( n17603 , n17434 , n17595 );
xor ( n17604 , n17603 , n17598 );
and ( n17605 , n16279 , n16750 );
and ( n17606 , n16247 , n16748 );
nor ( n17607 , n17605 , n17606 );
xnor ( n17608 , n17607 , n16647 );
and ( n17609 , n17045 , n16158 );
and ( n17610 , n16936 , n16156 );
nor ( n17611 , n17609 , n17610 );
xnor ( n17612 , n17611 , n16127 );
and ( n17613 , n17608 , n17612 );
and ( n17614 , n17240 , n16076 );
and ( n17615 , n17107 , n16074 );
nor ( n17616 , n17614 , n17615 );
xnor ( n17617 , n17616 , n16081 );
and ( n17618 , n17612 , n17617 );
and ( n17619 , n17608 , n17617 );
or ( n17620 , n17613 , n17618 , n17619 );
and ( n17621 , n16085 , n17317 );
and ( n17622 , n16096 , n17315 );
nor ( n17623 , n17621 , n17622 );
xnor ( n17624 , n17623 , n17215 );
buf ( n17625 , n17624 );
and ( n17626 , n17620 , n17625 );
and ( n17627 , n16472 , n16450 );
and ( n17628 , n16457 , n16448 );
nor ( n17629 , n17627 , n17628 );
xnor ( n17630 , n17629 , n16395 );
and ( n17631 , n17625 , n17630 );
and ( n17632 , n17620 , n17630 );
or ( n17633 , n17626 , n17631 , n17632 );
xor ( n17634 , n17438 , n17442 );
xor ( n17635 , n17634 , n17447 );
xor ( n17636 , n17493 , n17497 );
xor ( n17637 , n17636 , n17502 );
and ( n17638 , n17635 , n17637 );
xor ( n17639 , n17458 , n17462 );
xor ( n17640 , n17639 , n17467 );
and ( n17641 , n17637 , n17640 );
and ( n17642 , n17635 , n17640 );
or ( n17643 , n17638 , n17641 , n17642 );
and ( n17644 , n17633 , n17643 );
xor ( n17645 , n17450 , n17470 );
xor ( n17646 , n17645 , n17486 );
and ( n17647 , n17643 , n17646 );
and ( n17648 , n17633 , n17646 );
or ( n17649 , n17644 , n17647 , n17648 );
and ( n17650 , n16247 , n16913 );
and ( n17651 , n16229 , n16911 );
nor ( n17652 , n17650 , n17651 );
xnor ( n17653 , n17652 , n16848 );
and ( n17654 , n16611 , n16450 );
and ( n17655 , n16510 , n16448 );
nor ( n17656 , n17654 , n17655 );
xnor ( n17657 , n17656 , n16395 );
and ( n17658 , n17653 , n17657 );
and ( n17659 , n16725 , n16331 );
and ( n17660 , n16688 , n16329 );
nor ( n17661 , n17659 , n17660 );
xnor ( n17662 , n17661 , n16299 );
and ( n17663 , n17657 , n17662 );
and ( n17664 , n17653 , n17662 );
or ( n17665 , n17658 , n17663 , n17664 );
and ( n17666 , n16105 , n17317 );
and ( n17667 , n16085 , n17315 );
nor ( n17668 , n17666 , n17667 );
xnor ( n17669 , n17668 , n17215 );
and ( n17670 , n16936 , n16237 );
and ( n17671 , n16820 , n16235 );
nor ( n17672 , n17670 , n17671 );
xnor ( n17673 , n17672 , n16186 );
and ( n17674 , n17669 , n17673 );
and ( n17675 , n17107 , n16158 );
and ( n17676 , n17045 , n16156 );
nor ( n17677 , n17675 , n17676 );
xnor ( n17678 , n17677 , n16127 );
and ( n17679 , n17673 , n17678 );
and ( n17680 , n17669 , n17678 );
or ( n17681 , n17674 , n17679 , n17680 );
and ( n17682 , n17665 , n17681 );
not ( n17683 , n17624 );
and ( n17684 , n17681 , n17683 );
and ( n17685 , n17665 , n17683 );
or ( n17686 , n17682 , n17684 , n17685 );
xor ( n17687 , n17475 , n17479 );
xor ( n17688 , n17687 , n17483 );
and ( n17689 , n17686 , n17688 );
xor ( n17690 , n17620 , n17625 );
xor ( n17691 , n17690 , n17630 );
and ( n17692 , n17688 , n17691 );
and ( n17693 , n17686 , n17691 );
or ( n17694 , n17689 , n17692 , n17693 );
xor ( n17695 , n17505 , n17507 );
xor ( n17696 , n17695 , n17510 );
and ( n17697 , n17694 , n17696 );
xor ( n17698 , n17573 , n17575 );
xor ( n17699 , n17698 , n17578 );
and ( n17700 , n17696 , n17699 );
and ( n17701 , n17694 , n17699 );
or ( n17702 , n17697 , n17700 , n17701 );
and ( n17703 , n17649 , n17702 );
xor ( n17704 , n17489 , n17513 );
xor ( n17705 , n17704 , n17516 );
and ( n17706 , n17702 , n17705 );
and ( n17707 , n17649 , n17705 );
or ( n17708 , n17703 , n17706 , n17707 );
xor ( n17709 , n17404 , n17428 );
xor ( n17710 , n17709 , n17431 );
and ( n17711 , n17708 , n17710 );
xor ( n17712 , n17519 , n17589 );
xor ( n17713 , n17712 , n17592 );
and ( n17714 , n17710 , n17713 );
and ( n17715 , n17708 , n17713 );
or ( n17716 , n17711 , n17714 , n17715 );
and ( n17717 , n17604 , n17716 );
xor ( n17718 , n17708 , n17710 );
xor ( n17719 , n17718 , n17713 );
buf ( n544980 , n1179 );
buf ( n17721 , n544980 );
buf ( n544982 , n1180 );
buf ( n17723 , n544982 );
and ( n17724 , n17721 , n17723 );
not ( n17725 , n17724 );
and ( n17726 , n17454 , n17725 );
not ( n17727 , n17726 );
and ( n17728 , n16096 , n17555 );
and ( n17729 , n16066 , n17553 );
nor ( n17730 , n17728 , n17729 );
xnor ( n17731 , n17730 , n17457 );
and ( n17732 , n17727 , n17731 );
and ( n17733 , n16150 , n17116 );
and ( n17734 , n16135 , n17114 );
nor ( n17735 , n17733 , n17734 );
xnor ( n17736 , n17735 , n17000 );
and ( n17737 , n17731 , n17736 );
and ( n17738 , n17727 , n17736 );
or ( n17739 , n17732 , n17737 , n17738 );
and ( n17740 , n16365 , n16750 );
and ( n17741 , n16279 , n16748 );
nor ( n17742 , n17740 , n17741 );
xnor ( n17743 , n17742 , n16647 );
and ( n17744 , n17327 , n16076 );
and ( n17745 , n17240 , n16074 );
nor ( n17746 , n17744 , n17745 );
xnor ( n17747 , n17746 , n16081 );
and ( n17748 , n17743 , n17747 );
and ( n17749 , n17530 , n16093 );
and ( n17750 , n17482 , n16091 );
nor ( n17751 , n17749 , n17750 );
xnor ( n17752 , n17751 , n16101 );
and ( n17753 , n17747 , n17752 );
and ( n17754 , n17743 , n17752 );
or ( n17755 , n17748 , n17753 , n17754 );
and ( n17756 , n17739 , n17755 );
xor ( n17757 , n17523 , n17527 );
xor ( n17758 , n17757 , n17531 );
and ( n17759 , n17755 , n17758 );
and ( n17760 , n17739 , n17758 );
or ( n17761 , n17756 , n17759 , n17760 );
xor ( n17762 , n17538 , n17542 );
xor ( n17763 , n17762 , n17547 );
xor ( n17764 , n17558 , n17562 );
xor ( n17765 , n17764 , n17567 );
and ( n17766 , n17763 , n17765 );
xor ( n17767 , n17608 , n17612 );
xor ( n17768 , n17767 , n17617 );
and ( n17769 , n17765 , n17768 );
and ( n17770 , n17763 , n17768 );
or ( n17771 , n17766 , n17769 , n17770 );
and ( n17772 , n17761 , n17771 );
xor ( n17773 , n17534 , n17550 );
xor ( n17774 , n17773 , n17570 );
and ( n17775 , n17771 , n17774 );
and ( n17776 , n17761 , n17774 );
or ( n17777 , n17772 , n17775 , n17776 );
and ( n17778 , n16229 , n17116 );
and ( n17779 , n16150 , n17114 );
nor ( n17780 , n17778 , n17779 );
xnor ( n17781 , n17780 , n17000 );
and ( n17782 , n16688 , n16450 );
and ( n17783 , n16611 , n16448 );
nor ( n17784 , n17782 , n17783 );
xnor ( n17785 , n17784 , n16395 );
and ( n17786 , n17781 , n17785 );
and ( n17787 , n16820 , n16331 );
and ( n17788 , n16725 , n16329 );
nor ( n17789 , n17787 , n17788 );
xnor ( n17790 , n17789 , n16299 );
and ( n17791 , n17785 , n17790 );
and ( n17792 , n17781 , n17790 );
or ( n17793 , n17786 , n17791 , n17792 );
xor ( n17794 , n17454 , n17721 );
xor ( n17795 , n17721 , n17723 );
not ( n17796 , n17795 );
and ( n17797 , n17794 , n17796 );
and ( n17798 , n16066 , n17797 );
not ( n17799 , n17798 );
xnor ( n17800 , n17799 , n17726 );
and ( n17801 , n16457 , n16750 );
and ( n17802 , n16365 , n16748 );
nor ( n17803 , n17801 , n17802 );
xnor ( n17804 , n17803 , n16647 );
and ( n17805 , n17800 , n17804 );
and ( n17806 , n17482 , n16076 );
and ( n17807 , n17327 , n16074 );
nor ( n17808 , n17806 , n17807 );
xnor ( n17809 , n17808 , n16081 );
and ( n17810 , n17804 , n17809 );
and ( n17811 , n17800 , n17809 );
or ( n17812 , n17805 , n17810 , n17811 );
and ( n17813 , n17793 , n17812 );
and ( n17814 , n16279 , n16913 );
and ( n17815 , n16247 , n16911 );
nor ( n17816 , n17814 , n17815 );
xnor ( n17817 , n17816 , n16848 );
and ( n17818 , n17045 , n16237 );
and ( n17819 , n16936 , n16235 );
nor ( n17820 , n17818 , n17819 );
xnor ( n17821 , n17820 , n16186 );
and ( n17822 , n17817 , n17821 );
and ( n17823 , n17240 , n16158 );
and ( n17824 , n17107 , n16156 );
nor ( n17825 , n17823 , n17824 );
xnor ( n17826 , n17825 , n16127 );
and ( n17827 , n17821 , n17826 );
and ( n17828 , n17817 , n17826 );
or ( n17829 , n17822 , n17827 , n17828 );
and ( n17830 , n17812 , n17829 );
and ( n17831 , n17793 , n17829 );
or ( n17832 , n17813 , n17830 , n17831 );
and ( n17833 , n16085 , n17555 );
and ( n17834 , n16096 , n17553 );
nor ( n17835 , n17833 , n17834 );
xnor ( n17836 , n17835 , n17457 );
buf ( n17837 , n17836 );
and ( n17838 , n16472 , n16543 );
and ( n17839 , n16457 , n16541 );
nor ( n17840 , n17838 , n17839 );
xnor ( n17841 , n17840 , n16521 );
and ( n17842 , n17837 , n17841 );
buf ( n545103 , n1114 );
buf ( n17844 , n545103 );
and ( n17845 , n17844 , n16087 );
and ( n17846 , n17841 , n17845 );
and ( n17847 , n17837 , n17845 );
or ( n17848 , n17842 , n17846 , n17847 );
and ( n17849 , n17832 , n17848 );
xor ( n17850 , n17665 , n17681 );
xor ( n17851 , n17850 , n17683 );
and ( n17852 , n17848 , n17851 );
and ( n17853 , n17832 , n17851 );
or ( n17854 , n17849 , n17852 , n17853 );
xor ( n17855 , n17635 , n17637 );
xor ( n17856 , n17855 , n17640 );
and ( n17857 , n17854 , n17856 );
xor ( n17858 , n17686 , n17688 );
xor ( n17859 , n17858 , n17691 );
and ( n17860 , n17856 , n17859 );
and ( n17861 , n17854 , n17859 );
or ( n17862 , n17857 , n17860 , n17861 );
and ( n17863 , n17777 , n17862 );
xor ( n17864 , n17633 , n17643 );
xor ( n17865 , n17864 , n17646 );
and ( n17866 , n17862 , n17865 );
and ( n17867 , n17777 , n17865 );
or ( n17868 , n17863 , n17866 , n17867 );
xor ( n17869 , n17581 , n17583 );
xor ( n17870 , n17869 , n17586 );
and ( n17871 , n17868 , n17870 );
xor ( n17872 , n17649 , n17702 );
xor ( n17873 , n17872 , n17705 );
and ( n17874 , n17870 , n17873 );
and ( n17875 , n17868 , n17873 );
or ( n17876 , n17871 , n17874 , n17875 );
and ( n17877 , n17719 , n17876 );
xor ( n17878 , n17868 , n17870 );
xor ( n17879 , n17878 , n17873 );
and ( n17880 , n16247 , n17116 );
and ( n17881 , n16229 , n17114 );
nor ( n17882 , n17880 , n17881 );
xnor ( n17883 , n17882 , n17000 );
and ( n17884 , n16611 , n16543 );
and ( n17885 , n16510 , n16541 );
nor ( n17886 , n17884 , n17885 );
xnor ( n17887 , n17886 , n16521 );
and ( n17888 , n17883 , n17887 );
and ( n17889 , n16725 , n16450 );
and ( n17890 , n16688 , n16448 );
nor ( n17891 , n17889 , n17890 );
xnor ( n17892 , n17891 , n16395 );
and ( n17893 , n17887 , n17892 );
and ( n17894 , n17883 , n17892 );
or ( n17895 , n17888 , n17893 , n17894 );
and ( n17896 , n16105 , n17555 );
and ( n17897 , n16085 , n17553 );
nor ( n17898 , n17896 , n17897 );
xnor ( n17899 , n17898 , n17457 );
and ( n17900 , n16936 , n16331 );
and ( n17901 , n16820 , n16329 );
nor ( n17902 , n17900 , n17901 );
xnor ( n17903 , n17902 , n16299 );
and ( n17904 , n17899 , n17903 );
and ( n17905 , n17107 , n16237 );
and ( n17906 , n17045 , n16235 );
nor ( n17907 , n17905 , n17906 );
xnor ( n17908 , n17907 , n16186 );
and ( n17909 , n17903 , n17908 );
and ( n17910 , n17899 , n17908 );
or ( n17911 , n17904 , n17909 , n17910 );
and ( n17912 , n17895 , n17911 );
buf ( n545173 , n1181 );
buf ( n17914 , n545173 );
buf ( n545175 , n1182 );
buf ( n17916 , n545175 );
and ( n17917 , n17914 , n17916 );
not ( n17918 , n17917 );
and ( n17919 , n17723 , n17918 );
not ( n17920 , n17919 );
and ( n17921 , n16096 , n17797 );
and ( n17922 , n16066 , n17795 );
nor ( n17923 , n17921 , n17922 );
xnor ( n17924 , n17923 , n17726 );
and ( n17925 , n17920 , n17924 );
and ( n17926 , n16150 , n17317 );
and ( n17927 , n16135 , n17315 );
nor ( n17928 , n17926 , n17927 );
xnor ( n17929 , n17928 , n17215 );
and ( n17930 , n17924 , n17929 );
and ( n17931 , n17920 , n17929 );
or ( n17932 , n17925 , n17930 , n17931 );
and ( n17933 , n17911 , n17932 );
and ( n17934 , n17895 , n17932 );
or ( n17935 , n17912 , n17933 , n17934 );
and ( n17936 , n16365 , n16913 );
and ( n17937 , n16279 , n16911 );
nor ( n17938 , n17936 , n17937 );
xnor ( n17939 , n17938 , n16848 );
and ( n17940 , n17327 , n16158 );
and ( n17941 , n17240 , n16156 );
nor ( n17942 , n17940 , n17941 );
xnor ( n17943 , n17942 , n16127 );
and ( n17944 , n17939 , n17943 );
and ( n17945 , n17530 , n16076 );
and ( n17946 , n17482 , n16074 );
nor ( n17947 , n17945 , n17946 );
xnor ( n17948 , n17947 , n16081 );
and ( n17949 , n17943 , n17948 );
and ( n17950 , n17939 , n17948 );
or ( n17951 , n17944 , n17949 , n17950 );
not ( n17952 , n17836 );
and ( n17953 , n17951 , n17952 );
and ( n17954 , n16510 , n16543 );
and ( n17955 , n16472 , n16541 );
nor ( n17956 , n17954 , n17955 );
xnor ( n17957 , n17956 , n16521 );
and ( n17958 , n17952 , n17957 );
and ( n17959 , n17951 , n17957 );
or ( n17960 , n17953 , n17958 , n17959 );
and ( n17961 , n17935 , n17960 );
xor ( n17962 , n17793 , n17812 );
xor ( n17963 , n17962 , n17829 );
and ( n17964 , n17960 , n17963 );
and ( n17965 , n17935 , n17963 );
or ( n17966 , n17961 , n17964 , n17965 );
xor ( n17967 , n17763 , n17765 );
xor ( n17968 , n17967 , n17768 );
and ( n17969 , n17966 , n17968 );
xor ( n17970 , n17832 , n17848 );
xor ( n17971 , n17970 , n17851 );
and ( n17972 , n17968 , n17971 );
and ( n17973 , n17966 , n17971 );
or ( n17974 , n17969 , n17972 , n17973 );
and ( n17975 , n16135 , n17317 );
and ( n17976 , n16105 , n17315 );
nor ( n17977 , n17975 , n17976 );
xnor ( n17978 , n17977 , n17215 );
and ( n17979 , n17844 , n16093 );
and ( n17980 , n17530 , n16091 );
nor ( n17981 , n17979 , n17980 );
xnor ( n17982 , n17981 , n16101 );
and ( n17983 , n17978 , n17982 );
buf ( n545244 , n1115 );
buf ( n17985 , n545244 );
and ( n17986 , n17985 , n16087 );
and ( n17987 , n17982 , n17986 );
and ( n17988 , n17978 , n17986 );
or ( n17989 , n17983 , n17987 , n17988 );
xor ( n17990 , n17653 , n17657 );
xor ( n17991 , n17990 , n17662 );
and ( n17992 , n17989 , n17991 );
xor ( n17993 , n17727 , n17731 );
xor ( n17994 , n17993 , n17736 );
and ( n17995 , n17991 , n17994 );
and ( n17996 , n17989 , n17994 );
or ( n17997 , n17992 , n17995 , n17996 );
xor ( n17998 , n17669 , n17673 );
xor ( n17999 , n17998 , n17678 );
xor ( n18000 , n17743 , n17747 );
xor ( n18001 , n18000 , n17752 );
and ( n18002 , n17999 , n18001 );
xor ( n18003 , n17837 , n17841 );
xor ( n18004 , n18003 , n17845 );
and ( n18005 , n18001 , n18004 );
and ( n18006 , n17999 , n18004 );
or ( n18007 , n18002 , n18005 , n18006 );
and ( n18008 , n17997 , n18007 );
xor ( n18009 , n17739 , n17755 );
xor ( n18010 , n18009 , n17758 );
and ( n18011 , n18007 , n18010 );
and ( n18012 , n17997 , n18010 );
or ( n18013 , n18008 , n18011 , n18012 );
and ( n18014 , n17974 , n18013 );
xor ( n18015 , n17761 , n17771 );
xor ( n18016 , n18015 , n17774 );
and ( n18017 , n18013 , n18016 );
and ( n18018 , n17974 , n18016 );
or ( n18019 , n18014 , n18017 , n18018 );
xor ( n18020 , n17694 , n17696 );
xor ( n18021 , n18020 , n17699 );
and ( n18022 , n18019 , n18021 );
xor ( n18023 , n17777 , n17862 );
xor ( n18024 , n18023 , n17865 );
and ( n18025 , n18021 , n18024 );
and ( n18026 , n18019 , n18024 );
or ( n18027 , n18022 , n18025 , n18026 );
and ( n18028 , n17879 , n18027 );
xor ( n18029 , n18019 , n18021 );
xor ( n18030 , n18029 , n18024 );
xor ( n18031 , n17800 , n17804 );
xor ( n18032 , n18031 , n17809 );
xor ( n18033 , n17817 , n17821 );
xor ( n18034 , n18033 , n17826 );
and ( n18035 , n18032 , n18034 );
xor ( n18036 , n17951 , n17952 );
xor ( n18037 , n18036 , n17957 );
and ( n18038 , n18034 , n18037 );
and ( n18039 , n18032 , n18037 );
or ( n18040 , n18035 , n18038 , n18039 );
and ( n18041 , n16279 , n17116 );
and ( n18042 , n16247 , n17114 );
nor ( n18043 , n18041 , n18042 );
xnor ( n18044 , n18043 , n17000 );
and ( n18045 , n16820 , n16450 );
and ( n18046 , n16725 , n16448 );
nor ( n18047 , n18045 , n18046 );
xnor ( n18048 , n18047 , n16395 );
and ( n18049 , n18044 , n18048 );
and ( n18050 , n17045 , n16331 );
and ( n18051 , n16936 , n16329 );
nor ( n18052 , n18050 , n18051 );
xnor ( n18053 , n18052 , n16299 );
and ( n18054 , n18048 , n18053 );
and ( n18055 , n18044 , n18053 );
or ( n18056 , n18049 , n18054 , n18055 );
and ( n18057 , n16085 , n17797 );
and ( n18058 , n16096 , n17795 );
nor ( n18059 , n18057 , n18058 );
xnor ( n18060 , n18059 , n17726 );
and ( n18061 , n16229 , n17317 );
and ( n18062 , n16150 , n17315 );
nor ( n18063 , n18061 , n18062 );
xnor ( n18064 , n18063 , n17215 );
and ( n18065 , n18060 , n18064 );
and ( n18066 , n16688 , n16543 );
and ( n18067 , n16611 , n16541 );
nor ( n18068 , n18066 , n18067 );
xnor ( n18069 , n18068 , n16521 );
and ( n18070 , n18064 , n18069 );
and ( n18071 , n18060 , n18069 );
or ( n18072 , n18065 , n18070 , n18071 );
and ( n18073 , n18056 , n18072 );
xor ( n18074 , n17723 , n17914 );
xor ( n18075 , n17914 , n17916 );
not ( n18076 , n18075 );
and ( n18077 , n18074 , n18076 );
and ( n18078 , n16066 , n18077 );
not ( n18079 , n18078 );
xnor ( n18080 , n18079 , n17919 );
buf ( n18081 , n18080 );
and ( n18082 , n18072 , n18081 );
and ( n18083 , n18056 , n18081 );
or ( n18084 , n18073 , n18082 , n18083 );
and ( n18085 , n16510 , n16750 );
and ( n18086 , n16472 , n16748 );
nor ( n18087 , n18085 , n18086 );
xnor ( n18088 , n18087 , n16647 );
and ( n18089 , n17482 , n16158 );
and ( n18090 , n17327 , n16156 );
nor ( n18091 , n18089 , n18090 );
xnor ( n18092 , n18091 , n16127 );
and ( n18093 , n18088 , n18092 );
and ( n18094 , n17844 , n16076 );
and ( n18095 , n17530 , n16074 );
nor ( n18096 , n18094 , n18095 );
xnor ( n18097 , n18096 , n16081 );
and ( n18098 , n18092 , n18097 );
and ( n18099 , n18088 , n18097 );
or ( n18100 , n18093 , n18098 , n18099 );
and ( n18101 , n16135 , n17555 );
and ( n18102 , n16105 , n17553 );
nor ( n18103 , n18101 , n18102 );
xnor ( n18104 , n18103 , n17457 );
and ( n18105 , n16457 , n16913 );
and ( n18106 , n16365 , n16911 );
nor ( n18107 , n18105 , n18106 );
xnor ( n18108 , n18107 , n16848 );
and ( n18109 , n18104 , n18108 );
and ( n18110 , n17240 , n16237 );
and ( n18111 , n17107 , n16235 );
nor ( n18112 , n18110 , n18111 );
xnor ( n18113 , n18112 , n16186 );
and ( n18114 , n18108 , n18113 );
and ( n18115 , n18104 , n18113 );
or ( n18116 , n18109 , n18114 , n18115 );
and ( n18117 , n18100 , n18116 );
xor ( n18118 , n17883 , n17887 );
xor ( n18119 , n18118 , n17892 );
and ( n18120 , n18116 , n18119 );
and ( n18121 , n18100 , n18119 );
or ( n18122 , n18117 , n18120 , n18121 );
and ( n18123 , n18084 , n18122 );
xor ( n18124 , n17895 , n17911 );
xor ( n18125 , n18124 , n17932 );
and ( n18126 , n18122 , n18125 );
and ( n18127 , n18084 , n18125 );
or ( n18128 , n18123 , n18126 , n18127 );
and ( n18129 , n18040 , n18128 );
xor ( n18130 , n17935 , n17960 );
xor ( n18131 , n18130 , n17963 );
and ( n18132 , n18128 , n18131 );
and ( n18133 , n18040 , n18131 );
or ( n18134 , n18129 , n18132 , n18133 );
and ( n18135 , n16472 , n16750 );
and ( n18136 , n16457 , n16748 );
nor ( n18137 , n18135 , n18136 );
xnor ( n18138 , n18137 , n16647 );
and ( n18139 , n17985 , n16093 );
and ( n18140 , n17844 , n16091 );
nor ( n18141 , n18139 , n18140 );
xnor ( n18142 , n18141 , n16101 );
and ( n18143 , n18138 , n18142 );
buf ( n545404 , n1116 );
buf ( n18145 , n545404 );
and ( n18146 , n18145 , n16087 );
and ( n18147 , n18142 , n18146 );
and ( n18148 , n18138 , n18146 );
or ( n18149 , n18143 , n18147 , n18148 );
xor ( n18150 , n17978 , n17982 );
xor ( n18151 , n18150 , n17986 );
and ( n18152 , n18149 , n18151 );
xor ( n18153 , n17781 , n17785 );
xor ( n18154 , n18153 , n17790 );
and ( n18155 , n18151 , n18154 );
and ( n18156 , n18149 , n18154 );
or ( n18157 , n18152 , n18155 , n18156 );
xor ( n18158 , n17989 , n17991 );
xor ( n18159 , n18158 , n17994 );
and ( n18160 , n18157 , n18159 );
xor ( n18161 , n17999 , n18001 );
xor ( n18162 , n18161 , n18004 );
and ( n18163 , n18159 , n18162 );
and ( n18164 , n18157 , n18162 );
or ( n18165 , n18160 , n18163 , n18164 );
and ( n18166 , n18134 , n18165 );
xor ( n18167 , n17997 , n18007 );
xor ( n18168 , n18167 , n18010 );
and ( n18169 , n18165 , n18168 );
and ( n18170 , n18134 , n18168 );
or ( n18171 , n18166 , n18169 , n18170 );
xor ( n18172 , n17854 , n17856 );
xor ( n18173 , n18172 , n17859 );
and ( n18174 , n18171 , n18173 );
xor ( n18175 , n17974 , n18013 );
xor ( n18176 , n18175 , n18016 );
and ( n18177 , n18173 , n18176 );
and ( n18178 , n18171 , n18176 );
or ( n18179 , n18174 , n18177 , n18178 );
and ( n18180 , n18030 , n18179 );
xor ( n18181 , n18171 , n18173 );
xor ( n18182 , n18181 , n18176 );
xor ( n18183 , n17920 , n17924 );
xor ( n18184 , n18183 , n17929 );
xor ( n18185 , n18138 , n18142 );
xor ( n18186 , n18185 , n18146 );
and ( n18187 , n18184 , n18186 );
xor ( n18188 , n17939 , n17943 );
xor ( n18189 , n18188 , n17948 );
and ( n18190 , n18186 , n18189 );
and ( n18191 , n18184 , n18189 );
or ( n18192 , n18187 , n18190 , n18191 );
and ( n18193 , n16611 , n16750 );
and ( n18194 , n16510 , n16748 );
nor ( n18195 , n18193 , n18194 );
xnor ( n18196 , n18195 , n16647 );
and ( n18197 , n16725 , n16543 );
and ( n18198 , n16688 , n16541 );
nor ( n18199 , n18197 , n18198 );
xnor ( n18200 , n18199 , n16521 );
and ( n18201 , n18196 , n18200 );
buf ( n545462 , n1118 );
buf ( n18203 , n545462 );
and ( n18204 , n18203 , n16087 );
and ( n18205 , n18200 , n18204 );
and ( n18206 , n18196 , n18204 );
or ( n18207 , n18201 , n18205 , n18206 );
buf ( n545468 , n1183 );
buf ( n18209 , n545468 );
buf ( n545470 , n1184 );
buf ( n18211 , n545470 );
and ( n18212 , n18209 , n18211 );
not ( n18213 , n18212 );
and ( n18214 , n17916 , n18213 );
not ( n18215 , n18214 );
and ( n18216 , n16096 , n18077 );
and ( n18217 , n16066 , n18075 );
nor ( n18218 , n18216 , n18217 );
xnor ( n18219 , n18218 , n17919 );
and ( n18220 , n18215 , n18219 );
and ( n18221 , n16150 , n17555 );
and ( n18222 , n16135 , n17553 );
nor ( n18223 , n18221 , n18222 );
xnor ( n18224 , n18223 , n17457 );
and ( n18225 , n18219 , n18224 );
and ( n18226 , n18215 , n18224 );
or ( n18227 , n18220 , n18225 , n18226 );
and ( n18228 , n18207 , n18227 );
and ( n18229 , n16247 , n17317 );
and ( n18230 , n16229 , n17315 );
nor ( n18231 , n18229 , n18230 );
xnor ( n18232 , n18231 , n17215 );
and ( n18233 , n16936 , n16450 );
and ( n18234 , n16820 , n16448 );
nor ( n18235 , n18233 , n18234 );
xnor ( n18236 , n18235 , n16395 );
and ( n18237 , n18232 , n18236 );
and ( n18238 , n17107 , n16331 );
and ( n18239 , n17045 , n16329 );
nor ( n18240 , n18238 , n18239 );
xnor ( n18241 , n18240 , n16299 );
and ( n18242 , n18236 , n18241 );
and ( n18243 , n18232 , n18241 );
or ( n18244 , n18237 , n18242 , n18243 );
and ( n18245 , n18227 , n18244 );
and ( n18246 , n18207 , n18244 );
or ( n18247 , n18228 , n18245 , n18246 );
not ( n18248 , n18080 );
and ( n18249 , n18145 , n16093 );
and ( n18250 , n17985 , n16091 );
nor ( n18251 , n18249 , n18250 );
xnor ( n18252 , n18251 , n16101 );
and ( n18253 , n18248 , n18252 );
buf ( n545514 , n1117 );
buf ( n18255 , n545514 );
and ( n18256 , n18255 , n16087 );
and ( n18257 , n18252 , n18256 );
and ( n18258 , n18248 , n18256 );
or ( n18259 , n18253 , n18257 , n18258 );
and ( n18260 , n18247 , n18259 );
xor ( n18261 , n17899 , n17903 );
xor ( n18262 , n18261 , n17908 );
and ( n18263 , n18259 , n18262 );
and ( n18264 , n18247 , n18262 );
or ( n18265 , n18260 , n18263 , n18264 );
and ( n18266 , n18192 , n18265 );
xor ( n18267 , n18149 , n18151 );
xor ( n18268 , n18267 , n18154 );
and ( n18269 , n18265 , n18268 );
and ( n18270 , n18192 , n18268 );
or ( n18271 , n18266 , n18269 , n18270 );
xor ( n18272 , n18040 , n18128 );
xor ( n18273 , n18272 , n18131 );
and ( n18274 , n18271 , n18273 );
xor ( n18275 , n18157 , n18159 );
xor ( n18276 , n18275 , n18162 );
and ( n18277 , n18273 , n18276 );
and ( n18278 , n18271 , n18276 );
or ( n18279 , n18274 , n18277 , n18278 );
xor ( n18280 , n17966 , n17968 );
xor ( n18281 , n18280 , n17971 );
and ( n18282 , n18279 , n18281 );
xor ( n18283 , n18134 , n18165 );
xor ( n18284 , n18283 , n18168 );
and ( n18285 , n18281 , n18284 );
and ( n18286 , n18279 , n18284 );
or ( n18287 , n18282 , n18285 , n18286 );
and ( n18288 , n18182 , n18287 );
xor ( n18289 , n18279 , n18281 );
xor ( n18290 , n18289 , n18284 );
and ( n18291 , n16472 , n16913 );
and ( n18292 , n16457 , n16911 );
nor ( n18293 , n18291 , n18292 );
xnor ( n18294 , n18293 , n16848 );
and ( n18295 , n17530 , n16158 );
and ( n18296 , n17482 , n16156 );
nor ( n18297 , n18295 , n18296 );
xnor ( n18298 , n18297 , n16127 );
and ( n18299 , n18294 , n18298 );
and ( n18300 , n17985 , n16076 );
and ( n18301 , n17844 , n16074 );
nor ( n18302 , n18300 , n18301 );
xnor ( n18303 , n18302 , n16081 );
and ( n18304 , n18298 , n18303 );
and ( n18305 , n18294 , n18303 );
or ( n18306 , n18299 , n18304 , n18305 );
and ( n18307 , n16105 , n17797 );
and ( n18308 , n16085 , n17795 );
nor ( n18309 , n18307 , n18308 );
xnor ( n18310 , n18309 , n17726 );
and ( n18311 , n16365 , n17116 );
and ( n18312 , n16279 , n17114 );
nor ( n18313 , n18311 , n18312 );
xnor ( n18314 , n18313 , n17000 );
and ( n18315 , n18310 , n18314 );
and ( n18316 , n17327 , n16237 );
and ( n18317 , n17240 , n16235 );
nor ( n18318 , n18316 , n18317 );
xnor ( n18319 , n18318 , n16186 );
and ( n18320 , n18314 , n18319 );
and ( n18321 , n18310 , n18319 );
or ( n18322 , n18315 , n18320 , n18321 );
and ( n18323 , n18306 , n18322 );
xor ( n18324 , n18060 , n18064 );
xor ( n18325 , n18324 , n18069 );
and ( n18326 , n18322 , n18325 );
and ( n18327 , n18306 , n18325 );
or ( n18328 , n18323 , n18326 , n18327 );
xor ( n18329 , n18056 , n18072 );
xor ( n18330 , n18329 , n18081 );
and ( n18331 , n18328 , n18330 );
xor ( n18332 , n18100 , n18116 );
xor ( n18333 , n18332 , n18119 );
and ( n18334 , n18330 , n18333 );
and ( n18335 , n18328 , n18333 );
or ( n18336 , n18331 , n18334 , n18335 );
xor ( n18337 , n18032 , n18034 );
xor ( n18338 , n18337 , n18037 );
and ( n18339 , n18336 , n18338 );
xor ( n18340 , n18084 , n18122 );
xor ( n18341 , n18340 , n18125 );
and ( n18342 , n18338 , n18341 );
and ( n18343 , n18336 , n18341 );
or ( n18344 , n18339 , n18342 , n18343 );
xor ( n18345 , n18088 , n18092 );
xor ( n18346 , n18345 , n18097 );
xor ( n18347 , n18044 , n18048 );
xor ( n18348 , n18347 , n18053 );
and ( n18349 , n18346 , n18348 );
xor ( n18350 , n18104 , n18108 );
xor ( n18351 , n18350 , n18113 );
and ( n18352 , n18348 , n18351 );
and ( n18353 , n18346 , n18351 );
or ( n18354 , n18349 , n18352 , n18353 );
xor ( n18355 , n18184 , n18186 );
xor ( n18356 , n18355 , n18189 );
and ( n18357 , n18354 , n18356 );
xor ( n18358 , n18247 , n18259 );
xor ( n18359 , n18358 , n18262 );
and ( n18360 , n18356 , n18359 );
and ( n18361 , n18354 , n18359 );
or ( n18362 , n18357 , n18360 , n18361 );
xor ( n18363 , n18192 , n18265 );
xor ( n18364 , n18363 , n18268 );
and ( n18365 , n18362 , n18364 );
xor ( n18366 , n18336 , n18338 );
xor ( n18367 , n18366 , n18341 );
and ( n18368 , n18364 , n18367 );
and ( n18369 , n18362 , n18367 );
or ( n18370 , n18365 , n18368 , n18369 );
and ( n18371 , n18344 , n18370 );
xor ( n18372 , n18271 , n18273 );
xor ( n18373 , n18372 , n18276 );
and ( n18374 , n18370 , n18373 );
and ( n18375 , n18344 , n18373 );
or ( n18376 , n18371 , n18374 , n18375 );
and ( n18377 , n18290 , n18376 );
xor ( n18378 , n18328 , n18330 );
xor ( n18379 , n18378 , n18333 );
and ( n18380 , n16510 , n16913 );
and ( n18381 , n16472 , n16911 );
nor ( n18382 , n18380 , n18381 );
xnor ( n18383 , n18382 , n16848 );
and ( n18384 , n18145 , n16076 );
and ( n18385 , n17985 , n16074 );
nor ( n18386 , n18384 , n18385 );
xnor ( n18387 , n18386 , n16081 );
and ( n18388 , n18383 , n18387 );
and ( n18389 , n18203 , n16093 );
and ( n18390 , n18255 , n16091 );
nor ( n18391 , n18389 , n18390 );
xnor ( n18392 , n18391 , n16101 );
and ( n18393 , n18387 , n18392 );
and ( n18394 , n18383 , n18392 );
or ( n18395 , n18388 , n18393 , n18394 );
xor ( n18396 , n18196 , n18200 );
xor ( n18397 , n18396 , n18204 );
and ( n18398 , n18395 , n18397 );
xor ( n18399 , n18215 , n18219 );
xor ( n18400 , n18399 , n18224 );
and ( n18401 , n18397 , n18400 );
and ( n18402 , n18395 , n18400 );
or ( n18403 , n18398 , n18401 , n18402 );
xor ( n18404 , n18207 , n18227 );
xor ( n18405 , n18404 , n18244 );
and ( n18406 , n18403 , n18405 );
xor ( n18407 , n18306 , n18322 );
xor ( n18408 , n18407 , n18325 );
and ( n18409 , n18405 , n18408 );
and ( n18410 , n18403 , n18408 );
or ( n18411 , n18406 , n18409 , n18410 );
and ( n18412 , n18379 , n18411 );
xor ( n18413 , n18294 , n18298 );
xor ( n18414 , n18413 , n18303 );
xor ( n18415 , n18232 , n18236 );
xor ( n18416 , n18415 , n18241 );
and ( n18417 , n18414 , n18416 );
xor ( n18418 , n18310 , n18314 );
xor ( n18419 , n18418 , n18319 );
and ( n18420 , n18416 , n18419 );
and ( n18421 , n18414 , n18419 );
or ( n18422 , n18417 , n18420 , n18421 );
xor ( n18423 , n18346 , n18348 );
xor ( n18424 , n18423 , n18351 );
and ( n18425 , n18422 , n18424 );
and ( n18426 , n18411 , n18425 );
and ( n18427 , n18379 , n18425 );
or ( n18428 , n18412 , n18426 , n18427 );
xor ( n18429 , n18362 , n18364 );
xor ( n18430 , n18429 , n18367 );
and ( n18431 , n18428 , n18430 );
xor ( n18432 , n18354 , n18356 );
xor ( n18433 , n18432 , n18359 );
xor ( n18434 , n18248 , n18252 );
xor ( n18435 , n18434 , n18256 );
and ( n18436 , n16135 , n17797 );
and ( n18437 , n16105 , n17795 );
nor ( n18438 , n18436 , n18437 );
xnor ( n18439 , n18438 , n17726 );
and ( n18440 , n17045 , n16450 );
and ( n18441 , n16936 , n16448 );
nor ( n18442 , n18440 , n18441 );
xnor ( n18443 , n18442 , n16395 );
and ( n18444 , n18439 , n18443 );
and ( n18445 , n17240 , n16331 );
and ( n18446 , n17107 , n16329 );
nor ( n18447 , n18445 , n18446 );
xnor ( n18448 , n18447 , n16299 );
and ( n18449 , n18443 , n18448 );
and ( n18450 , n18439 , n18448 );
or ( n18451 , n18444 , n18449 , n18450 );
and ( n18452 , n16457 , n17116 );
and ( n18453 , n16365 , n17114 );
nor ( n18454 , n18452 , n18453 );
xnor ( n18455 , n18454 , n17000 );
and ( n18456 , n17482 , n16237 );
and ( n18457 , n17327 , n16235 );
nor ( n18458 , n18456 , n18457 );
xnor ( n18459 , n18458 , n16186 );
and ( n18460 , n18455 , n18459 );
and ( n18461 , n17844 , n16158 );
and ( n18462 , n17530 , n16156 );
nor ( n18463 , n18461 , n18462 );
xnor ( n18464 , n18463 , n16127 );
and ( n18465 , n18459 , n18464 );
and ( n18466 , n18455 , n18464 );
or ( n18467 , n18460 , n18465 , n18466 );
and ( n18468 , n18451 , n18467 );
and ( n18469 , n16279 , n17317 );
and ( n18470 , n16247 , n17315 );
nor ( n18471 , n18469 , n18470 );
xnor ( n18472 , n18471 , n17215 );
and ( n18473 , n16688 , n16750 );
and ( n18474 , n16611 , n16748 );
nor ( n18475 , n18473 , n18474 );
xnor ( n18476 , n18475 , n16647 );
and ( n18477 , n18472 , n18476 );
and ( n18478 , n16820 , n16543 );
and ( n18479 , n16725 , n16541 );
nor ( n18480 , n18478 , n18479 );
xnor ( n18481 , n18480 , n16521 );
and ( n18482 , n18476 , n18481 );
and ( n18483 , n18472 , n18481 );
or ( n18484 , n18477 , n18482 , n18483 );
and ( n18485 , n18467 , n18484 );
and ( n18486 , n18451 , n18484 );
or ( n18487 , n18468 , n18485 , n18486 );
and ( n18488 , n18435 , n18487 );
xor ( n18489 , n18403 , n18405 );
xor ( n18490 , n18489 , n18408 );
and ( n18491 , n18487 , n18490 );
and ( n18492 , n18435 , n18490 );
or ( n18493 , n18488 , n18491 , n18492 );
and ( n18494 , n18433 , n18493 );
xor ( n18495 , n18422 , n18424 );
and ( n18496 , n16085 , n18077 );
and ( n18497 , n16096 , n18075 );
nor ( n18498 , n18496 , n18497 );
xnor ( n18499 , n18498 , n17919 );
and ( n18500 , n16229 , n17555 );
and ( n18501 , n16150 , n17553 );
nor ( n18502 , n18500 , n18501 );
xnor ( n18503 , n18502 , n17457 );
xor ( n18504 , n18499 , n18503 );
buf ( n545765 , n1119 );
buf ( n18506 , n545765 );
and ( n18507 , n18506 , n16087 );
xor ( n18508 , n18504 , n18507 );
xor ( n18509 , n18439 , n18443 );
xor ( n18510 , n18509 , n18448 );
and ( n18511 , n18508 , n18510 );
xor ( n18512 , n18455 , n18459 );
xor ( n18513 , n18512 , n18464 );
and ( n18514 , n18510 , n18513 );
and ( n18515 , n18508 , n18513 );
or ( n18516 , n18511 , n18514 , n18515 );
and ( n18517 , n16472 , n17116 );
and ( n18518 , n16457 , n17114 );
nor ( n18519 , n18517 , n18518 );
xnor ( n18520 , n18519 , n17000 );
and ( n18521 , n17530 , n16237 );
and ( n18522 , n17482 , n16235 );
nor ( n18523 , n18521 , n18522 );
xnor ( n18524 , n18523 , n16186 );
and ( n18525 , n18520 , n18524 );
and ( n18526 , n17985 , n16158 );
and ( n18527 , n17844 , n16156 );
nor ( n18528 , n18526 , n18527 );
xnor ( n18529 , n18528 , n16127 );
and ( n18530 , n18524 , n18529 );
and ( n18531 , n18520 , n18529 );
or ( n18532 , n18525 , n18530 , n18531 );
xor ( n18533 , n18383 , n18387 );
xor ( n18534 , n18533 , n18392 );
and ( n18535 , n18532 , n18534 );
xor ( n18536 , n18472 , n18476 );
xor ( n18537 , n18536 , n18481 );
and ( n18538 , n18534 , n18537 );
and ( n18539 , n18532 , n18537 );
or ( n18540 , n18535 , n18538 , n18539 );
and ( n18541 , n18516 , n18540 );
xor ( n18542 , n18451 , n18467 );
xor ( n18543 , n18542 , n18484 );
and ( n18544 , n18540 , n18543 );
and ( n18545 , n18516 , n18543 );
or ( n18546 , n18541 , n18544 , n18545 );
and ( n18547 , n18495 , n18546 );
xor ( n18548 , n18395 , n18397 );
xor ( n18549 , n18548 , n18400 );
xor ( n18550 , n18414 , n18416 );
xor ( n18551 , n18550 , n18419 );
and ( n18552 , n18549 , n18551 );
and ( n18553 , n18546 , n18552 );
and ( n18554 , n18495 , n18552 );
or ( n18555 , n18547 , n18553 , n18554 );
and ( n18556 , n18493 , n18555 );
and ( n18557 , n18433 , n18555 );
or ( n18558 , n18494 , n18556 , n18557 );
and ( n18559 , n18430 , n18558 );
and ( n18560 , n18428 , n18558 );
or ( n18561 , n18431 , n18559 , n18560 );
xor ( n18562 , n18344 , n18370 );
xor ( n18563 , n18562 , n18373 );
and ( n18564 , n18561 , n18563 );
xor ( n18565 , n18379 , n18411 );
xor ( n18566 , n18565 , n18425 );
xor ( n18567 , n17916 , n18209 );
xor ( n18568 , n18209 , n18211 );
not ( n18569 , n18568 );
and ( n18570 , n18567 , n18569 );
and ( n18571 , n16066 , n18570 );
not ( n18572 , n18571 );
xnor ( n18573 , n18572 , n18214 );
buf ( n18574 , n18573 );
and ( n18575 , n18255 , n16093 );
and ( n18576 , n18145 , n16091 );
nor ( n18577 , n18575 , n18576 );
xnor ( n18578 , n18577 , n16101 );
and ( n18579 , n18574 , n18578 );
and ( n18580 , n18499 , n18503 );
and ( n18581 , n18503 , n18507 );
and ( n18582 , n18499 , n18507 );
or ( n18583 , n18580 , n18581 , n18582 );
and ( n18584 , n16105 , n18077 );
and ( n18585 , n16085 , n18075 );
nor ( n18586 , n18584 , n18585 );
xnor ( n18587 , n18586 , n17919 );
and ( n18588 , n16365 , n17317 );
and ( n18589 , n16279 , n17315 );
nor ( n18590 , n18588 , n18589 );
xnor ( n18591 , n18590 , n17215 );
and ( n18592 , n18587 , n18591 );
and ( n18593 , n17327 , n16331 );
and ( n18594 , n17240 , n16329 );
nor ( n18595 , n18593 , n18594 );
xnor ( n18596 , n18595 , n16299 );
and ( n18597 , n18591 , n18596 );
and ( n18598 , n18587 , n18596 );
or ( n18599 , n18592 , n18597 , n18598 );
and ( n18600 , n16096 , n18570 );
and ( n18601 , n16066 , n18568 );
nor ( n18602 , n18600 , n18601 );
xnor ( n18603 , n18602 , n18214 );
and ( n18604 , n16150 , n17797 );
and ( n18605 , n16135 , n17795 );
nor ( n18606 , n18604 , n18605 );
xnor ( n18607 , n18606 , n17726 );
and ( n18608 , n18603 , n18607 );
and ( n18609 , n16725 , n16750 );
and ( n18610 , n16688 , n16748 );
nor ( n18611 , n18609 , n18610 );
xnor ( n18612 , n18611 , n16647 );
and ( n18613 , n18607 , n18612 );
and ( n18614 , n18603 , n18612 );
or ( n18615 , n18608 , n18613 , n18614 );
and ( n18616 , n18599 , n18615 );
and ( n18617 , n16247 , n17555 );
and ( n18618 , n16229 , n17553 );
nor ( n18619 , n18617 , n18618 );
xnor ( n18620 , n18619 , n17457 );
and ( n18621 , n16936 , n16543 );
and ( n18622 , n16820 , n16541 );
nor ( n18623 , n18621 , n18622 );
xnor ( n18624 , n18623 , n16521 );
and ( n18625 , n18620 , n18624 );
and ( n18626 , n17107 , n16450 );
and ( n18627 , n17045 , n16448 );
nor ( n18628 , n18626 , n18627 );
xnor ( n18629 , n18628 , n16395 );
and ( n18630 , n18624 , n18629 );
and ( n18631 , n18620 , n18629 );
or ( n18632 , n18625 , n18630 , n18631 );
and ( n18633 , n18615 , n18632 );
and ( n18634 , n18599 , n18632 );
or ( n18635 , n18616 , n18633 , n18634 );
and ( n18636 , n18583 , n18635 );
xor ( n18637 , n18516 , n18540 );
xor ( n18638 , n18637 , n18543 );
and ( n18639 , n18635 , n18638 );
and ( n18640 , n18583 , n18638 );
or ( n18641 , n18636 , n18639 , n18640 );
and ( n18642 , n18579 , n18641 );
xor ( n18643 , n18549 , n18551 );
and ( n18644 , n16611 , n16913 );
and ( n18645 , n16510 , n16911 );
nor ( n18646 , n18644 , n18645 );
xnor ( n18647 , n18646 , n16848 );
and ( n18648 , n18506 , n16093 );
and ( n18649 , n18203 , n16091 );
nor ( n18650 , n18648 , n18649 );
xnor ( n18651 , n18650 , n16101 );
and ( n18652 , n18647 , n18651 );
buf ( n545913 , n1120 );
buf ( n18654 , n545913 );
and ( n18655 , n18654 , n16087 );
and ( n18656 , n18651 , n18655 );
and ( n18657 , n18647 , n18655 );
or ( n18658 , n18652 , n18656 , n18657 );
not ( n18659 , n18211 );
buf ( n18660 , n18659 );
and ( n18661 , n18658 , n18660 );
not ( n18662 , n18573 );
and ( n18663 , n18660 , n18662 );
and ( n18664 , n18658 , n18662 );
or ( n18665 , n18661 , n18663 , n18664 );
and ( n18666 , n18643 , n18665 );
xor ( n18667 , n18508 , n18510 );
xor ( n18668 , n18667 , n18513 );
xor ( n18669 , n18532 , n18534 );
xor ( n18670 , n18669 , n18537 );
and ( n18671 , n18668 , n18670 );
and ( n18672 , n18665 , n18671 );
and ( n18673 , n18643 , n18671 );
or ( n18674 , n18666 , n18672 , n18673 );
and ( n18675 , n18641 , n18674 );
and ( n18676 , n18579 , n18674 );
or ( n18677 , n18642 , n18675 , n18676 );
and ( n18678 , n18566 , n18677 );
xor ( n18679 , n18433 , n18493 );
xor ( n18680 , n18679 , n18555 );
and ( n18681 , n18677 , n18680 );
and ( n18682 , n18566 , n18680 );
or ( n18683 , n18678 , n18681 , n18682 );
xor ( n18684 , n18428 , n18430 );
xor ( n18685 , n18684 , n18558 );
and ( n18686 , n18683 , n18685 );
xor ( n18687 , n18435 , n18487 );
xor ( n18688 , n18687 , n18490 );
xor ( n18689 , n18495 , n18546 );
xor ( n18690 , n18689 , n18552 );
and ( n18691 , n18688 , n18690 );
xor ( n18692 , n18599 , n18615 );
xor ( n18693 , n18692 , n18632 );
buf ( n545954 , n1185 );
buf ( n18695 , n545954 );
xor ( n18696 , n18211 , n18695 );
not ( n18697 , n18695 );
and ( n18698 , n18696 , n18697 );
and ( n18699 , n16066 , n18698 );
not ( n18700 , n18699 );
xnor ( n18701 , n18700 , n18211 );
and ( n18702 , n16085 , n18570 );
and ( n18703 , n16096 , n18568 );
nor ( n18704 , n18702 , n18703 );
xnor ( n18705 , n18704 , n18214 );
and ( n18706 , n18701 , n18705 );
buf ( n545967 , n1121 );
buf ( n18708 , n545967 );
and ( n18709 , n18708 , n16087 );
and ( n18710 , n18705 , n18709 );
and ( n18711 , n18701 , n18709 );
or ( n18712 , n18706 , n18710 , n18711 );
and ( n18713 , n18712 , n18211 );
and ( n18714 , n18255 , n16076 );
and ( n18715 , n18145 , n16074 );
nor ( n18716 , n18714 , n18715 );
xnor ( n18717 , n18716 , n16081 );
and ( n18718 , n18211 , n18717 );
and ( n18719 , n18712 , n18717 );
or ( n18720 , n18713 , n18718 , n18719 );
and ( n18721 , n18693 , n18720 );
and ( n18722 , n16279 , n17555 );
and ( n18723 , n16247 , n17553 );
nor ( n18724 , n18722 , n18723 );
xnor ( n18725 , n18724 , n17457 );
and ( n18726 , n16820 , n16750 );
and ( n18727 , n16725 , n16748 );
nor ( n18728 , n18726 , n18727 );
xnor ( n18729 , n18728 , n16647 );
and ( n18730 , n18725 , n18729 );
and ( n18731 , n17045 , n16543 );
and ( n18732 , n16936 , n16541 );
nor ( n18733 , n18731 , n18732 );
xnor ( n18734 , n18733 , n16521 );
and ( n18735 , n18729 , n18734 );
and ( n18736 , n18725 , n18734 );
or ( n18737 , n18730 , n18735 , n18736 );
and ( n18738 , n16229 , n17797 );
and ( n18739 , n16150 , n17795 );
nor ( n18740 , n18738 , n18739 );
xnor ( n18741 , n18740 , n17726 );
and ( n18742 , n16688 , n16913 );
and ( n18743 , n16611 , n16911 );
nor ( n18744 , n18742 , n18743 );
xnor ( n18745 , n18744 , n16848 );
and ( n18746 , n18741 , n18745 );
and ( n18747 , n18654 , n16093 );
and ( n18748 , n18506 , n16091 );
nor ( n18749 , n18747 , n18748 );
xnor ( n18750 , n18749 , n16101 );
and ( n18751 , n18745 , n18750 );
and ( n18752 , n18741 , n18750 );
or ( n18753 , n18746 , n18751 , n18752 );
and ( n18754 , n18737 , n18753 );
and ( n18755 , n16510 , n17116 );
and ( n18756 , n16472 , n17114 );
nor ( n18757 , n18755 , n18756 );
xnor ( n18758 , n18757 , n17000 );
and ( n18759 , n17482 , n16331 );
and ( n18760 , n17327 , n16329 );
nor ( n18761 , n18759 , n18760 );
xnor ( n18762 , n18761 , n16299 );
and ( n18763 , n18758 , n18762 );
and ( n18764 , n17844 , n16237 );
and ( n18765 , n17530 , n16235 );
nor ( n18766 , n18764 , n18765 );
xnor ( n18767 , n18766 , n16186 );
and ( n18768 , n18762 , n18767 );
and ( n18769 , n18758 , n18767 );
or ( n18770 , n18763 , n18768 , n18769 );
and ( n18771 , n18753 , n18770 );
and ( n18772 , n18737 , n18770 );
or ( n18773 , n18754 , n18771 , n18772 );
and ( n18774 , n18720 , n18773 );
and ( n18775 , n18693 , n18773 );
or ( n18776 , n18721 , n18774 , n18775 );
xor ( n18777 , n18574 , n18578 );
and ( n18778 , n18776 , n18777 );
xor ( n18779 , n18587 , n18591 );
xor ( n18780 , n18779 , n18596 );
xor ( n18781 , n18603 , n18607 );
xor ( n18782 , n18781 , n18612 );
and ( n18783 , n18780 , n18782 );
xor ( n18784 , n18620 , n18624 );
xor ( n18785 , n18784 , n18629 );
and ( n18786 , n18782 , n18785 );
and ( n18787 , n18780 , n18785 );
or ( n18788 , n18783 , n18786 , n18787 );
and ( n18789 , n16135 , n18077 );
and ( n18790 , n16105 , n18075 );
nor ( n18791 , n18789 , n18790 );
xnor ( n18792 , n18791 , n17919 );
and ( n18793 , n16457 , n17317 );
and ( n18794 , n16365 , n17315 );
nor ( n18795 , n18793 , n18794 );
xnor ( n18796 , n18795 , n17215 );
and ( n18797 , n18792 , n18796 );
and ( n18798 , n17240 , n16450 );
and ( n18799 , n17107 , n16448 );
nor ( n18800 , n18798 , n18799 );
xnor ( n18801 , n18800 , n16395 );
and ( n18802 , n18796 , n18801 );
and ( n18803 , n18792 , n18801 );
or ( n18804 , n18797 , n18802 , n18803 );
xor ( n18805 , n18520 , n18524 );
xor ( n18806 , n18805 , n18529 );
and ( n18807 , n18804 , n18806 );
xor ( n18808 , n18647 , n18651 );
xor ( n18809 , n18808 , n18655 );
and ( n18810 , n18806 , n18809 );
and ( n18811 , n18804 , n18809 );
or ( n18812 , n18807 , n18810 , n18811 );
and ( n18813 , n18788 , n18812 );
xor ( n18814 , n18658 , n18660 );
xor ( n18815 , n18814 , n18662 );
and ( n18816 , n18812 , n18815 );
and ( n18817 , n18788 , n18815 );
or ( n18818 , n18813 , n18816 , n18817 );
and ( n18819 , n18777 , n18818 );
and ( n18820 , n18776 , n18818 );
or ( n18821 , n18778 , n18819 , n18820 );
and ( n18822 , n18690 , n18821 );
and ( n18823 , n18688 , n18821 );
or ( n18824 , n18691 , n18822 , n18823 );
xor ( n18825 , n18566 , n18677 );
xor ( n18826 , n18825 , n18680 );
and ( n18827 , n18824 , n18826 );
xor ( n18828 , n18668 , n18670 );
and ( n18829 , n16096 , n18698 );
and ( n18830 , n16066 , n18695 );
nor ( n18831 , n18829 , n18830 );
xnor ( n18832 , n18831 , n18211 );
and ( n18833 , n18708 , n16091 );
not ( n18834 , n18833 );
and ( n18835 , n18834 , n16101 );
and ( n18836 , n18832 , n18835 );
and ( n18837 , n18145 , n16158 );
and ( n18838 , n17985 , n16156 );
nor ( n18839 , n18837 , n18838 );
xnor ( n18840 , n18839 , n16127 );
and ( n18841 , n18836 , n18840 );
and ( n18842 , n18203 , n16076 );
and ( n18843 , n18255 , n16074 );
nor ( n18844 , n18842 , n18843 );
xnor ( n18845 , n18844 , n16081 );
and ( n18846 , n18840 , n18845 );
and ( n18847 , n18836 , n18845 );
or ( n18848 , n18841 , n18846 , n18847 );
and ( n18849 , n16365 , n17555 );
and ( n18850 , n16279 , n17553 );
nor ( n18851 , n18849 , n18850 );
xnor ( n18852 , n18851 , n17457 );
and ( n18853 , n16725 , n16913 );
and ( n18854 , n16688 , n16911 );
nor ( n18855 , n18853 , n18854 );
xnor ( n18856 , n18855 , n16848 );
and ( n18857 , n18852 , n18856 );
and ( n18858 , n16936 , n16750 );
and ( n18859 , n16820 , n16748 );
nor ( n18860 , n18858 , n18859 );
xnor ( n18861 , n18860 , n16647 );
and ( n18862 , n18856 , n18861 );
and ( n18863 , n18852 , n18861 );
or ( n18864 , n18857 , n18862 , n18863 );
and ( n18865 , n16105 , n18570 );
and ( n18866 , n16085 , n18568 );
nor ( n18867 , n18865 , n18866 );
xnor ( n18868 , n18867 , n18214 );
and ( n18869 , n16247 , n17797 );
and ( n18870 , n16229 , n17795 );
nor ( n18871 , n18869 , n18870 );
xnor ( n18872 , n18871 , n17726 );
and ( n18873 , n18868 , n18872 );
and ( n18874 , n18708 , n16093 );
and ( n18875 , n18654 , n16091 );
nor ( n18876 , n18874 , n18875 );
xnor ( n18877 , n18876 , n16101 );
and ( n18878 , n18872 , n18877 );
and ( n18879 , n18868 , n18877 );
or ( n18880 , n18873 , n18878 , n18879 );
and ( n18881 , n18864 , n18880 );
and ( n18882 , n16150 , n18077 );
and ( n18883 , n16135 , n18075 );
nor ( n18884 , n18882 , n18883 );
xnor ( n18885 , n18884 , n17919 );
and ( n18886 , n17107 , n16543 );
and ( n18887 , n17045 , n16541 );
nor ( n18888 , n18886 , n18887 );
xnor ( n18889 , n18888 , n16521 );
and ( n18890 , n18885 , n18889 );
and ( n18891 , n17327 , n16450 );
and ( n18892 , n17240 , n16448 );
nor ( n18893 , n18891 , n18892 );
xnor ( n18894 , n18893 , n16395 );
and ( n18895 , n18889 , n18894 );
and ( n18896 , n18885 , n18894 );
or ( n18897 , n18890 , n18895 , n18896 );
and ( n18898 , n18880 , n18897 );
and ( n18899 , n18864 , n18897 );
or ( n18900 , n18881 , n18898 , n18899 );
and ( n18901 , n18848 , n18900 );
and ( n18902 , n16611 , n17116 );
and ( n18903 , n16510 , n17114 );
nor ( n18904 , n18902 , n18903 );
xnor ( n18905 , n18904 , n17000 );
and ( n18906 , n18255 , n16158 );
and ( n18907 , n18145 , n16156 );
nor ( n18908 , n18906 , n18907 );
xnor ( n18909 , n18908 , n16127 );
and ( n18910 , n18905 , n18909 );
and ( n18911 , n18506 , n16076 );
and ( n18912 , n18203 , n16074 );
nor ( n18913 , n18911 , n18912 );
xnor ( n18914 , n18913 , n16081 );
and ( n18915 , n18909 , n18914 );
and ( n18916 , n18905 , n18914 );
or ( n18917 , n18910 , n18915 , n18916 );
and ( n18918 , n16472 , n17317 );
and ( n18919 , n16457 , n17315 );
nor ( n18920 , n18918 , n18919 );
xnor ( n18921 , n18920 , n17215 );
and ( n18922 , n17530 , n16331 );
and ( n18923 , n17482 , n16329 );
nor ( n18924 , n18922 , n18923 );
xnor ( n18925 , n18924 , n16299 );
and ( n18926 , n18921 , n18925 );
and ( n18927 , n17985 , n16237 );
and ( n18928 , n17844 , n16235 );
nor ( n18929 , n18927 , n18928 );
xnor ( n18930 , n18929 , n16186 );
and ( n18931 , n18925 , n18930 );
and ( n18932 , n18921 , n18930 );
or ( n18933 , n18926 , n18931 , n18932 );
and ( n18934 , n18917 , n18933 );
xor ( n18935 , n18701 , n18705 );
xor ( n18936 , n18935 , n18709 );
and ( n18937 , n18933 , n18936 );
and ( n18938 , n18917 , n18936 );
or ( n18939 , n18934 , n18937 , n18938 );
and ( n18940 , n18900 , n18939 );
and ( n18941 , n18848 , n18939 );
or ( n18942 , n18901 , n18940 , n18941 );
and ( n18943 , n18828 , n18942 );
xor ( n18944 , n18712 , n18211 );
xor ( n18945 , n18944 , n18717 );
xor ( n18946 , n18725 , n18729 );
xor ( n18947 , n18946 , n18734 );
xor ( n18948 , n18792 , n18796 );
xor ( n18949 , n18948 , n18801 );
and ( n18950 , n18947 , n18949 );
xor ( n18951 , n18758 , n18762 );
xor ( n18952 , n18951 , n18767 );
and ( n18953 , n18949 , n18952 );
and ( n18954 , n18947 , n18952 );
or ( n18955 , n18950 , n18953 , n18954 );
and ( n18956 , n18945 , n18955 );
xor ( n18957 , n18737 , n18753 );
xor ( n18958 , n18957 , n18770 );
and ( n18959 , n18955 , n18958 );
and ( n18960 , n18945 , n18958 );
or ( n18961 , n18956 , n18959 , n18960 );
and ( n18962 , n18942 , n18961 );
and ( n18963 , n18828 , n18961 );
or ( n18964 , n18943 , n18962 , n18963 );
xor ( n18965 , n18583 , n18635 );
xor ( n18966 , n18965 , n18638 );
and ( n18967 , n18964 , n18966 );
xor ( n18968 , n18643 , n18665 );
xor ( n18969 , n18968 , n18671 );
and ( n18970 , n18966 , n18969 );
and ( n18971 , n18964 , n18969 );
or ( n18972 , n18967 , n18970 , n18971 );
xor ( n18973 , n18579 , n18641 );
xor ( n18974 , n18973 , n18674 );
and ( n18975 , n18972 , n18974 );
xor ( n18976 , n18693 , n18720 );
xor ( n18977 , n18976 , n18773 );
xor ( n18978 , n18788 , n18812 );
xor ( n18979 , n18978 , n18815 );
and ( n18980 , n18977 , n18979 );
and ( n18981 , n16229 , n18077 );
and ( n18982 , n16150 , n18075 );
nor ( n18983 , n18981 , n18982 );
xnor ( n18984 , n18983 , n17919 );
and ( n18985 , n16510 , n17317 );
and ( n18986 , n16472 , n17315 );
nor ( n18987 , n18985 , n18986 );
xnor ( n18988 , n18987 , n17215 );
and ( n18989 , n18984 , n18988 );
and ( n18990 , n17844 , n16331 );
and ( n18991 , n17530 , n16329 );
nor ( n18992 , n18990 , n18991 );
xnor ( n18993 , n18992 , n16299 );
and ( n18994 , n18988 , n18993 );
and ( n18995 , n18984 , n18993 );
or ( n18996 , n18989 , n18994 , n18995 );
and ( n18997 , n16688 , n17116 );
and ( n18998 , n16611 , n17114 );
nor ( n18999 , n18997 , n18998 );
xnor ( n19000 , n18999 , n17000 );
and ( n19001 , n18145 , n16237 );
and ( n19002 , n17985 , n16235 );
nor ( n19003 , n19001 , n19002 );
xnor ( n19004 , n19003 , n16186 );
and ( n19005 , n19000 , n19004 );
and ( n19006 , n18203 , n16158 );
and ( n19007 , n18255 , n16156 );
nor ( n19008 , n19006 , n19007 );
xnor ( n19009 , n19008 , n16127 );
and ( n19010 , n19004 , n19009 );
and ( n19011 , n19000 , n19009 );
or ( n19012 , n19005 , n19010 , n19011 );
and ( n19013 , n18996 , n19012 );
and ( n19014 , n16457 , n17555 );
and ( n19015 , n16365 , n17553 );
nor ( n19016 , n19014 , n19015 );
xnor ( n19017 , n19016 , n17457 );
and ( n19018 , n17240 , n16543 );
and ( n19019 , n17107 , n16541 );
nor ( n19020 , n19018 , n19019 );
xnor ( n19021 , n19020 , n16521 );
and ( n19022 , n19017 , n19021 );
and ( n19023 , n17482 , n16450 );
and ( n19024 , n17327 , n16448 );
nor ( n19025 , n19023 , n19024 );
xnor ( n19026 , n19025 , n16395 );
and ( n19027 , n19021 , n19026 );
and ( n19028 , n19017 , n19026 );
or ( n19029 , n19022 , n19027 , n19028 );
and ( n19030 , n19012 , n19029 );
and ( n19031 , n18996 , n19029 );
or ( n19032 , n19013 , n19030 , n19031 );
xor ( n19033 , n18741 , n18745 );
xor ( n19034 , n19033 , n18750 );
and ( n19035 , n19032 , n19034 );
xor ( n19036 , n18836 , n18840 );
xor ( n19037 , n19036 , n18845 );
and ( n19038 , n19034 , n19037 );
and ( n19039 , n19032 , n19037 );
or ( n19040 , n19035 , n19038 , n19039 );
xor ( n19041 , n18780 , n18782 );
xor ( n19042 , n19041 , n18785 );
and ( n19043 , n19040 , n19042 );
xor ( n19044 , n18804 , n18806 );
xor ( n19045 , n19044 , n18809 );
and ( n19046 , n19042 , n19045 );
and ( n19047 , n19040 , n19045 );
or ( n19048 , n19043 , n19046 , n19047 );
and ( n19049 , n18979 , n19048 );
and ( n19050 , n18977 , n19048 );
or ( n19051 , n18980 , n19049 , n19050 );
xor ( n19052 , n18776 , n18777 );
xor ( n19053 , n19052 , n18818 );
and ( n19054 , n19051 , n19053 );
xor ( n19055 , n18964 , n18966 );
xor ( n19056 , n19055 , n18969 );
and ( n19057 , n19053 , n19056 );
and ( n19058 , n19051 , n19056 );
or ( n19059 , n19054 , n19057 , n19058 );
and ( n19060 , n18974 , n19059 );
and ( n19061 , n18972 , n19059 );
or ( n19062 , n18975 , n19060 , n19061 );
and ( n19063 , n18826 , n19062 );
and ( n19064 , n18824 , n19062 );
or ( n19065 , n18827 , n19063 , n19064 );
and ( n19066 , n18685 , n19065 );
and ( n19067 , n18683 , n19065 );
or ( n19068 , n18686 , n19066 , n19067 );
and ( n19069 , n18563 , n19068 );
and ( n19070 , n18561 , n19068 );
or ( n19071 , n18564 , n19069 , n19070 );
and ( n19072 , n18376 , n19071 );
and ( n19073 , n18290 , n19071 );
or ( n19074 , n18377 , n19072 , n19073 );
and ( n19075 , n18287 , n19074 );
and ( n19076 , n18182 , n19074 );
or ( n19077 , n18288 , n19075 , n19076 );
and ( n19078 , n18179 , n19077 );
and ( n19079 , n18030 , n19077 );
or ( n19080 , n18180 , n19078 , n19079 );
and ( n19081 , n18027 , n19080 );
and ( n19082 , n17879 , n19080 );
or ( n19083 , n18028 , n19081 , n19082 );
and ( n19084 , n17876 , n19083 );
and ( n19085 , n17719 , n19083 );
or ( n19086 , n17877 , n19084 , n19085 );
and ( n19087 , n17716 , n19086 );
and ( n19088 , n17604 , n19086 );
or ( n19089 , n17717 , n19087 , n19088 );
and ( n19090 , n17601 , n19089 );
and ( n19091 , n17383 , n19089 );
or ( n19092 , n17602 , n19090 , n19091 );
and ( n19093 , n17380 , n19092 );
and ( n19094 , n17313 , n19092 );
or ( n19095 , n17381 , n19093 , n19094 );
and ( n19096 , n17310 , n19095 );
and ( n19097 , n17192 , n19095 );
or ( n19098 , n17311 , n19096 , n19097 );
and ( n19099 , n17189 , n19098 );
and ( n19100 , n17080 , n19098 );
or ( n19101 , n17190 , n19099 , n19100 );
and ( n19102 , n17077 , n19101 );
and ( n19103 , n16983 , n19101 );
or ( n19104 , n17078 , n19102 , n19103 );
and ( n19105 , n16980 , n19104 );
and ( n19106 , n16809 , n19104 );
or ( n19107 , n16981 , n19105 , n19106 );
and ( n19108 , n16806 , n19107 );
and ( n19109 , n16804 , n19107 );
or ( n19110 , n16807 , n19108 , n19109 );
and ( n19111 , n16777 , n19110 );
and ( n19112 , n16640 , n19110 );
or ( n19113 , n16778 , n19111 , n19112 );
and ( n19114 , n16637 , n19113 );
and ( n19115 , n16584 , n19113 );
or ( n19116 , n16638 , n19114 , n19115 );
and ( n19117 , n16581 , n19116 );
and ( n19118 , n16499 , n19116 );
or ( n19119 , n16582 , n19117 , n19118 );
and ( n19120 , n16496 , n19119 );
and ( n19121 , n16388 , n19119 );
or ( n19122 , n16497 , n19120 , n19121 );
and ( n19123 , n16385 , n19122 );
and ( n19124 , n16383 , n19122 );
or ( n19125 , n16386 , n19123 , n19124 );
and ( n19126 , n16326 , n19125 );
and ( n19127 , n16268 , n19125 );
or ( n19128 , n16327 , n19126 , n19127 );
and ( n19129 , n16265 , n19128 );
and ( n19130 , n16217 , n19128 );
or ( n19131 , n16266 , n19129 , n19130 );
and ( n19132 , n16214 , n19131 );
and ( n19133 , n16179 , n19131 );
or ( n19134 , n16215 , n19132 , n19133 );
xor ( n19135 , n16177 , n19134 );
xor ( n19136 , n16179 , n16214 );
xor ( n19137 , n19136 , n19131 );
xor ( n19138 , n16217 , n16265 );
xor ( n19139 , n19138 , n19128 );
xor ( n19140 , n16268 , n16326 );
xor ( n19141 , n19140 , n19125 );
xor ( n19142 , n16383 , n16385 );
xor ( n19143 , n19142 , n19122 );
xor ( n19144 , n16388 , n16496 );
xor ( n19145 , n19144 , n19119 );
xor ( n19146 , n16499 , n16581 );
xor ( n19147 , n19146 , n19116 );
xor ( n19148 , n16584 , n16637 );
xor ( n19149 , n19148 , n19113 );
xor ( n19150 , n16640 , n16777 );
xor ( n19151 , n19150 , n19110 );
xor ( n19152 , n16804 , n16806 );
xor ( n19153 , n19152 , n19107 );
xor ( n19154 , n16809 , n16980 );
xor ( n19155 , n19154 , n19104 );
xor ( n19156 , n16983 , n17077 );
xor ( n19157 , n19156 , n19101 );
xor ( n19158 , n17080 , n17189 );
xor ( n19159 , n19158 , n19098 );
xor ( n19160 , n17192 , n17310 );
xor ( n19161 , n19160 , n19095 );
xor ( n19162 , n17313 , n17380 );
xor ( n19163 , n19162 , n19092 );
xor ( n19164 , n17383 , n17601 );
xor ( n19165 , n19164 , n19089 );
xor ( n19166 , n17604 , n17716 );
xor ( n19167 , n19166 , n19086 );
xor ( n19168 , n17719 , n17876 );
xor ( n19169 , n19168 , n19083 );
xor ( n19170 , n17879 , n18027 );
xor ( n19171 , n19170 , n19080 );
xor ( n19172 , n18030 , n18179 );
xor ( n19173 , n19172 , n19077 );
xor ( n19174 , n18182 , n18287 );
xor ( n19175 , n19174 , n19074 );
xor ( n19176 , n18290 , n18376 );
xor ( n19177 , n19176 , n19071 );
xor ( n19178 , n18561 , n18563 );
xor ( n19179 , n19178 , n19068 );
xor ( n19180 , n18683 , n18685 );
xor ( n19181 , n19180 , n19065 );
xor ( n19182 , n18824 , n18826 );
xor ( n19183 , n19182 , n19062 );
xor ( n19184 , n18688 , n18690 );
xor ( n19185 , n19184 , n18821 );
xor ( n19186 , n18972 , n18974 );
xor ( n19187 , n19186 , n19059 );
and ( n19188 , n19185 , n19187 );
xor ( n19189 , n18832 , n18835 );
and ( n19190 , n16085 , n18698 );
and ( n19191 , n16096 , n18695 );
nor ( n19192 , n19190 , n19191 );
xnor ( n19193 , n19192 , n18211 );
and ( n19194 , n16135 , n18570 );
and ( n19195 , n16105 , n18568 );
nor ( n19196 , n19194 , n19195 );
xnor ( n19197 , n19196 , n18214 );
and ( n19198 , n19193 , n19197 );
and ( n19199 , n19197 , n18833 );
and ( n19200 , n19193 , n18833 );
or ( n19201 , n19198 , n19199 , n19200 );
and ( n19202 , n19189 , n19201 );
and ( n19203 , n16279 , n17797 );
and ( n19204 , n16247 , n17795 );
nor ( n19205 , n19203 , n19204 );
xnor ( n19206 , n19205 , n17726 );
and ( n19207 , n16820 , n16913 );
and ( n19208 , n16725 , n16911 );
nor ( n19209 , n19207 , n19208 );
xnor ( n19210 , n19209 , n16848 );
and ( n19211 , n19206 , n19210 );
and ( n19212 , n17045 , n16750 );
and ( n19213 , n16936 , n16748 );
nor ( n19214 , n19212 , n19213 );
xnor ( n19215 , n19214 , n16647 );
and ( n19216 , n19210 , n19215 );
and ( n19217 , n19206 , n19215 );
or ( n19218 , n19211 , n19216 , n19217 );
and ( n19219 , n19201 , n19218 );
and ( n19220 , n19189 , n19218 );
or ( n19221 , n19202 , n19219 , n19220 );
xor ( n19222 , n18905 , n18909 );
xor ( n19223 , n19222 , n18914 );
xor ( n19224 , n18852 , n18856 );
xor ( n19225 , n19224 , n18861 );
and ( n19226 , n19223 , n19225 );
xor ( n19227 , n18868 , n18872 );
xor ( n19228 , n19227 , n18877 );
and ( n19229 , n19225 , n19228 );
and ( n19230 , n19223 , n19228 );
or ( n19231 , n19226 , n19229 , n19230 );
and ( n19232 , n19221 , n19231 );
xor ( n19233 , n18917 , n18933 );
xor ( n19234 , n19233 , n18936 );
and ( n19235 , n19231 , n19234 );
and ( n19236 , n19221 , n19234 );
or ( n19237 , n19232 , n19235 , n19236 );
xor ( n19238 , n18848 , n18900 );
xor ( n19239 , n19238 , n18939 );
and ( n19240 , n19237 , n19239 );
xor ( n19241 , n18828 , n18942 );
xor ( n19242 , n19241 , n18961 );
and ( n19243 , n19240 , n19242 );
xor ( n19244 , n18945 , n18955 );
xor ( n19245 , n19244 , n18958 );
xor ( n19246 , n19040 , n19042 );
xor ( n19247 , n19246 , n19045 );
and ( n19248 , n19245 , n19247 );
xor ( n19249 , n19237 , n19239 );
and ( n19250 , n19247 , n19249 );
and ( n19251 , n19245 , n19249 );
or ( n19252 , n19248 , n19250 , n19251 );
and ( n19253 , n19242 , n19252 );
and ( n19254 , n19240 , n19252 );
or ( n19255 , n19243 , n19253 , n19254 );
xor ( n19256 , n19051 , n19053 );
xor ( n19257 , n19256 , n19056 );
and ( n19258 , n19255 , n19257 );
xor ( n19259 , n18977 , n18979 );
xor ( n19260 , n19259 , n19048 );
xor ( n19261 , n18864 , n18880 );
xor ( n19262 , n19261 , n18897 );
xor ( n19263 , n18947 , n18949 );
xor ( n19264 , n19263 , n18952 );
and ( n19265 , n19262 , n19264 );
xor ( n19266 , n19221 , n19231 );
xor ( n19267 , n19266 , n19234 );
and ( n19268 , n19264 , n19267 );
and ( n19269 , n19262 , n19267 );
or ( n19270 , n19265 , n19268 , n19269 );
and ( n19271 , n16150 , n18570 );
and ( n19272 , n16135 , n18568 );
nor ( n19273 , n19271 , n19272 );
xnor ( n19274 , n19273 , n18214 );
and ( n19275 , n16365 , n17797 );
and ( n19276 , n16279 , n17795 );
nor ( n19277 , n19275 , n19276 );
xnor ( n19278 , n19277 , n17726 );
and ( n19279 , n19274 , n19278 );
and ( n19280 , n16936 , n16913 );
and ( n19281 , n16820 , n16911 );
nor ( n19282 , n19280 , n19281 );
xnor ( n19283 , n19282 , n16848 );
and ( n19284 , n19278 , n19283 );
and ( n19285 , n19274 , n19283 );
or ( n19286 , n19279 , n19284 , n19285 );
and ( n19287 , n16105 , n18698 );
and ( n19288 , n16085 , n18695 );
nor ( n19289 , n19287 , n19288 );
xnor ( n19290 , n19289 , n18211 );
and ( n19291 , n18708 , n16074 );
not ( n19292 , n19291 );
and ( n19293 , n19292 , n16081 );
and ( n19294 , n19290 , n19293 );
and ( n19295 , n19286 , n19294 );
and ( n19296 , n18654 , n16076 );
and ( n19297 , n18506 , n16074 );
nor ( n19298 , n19296 , n19297 );
xnor ( n19299 , n19298 , n16081 );
and ( n19300 , n19294 , n19299 );
and ( n19301 , n19286 , n19299 );
or ( n19302 , n19295 , n19300 , n19301 );
xor ( n19303 , n18996 , n19012 );
xor ( n19304 , n19303 , n19029 );
and ( n19305 , n19302 , n19304 );
xor ( n19306 , n19189 , n19201 );
xor ( n19307 , n19306 , n19218 );
and ( n19308 , n19304 , n19307 );
and ( n19309 , n19302 , n19307 );
or ( n19310 , n19305 , n19308 , n19309 );
xor ( n19311 , n19193 , n19197 );
xor ( n19312 , n19311 , n18833 );
xor ( n19313 , n18984 , n18988 );
xor ( n19314 , n19313 , n18993 );
and ( n19315 , n19312 , n19314 );
xor ( n19316 , n19000 , n19004 );
xor ( n19317 , n19316 , n19009 );
and ( n19318 , n19314 , n19317 );
and ( n19319 , n19312 , n19317 );
or ( n19320 , n19315 , n19318 , n19319 );
xor ( n19321 , n19290 , n19293 );
and ( n19322 , n18506 , n16158 );
and ( n19323 , n18203 , n16156 );
nor ( n19324 , n19322 , n19323 );
xnor ( n19325 , n19324 , n16127 );
and ( n19326 , n19321 , n19325 );
and ( n19327 , n18708 , n16076 );
and ( n19328 , n18654 , n16074 );
nor ( n19329 , n19327 , n19328 );
xnor ( n19330 , n19329 , n16081 );
and ( n19331 , n19325 , n19330 );
and ( n19332 , n19321 , n19330 );
or ( n19333 , n19326 , n19331 , n19332 );
xor ( n19334 , n19206 , n19210 );
xor ( n19335 , n19334 , n19215 );
and ( n19336 , n19333 , n19335 );
xor ( n19337 , n19017 , n19021 );
xor ( n19338 , n19337 , n19026 );
and ( n19339 , n19335 , n19338 );
and ( n19340 , n19333 , n19338 );
or ( n19341 , n19336 , n19339 , n19340 );
and ( n19342 , n19320 , n19341 );
xor ( n19343 , n19223 , n19225 );
xor ( n19344 , n19343 , n19228 );
and ( n19345 , n19341 , n19344 );
and ( n19346 , n19320 , n19344 );
or ( n19347 , n19342 , n19345 , n19346 );
and ( n19348 , n19310 , n19347 );
xor ( n19349 , n19032 , n19034 );
xor ( n19350 , n19349 , n19037 );
and ( n19351 , n19347 , n19350 );
and ( n19352 , n19310 , n19350 );
or ( n19353 , n19348 , n19351 , n19352 );
and ( n19354 , n19270 , n19353 );
xor ( n19355 , n19245 , n19247 );
xor ( n19356 , n19355 , n19249 );
and ( n19357 , n19353 , n19356 );
and ( n19358 , n19270 , n19356 );
or ( n19359 , n19354 , n19357 , n19358 );
and ( n19360 , n19260 , n19359 );
xor ( n19361 , n19240 , n19242 );
xor ( n19362 , n19361 , n19252 );
and ( n19363 , n19359 , n19362 );
and ( n19364 , n19260 , n19362 );
or ( n19365 , n19360 , n19363 , n19364 );
and ( n19366 , n19257 , n19365 );
and ( n19367 , n19255 , n19365 );
or ( n19368 , n19258 , n19366 , n19367 );
and ( n19369 , n19187 , n19368 );
and ( n19370 , n19185 , n19368 );
or ( n19371 , n19188 , n19369 , n19370 );
and ( n19372 , n19183 , n19371 );
xor ( n19373 , n19183 , n19371 );
xor ( n19374 , n19185 , n19187 );
xor ( n19375 , n19374 , n19368 );
xor ( n19376 , n19255 , n19257 );
xor ( n19377 , n19376 , n19365 );
and ( n19378 , n16229 , n18570 );
and ( n19379 , n16150 , n18568 );
nor ( n19380 , n19378 , n19379 );
xnor ( n19381 , n19380 , n18214 );
and ( n19382 , n16457 , n17797 );
and ( n19383 , n16365 , n17795 );
nor ( n19384 , n19382 , n19383 );
xnor ( n19385 , n19384 , n17726 );
and ( n19386 , n19381 , n19385 );
and ( n19387 , n19385 , n19291 );
and ( n19388 , n19381 , n19291 );
or ( n19389 , n19386 , n19387 , n19388 );
and ( n19390 , n16135 , n18698 );
and ( n19391 , n16105 , n18695 );
nor ( n19392 , n19390 , n19391 );
xnor ( n19393 , n19392 , n18211 );
and ( n19394 , n17482 , n16543 );
and ( n19395 , n17327 , n16541 );
nor ( n19396 , n19394 , n19395 );
xnor ( n19397 , n19396 , n16521 );
and ( n19398 , n19393 , n19397 );
and ( n19399 , n17844 , n16450 );
and ( n19400 , n17530 , n16448 );
nor ( n19401 , n19399 , n19400 );
xnor ( n19402 , n19401 , n16395 );
and ( n19403 , n19397 , n19402 );
and ( n19404 , n19393 , n19402 );
or ( n19405 , n19398 , n19403 , n19404 );
and ( n19406 , n19389 , n19405 );
and ( n19407 , n16510 , n17555 );
and ( n19408 , n16472 , n17553 );
nor ( n19409 , n19407 , n19408 );
xnor ( n19410 , n19409 , n17457 );
and ( n19411 , n17045 , n16913 );
and ( n19412 , n16936 , n16911 );
nor ( n19413 , n19411 , n19412 );
xnor ( n19414 , n19413 , n16848 );
and ( n19415 , n19410 , n19414 );
and ( n19416 , n17240 , n16750 );
and ( n19417 , n17107 , n16748 );
nor ( n19418 , n19416 , n19417 );
xnor ( n19419 , n19418 , n16647 );
and ( n19420 , n19414 , n19419 );
and ( n19421 , n19410 , n19419 );
or ( n19422 , n19415 , n19420 , n19421 );
and ( n19423 , n19405 , n19422 );
and ( n19424 , n19389 , n19422 );
or ( n19425 , n19406 , n19423 , n19424 );
and ( n19426 , n16472 , n17555 );
and ( n19427 , n16457 , n17553 );
nor ( n19428 , n19426 , n19427 );
xnor ( n19429 , n19428 , n17457 );
and ( n19430 , n17107 , n16750 );
and ( n19431 , n17045 , n16748 );
nor ( n19432 , n19430 , n19431 );
xnor ( n19433 , n19432 , n16647 );
xor ( n19434 , n19429 , n19433 );
and ( n19435 , n17327 , n16543 );
and ( n19436 , n17240 , n16541 );
nor ( n19437 , n19435 , n19436 );
xnor ( n19438 , n19437 , n16521 );
xor ( n19439 , n19434 , n19438 );
and ( n19440 , n16725 , n17116 );
and ( n19441 , n16688 , n17114 );
nor ( n19442 , n19440 , n19441 );
xnor ( n19443 , n19442 , n17000 );
and ( n19444 , n17985 , n16331 );
and ( n19445 , n17844 , n16329 );
nor ( n19446 , n19444 , n19445 );
xnor ( n19447 , n19446 , n16299 );
xor ( n19448 , n19443 , n19447 );
and ( n19449 , n18255 , n16237 );
and ( n19450 , n18145 , n16235 );
nor ( n19451 , n19449 , n19450 );
xnor ( n19452 , n19451 , n16186 );
xor ( n19453 , n19448 , n19452 );
and ( n19454 , n19439 , n19453 );
and ( n19455 , n16247 , n18077 );
and ( n19456 , n16229 , n18075 );
nor ( n19457 , n19455 , n19456 );
xnor ( n19458 , n19457 , n17919 );
and ( n19459 , n16611 , n17317 );
and ( n19460 , n16510 , n17315 );
nor ( n19461 , n19459 , n19460 );
xnor ( n19462 , n19461 , n17215 );
xor ( n19463 , n19458 , n19462 );
and ( n19464 , n17530 , n16450 );
and ( n19465 , n17482 , n16448 );
nor ( n19466 , n19464 , n19465 );
xnor ( n19467 , n19466 , n16395 );
xor ( n19468 , n19463 , n19467 );
and ( n19469 , n19453 , n19468 );
and ( n19470 , n19439 , n19468 );
or ( n19471 , n19454 , n19469 , n19470 );
and ( n19472 , n19425 , n19471 );
xor ( n19473 , n19286 , n19294 );
xor ( n19474 , n19473 , n19299 );
and ( n19475 , n19471 , n19474 );
and ( n19476 , n19425 , n19474 );
or ( n19477 , n19472 , n19475 , n19476 );
and ( n19478 , n16279 , n18077 );
and ( n19479 , n16247 , n18075 );
nor ( n19480 , n19478 , n19479 );
xnor ( n19481 , n19480 , n17919 );
and ( n19482 , n16820 , n17116 );
and ( n19483 , n16725 , n17114 );
nor ( n19484 , n19482 , n19483 );
xnor ( n19485 , n19484 , n17000 );
and ( n19486 , n19481 , n19485 );
and ( n19487 , n18654 , n16158 );
and ( n19488 , n18506 , n16156 );
nor ( n19489 , n19487 , n19488 );
xnor ( n19490 , n19489 , n16127 );
and ( n19491 , n19485 , n19490 );
and ( n19492 , n19481 , n19490 );
or ( n19493 , n19486 , n19491 , n19492 );
and ( n19494 , n16688 , n17317 );
and ( n19495 , n16611 , n17315 );
nor ( n19496 , n19494 , n19495 );
xnor ( n19497 , n19496 , n17215 );
and ( n19498 , n18145 , n16331 );
and ( n19499 , n17985 , n16329 );
nor ( n19500 , n19498 , n19499 );
xnor ( n19501 , n19500 , n16299 );
and ( n19502 , n19497 , n19501 );
and ( n19503 , n18203 , n16237 );
and ( n19504 , n18255 , n16235 );
nor ( n19505 , n19503 , n19504 );
xnor ( n19506 , n19505 , n16186 );
and ( n19507 , n19501 , n19506 );
and ( n19508 , n19497 , n19506 );
or ( n19509 , n19502 , n19507 , n19508 );
and ( n19510 , n19493 , n19509 );
xor ( n19511 , n19274 , n19278 );
xor ( n19512 , n19511 , n19283 );
and ( n19513 , n19509 , n19512 );
and ( n19514 , n19493 , n19512 );
or ( n19515 , n19510 , n19513 , n19514 );
and ( n19516 , n19429 , n19433 );
and ( n19517 , n19433 , n19438 );
and ( n19518 , n19429 , n19438 );
or ( n19519 , n19516 , n19517 , n19518 );
and ( n19520 , n19443 , n19447 );
and ( n19521 , n19447 , n19452 );
and ( n19522 , n19443 , n19452 );
or ( n19523 , n19520 , n19521 , n19522 );
xor ( n19524 , n19519 , n19523 );
and ( n19525 , n19458 , n19462 );
and ( n19526 , n19462 , n19467 );
and ( n19527 , n19458 , n19467 );
or ( n19528 , n19525 , n19526 , n19527 );
xor ( n19529 , n19524 , n19528 );
and ( n19530 , n19515 , n19529 );
xor ( n19531 , n19333 , n19335 );
xor ( n19532 , n19531 , n19338 );
and ( n19533 , n19529 , n19532 );
and ( n19534 , n19515 , n19532 );
or ( n19535 , n19530 , n19533 , n19534 );
and ( n19536 , n19477 , n19535 );
and ( n19537 , n19519 , n19523 );
and ( n19538 , n19523 , n19528 );
and ( n19539 , n19519 , n19528 );
or ( n19540 , n19537 , n19538 , n19539 );
xor ( n19541 , n18885 , n18889 );
xor ( n19542 , n19541 , n18894 );
xor ( n19543 , n19540 , n19542 );
xor ( n19544 , n18921 , n18925 );
xor ( n19545 , n19544 , n18930 );
xor ( n19546 , n19543 , n19545 );
and ( n19547 , n19535 , n19546 );
and ( n19548 , n19477 , n19546 );
or ( n19549 , n19536 , n19547 , n19548 );
and ( n19550 , n16472 , n17797 );
and ( n19551 , n16457 , n17795 );
nor ( n19552 , n19550 , n19551 );
xnor ( n19553 , n19552 , n17726 );
and ( n19554 , n17107 , n16913 );
and ( n19555 , n17045 , n16911 );
nor ( n19556 , n19554 , n19555 );
xnor ( n19557 , n19556 , n16848 );
and ( n19558 , n19553 , n19557 );
and ( n19559 , n17327 , n16750 );
and ( n19560 , n17240 , n16748 );
nor ( n19561 , n19559 , n19560 );
xnor ( n19562 , n19561 , n16647 );
and ( n19563 , n19557 , n19562 );
and ( n19564 , n19553 , n19562 );
or ( n19565 , n19558 , n19563 , n19564 );
and ( n19566 , n16611 , n17555 );
and ( n19567 , n16510 , n17553 );
nor ( n19568 , n19566 , n19567 );
xnor ( n19569 , n19568 , n17457 );
and ( n19570 , n17530 , n16543 );
and ( n19571 , n17482 , n16541 );
nor ( n19572 , n19570 , n19571 );
xnor ( n19573 , n19572 , n16521 );
and ( n19574 , n19569 , n19573 );
and ( n19575 , n17985 , n16450 );
and ( n19576 , n17844 , n16448 );
nor ( n19577 , n19575 , n19576 );
xnor ( n19578 , n19577 , n16395 );
and ( n19579 , n19573 , n19578 );
and ( n19580 , n19569 , n19578 );
or ( n19581 , n19574 , n19579 , n19580 );
and ( n19582 , n19565 , n19581 );
and ( n19583 , n16247 , n18570 );
and ( n19584 , n16229 , n18568 );
nor ( n19585 , n19583 , n19584 );
xnor ( n19586 , n19585 , n18214 );
and ( n19587 , n18708 , n16156 );
not ( n19588 , n19587 );
and ( n19589 , n19588 , n16127 );
and ( n19590 , n19586 , n19589 );
and ( n19591 , n19581 , n19590 );
and ( n19592 , n19565 , n19590 );
or ( n19593 , n19582 , n19591 , n19592 );
xor ( n19594 , n19381 , n19385 );
xor ( n19595 , n19594 , n19291 );
xor ( n19596 , n19481 , n19485 );
xor ( n19597 , n19596 , n19490 );
and ( n19598 , n19595 , n19597 );
xor ( n19599 , n19393 , n19397 );
xor ( n19600 , n19599 , n19402 );
and ( n19601 , n19597 , n19600 );
and ( n19602 , n19595 , n19600 );
or ( n19603 , n19598 , n19601 , n19602 );
and ( n19604 , n19593 , n19603 );
xor ( n19605 , n19321 , n19325 );
xor ( n19606 , n19605 , n19330 );
and ( n19607 , n19603 , n19606 );
and ( n19608 , n19593 , n19606 );
or ( n19609 , n19604 , n19607 , n19608 );
and ( n19610 , n16365 , n18077 );
and ( n19611 , n16279 , n18075 );
nor ( n19612 , n19610 , n19611 );
xnor ( n19613 , n19612 , n17919 );
and ( n19614 , n18506 , n16237 );
and ( n19615 , n18203 , n16235 );
nor ( n19616 , n19614 , n19615 );
xnor ( n19617 , n19616 , n16186 );
and ( n19618 , n19613 , n19617 );
and ( n19619 , n18708 , n16158 );
and ( n19620 , n18654 , n16156 );
nor ( n19621 , n19619 , n19620 );
xnor ( n19622 , n19621 , n16127 );
and ( n19623 , n19617 , n19622 );
and ( n19624 , n19613 , n19622 );
or ( n19625 , n19618 , n19623 , n19624 );
and ( n19626 , n16150 , n18698 );
and ( n19627 , n16135 , n18695 );
nor ( n19628 , n19626 , n19627 );
xnor ( n19629 , n19628 , n18211 );
and ( n19630 , n16725 , n17317 );
and ( n19631 , n16688 , n17315 );
nor ( n19632 , n19630 , n19631 );
xnor ( n19633 , n19632 , n17215 );
and ( n19634 , n19629 , n19633 );
and ( n19635 , n18255 , n16331 );
and ( n19636 , n18145 , n16329 );
nor ( n19637 , n19635 , n19636 );
xnor ( n19638 , n19637 , n16299 );
and ( n19639 , n19633 , n19638 );
and ( n19640 , n19629 , n19638 );
or ( n19641 , n19634 , n19639 , n19640 );
and ( n19642 , n19625 , n19641 );
xor ( n19643 , n19410 , n19414 );
xor ( n19644 , n19643 , n19419 );
and ( n19645 , n19641 , n19644 );
and ( n19646 , n19625 , n19644 );
or ( n19647 , n19642 , n19645 , n19646 );
xor ( n19648 , n19389 , n19405 );
xor ( n19649 , n19648 , n19422 );
and ( n19650 , n19647 , n19649 );
xor ( n19651 , n19493 , n19509 );
xor ( n19652 , n19651 , n19512 );
and ( n19653 , n19649 , n19652 );
and ( n19654 , n19647 , n19652 );
or ( n19655 , n19650 , n19653 , n19654 );
and ( n19656 , n19609 , n19655 );
xor ( n19657 , n19312 , n19314 );
xor ( n19658 , n19657 , n19317 );
and ( n19659 , n19655 , n19658 );
and ( n19660 , n19609 , n19658 );
or ( n19661 , n19656 , n19659 , n19660 );
xor ( n19662 , n19302 , n19304 );
xor ( n19663 , n19662 , n19307 );
and ( n19664 , n19661 , n19663 );
xor ( n19665 , n19320 , n19341 );
xor ( n19666 , n19665 , n19344 );
and ( n19667 , n19663 , n19666 );
and ( n19668 , n19661 , n19666 );
or ( n19669 , n19664 , n19667 , n19668 );
and ( n19670 , n19549 , n19669 );
and ( n19671 , n19540 , n19542 );
and ( n19672 , n19542 , n19545 );
and ( n19673 , n19540 , n19545 );
or ( n19674 , n19671 , n19672 , n19673 );
xor ( n19675 , n19262 , n19264 );
xor ( n19676 , n19675 , n19267 );
and ( n19677 , n19674 , n19676 );
xor ( n19678 , n19310 , n19347 );
xor ( n19679 , n19678 , n19350 );
and ( n19680 , n19676 , n19679 );
and ( n19681 , n19674 , n19679 );
or ( n19682 , n19677 , n19680 , n19681 );
and ( n19683 , n19670 , n19682 );
xor ( n19684 , n19270 , n19353 );
xor ( n19685 , n19684 , n19356 );
and ( n19686 , n19682 , n19685 );
and ( n19687 , n19670 , n19685 );
or ( n19688 , n19683 , n19686 , n19687 );
xor ( n19689 , n19260 , n19359 );
xor ( n19690 , n19689 , n19362 );
and ( n19691 , n19688 , n19690 );
xor ( n19692 , n19688 , n19690 );
xor ( n19693 , n19549 , n19669 );
and ( n19694 , n16820 , n17317 );
and ( n19695 , n16725 , n17315 );
nor ( n19696 , n19694 , n19695 );
xnor ( n19697 , n19696 , n17215 );
and ( n19698 , n18203 , n16331 );
and ( n19699 , n18255 , n16329 );
nor ( n19700 , n19698 , n19699 );
xnor ( n19701 , n19700 , n16299 );
and ( n19702 , n19697 , n19701 );
and ( n19703 , n18654 , n16237 );
and ( n19704 , n18506 , n16235 );
nor ( n19705 , n19703 , n19704 );
xnor ( n19706 , n19705 , n16186 );
and ( n19707 , n19701 , n19706 );
and ( n19708 , n19697 , n19706 );
or ( n19709 , n19702 , n19707 , n19708 );
and ( n19710 , n16688 , n17555 );
and ( n19711 , n16611 , n17553 );
nor ( n19712 , n19710 , n19711 );
xnor ( n19713 , n19712 , n17457 );
and ( n19714 , n17240 , n16913 );
and ( n19715 , n17107 , n16911 );
nor ( n19716 , n19714 , n19715 );
xnor ( n19717 , n19716 , n16848 );
and ( n19718 , n19713 , n19717 );
and ( n19719 , n17482 , n16750 );
and ( n19720 , n17327 , n16748 );
nor ( n19721 , n19719 , n19720 );
xnor ( n19722 , n19721 , n16647 );
and ( n19723 , n19717 , n19722 );
and ( n19724 , n19713 , n19722 );
or ( n19725 , n19718 , n19723 , n19724 );
and ( n19726 , n19709 , n19725 );
and ( n19727 , n16229 , n18698 );
and ( n19728 , n16150 , n18695 );
nor ( n19729 , n19727 , n19728 );
xnor ( n19730 , n19729 , n18211 );
and ( n19731 , n17844 , n16543 );
and ( n19732 , n17530 , n16541 );
nor ( n19733 , n19731 , n19732 );
xnor ( n19734 , n19733 , n16521 );
and ( n19735 , n19730 , n19734 );
and ( n19736 , n18145 , n16450 );
and ( n19737 , n17985 , n16448 );
nor ( n19738 , n19736 , n19737 );
xnor ( n19739 , n19738 , n16395 );
and ( n19740 , n19734 , n19739 );
and ( n19741 , n19730 , n19739 );
or ( n19742 , n19735 , n19740 , n19741 );
and ( n19743 , n19725 , n19742 );
and ( n19744 , n19709 , n19742 );
or ( n19745 , n19726 , n19743 , n19744 );
xor ( n19746 , n19586 , n19589 );
and ( n19747 , n16279 , n18570 );
and ( n19748 , n16247 , n18568 );
nor ( n19749 , n19747 , n19748 );
xnor ( n19750 , n19749 , n18214 );
and ( n19751 , n16510 , n17797 );
and ( n19752 , n16472 , n17795 );
nor ( n19753 , n19751 , n19752 );
xnor ( n19754 , n19753 , n17726 );
and ( n19755 , n19750 , n19754 );
and ( n19756 , n19754 , n19587 );
and ( n19757 , n19750 , n19587 );
or ( n19758 , n19755 , n19756 , n19757 );
and ( n19759 , n19746 , n19758 );
and ( n19760 , n16936 , n17116 );
and ( n19761 , n16820 , n17114 );
nor ( n19762 , n19760 , n19761 );
xnor ( n19763 , n19762 , n17000 );
and ( n19764 , n19758 , n19763 );
and ( n19765 , n19746 , n19763 );
or ( n19766 , n19759 , n19764 , n19765 );
and ( n19767 , n19745 , n19766 );
xor ( n19768 , n19497 , n19501 );
xor ( n19769 , n19768 , n19506 );
and ( n19770 , n19766 , n19769 );
and ( n19771 , n19745 , n19769 );
or ( n19772 , n19767 , n19770 , n19771 );
xor ( n19773 , n19613 , n19617 );
xor ( n19774 , n19773 , n19622 );
xor ( n19775 , n19553 , n19557 );
xor ( n19776 , n19775 , n19562 );
and ( n19777 , n19774 , n19776 );
xor ( n19778 , n19629 , n19633 );
xor ( n19779 , n19778 , n19638 );
and ( n19780 , n19776 , n19779 );
and ( n19781 , n19774 , n19779 );
or ( n19782 , n19777 , n19780 , n19781 );
xor ( n19783 , n19565 , n19581 );
xor ( n19784 , n19783 , n19590 );
and ( n19785 , n19782 , n19784 );
xor ( n19786 , n19625 , n19641 );
xor ( n19787 , n19786 , n19644 );
and ( n19788 , n19784 , n19787 );
and ( n19789 , n19782 , n19787 );
or ( n19790 , n19785 , n19788 , n19789 );
and ( n19791 , n19772 , n19790 );
xor ( n19792 , n19439 , n19453 );
xor ( n19793 , n19792 , n19468 );
and ( n19794 , n19790 , n19793 );
and ( n19795 , n19772 , n19793 );
or ( n19796 , n19791 , n19794 , n19795 );
xor ( n19797 , n19425 , n19471 );
xor ( n19798 , n19797 , n19474 );
and ( n19799 , n19796 , n19798 );
xor ( n19800 , n19515 , n19529 );
xor ( n19801 , n19800 , n19532 );
and ( n19802 , n19798 , n19801 );
and ( n19803 , n19796 , n19801 );
or ( n19804 , n19799 , n19802 , n19803 );
xor ( n19805 , n19477 , n19535 );
xor ( n19806 , n19805 , n19546 );
and ( n19807 , n19804 , n19806 );
xor ( n19808 , n19661 , n19663 );
xor ( n19809 , n19808 , n19666 );
and ( n19810 , n19806 , n19809 );
and ( n19811 , n19804 , n19809 );
or ( n19812 , n19807 , n19810 , n19811 );
and ( n19813 , n19693 , n19812 );
xor ( n19814 , n19674 , n19676 );
xor ( n19815 , n19814 , n19679 );
and ( n19816 , n19812 , n19815 );
and ( n19817 , n19693 , n19815 );
or ( n19818 , n19813 , n19816 , n19817 );
xor ( n19819 , n19670 , n19682 );
xor ( n19820 , n19819 , n19685 );
and ( n19821 , n19818 , n19820 );
xor ( n19822 , n19818 , n19820 );
xor ( n19823 , n19693 , n19812 );
xor ( n19824 , n19823 , n19815 );
xor ( n19825 , n19804 , n19806 );
xor ( n19826 , n19825 , n19809 );
xor ( n19827 , n19593 , n19603 );
xor ( n19828 , n19827 , n19606 );
xor ( n19829 , n19647 , n19649 );
xor ( n19830 , n19829 , n19652 );
and ( n19831 , n19828 , n19830 );
xor ( n19832 , n19772 , n19790 );
xor ( n19833 , n19832 , n19793 );
and ( n19834 , n19830 , n19833 );
and ( n19835 , n19828 , n19833 );
or ( n19836 , n19831 , n19834 , n19835 );
xor ( n19837 , n19609 , n19655 );
xor ( n19838 , n19837 , n19658 );
and ( n19839 , n19836 , n19838 );
xor ( n19840 , n19796 , n19798 );
xor ( n19841 , n19840 , n19801 );
and ( n19842 , n19838 , n19841 );
and ( n19843 , n19836 , n19841 );
or ( n19844 , n19839 , n19842 , n19843 );
and ( n19845 , n19826 , n19844 );
xor ( n19846 , n19836 , n19838 );
xor ( n19847 , n19846 , n19841 );
and ( n19848 , n16365 , n18570 );
and ( n19849 , n16279 , n18568 );
nor ( n19850 , n19848 , n19849 );
xnor ( n19851 , n19850 , n18214 );
and ( n19852 , n18708 , n16235 );
not ( n19853 , n19852 );
and ( n19854 , n19853 , n16186 );
and ( n19855 , n19851 , n19854 );
and ( n19856 , n16457 , n18077 );
and ( n19857 , n16365 , n18075 );
nor ( n19858 , n19856 , n19857 );
xnor ( n19859 , n19858 , n17919 );
and ( n19860 , n19855 , n19859 );
and ( n19861 , n17045 , n17116 );
and ( n19862 , n16936 , n17114 );
nor ( n19863 , n19861 , n19862 );
xnor ( n19864 , n19863 , n17000 );
and ( n19865 , n19859 , n19864 );
and ( n19866 , n19855 , n19864 );
or ( n19867 , n19860 , n19865 , n19866 );
xor ( n19868 , n19569 , n19573 );
xor ( n19869 , n19868 , n19578 );
and ( n19870 , n19867 , n19869 );
xor ( n19871 , n19746 , n19758 );
xor ( n19872 , n19871 , n19763 );
and ( n19873 , n19869 , n19872 );
and ( n19874 , n19867 , n19872 );
or ( n19875 , n19870 , n19873 , n19874 );
xor ( n19876 , n19595 , n19597 );
xor ( n19877 , n19876 , n19600 );
and ( n19878 , n19875 , n19877 );
xor ( n19879 , n19828 , n19830 );
xor ( n19880 , n19879 , n19833 );
and ( n19881 , n19878 , n19880 );
xor ( n19882 , n19697 , n19701 );
xor ( n19883 , n19882 , n19706 );
xor ( n19884 , n19713 , n19717 );
xor ( n19885 , n19884 , n19722 );
and ( n19886 , n19883 , n19885 );
xor ( n19887 , n19855 , n19859 );
xor ( n19888 , n19887 , n19864 );
and ( n19889 , n19885 , n19888 );
and ( n19890 , n19883 , n19888 );
or ( n19891 , n19886 , n19889 , n19890 );
xor ( n19892 , n19774 , n19776 );
xor ( n19893 , n19892 , n19779 );
and ( n19894 , n19891 , n19893 );
xor ( n19895 , n19867 , n19869 );
xor ( n19896 , n19895 , n19872 );
and ( n19897 , n19893 , n19896 );
and ( n19898 , n19891 , n19896 );
or ( n19899 , n19894 , n19897 , n19898 );
xor ( n19900 , n19745 , n19766 );
xor ( n19901 , n19900 , n19769 );
and ( n19902 , n19899 , n19901 );
xor ( n19903 , n19782 , n19784 );
xor ( n19904 , n19903 , n19787 );
and ( n19905 , n19901 , n19904 );
and ( n19906 , n19899 , n19904 );
or ( n19907 , n19902 , n19905 , n19906 );
and ( n19908 , n19880 , n19907 );
and ( n19909 , n19878 , n19907 );
or ( n19910 , n19881 , n19908 , n19909 );
and ( n19911 , n19847 , n19910 );
xor ( n19912 , n19709 , n19725 );
xor ( n19913 , n19912 , n19742 );
and ( n19914 , n16472 , n18077 );
and ( n19915 , n16457 , n18075 );
nor ( n19916 , n19914 , n19915 );
xnor ( n19917 , n19916 , n17919 );
and ( n19918 , n17107 , n17116 );
and ( n19919 , n17045 , n17114 );
nor ( n19920 , n19918 , n19919 );
xnor ( n19921 , n19920 , n17000 );
and ( n19922 , n19917 , n19921 );
and ( n19923 , n18708 , n16237 );
and ( n19924 , n18654 , n16235 );
nor ( n19925 , n19923 , n19924 );
xnor ( n19926 , n19925 , n16186 );
and ( n19927 , n19921 , n19926 );
and ( n19928 , n19917 , n19926 );
or ( n19929 , n19922 , n19927 , n19928 );
xor ( n19930 , n19750 , n19754 );
xor ( n19931 , n19930 , n19587 );
and ( n19932 , n19929 , n19931 );
xor ( n19933 , n19730 , n19734 );
xor ( n19934 , n19933 , n19739 );
and ( n19935 , n19931 , n19934 );
and ( n19936 , n19929 , n19934 );
or ( n19937 , n19932 , n19935 , n19936 );
and ( n19938 , n19913 , n19937 );
and ( n19939 , n16247 , n18698 );
and ( n19940 , n16229 , n18695 );
nor ( n19941 , n19939 , n19940 );
xnor ( n19942 , n19941 , n18211 );
and ( n19943 , n16936 , n17317 );
and ( n19944 , n16820 , n17315 );
nor ( n19945 , n19943 , n19944 );
xnor ( n19946 , n19945 , n17215 );
and ( n19947 , n19942 , n19946 );
and ( n19948 , n18506 , n16331 );
and ( n19949 , n18203 , n16329 );
nor ( n19950 , n19948 , n19949 );
xnor ( n19951 , n19950 , n16299 );
and ( n19952 , n19946 , n19951 );
and ( n19953 , n19942 , n19951 );
or ( n19954 , n19947 , n19952 , n19953 );
and ( n19955 , n16611 , n17797 );
and ( n19956 , n16510 , n17795 );
nor ( n19957 , n19955 , n19956 );
xnor ( n19958 , n19957 , n17726 );
and ( n19959 , n17327 , n16913 );
and ( n19960 , n17240 , n16911 );
nor ( n19961 , n19959 , n19960 );
xnor ( n19962 , n19961 , n16848 );
and ( n19963 , n19958 , n19962 );
and ( n19964 , n17530 , n16750 );
and ( n19965 , n17482 , n16748 );
nor ( n19966 , n19964 , n19965 );
xnor ( n19967 , n19966 , n16647 );
and ( n19968 , n19962 , n19967 );
and ( n19969 , n19958 , n19967 );
or ( n19970 , n19963 , n19968 , n19969 );
and ( n19971 , n19954 , n19970 );
and ( n19972 , n16725 , n17555 );
and ( n19973 , n16688 , n17553 );
nor ( n19974 , n19972 , n19973 );
xnor ( n19975 , n19974 , n17457 );
and ( n19976 , n17985 , n16543 );
and ( n19977 , n17844 , n16541 );
nor ( n19978 , n19976 , n19977 );
xnor ( n19979 , n19978 , n16521 );
and ( n19980 , n19975 , n19979 );
and ( n19981 , n18255 , n16450 );
and ( n19982 , n18145 , n16448 );
nor ( n19983 , n19981 , n19982 );
xnor ( n19984 , n19983 , n16395 );
and ( n19985 , n19979 , n19984 );
and ( n19986 , n19975 , n19984 );
or ( n19987 , n19980 , n19985 , n19986 );
and ( n19988 , n19970 , n19987 );
and ( n19989 , n19954 , n19987 );
or ( n19990 , n19971 , n19988 , n19989 );
and ( n19991 , n19937 , n19990 );
and ( n19992 , n19913 , n19990 );
or ( n19993 , n19938 , n19991 , n19992 );
xor ( n19994 , n19875 , n19877 );
and ( n19995 , n19993 , n19994 );
xor ( n19996 , n19851 , n19854 );
and ( n19997 , n16279 , n18698 );
and ( n19998 , n16247 , n18695 );
nor ( n19999 , n19997 , n19998 );
xnor ( n20000 , n19999 , n18211 );
and ( n20001 , n18145 , n16543 );
and ( n20002 , n17985 , n16541 );
nor ( n20003 , n20001 , n20002 );
xnor ( n20004 , n20003 , n16521 );
and ( n20005 , n20000 , n20004 );
and ( n20006 , n18203 , n16450 );
and ( n20007 , n18255 , n16448 );
nor ( n20008 , n20006 , n20007 );
xnor ( n20009 , n20008 , n16395 );
and ( n20010 , n20004 , n20009 );
and ( n20011 , n20000 , n20009 );
or ( n20012 , n20005 , n20010 , n20011 );
and ( n20013 , n19996 , n20012 );
and ( n20014 , n16820 , n17555 );
and ( n20015 , n16725 , n17553 );
nor ( n20016 , n20014 , n20015 );
xnor ( n20017 , n20016 , n17457 );
and ( n20018 , n17482 , n16913 );
and ( n20019 , n17327 , n16911 );
nor ( n20020 , n20018 , n20019 );
xnor ( n20021 , n20020 , n16848 );
and ( n20022 , n20017 , n20021 );
and ( n20023 , n17844 , n16750 );
and ( n20024 , n17530 , n16748 );
nor ( n20025 , n20023 , n20024 );
xnor ( n20026 , n20025 , n16647 );
and ( n20027 , n20021 , n20026 );
and ( n20028 , n20017 , n20026 );
or ( n20029 , n20022 , n20027 , n20028 );
and ( n20030 , n20012 , n20029 );
and ( n20031 , n19996 , n20029 );
or ( n20032 , n20013 , n20030 , n20031 );
and ( n20033 , n16510 , n18077 );
and ( n20034 , n16472 , n18075 );
nor ( n20035 , n20033 , n20034 );
xnor ( n20036 , n20035 , n17919 );
and ( n20037 , n17045 , n17317 );
and ( n20038 , n16936 , n17315 );
nor ( n20039 , n20037 , n20038 );
xnor ( n20040 , n20039 , n17215 );
and ( n20041 , n20036 , n20040 );
and ( n20042 , n18654 , n16331 );
and ( n20043 , n18506 , n16329 );
nor ( n20044 , n20042 , n20043 );
xnor ( n20045 , n20044 , n16299 );
and ( n20046 , n20040 , n20045 );
and ( n20047 , n20036 , n20045 );
or ( n20048 , n20041 , n20046 , n20047 );
and ( n20049 , n16457 , n18570 );
and ( n20050 , n16365 , n18568 );
nor ( n20051 , n20049 , n20050 );
xnor ( n20052 , n20051 , n18214 );
and ( n20053 , n16688 , n17797 );
and ( n20054 , n16611 , n17795 );
nor ( n20055 , n20053 , n20054 );
xnor ( n20056 , n20055 , n17726 );
and ( n20057 , n20052 , n20056 );
and ( n20058 , n20056 , n19852 );
and ( n20059 , n20052 , n19852 );
or ( n20060 , n20057 , n20058 , n20059 );
and ( n20061 , n20048 , n20060 );
xor ( n20062 , n19917 , n19921 );
xor ( n20063 , n20062 , n19926 );
and ( n20064 , n20060 , n20063 );
and ( n20065 , n20048 , n20063 );
or ( n20066 , n20061 , n20064 , n20065 );
and ( n20067 , n20032 , n20066 );
xor ( n20068 , n19929 , n19931 );
xor ( n20069 , n20068 , n19934 );
xor ( n20070 , n19942 , n19946 );
xor ( n20071 , n20070 , n19951 );
xor ( n20072 , n19958 , n19962 );
xor ( n20073 , n20072 , n19967 );
and ( n20074 , n20071 , n20073 );
xor ( n20075 , n19975 , n19979 );
xor ( n20076 , n20075 , n19984 );
and ( n20077 , n20073 , n20076 );
and ( n20078 , n20071 , n20076 );
or ( n20079 , n20074 , n20077 , n20078 );
and ( n20080 , n20069 , n20079 );
xor ( n20081 , n19954 , n19970 );
xor ( n20082 , n20081 , n19987 );
and ( n20083 , n20079 , n20082 );
and ( n20084 , n20069 , n20082 );
or ( n20085 , n20080 , n20083 , n20084 );
and ( n20086 , n20067 , n20085 );
xor ( n20087 , n19913 , n19937 );
xor ( n20088 , n20087 , n19990 );
and ( n20089 , n20085 , n20088 );
and ( n20090 , n20067 , n20088 );
or ( n20091 , n20086 , n20089 , n20090 );
and ( n20092 , n19994 , n20091 );
and ( n20093 , n19993 , n20091 );
or ( n20094 , n19995 , n20092 , n20093 );
xor ( n20095 , n19899 , n19901 );
xor ( n20096 , n20095 , n19904 );
xor ( n20097 , n19891 , n19893 );
xor ( n20098 , n20097 , n19896 );
xor ( n20099 , n19883 , n19885 );
xor ( n20100 , n20099 , n19888 );
xor ( n20101 , n20032 , n20066 );
and ( n20102 , n20100 , n20101 );
and ( n20103 , n16936 , n17555 );
and ( n20104 , n16820 , n17553 );
nor ( n20105 , n20103 , n20104 );
xnor ( n20106 , n20105 , n17457 );
and ( n20107 , n18255 , n16543 );
and ( n20108 , n18145 , n16541 );
nor ( n20109 , n20107 , n20108 );
xnor ( n20110 , n20109 , n16521 );
and ( n20111 , n20106 , n20110 );
and ( n20112 , n18506 , n16450 );
and ( n20113 , n18203 , n16448 );
nor ( n20114 , n20112 , n20113 );
xnor ( n20115 , n20114 , n16395 );
and ( n20116 , n20110 , n20115 );
and ( n20117 , n20106 , n20115 );
or ( n20118 , n20111 , n20116 , n20117 );
and ( n20119 , n16472 , n18570 );
and ( n20120 , n16457 , n18568 );
nor ( n20121 , n20119 , n20120 );
xnor ( n20122 , n20121 , n18214 );
and ( n20123 , n18708 , n16329 );
not ( n20124 , n20123 );
and ( n20125 , n20124 , n16299 );
and ( n20126 , n20122 , n20125 );
and ( n20127 , n20118 , n20126 );
and ( n20128 , n17240 , n17116 );
and ( n20129 , n17107 , n17114 );
nor ( n20130 , n20128 , n20129 );
xnor ( n20131 , n20130 , n17000 );
and ( n20132 , n20126 , n20131 );
and ( n20133 , n20118 , n20131 );
or ( n20134 , n20127 , n20132 , n20133 );
xor ( n20135 , n20000 , n20004 );
xor ( n20136 , n20135 , n20009 );
xor ( n20137 , n20052 , n20056 );
xor ( n20138 , n20137 , n19852 );
and ( n20139 , n20136 , n20138 );
xor ( n20140 , n20017 , n20021 );
xor ( n20141 , n20140 , n20026 );
and ( n20142 , n20138 , n20141 );
and ( n20143 , n20136 , n20141 );
or ( n20144 , n20139 , n20142 , n20143 );
and ( n20145 , n20134 , n20144 );
xor ( n20146 , n20048 , n20060 );
xor ( n20147 , n20146 , n20063 );
and ( n20148 , n20144 , n20147 );
and ( n20149 , n20134 , n20147 );
or ( n20150 , n20145 , n20148 , n20149 );
and ( n20151 , n20101 , n20150 );
and ( n20152 , n20100 , n20150 );
or ( n20153 , n20102 , n20151 , n20152 );
and ( n20154 , n20098 , n20153 );
xor ( n20155 , n20067 , n20085 );
xor ( n20156 , n20155 , n20088 );
and ( n20157 , n20153 , n20156 );
and ( n20158 , n20098 , n20156 );
or ( n20159 , n20154 , n20157 , n20158 );
and ( n20160 , n20096 , n20159 );
xor ( n20161 , n19993 , n19994 );
xor ( n20162 , n20161 , n20091 );
and ( n20163 , n20159 , n20162 );
and ( n20164 , n20096 , n20162 );
or ( n20165 , n20160 , n20163 , n20164 );
and ( n20166 , n20094 , n20165 );
xor ( n20167 , n19878 , n19880 );
xor ( n20168 , n20167 , n19907 );
and ( n20169 , n20165 , n20168 );
and ( n20170 , n20094 , n20168 );
or ( n20171 , n20166 , n20169 , n20170 );
and ( n20172 , n19910 , n20171 );
and ( n20173 , n19847 , n20171 );
or ( n20174 , n19911 , n20172 , n20173 );
and ( n20175 , n19844 , n20174 );
and ( n20176 , n19826 , n20174 );
or ( n20177 , n19845 , n20175 , n20176 );
and ( n20178 , n19824 , n20177 );
xor ( n20179 , n19824 , n20177 );
xor ( n20180 , n19826 , n19844 );
xor ( n20181 , n20180 , n20174 );
xor ( n20182 , n19847 , n19910 );
xor ( n20183 , n20182 , n20171 );
xor ( n20184 , n20094 , n20165 );
xor ( n20185 , n20184 , n20168 );
xor ( n20186 , n20096 , n20159 );
xor ( n20187 , n20186 , n20162 );
and ( n20188 , n16725 , n17797 );
and ( n20189 , n16688 , n17795 );
nor ( n20190 , n20188 , n20189 );
xnor ( n20191 , n20190 , n17726 );
and ( n20192 , n17530 , n16913 );
and ( n20193 , n17482 , n16911 );
nor ( n20194 , n20192 , n20193 );
xnor ( n20195 , n20194 , n16848 );
and ( n20196 , n20191 , n20195 );
and ( n20197 , n17985 , n16750 );
and ( n20198 , n17844 , n16748 );
nor ( n20199 , n20197 , n20198 );
xnor ( n20200 , n20199 , n16647 );
and ( n20201 , n20195 , n20200 );
and ( n20202 , n20191 , n20200 );
or ( n20203 , n20196 , n20201 , n20202 );
and ( n20204 , n16365 , n18698 );
and ( n20205 , n16279 , n18695 );
nor ( n20206 , n20204 , n20205 );
xnor ( n20207 , n20206 , n18211 );
and ( n20208 , n16611 , n18077 );
and ( n20209 , n16510 , n18075 );
nor ( n20210 , n20208 , n20209 );
xnor ( n20211 , n20210 , n17919 );
and ( n20212 , n20207 , n20211 );
and ( n20213 , n18708 , n16331 );
and ( n20214 , n18654 , n16329 );
nor ( n20215 , n20213 , n20214 );
xnor ( n20216 , n20215 , n16299 );
and ( n20217 , n20211 , n20216 );
and ( n20218 , n20207 , n20216 );
or ( n20219 , n20212 , n20217 , n20218 );
and ( n20220 , n20203 , n20219 );
xor ( n20221 , n20036 , n20040 );
xor ( n20222 , n20221 , n20045 );
and ( n20223 , n20219 , n20222 );
and ( n20224 , n20203 , n20222 );
or ( n20225 , n20220 , n20223 , n20224 );
xor ( n20226 , n19996 , n20012 );
xor ( n20227 , n20226 , n20029 );
and ( n20228 , n20225 , n20227 );
xor ( n20229 , n20069 , n20079 );
xor ( n20230 , n20229 , n20082 );
and ( n20231 , n20228 , n20230 );
and ( n20232 , n16688 , n18077 );
and ( n20233 , n16611 , n18075 );
nor ( n20234 , n20232 , n20233 );
xnor ( n20235 , n20234 , n17919 );
and ( n20236 , n17240 , n17317 );
and ( n20237 , n17107 , n17315 );
nor ( n20238 , n20236 , n20237 );
xnor ( n20239 , n20238 , n17215 );
and ( n20240 , n20235 , n20239 );
and ( n20241 , n17482 , n17116 );
and ( n20242 , n17327 , n17114 );
nor ( n20243 , n20241 , n20242 );
xnor ( n20244 , n20243 , n17000 );
and ( n20245 , n20239 , n20244 );
and ( n20246 , n20235 , n20244 );
or ( n20247 , n20240 , n20245 , n20246 );
and ( n20248 , n16457 , n18698 );
and ( n20249 , n16365 , n18695 );
nor ( n20250 , n20248 , n20249 );
xnor ( n20251 , n20250 , n18211 );
and ( n20252 , n18203 , n16543 );
and ( n20253 , n18255 , n16541 );
nor ( n20254 , n20252 , n20253 );
xnor ( n20255 , n20254 , n16521 );
and ( n20256 , n20251 , n20255 );
and ( n20257 , n18654 , n16450 );
and ( n20258 , n18506 , n16448 );
nor ( n20259 , n20257 , n20258 );
xnor ( n20260 , n20259 , n16395 );
and ( n20261 , n20255 , n20260 );
and ( n20262 , n20251 , n20260 );
or ( n20263 , n20256 , n20261 , n20262 );
and ( n20264 , n20247 , n20263 );
and ( n20265 , n16510 , n18570 );
and ( n20266 , n16472 , n18568 );
nor ( n20267 , n20265 , n20266 );
xnor ( n20268 , n20267 , n18214 );
and ( n20269 , n16820 , n17797 );
and ( n20270 , n16725 , n17795 );
nor ( n20271 , n20269 , n20270 );
xnor ( n20272 , n20271 , n17726 );
and ( n20273 , n20268 , n20272 );
and ( n20274 , n20272 , n20123 );
and ( n20275 , n20268 , n20123 );
or ( n20276 , n20273 , n20274 , n20275 );
and ( n20277 , n20263 , n20276 );
and ( n20278 , n20247 , n20276 );
or ( n20279 , n20264 , n20277 , n20278 );
xor ( n20280 , n20122 , n20125 );
and ( n20281 , n17107 , n17317 );
and ( n20282 , n17045 , n17315 );
nor ( n20283 , n20281 , n20282 );
xnor ( n20284 , n20283 , n17215 );
and ( n20285 , n20280 , n20284 );
and ( n20286 , n17327 , n17116 );
and ( n20287 , n17240 , n17114 );
nor ( n20288 , n20286 , n20287 );
xnor ( n20289 , n20288 , n17000 );
and ( n20290 , n20284 , n20289 );
and ( n20291 , n20280 , n20289 );
or ( n20292 , n20285 , n20290 , n20291 );
and ( n20293 , n20279 , n20292 );
xor ( n20294 , n20118 , n20126 );
xor ( n20295 , n20294 , n20131 );
and ( n20296 , n20292 , n20295 );
and ( n20297 , n20279 , n20295 );
or ( n20298 , n20293 , n20296 , n20297 );
and ( n20299 , n17045 , n17555 );
and ( n20300 , n16936 , n17553 );
nor ( n20301 , n20299 , n20300 );
xnor ( n20302 , n20301 , n17457 );
and ( n20303 , n17844 , n16913 );
and ( n20304 , n17530 , n16911 );
nor ( n20305 , n20303 , n20304 );
xnor ( n20306 , n20305 , n16848 );
and ( n20307 , n20302 , n20306 );
and ( n20308 , n18145 , n16750 );
and ( n20309 , n17985 , n16748 );
nor ( n20310 , n20308 , n20309 );
xnor ( n20311 , n20310 , n16647 );
and ( n20312 , n20306 , n20311 );
and ( n20313 , n20302 , n20311 );
or ( n20314 , n20307 , n20312 , n20313 );
xor ( n20315 , n20207 , n20211 );
xor ( n20316 , n20315 , n20216 );
and ( n20317 , n20314 , n20316 );
xor ( n20318 , n20106 , n20110 );
xor ( n20319 , n20318 , n20115 );
and ( n20320 , n20316 , n20319 );
and ( n20321 , n20314 , n20319 );
or ( n20322 , n20317 , n20320 , n20321 );
xor ( n20323 , n20203 , n20219 );
xor ( n20324 , n20323 , n20222 );
and ( n20325 , n20322 , n20324 );
xor ( n20326 , n20136 , n20138 );
xor ( n20327 , n20326 , n20141 );
and ( n20328 , n20324 , n20327 );
and ( n20329 , n20322 , n20327 );
or ( n20330 , n20325 , n20328 , n20329 );
and ( n20331 , n20298 , n20330 );
xor ( n20332 , n20134 , n20144 );
xor ( n20333 , n20332 , n20147 );
and ( n20334 , n20330 , n20333 );
and ( n20335 , n20298 , n20333 );
or ( n20336 , n20331 , n20334 , n20335 );
and ( n20337 , n20230 , n20336 );
and ( n20338 , n20228 , n20336 );
or ( n20339 , n20231 , n20337 , n20338 );
xor ( n20340 , n20098 , n20153 );
xor ( n20341 , n20340 , n20156 );
and ( n20342 , n20339 , n20341 );
xor ( n20343 , n20100 , n20101 );
xor ( n20344 , n20343 , n20150 );
xor ( n20345 , n20071 , n20073 );
xor ( n20346 , n20345 , n20076 );
xor ( n20347 , n20225 , n20227 );
and ( n20348 , n20346 , n20347 );
xor ( n20349 , n20298 , n20330 );
xor ( n20350 , n20349 , n20333 );
and ( n20351 , n20347 , n20350 );
and ( n20352 , n20346 , n20350 );
or ( n20353 , n20348 , n20351 , n20352 );
and ( n20354 , n20344 , n20353 );
xor ( n20355 , n20228 , n20230 );
xor ( n20356 , n20355 , n20336 );
and ( n20357 , n20353 , n20356 );
and ( n20358 , n20344 , n20356 );
or ( n20359 , n20354 , n20357 , n20358 );
and ( n20360 , n20341 , n20359 );
and ( n20361 , n20339 , n20359 );
or ( n20362 , n20342 , n20360 , n20361 );
and ( n20363 , n20187 , n20362 );
xor ( n20364 , n20187 , n20362 );
xor ( n20365 , n20339 , n20341 );
xor ( n20366 , n20365 , n20359 );
xor ( n20367 , n20279 , n20292 );
xor ( n20368 , n20367 , n20295 );
xor ( n20369 , n20322 , n20324 );
xor ( n20370 , n20369 , n20327 );
and ( n20371 , n20368 , n20370 );
and ( n20372 , n16936 , n17797 );
and ( n20373 , n16820 , n17795 );
nor ( n20374 , n20372 , n20373 );
xnor ( n20375 , n20374 , n17726 );
and ( n20376 , n17985 , n16913 );
and ( n20377 , n17844 , n16911 );
nor ( n20378 , n20376 , n20377 );
xnor ( n20379 , n20378 , n16848 );
and ( n20380 , n20375 , n20379 );
and ( n20381 , n18255 , n16750 );
and ( n20382 , n18145 , n16748 );
nor ( n20383 , n20381 , n20382 );
xnor ( n20384 , n20383 , n16647 );
and ( n20385 , n20379 , n20384 );
and ( n20386 , n20375 , n20384 );
or ( n20387 , n20380 , n20385 , n20386 );
xor ( n20388 , n20235 , n20239 );
xor ( n20389 , n20388 , n20244 );
and ( n20390 , n20387 , n20389 );
xor ( n20391 , n20302 , n20306 );
xor ( n20392 , n20391 , n20311 );
and ( n20393 , n20389 , n20392 );
and ( n20394 , n20387 , n20392 );
or ( n20395 , n20390 , n20393 , n20394 );
xor ( n20396 , n20247 , n20263 );
xor ( n20397 , n20396 , n20276 );
and ( n20398 , n20395 , n20397 );
xor ( n20399 , n20314 , n20316 );
xor ( n20400 , n20399 , n20319 );
and ( n20401 , n20397 , n20400 );
and ( n20402 , n20395 , n20400 );
or ( n20403 , n20398 , n20401 , n20402 );
and ( n20404 , n20370 , n20403 );
and ( n20405 , n20368 , n20403 );
or ( n20406 , n20371 , n20404 , n20405 );
xor ( n20407 , n20191 , n20195 );
xor ( n20408 , n20407 , n20200 );
xor ( n20409 , n20280 , n20284 );
xor ( n20410 , n20409 , n20289 );
and ( n20411 , n20408 , n20410 );
and ( n20412 , n16472 , n18698 );
and ( n20413 , n16457 , n18695 );
nor ( n20414 , n20412 , n20413 );
xnor ( n20415 , n20414 , n18211 );
and ( n20416 , n16725 , n18077 );
and ( n20417 , n16688 , n18075 );
nor ( n20418 , n20416 , n20417 );
xnor ( n20419 , n20418 , n17919 );
and ( n20420 , n20415 , n20419 );
and ( n20421 , n17327 , n17317 );
and ( n20422 , n17240 , n17315 );
nor ( n20423 , n20421 , n20422 );
xnor ( n20424 , n20423 , n17215 );
and ( n20425 , n20419 , n20424 );
and ( n20426 , n20415 , n20424 );
or ( n20427 , n20420 , n20425 , n20426 );
and ( n20428 , n16611 , n18570 );
and ( n20429 , n16510 , n18568 );
nor ( n20430 , n20428 , n20429 );
xnor ( n20431 , n20430 , n18214 );
and ( n20432 , n18708 , n16448 );
not ( n20433 , n20432 );
and ( n20434 , n20433 , n16395 );
and ( n20435 , n20431 , n20434 );
and ( n20436 , n20427 , n20435 );
and ( n20437 , n18506 , n16543 );
and ( n20438 , n18203 , n16541 );
nor ( n20439 , n20437 , n20438 );
xnor ( n20440 , n20439 , n16521 );
and ( n20441 , n18708 , n16450 );
and ( n20442 , n18654 , n16448 );
nor ( n20443 , n20441 , n20442 );
xnor ( n20444 , n20443 , n16395 );
and ( n20445 , n20440 , n20444 );
and ( n20446 , n20435 , n20445 );
and ( n20447 , n20427 , n20445 );
or ( n20448 , n20436 , n20446 , n20447 );
xor ( n20449 , n20395 , n20397 );
xor ( n20450 , n20449 , n20400 );
and ( n20451 , n20448 , n20450 );
xor ( n20452 , n20408 , n20410 );
and ( n20453 , n20450 , n20452 );
and ( n20454 , n20448 , n20452 );
or ( n20455 , n20451 , n20453 , n20454 );
and ( n20456 , n20411 , n20455 );
xor ( n20457 , n20368 , n20370 );
xor ( n20458 , n20457 , n20403 );
and ( n20459 , n20455 , n20458 );
and ( n20460 , n20411 , n20458 );
or ( n20461 , n20456 , n20459 , n20460 );
and ( n20462 , n20406 , n20461 );
xor ( n20463 , n20346 , n20347 );
xor ( n20464 , n20463 , n20350 );
and ( n20465 , n20461 , n20464 );
and ( n20466 , n20406 , n20464 );
or ( n20467 , n20462 , n20465 , n20466 );
xor ( n20468 , n20344 , n20353 );
xor ( n20469 , n20468 , n20356 );
and ( n20470 , n20467 , n20469 );
xor ( n20471 , n20467 , n20469 );
xor ( n20472 , n20406 , n20461 );
xor ( n20473 , n20472 , n20464 );
xor ( n20474 , n20431 , n20434 );
and ( n20475 , n16688 , n18570 );
and ( n20476 , n16611 , n18568 );
nor ( n20477 , n20475 , n20476 );
xnor ( n20478 , n20477 , n18214 );
and ( n20479 , n18145 , n16913 );
and ( n20480 , n17985 , n16911 );
nor ( n20481 , n20479 , n20480 );
xnor ( n20482 , n20481 , n16848 );
and ( n20483 , n20478 , n20482 );
and ( n20484 , n18203 , n16750 );
and ( n20485 , n18255 , n16748 );
nor ( n20486 , n20484 , n20485 );
xnor ( n20487 , n20486 , n16647 );
and ( n20488 , n20482 , n20487 );
and ( n20489 , n20478 , n20487 );
or ( n20490 , n20483 , n20488 , n20489 );
and ( n20491 , n20474 , n20490 );
and ( n20492 , n17530 , n17116 );
and ( n20493 , n17482 , n17114 );
nor ( n20494 , n20492 , n20493 );
xnor ( n20495 , n20494 , n17000 );
and ( n20496 , n20490 , n20495 );
and ( n20497 , n20474 , n20495 );
or ( n20498 , n20491 , n20496 , n20497 );
xor ( n20499 , n20251 , n20255 );
xor ( n20500 , n20499 , n20260 );
and ( n20501 , n20498 , n20500 );
xor ( n20502 , n20268 , n20272 );
xor ( n20503 , n20502 , n20123 );
and ( n20504 , n20500 , n20503 );
and ( n20505 , n20498 , n20503 );
or ( n20506 , n20501 , n20504 , n20505 );
and ( n20507 , n16510 , n18698 );
and ( n20508 , n16472 , n18695 );
nor ( n20509 , n20507 , n20508 );
xnor ( n20510 , n20509 , n18211 );
and ( n20511 , n17045 , n17797 );
and ( n20512 , n16936 , n17795 );
nor ( n20513 , n20511 , n20512 );
xnor ( n20514 , n20513 , n17726 );
and ( n20515 , n20510 , n20514 );
and ( n20516 , n20514 , n20432 );
and ( n20517 , n20510 , n20432 );
or ( n20518 , n20515 , n20516 , n20517 );
and ( n20519 , n16820 , n18077 );
and ( n20520 , n16725 , n18075 );
nor ( n20521 , n20519 , n20520 );
xnor ( n20522 , n20521 , n17919 );
and ( n20523 , n17240 , n17555 );
and ( n20524 , n17107 , n17553 );
nor ( n20525 , n20523 , n20524 );
xnor ( n20526 , n20525 , n17457 );
and ( n20527 , n20522 , n20526 );
and ( n20528 , n18654 , n16543 );
and ( n20529 , n18506 , n16541 );
nor ( n20530 , n20528 , n20529 );
xnor ( n20531 , n20530 , n16521 );
and ( n20532 , n20526 , n20531 );
and ( n20533 , n20522 , n20531 );
or ( n20534 , n20527 , n20532 , n20533 );
and ( n20535 , n20518 , n20534 );
xor ( n20536 , n20415 , n20419 );
xor ( n20537 , n20536 , n20424 );
and ( n20538 , n20534 , n20537 );
and ( n20539 , n20518 , n20537 );
or ( n20540 , n20535 , n20538 , n20539 );
and ( n20541 , n17107 , n17555 );
and ( n20542 , n17045 , n17553 );
nor ( n20543 , n20541 , n20542 );
xnor ( n20544 , n20543 , n17457 );
xor ( n20545 , n20375 , n20379 );
xor ( n20546 , n20545 , n20384 );
and ( n20547 , n20544 , n20546 );
xor ( n20548 , n20440 , n20444 );
and ( n20549 , n20546 , n20548 );
and ( n20550 , n20544 , n20548 );
or ( n20551 , n20547 , n20549 , n20550 );
and ( n20552 , n20540 , n20551 );
xor ( n20553 , n20427 , n20435 );
xor ( n20554 , n20553 , n20445 );
and ( n20555 , n20551 , n20554 );
and ( n20556 , n20540 , n20554 );
or ( n20557 , n20552 , n20555 , n20556 );
and ( n20558 , n20506 , n20557 );
and ( n20559 , n16936 , n18077 );
and ( n20560 , n16820 , n18075 );
nor ( n20561 , n20559 , n20560 );
xnor ( n20562 , n20561 , n17919 );
and ( n20563 , n17530 , n17317 );
and ( n20564 , n17482 , n17315 );
nor ( n20565 , n20563 , n20564 );
xnor ( n20566 , n20565 , n17215 );
and ( n20567 , n20562 , n20566 );
and ( n20568 , n17985 , n17116 );
and ( n20569 , n17844 , n17114 );
nor ( n20570 , n20568 , n20569 );
xnor ( n20571 , n20570 , n17000 );
and ( n20572 , n20566 , n20571 );
and ( n20573 , n20562 , n20571 );
or ( n20574 , n20567 , n20572 , n20573 );
and ( n20575 , n17107 , n17797 );
and ( n20576 , n17045 , n17795 );
nor ( n20577 , n20575 , n20576 );
xnor ( n20578 , n20577 , n17726 );
and ( n20579 , n18255 , n16913 );
and ( n20580 , n18145 , n16911 );
nor ( n20581 , n20579 , n20580 );
xnor ( n20582 , n20581 , n16848 );
and ( n20583 , n20578 , n20582 );
and ( n20584 , n18506 , n16750 );
and ( n20585 , n18203 , n16748 );
nor ( n20586 , n20584 , n20585 );
xnor ( n20587 , n20586 , n16647 );
and ( n20588 , n20582 , n20587 );
and ( n20589 , n20578 , n20587 );
or ( n20590 , n20583 , n20588 , n20589 );
and ( n20591 , n20574 , n20590 );
and ( n20592 , n16725 , n18570 );
and ( n20593 , n16688 , n18568 );
nor ( n20594 , n20592 , n20593 );
xnor ( n20595 , n20594 , n18214 );
and ( n20596 , n17327 , n17555 );
and ( n20597 , n17240 , n17553 );
nor ( n20598 , n20596 , n20597 );
xnor ( n20599 , n20598 , n17457 );
and ( n20600 , n20595 , n20599 );
and ( n20601 , n18708 , n16543 );
and ( n20602 , n18654 , n16541 );
nor ( n20603 , n20601 , n20602 );
xnor ( n20604 , n20603 , n16521 );
and ( n20605 , n20599 , n20604 );
and ( n20606 , n20595 , n20604 );
or ( n20607 , n20600 , n20605 , n20606 );
and ( n20608 , n20590 , n20607 );
and ( n20609 , n20574 , n20607 );
or ( n20610 , n20591 , n20608 , n20609 );
xor ( n20611 , n20474 , n20490 );
xor ( n20612 , n20611 , n20495 );
and ( n20613 , n20610 , n20612 );
xor ( n20614 , n20518 , n20534 );
xor ( n20615 , n20614 , n20537 );
and ( n20616 , n20612 , n20615 );
and ( n20617 , n20610 , n20615 );
or ( n20618 , n20613 , n20616 , n20617 );
xor ( n20619 , n20387 , n20389 );
xor ( n20620 , n20619 , n20392 );
and ( n20621 , n20618 , n20620 );
xor ( n20622 , n20498 , n20500 );
xor ( n20623 , n20622 , n20503 );
and ( n20624 , n20620 , n20623 );
and ( n20625 , n20618 , n20623 );
or ( n20626 , n20621 , n20624 , n20625 );
and ( n20627 , n20557 , n20626 );
and ( n20628 , n20506 , n20626 );
or ( n20629 , n20558 , n20627 , n20628 );
xor ( n20630 , n20411 , n20455 );
xor ( n20631 , n20630 , n20458 );
and ( n20632 , n20629 , n20631 );
xor ( n20633 , n20448 , n20450 );
xor ( n20634 , n20633 , n20452 );
and ( n20635 , n16611 , n18698 );
and ( n20636 , n16510 , n18695 );
nor ( n20637 , n20635 , n20636 );
xnor ( n20638 , n20637 , n18211 );
and ( n20639 , n18708 , n16541 );
not ( n20640 , n20639 );
and ( n20641 , n20640 , n16521 );
and ( n20642 , n20638 , n20641 );
and ( n20643 , n17482 , n17317 );
and ( n20644 , n17327 , n17315 );
nor ( n20645 , n20643 , n20644 );
xnor ( n20646 , n20645 , n17215 );
and ( n20647 , n20642 , n20646 );
and ( n20648 , n17844 , n17116 );
and ( n20649 , n17530 , n17114 );
nor ( n20650 , n20648 , n20649 );
xnor ( n20651 , n20650 , n17000 );
and ( n20652 , n20646 , n20651 );
and ( n20653 , n20642 , n20651 );
or ( n20654 , n20647 , n20652 , n20653 );
xor ( n20655 , n20510 , n20514 );
xor ( n20656 , n20655 , n20432 );
xor ( n20657 , n20478 , n20482 );
xor ( n20658 , n20657 , n20487 );
and ( n20659 , n20656 , n20658 );
xor ( n20660 , n20522 , n20526 );
xor ( n20661 , n20660 , n20531 );
and ( n20662 , n20658 , n20661 );
and ( n20663 , n20656 , n20661 );
or ( n20664 , n20659 , n20662 , n20663 );
and ( n20665 , n20654 , n20664 );
xor ( n20666 , n20544 , n20546 );
xor ( n20667 , n20666 , n20548 );
and ( n20668 , n20664 , n20667 );
and ( n20669 , n20654 , n20667 );
or ( n20670 , n20665 , n20668 , n20669 );
xor ( n20671 , n20540 , n20551 );
xor ( n20672 , n20671 , n20554 );
and ( n20673 , n20670 , n20672 );
xor ( n20674 , n20618 , n20620 );
xor ( n20675 , n20674 , n20623 );
and ( n20676 , n20672 , n20675 );
and ( n20677 , n20670 , n20675 );
or ( n20678 , n20673 , n20676 , n20677 );
and ( n20679 , n20634 , n20678 );
xor ( n20680 , n20506 , n20557 );
xor ( n20681 , n20680 , n20626 );
and ( n20682 , n20678 , n20681 );
and ( n20683 , n20634 , n20681 );
or ( n20684 , n20679 , n20682 , n20683 );
and ( n20685 , n20631 , n20684 );
and ( n20686 , n20629 , n20684 );
or ( n20687 , n20632 , n20685 , n20686 );
and ( n20688 , n20473 , n20687 );
xor ( n20689 , n20473 , n20687 );
xor ( n20690 , n20629 , n20631 );
xor ( n20691 , n20690 , n20684 );
xor ( n20692 , n20634 , n20678 );
xor ( n20693 , n20692 , n20681 );
xor ( n20694 , n20610 , n20612 );
xor ( n20695 , n20694 , n20615 );
xor ( n20696 , n20638 , n20641 );
and ( n20697 , n16688 , n18698 );
and ( n20698 , n16611 , n18695 );
nor ( n20699 , n20697 , n20698 );
xnor ( n20700 , n20699 , n18211 );
and ( n20701 , n17240 , n17797 );
and ( n20702 , n17107 , n17795 );
nor ( n20703 , n20701 , n20702 );
xnor ( n20704 , n20703 , n17726 );
and ( n20705 , n20700 , n20704 );
and ( n20706 , n20704 , n20639 );
and ( n20707 , n20700 , n20639 );
or ( n20708 , n20705 , n20706 , n20707 );
and ( n20709 , n20696 , n20708 );
and ( n20710 , n16820 , n18570 );
and ( n20711 , n16725 , n18568 );
nor ( n20712 , n20710 , n20711 );
xnor ( n20713 , n20712 , n18214 );
and ( n20714 , n18203 , n16913 );
and ( n20715 , n18255 , n16911 );
nor ( n20716 , n20714 , n20715 );
xnor ( n20717 , n20716 , n16848 );
and ( n20718 , n20713 , n20717 );
and ( n20719 , n18654 , n16750 );
and ( n20720 , n18506 , n16748 );
nor ( n20721 , n20719 , n20720 );
xnor ( n20722 , n20721 , n16647 );
and ( n20723 , n20717 , n20722 );
and ( n20724 , n20713 , n20722 );
or ( n20725 , n20718 , n20723 , n20724 );
and ( n20726 , n20708 , n20725 );
and ( n20727 , n20696 , n20725 );
or ( n20728 , n20709 , n20726 , n20727 );
and ( n20729 , n17045 , n18077 );
and ( n20730 , n16936 , n18075 );
nor ( n20731 , n20729 , n20730 );
xnor ( n20732 , n20731 , n17919 );
and ( n20733 , n17482 , n17555 );
and ( n20734 , n17327 , n17553 );
nor ( n20735 , n20733 , n20734 );
xnor ( n20736 , n20735 , n17457 );
and ( n20737 , n20732 , n20736 );
and ( n20738 , n17844 , n17317 );
and ( n20739 , n17530 , n17315 );
nor ( n20740 , n20738 , n20739 );
xnor ( n20741 , n20740 , n17215 );
and ( n20742 , n20736 , n20741 );
and ( n20743 , n20732 , n20741 );
or ( n20744 , n20737 , n20742 , n20743 );
xor ( n20745 , n20562 , n20566 );
xor ( n20746 , n20745 , n20571 );
and ( n20747 , n20744 , n20746 );
xor ( n20748 , n20578 , n20582 );
xor ( n20749 , n20748 , n20587 );
and ( n20750 , n20746 , n20749 );
and ( n20751 , n20744 , n20749 );
or ( n20752 , n20747 , n20750 , n20751 );
and ( n20753 , n20728 , n20752 );
xor ( n20754 , n20642 , n20646 );
xor ( n20755 , n20754 , n20651 );
and ( n20756 , n20752 , n20755 );
and ( n20757 , n20728 , n20755 );
or ( n20758 , n20753 , n20756 , n20757 );
and ( n20759 , n20695 , n20758 );
xor ( n20760 , n20654 , n20664 );
xor ( n20761 , n20760 , n20667 );
and ( n20762 , n20758 , n20761 );
and ( n20763 , n20695 , n20761 );
or ( n20764 , n20759 , n20762 , n20763 );
xor ( n20765 , n20670 , n20672 );
xor ( n20766 , n20765 , n20675 );
and ( n20767 , n20764 , n20766 );
xor ( n20768 , n20574 , n20590 );
xor ( n20769 , n20768 , n20607 );
xor ( n20770 , n20656 , n20658 );
xor ( n20771 , n20770 , n20661 );
and ( n20772 , n20769 , n20771 );
xor ( n20773 , n20728 , n20752 );
xor ( n20774 , n20773 , n20755 );
and ( n20775 , n20771 , n20774 );
and ( n20776 , n20769 , n20774 );
or ( n20777 , n20772 , n20775 , n20776 );
xor ( n20778 , n20695 , n20758 );
xor ( n20779 , n20778 , n20761 );
and ( n20780 , n20777 , n20779 );
xor ( n20781 , n20595 , n20599 );
xor ( n20782 , n20781 , n20604 );
xor ( n20783 , n20696 , n20708 );
xor ( n20784 , n20783 , n20725 );
and ( n20785 , n20782 , n20784 );
and ( n20786 , n17327 , n17797 );
and ( n20787 , n17240 , n17795 );
nor ( n20788 , n20786 , n20787 );
xnor ( n20789 , n20788 , n17726 );
and ( n20790 , n18506 , n16913 );
and ( n20791 , n18203 , n16911 );
nor ( n20792 , n20790 , n20791 );
xnor ( n20793 , n20792 , n16848 );
and ( n20794 , n20789 , n20793 );
and ( n20795 , n18708 , n16750 );
and ( n20796 , n18654 , n16748 );
nor ( n20797 , n20795 , n20796 );
xnor ( n20798 , n20797 , n16647 );
and ( n20799 , n20793 , n20798 );
and ( n20800 , n20789 , n20798 );
or ( n20801 , n20794 , n20799 , n20800 );
and ( n20802 , n16725 , n18698 );
and ( n20803 , n16688 , n18695 );
nor ( n20804 , n20802 , n20803 );
xnor ( n20805 , n20804 , n18211 );
and ( n20806 , n18708 , n16748 );
not ( n20807 , n20806 );
and ( n20808 , n20807 , n16647 );
and ( n20809 , n20805 , n20808 );
and ( n20810 , n20801 , n20809 );
and ( n20811 , n18145 , n17116 );
and ( n20812 , n17985 , n17114 );
nor ( n20813 , n20811 , n20812 );
xnor ( n20814 , n20813 , n17000 );
and ( n20815 , n20809 , n20814 );
and ( n20816 , n20801 , n20814 );
or ( n20817 , n20810 , n20815 , n20816 );
and ( n20818 , n20784 , n20817 );
and ( n20819 , n20782 , n20817 );
or ( n20820 , n20785 , n20818 , n20819 );
xor ( n20821 , n20769 , n20771 );
xor ( n20822 , n20821 , n20774 );
and ( n20823 , n20820 , n20822 );
and ( n20824 , n16936 , n18570 );
and ( n20825 , n16820 , n18568 );
nor ( n20826 , n20824 , n20825 );
xnor ( n20827 , n20826 , n18214 );
and ( n20828 , n17107 , n18077 );
and ( n20829 , n17045 , n18075 );
nor ( n20830 , n20828 , n20829 );
xnor ( n20831 , n20830 , n17919 );
and ( n20832 , n20827 , n20831 );
and ( n20833 , n17530 , n17555 );
and ( n20834 , n17482 , n17553 );
nor ( n20835 , n20833 , n20834 );
xnor ( n20836 , n20835 , n17457 );
and ( n20837 , n20831 , n20836 );
and ( n20838 , n20827 , n20836 );
or ( n20839 , n20832 , n20837 , n20838 );
xor ( n20840 , n20700 , n20704 );
xor ( n20841 , n20840 , n20639 );
and ( n20842 , n20839 , n20841 );
xor ( n20843 , n20732 , n20736 );
xor ( n20844 , n20843 , n20741 );
and ( n20845 , n20841 , n20844 );
and ( n20846 , n20839 , n20844 );
or ( n20847 , n20842 , n20845 , n20846 );
xor ( n20848 , n20805 , n20808 );
and ( n20849 , n17985 , n17317 );
and ( n20850 , n17844 , n17315 );
nor ( n20851 , n20849 , n20850 );
xnor ( n20852 , n20851 , n17215 );
and ( n20853 , n20848 , n20852 );
and ( n20854 , n18255 , n17116 );
and ( n20855 , n18145 , n17114 );
nor ( n20856 , n20854 , n20855 );
xnor ( n20857 , n20856 , n17000 );
and ( n20858 , n20852 , n20857 );
and ( n20859 , n20848 , n20857 );
or ( n20860 , n20853 , n20858 , n20859 );
xor ( n20861 , n20713 , n20717 );
xor ( n20862 , n20861 , n20722 );
and ( n20863 , n20860 , n20862 );
xor ( n20864 , n20801 , n20809 );
xor ( n20865 , n20864 , n20814 );
and ( n20866 , n20862 , n20865 );
and ( n20867 , n20860 , n20865 );
or ( n20868 , n20863 , n20866 , n20867 );
and ( n20869 , n20847 , n20868 );
xor ( n20870 , n20744 , n20746 );
xor ( n20871 , n20870 , n20749 );
and ( n20872 , n20868 , n20871 );
and ( n20873 , n20847 , n20871 );
or ( n20874 , n20869 , n20872 , n20873 );
and ( n20875 , n20822 , n20874 );
and ( n20876 , n20820 , n20874 );
or ( n20877 , n20823 , n20875 , n20876 );
and ( n20878 , n20779 , n20877 );
and ( n20879 , n20777 , n20877 );
or ( n20880 , n20780 , n20878 , n20879 );
and ( n20881 , n20766 , n20880 );
and ( n20882 , n20764 , n20880 );
or ( n20883 , n20767 , n20881 , n20882 );
and ( n20884 , n20693 , n20883 );
xor ( n20885 , n20693 , n20883 );
xor ( n20886 , n20764 , n20766 );
xor ( n20887 , n20886 , n20880 );
xor ( n20888 , n20777 , n20779 );
xor ( n20889 , n20888 , n20877 );
xor ( n20890 , n20782 , n20784 );
xor ( n20891 , n20890 , n20817 );
xor ( n20892 , n20847 , n20868 );
xor ( n20893 , n20892 , n20871 );
and ( n20894 , n20891 , n20893 );
and ( n20895 , n16820 , n18698 );
and ( n20896 , n16725 , n18695 );
nor ( n20897 , n20895 , n20896 );
xnor ( n20898 , n20897 , n18211 );
and ( n20899 , n17045 , n18570 );
and ( n20900 , n16936 , n18568 );
nor ( n20901 , n20899 , n20900 );
xnor ( n20902 , n20901 , n18214 );
and ( n20903 , n20898 , n20902 );
and ( n20904 , n20902 , n20806 );
and ( n20905 , n20898 , n20806 );
or ( n20906 , n20903 , n20904 , n20905 );
and ( n20907 , n17240 , n18077 );
and ( n20908 , n17107 , n18075 );
nor ( n20909 , n20907 , n20908 );
xnor ( n20910 , n20909 , n17919 );
and ( n20911 , n18145 , n17317 );
and ( n20912 , n17985 , n17315 );
nor ( n20913 , n20911 , n20912 );
xnor ( n20914 , n20913 , n17215 );
and ( n20915 , n20910 , n20914 );
and ( n20916 , n18203 , n17116 );
and ( n20917 , n18255 , n17114 );
nor ( n20918 , n20916 , n20917 );
xnor ( n20919 , n20918 , n17000 );
and ( n20920 , n20914 , n20919 );
and ( n20921 , n20910 , n20919 );
or ( n20922 , n20915 , n20920 , n20921 );
and ( n20923 , n20906 , n20922 );
and ( n20924 , n17482 , n17797 );
and ( n20925 , n17327 , n17795 );
nor ( n20926 , n20924 , n20925 );
xnor ( n20927 , n20926 , n17726 );
and ( n20928 , n17844 , n17555 );
and ( n20929 , n17530 , n17553 );
nor ( n20930 , n20928 , n20929 );
xnor ( n20931 , n20930 , n17457 );
and ( n20932 , n20927 , n20931 );
and ( n20933 , n18654 , n16913 );
and ( n20934 , n18506 , n16911 );
nor ( n20935 , n20933 , n20934 );
xnor ( n20936 , n20935 , n16848 );
and ( n20937 , n20931 , n20936 );
and ( n20938 , n20927 , n20936 );
or ( n20939 , n20932 , n20937 , n20938 );
and ( n20940 , n20922 , n20939 );
and ( n20941 , n20906 , n20939 );
or ( n20942 , n20923 , n20940 , n20941 );
xor ( n20943 , n20827 , n20831 );
xor ( n20944 , n20943 , n20836 );
xor ( n20945 , n20789 , n20793 );
xor ( n20946 , n20945 , n20798 );
and ( n20947 , n20944 , n20946 );
xor ( n20948 , n20848 , n20852 );
xor ( n20949 , n20948 , n20857 );
and ( n20950 , n20946 , n20949 );
and ( n20951 , n20944 , n20949 );
or ( n20952 , n20947 , n20950 , n20951 );
and ( n20953 , n20942 , n20952 );
xor ( n20954 , n20839 , n20841 );
xor ( n20955 , n20954 , n20844 );
and ( n20956 , n20952 , n20955 );
and ( n20957 , n20942 , n20955 );
or ( n20958 , n20953 , n20956 , n20957 );
and ( n20959 , n20893 , n20958 );
and ( n20960 , n20891 , n20958 );
or ( n20961 , n20894 , n20959 , n20960 );
xor ( n20962 , n20820 , n20822 );
xor ( n20963 , n20962 , n20874 );
and ( n20964 , n20961 , n20963 );
and ( n20965 , n17327 , n18077 );
and ( n20966 , n17240 , n18075 );
nor ( n20967 , n20965 , n20966 );
xnor ( n20968 , n20967 , n17919 );
and ( n20969 , n17985 , n17555 );
and ( n20970 , n17844 , n17553 );
nor ( n20971 , n20969 , n20970 );
xnor ( n20972 , n20971 , n17457 );
and ( n20973 , n20968 , n20972 );
and ( n20974 , n18255 , n17317 );
and ( n20975 , n18145 , n17315 );
nor ( n20976 , n20974 , n20975 );
xnor ( n20977 , n20976 , n17215 );
and ( n20978 , n20972 , n20977 );
and ( n20979 , n20968 , n20977 );
or ( n20980 , n20973 , n20978 , n20979 );
and ( n20981 , n17107 , n18570 );
and ( n20982 , n17045 , n18568 );
nor ( n20983 , n20981 , n20982 );
xnor ( n20984 , n20983 , n18214 );
and ( n20985 , n17530 , n17797 );
and ( n20986 , n17482 , n17795 );
nor ( n20987 , n20985 , n20986 );
xnor ( n20988 , n20987 , n17726 );
and ( n20989 , n20984 , n20988 );
and ( n20990 , n18708 , n16913 );
and ( n20991 , n18654 , n16911 );
nor ( n20992 , n20990 , n20991 );
xnor ( n20993 , n20992 , n16848 );
and ( n20994 , n20988 , n20993 );
and ( n20995 , n20984 , n20993 );
or ( n20996 , n20989 , n20994 , n20995 );
and ( n20997 , n20980 , n20996 );
and ( n20998 , n16936 , n18698 );
and ( n20999 , n16820 , n18695 );
nor ( n21000 , n20998 , n20999 );
xnor ( n21001 , n21000 , n18211 );
and ( n21002 , n18708 , n16911 );
not ( n21003 , n21002 );
and ( n21004 , n21003 , n16848 );
and ( n21005 , n21001 , n21004 );
and ( n21006 , n20996 , n21005 );
and ( n21007 , n20980 , n21005 );
or ( n21008 , n20997 , n21006 , n21007 );
xor ( n21009 , n20898 , n20902 );
xor ( n21010 , n21009 , n20806 );
xor ( n21011 , n20910 , n20914 );
xor ( n21012 , n21011 , n20919 );
and ( n21013 , n21010 , n21012 );
xor ( n21014 , n20927 , n20931 );
xor ( n21015 , n21014 , n20936 );
and ( n21016 , n21012 , n21015 );
and ( n21017 , n21010 , n21015 );
or ( n21018 , n21013 , n21016 , n21017 );
and ( n21019 , n21008 , n21018 );
xor ( n21020 , n20906 , n20922 );
xor ( n21021 , n21020 , n20939 );
and ( n21022 , n21018 , n21021 );
and ( n21023 , n21008 , n21021 );
or ( n21024 , n21019 , n21022 , n21023 );
xor ( n21025 , n20860 , n20862 );
xor ( n21026 , n21025 , n20865 );
and ( n21027 , n21024 , n21026 );
xor ( n21028 , n20942 , n20952 );
xor ( n21029 , n21028 , n20955 );
and ( n21030 , n21026 , n21029 );
and ( n21031 , n21024 , n21029 );
or ( n21032 , n21027 , n21030 , n21031 );
xor ( n21033 , n20891 , n20893 );
xor ( n21034 , n21033 , n20958 );
and ( n21035 , n21032 , n21034 );
xor ( n21036 , n21001 , n21004 );
and ( n21037 , n17045 , n18698 );
and ( n21038 , n16936 , n18695 );
nor ( n21039 , n21037 , n21038 );
xnor ( n21040 , n21039 , n18211 );
and ( n21041 , n17240 , n18570 );
and ( n21042 , n17107 , n18568 );
nor ( n21043 , n21041 , n21042 );
xnor ( n21044 , n21043 , n18214 );
and ( n21045 , n21040 , n21044 );
and ( n21046 , n21044 , n21002 );
and ( n21047 , n21040 , n21002 );
or ( n21048 , n21045 , n21046 , n21047 );
and ( n21049 , n21036 , n21048 );
and ( n21050 , n18506 , n17116 );
and ( n21051 , n18203 , n17114 );
nor ( n21052 , n21050 , n21051 );
xnor ( n21053 , n21052 , n17000 );
and ( n21054 , n21048 , n21053 );
and ( n21055 , n21036 , n21053 );
or ( n21056 , n21049 , n21054 , n21055 );
and ( n21057 , n17482 , n18077 );
and ( n21058 , n17327 , n18075 );
nor ( n21059 , n21057 , n21058 );
xnor ( n21060 , n21059 , n17919 );
and ( n21061 , n17844 , n17797 );
and ( n21062 , n17530 , n17795 );
nor ( n21063 , n21061 , n21062 );
xnor ( n21064 , n21063 , n17726 );
and ( n21065 , n21060 , n21064 );
and ( n21066 , n18145 , n17555 );
and ( n21067 , n17985 , n17553 );
nor ( n21068 , n21066 , n21067 );
xnor ( n21069 , n21068 , n17457 );
and ( n21070 , n21064 , n21069 );
and ( n21071 , n21060 , n21069 );
or ( n21072 , n21065 , n21070 , n21071 );
xor ( n21073 , n20968 , n20972 );
xor ( n21074 , n21073 , n20977 );
and ( n21075 , n21072 , n21074 );
xor ( n21076 , n20984 , n20988 );
xor ( n21077 , n21076 , n20993 );
and ( n21078 , n21074 , n21077 );
and ( n21079 , n21072 , n21077 );
or ( n21080 , n21075 , n21078 , n21079 );
and ( n21081 , n21056 , n21080 );
xor ( n21082 , n20980 , n20996 );
xor ( n21083 , n21082 , n21005 );
and ( n21084 , n21080 , n21083 );
and ( n21085 , n21056 , n21083 );
or ( n21086 , n21081 , n21084 , n21085 );
xor ( n21087 , n20944 , n20946 );
xor ( n21088 , n21087 , n20949 );
and ( n21089 , n21086 , n21088 );
xor ( n21090 , n21008 , n21018 );
xor ( n21091 , n21090 , n21021 );
and ( n21092 , n21088 , n21091 );
and ( n21093 , n21086 , n21091 );
or ( n21094 , n21089 , n21092 , n21093 );
xor ( n21095 , n21024 , n21026 );
xor ( n21096 , n21095 , n21029 );
and ( n21097 , n21094 , n21096 );
xor ( n21098 , n21086 , n21088 );
xor ( n21099 , n21098 , n21091 );
and ( n21100 , n17107 , n18698 );
and ( n21101 , n17045 , n18695 );
nor ( n21102 , n21100 , n21101 );
xnor ( n21103 , n21102 , n18211 );
and ( n21104 , n18708 , n17114 );
not ( n21105 , n21104 );
and ( n21106 , n21105 , n17000 );
and ( n21107 , n21103 , n21106 );
and ( n21108 , n18203 , n17317 );
and ( n21109 , n18255 , n17315 );
nor ( n21110 , n21108 , n21109 );
xnor ( n21111 , n21110 , n17215 );
and ( n21112 , n21107 , n21111 );
and ( n21113 , n18654 , n17116 );
and ( n21114 , n18506 , n17114 );
nor ( n21115 , n21113 , n21114 );
xnor ( n21116 , n21115 , n17000 );
and ( n21117 , n21111 , n21116 );
and ( n21118 , n21107 , n21116 );
or ( n21119 , n21112 , n21117 , n21118 );
and ( n21120 , n17530 , n18077 );
and ( n21121 , n17482 , n18075 );
nor ( n21122 , n21120 , n21121 );
xnor ( n21123 , n21122 , n17919 );
and ( n21124 , n18506 , n17317 );
and ( n21125 , n18203 , n17315 );
nor ( n21126 , n21124 , n21125 );
xnor ( n21127 , n21126 , n17215 );
and ( n21128 , n21123 , n21127 );
and ( n21129 , n18708 , n17116 );
and ( n21130 , n18654 , n17114 );
nor ( n21131 , n21129 , n21130 );
xnor ( n21132 , n21131 , n17000 );
and ( n21133 , n21127 , n21132 );
and ( n21134 , n21123 , n21132 );
or ( n21135 , n21128 , n21133 , n21134 );
and ( n21136 , n17327 , n18570 );
and ( n21137 , n17240 , n18568 );
nor ( n21138 , n21136 , n21137 );
xnor ( n21139 , n21138 , n18214 );
and ( n21140 , n17985 , n17797 );
and ( n21141 , n17844 , n17795 );
nor ( n21142 , n21140 , n21141 );
xnor ( n21143 , n21142 , n17726 );
and ( n21144 , n21139 , n21143 );
and ( n21145 , n18255 , n17555 );
and ( n21146 , n18145 , n17553 );
nor ( n21147 , n21145 , n21146 );
xnor ( n21148 , n21147 , n17457 );
and ( n21149 , n21143 , n21148 );
and ( n21150 , n21139 , n21148 );
or ( n21151 , n21144 , n21149 , n21150 );
and ( n21152 , n21135 , n21151 );
xor ( n21153 , n21040 , n21044 );
xor ( n21154 , n21153 , n21002 );
and ( n21155 , n21151 , n21154 );
and ( n21156 , n21135 , n21154 );
or ( n21157 , n21152 , n21155 , n21156 );
and ( n21158 , n21119 , n21157 );
xor ( n21159 , n21036 , n21048 );
xor ( n21160 , n21159 , n21053 );
and ( n21161 , n21157 , n21160 );
and ( n21162 , n21119 , n21160 );
or ( n21163 , n21158 , n21161 , n21162 );
xor ( n21164 , n21010 , n21012 );
xor ( n21165 , n21164 , n21015 );
and ( n21166 , n21163 , n21165 );
xor ( n21167 , n21056 , n21080 );
xor ( n21168 , n21167 , n21083 );
and ( n21169 , n21165 , n21168 );
and ( n21170 , n21163 , n21168 );
or ( n21171 , n21166 , n21169 , n21170 );
and ( n21172 , n21099 , n21171 );
xor ( n21173 , n21163 , n21165 );
xor ( n21174 , n21173 , n21168 );
xor ( n21175 , n21103 , n21106 );
and ( n21176 , n17240 , n18698 );
and ( n21177 , n17107 , n18695 );
nor ( n21178 , n21176 , n21177 );
xnor ( n21179 , n21178 , n18211 );
and ( n21180 , n18203 , n17555 );
and ( n21181 , n18255 , n17553 );
nor ( n21182 , n21180 , n21181 );
xnor ( n21183 , n21182 , n17457 );
and ( n21184 , n21179 , n21183 );
and ( n21185 , n18654 , n17317 );
and ( n21186 , n18506 , n17315 );
nor ( n21187 , n21185 , n21186 );
xnor ( n21188 , n21187 , n17215 );
and ( n21189 , n21183 , n21188 );
and ( n21190 , n21179 , n21188 );
or ( n21191 , n21184 , n21189 , n21190 );
and ( n21192 , n21175 , n21191 );
and ( n21193 , n17482 , n18570 );
and ( n21194 , n17327 , n18568 );
nor ( n21195 , n21193 , n21194 );
xnor ( n21196 , n21195 , n18214 );
and ( n21197 , n18145 , n17797 );
and ( n21198 , n17985 , n17795 );
nor ( n21199 , n21197 , n21198 );
xnor ( n21200 , n21199 , n17726 );
and ( n21201 , n21196 , n21200 );
and ( n21202 , n21200 , n21104 );
and ( n21203 , n21196 , n21104 );
or ( n21204 , n21201 , n21202 , n21203 );
and ( n21205 , n21191 , n21204 );
and ( n21206 , n21175 , n21204 );
or ( n21207 , n21192 , n21205 , n21206 );
xor ( n21208 , n21060 , n21064 );
xor ( n21209 , n21208 , n21069 );
and ( n21210 , n21207 , n21209 );
xor ( n21211 , n21107 , n21111 );
xor ( n21212 , n21211 , n21116 );
and ( n21213 , n21209 , n21212 );
and ( n21214 , n21207 , n21212 );
or ( n21215 , n21210 , n21213 , n21214 );
xor ( n21216 , n21072 , n21074 );
xor ( n21217 , n21216 , n21077 );
and ( n21218 , n21215 , n21217 );
xor ( n21219 , n21119 , n21157 );
xor ( n21220 , n21219 , n21160 );
and ( n21221 , n21217 , n21220 );
and ( n21222 , n21215 , n21220 );
or ( n21223 , n21218 , n21221 , n21222 );
and ( n21224 , n21174 , n21223 );
xor ( n21225 , n21215 , n21217 );
xor ( n21226 , n21225 , n21220 );
and ( n21227 , n17327 , n18698 );
and ( n21228 , n17240 , n18695 );
nor ( n21229 , n21227 , n21228 );
xnor ( n21230 , n21229 , n18211 );
and ( n21231 , n18255 , n17797 );
and ( n21232 , n18145 , n17795 );
nor ( n21233 , n21231 , n21232 );
xnor ( n21234 , n21233 , n17726 );
and ( n21235 , n21230 , n21234 );
and ( n21236 , n18506 , n17555 );
and ( n21237 , n18203 , n17553 );
nor ( n21238 , n21236 , n21237 );
xnor ( n21239 , n21238 , n17457 );
and ( n21240 , n21234 , n21239 );
and ( n21241 , n21230 , n21239 );
or ( n21242 , n21235 , n21240 , n21241 );
and ( n21243 , n17530 , n18570 );
and ( n21244 , n17482 , n18568 );
nor ( n21245 , n21243 , n21244 );
xnor ( n21246 , n21245 , n18214 );
and ( n21247 , n18708 , n17315 );
not ( n21248 , n21247 );
and ( n21249 , n21248 , n17215 );
and ( n21250 , n21246 , n21249 );
and ( n21251 , n21242 , n21250 );
and ( n21252 , n17844 , n18077 );
and ( n21253 , n17530 , n18075 );
nor ( n21254 , n21252 , n21253 );
xnor ( n21255 , n21254 , n17919 );
and ( n21256 , n21250 , n21255 );
and ( n21257 , n21242 , n21255 );
or ( n21258 , n21251 , n21256 , n21257 );
xor ( n21259 , n21123 , n21127 );
xor ( n21260 , n21259 , n21132 );
and ( n21261 , n21258 , n21260 );
xor ( n21262 , n21139 , n21143 );
xor ( n21263 , n21262 , n21148 );
and ( n21264 , n21260 , n21263 );
and ( n21265 , n21258 , n21263 );
or ( n21266 , n21261 , n21264 , n21265 );
xor ( n21267 , n21135 , n21151 );
xor ( n21268 , n21267 , n21154 );
and ( n21269 , n21266 , n21268 );
xor ( n21270 , n21207 , n21209 );
xor ( n21271 , n21270 , n21212 );
and ( n21272 , n21268 , n21271 );
and ( n21273 , n21266 , n21271 );
or ( n21274 , n21269 , n21272 , n21273 );
and ( n21275 , n21226 , n21274 );
xor ( n21276 , n21266 , n21268 );
xor ( n21277 , n21276 , n21271 );
xor ( n21278 , n21246 , n21249 );
and ( n21279 , n17985 , n18077 );
and ( n21280 , n17844 , n18075 );
nor ( n21281 , n21279 , n21280 );
xnor ( n21282 , n21281 , n17919 );
and ( n21283 , n21278 , n21282 );
and ( n21284 , n18708 , n17317 );
and ( n21285 , n18654 , n17315 );
nor ( n21286 , n21284 , n21285 );
xnor ( n21287 , n21286 , n17215 );
and ( n21288 , n21282 , n21287 );
and ( n21289 , n21278 , n21287 );
or ( n21290 , n21283 , n21288 , n21289 );
xor ( n21291 , n21179 , n21183 );
xor ( n21292 , n21291 , n21188 );
and ( n21293 , n21290 , n21292 );
xor ( n21294 , n21196 , n21200 );
xor ( n21295 , n21294 , n21104 );
and ( n21296 , n21292 , n21295 );
and ( n21297 , n21290 , n21295 );
or ( n21298 , n21293 , n21296 , n21297 );
xor ( n21299 , n21175 , n21191 );
xor ( n21300 , n21299 , n21204 );
and ( n21301 , n21298 , n21300 );
xor ( n21302 , n21258 , n21260 );
xor ( n21303 , n21302 , n21263 );
and ( n21304 , n21300 , n21303 );
and ( n21305 , n21298 , n21303 );
or ( n21306 , n21301 , n21304 , n21305 );
and ( n21307 , n21277 , n21306 );
xor ( n21308 , n21298 , n21300 );
xor ( n21309 , n21308 , n21303 );
and ( n21310 , n17482 , n18698 );
and ( n21311 , n17327 , n18695 );
nor ( n21312 , n21310 , n21311 );
xnor ( n21313 , n21312 , n18211 );
and ( n21314 , n18145 , n18077 );
and ( n21315 , n17985 , n18075 );
nor ( n21316 , n21314 , n21315 );
xnor ( n21317 , n21316 , n17919 );
and ( n21318 , n21313 , n21317 );
and ( n21319 , n18654 , n17555 );
and ( n21320 , n18506 , n17553 );
nor ( n21321 , n21319 , n21320 );
xnor ( n21322 , n21321 , n17457 );
and ( n21323 , n21317 , n21322 );
and ( n21324 , n21313 , n21322 );
or ( n21325 , n21318 , n21323 , n21324 );
and ( n21326 , n17844 , n18570 );
and ( n21327 , n17530 , n18568 );
nor ( n21328 , n21326 , n21327 );
xnor ( n21329 , n21328 , n18214 );
and ( n21330 , n18203 , n17797 );
and ( n21331 , n18255 , n17795 );
nor ( n21332 , n21330 , n21331 );
xnor ( n21333 , n21332 , n17726 );
and ( n21334 , n21329 , n21333 );
and ( n21335 , n21333 , n21247 );
and ( n21336 , n21329 , n21247 );
or ( n21337 , n21334 , n21335 , n21336 );
and ( n21338 , n21325 , n21337 );
xor ( n21339 , n21230 , n21234 );
xor ( n21340 , n21339 , n21239 );
and ( n21341 , n21337 , n21340 );
and ( n21342 , n21325 , n21340 );
or ( n21343 , n21338 , n21341 , n21342 );
xor ( n21344 , n21242 , n21250 );
xor ( n21345 , n21344 , n21255 );
and ( n21346 , n21343 , n21345 );
xor ( n21347 , n21290 , n21292 );
xor ( n21348 , n21347 , n21295 );
and ( n21349 , n21345 , n21348 );
and ( n21350 , n21343 , n21348 );
or ( n21351 , n21346 , n21349 , n21350 );
and ( n21352 , n21309 , n21351 );
xor ( n21353 , n21278 , n21282 );
xor ( n21354 , n21353 , n21287 );
xor ( n21355 , n21325 , n21337 );
xor ( n21356 , n21355 , n21340 );
and ( n21357 , n21354 , n21356 );
xor ( n21358 , n21329 , n21333 );
xor ( n21359 , n21358 , n21247 );
and ( n21360 , n17530 , n18698 );
and ( n21361 , n17482 , n18695 );
nor ( n21362 , n21360 , n21361 );
xnor ( n21363 , n21362 , n18211 );
and ( n21364 , n18506 , n17797 );
and ( n21365 , n18203 , n17795 );
nor ( n21366 , n21364 , n21365 );
xnor ( n21367 , n21366 , n17726 );
and ( n21368 , n21363 , n21367 );
and ( n21369 , n18708 , n17555 );
and ( n21370 , n18654 , n17553 );
nor ( n21371 , n21369 , n21370 );
xnor ( n21372 , n21371 , n17457 );
and ( n21373 , n21367 , n21372 );
and ( n21374 , n21363 , n21372 );
or ( n21375 , n21368 , n21373 , n21374 );
and ( n21376 , n21359 , n21375 );
and ( n21377 , n17985 , n18570 );
and ( n21378 , n17844 , n18568 );
nor ( n21379 , n21377 , n21378 );
xnor ( n21380 , n21379 , n18214 );
and ( n21381 , n18708 , n17553 );
not ( n21382 , n21381 );
and ( n21383 , n21382 , n17457 );
and ( n21384 , n21380 , n21383 );
and ( n21385 , n21375 , n21384 );
and ( n21386 , n21359 , n21384 );
or ( n21387 , n21376 , n21385 , n21386 );
and ( n21388 , n21356 , n21387 );
and ( n21389 , n21354 , n21387 );
or ( n21390 , n21357 , n21388 , n21389 );
xor ( n21391 , n21343 , n21345 );
xor ( n21392 , n21391 , n21348 );
and ( n21393 , n21390 , n21392 );
xor ( n21394 , n21380 , n21383 );
and ( n21395 , n17844 , n18698 );
and ( n21396 , n17530 , n18695 );
nor ( n21397 , n21395 , n21396 );
xnor ( n21398 , n21397 , n18211 );
and ( n21399 , n18654 , n17797 );
and ( n21400 , n18506 , n17795 );
nor ( n21401 , n21399 , n21400 );
xnor ( n21402 , n21401 , n17726 );
and ( n21403 , n21398 , n21402 );
and ( n21404 , n21402 , n21381 );
and ( n21405 , n21398 , n21381 );
or ( n21406 , n21403 , n21404 , n21405 );
and ( n21407 , n21394 , n21406 );
and ( n21408 , n18255 , n18077 );
and ( n21409 , n18145 , n18075 );
nor ( n21410 , n21408 , n21409 );
xnor ( n21411 , n21410 , n17919 );
and ( n21412 , n21406 , n21411 );
and ( n21413 , n21394 , n21411 );
or ( n21414 , n21407 , n21412 , n21413 );
xor ( n21415 , n21313 , n21317 );
xor ( n21416 , n21415 , n21322 );
and ( n21417 , n21414 , n21416 );
xor ( n21418 , n21354 , n21356 );
xor ( n21419 , n21418 , n21387 );
and ( n21420 , n21417 , n21419 );
xor ( n21421 , n21359 , n21375 );
xor ( n21422 , n21421 , n21384 );
xor ( n21423 , n21414 , n21416 );
and ( n21424 , n21422 , n21423 );
and ( n21425 , n17985 , n18698 );
and ( n21426 , n17844 , n18695 );
nor ( n21427 , n21425 , n21426 );
xnor ( n21428 , n21427 , n18211 );
and ( n21429 , n18708 , n17795 );
not ( n21430 , n21429 );
and ( n21431 , n21430 , n17726 );
and ( n21432 , n21428 , n21431 );
and ( n21433 , n18145 , n18570 );
and ( n21434 , n17985 , n18568 );
nor ( n21435 , n21433 , n21434 );
xnor ( n21436 , n21435 , n18214 );
and ( n21437 , n21432 , n21436 );
and ( n21438 , n18203 , n18077 );
and ( n21439 , n18255 , n18075 );
nor ( n21440 , n21438 , n21439 );
xnor ( n21441 , n21440 , n17919 );
and ( n21442 , n21436 , n21441 );
and ( n21443 , n21432 , n21441 );
or ( n21444 , n21437 , n21442 , n21443 );
xor ( n21445 , n21363 , n21367 );
xor ( n21446 , n21445 , n21372 );
and ( n21447 , n21444 , n21446 );
xor ( n21448 , n21394 , n21406 );
xor ( n21449 , n21448 , n21411 );
and ( n21450 , n21446 , n21449 );
and ( n21451 , n21444 , n21449 );
or ( n21452 , n21447 , n21450 , n21451 );
and ( n21453 , n21423 , n21452 );
and ( n21454 , n21422 , n21452 );
or ( n21455 , n21424 , n21453 , n21454 );
and ( n21456 , n21419 , n21455 );
and ( n21457 , n21417 , n21455 );
or ( n21458 , n21420 , n21456 , n21457 );
and ( n21459 , n21392 , n21458 );
and ( n21460 , n21390 , n21458 );
or ( n21461 , n21393 , n21459 , n21460 );
and ( n21462 , n21351 , n21461 );
and ( n21463 , n21309 , n21461 );
or ( n21464 , n21352 , n21462 , n21463 );
and ( n21465 , n21306 , n21464 );
and ( n21466 , n21277 , n21464 );
or ( n21467 , n21307 , n21465 , n21466 );
and ( n21468 , n21274 , n21467 );
and ( n21469 , n21226 , n21467 );
or ( n21470 , n21275 , n21468 , n21469 );
and ( n21471 , n21223 , n21470 );
and ( n21472 , n21174 , n21470 );
or ( n21473 , n21224 , n21471 , n21472 );
and ( n21474 , n21171 , n21473 );
and ( n21475 , n21099 , n21473 );
or ( n21476 , n21172 , n21474 , n21475 );
and ( n21477 , n21096 , n21476 );
and ( n21478 , n21094 , n21476 );
or ( n21479 , n21097 , n21477 , n21478 );
and ( n21480 , n21034 , n21479 );
and ( n21481 , n21032 , n21479 );
or ( n21482 , n21035 , n21480 , n21481 );
and ( n21483 , n20963 , n21482 );
and ( n21484 , n20961 , n21482 );
or ( n21485 , n20964 , n21483 , n21484 );
and ( n21486 , n20889 , n21485 );
xor ( n21487 , n20889 , n21485 );
xor ( n21488 , n20961 , n20963 );
xor ( n21489 , n21488 , n21482 );
xor ( n21490 , n21032 , n21034 );
xor ( n21491 , n21490 , n21479 );
xor ( n21492 , n21094 , n21096 );
xor ( n21493 , n21492 , n21476 );
xor ( n21494 , n21099 , n21171 );
xor ( n21495 , n21494 , n21473 );
xor ( n21496 , n21174 , n21223 );
xor ( n21497 , n21496 , n21470 );
xor ( n21498 , n21226 , n21274 );
xor ( n21499 , n21498 , n21467 );
xor ( n21500 , n21277 , n21306 );
xor ( n21501 , n21500 , n21464 );
xor ( n21502 , n21309 , n21351 );
xor ( n21503 , n21502 , n21461 );
xor ( n21504 , n21390 , n21392 );
xor ( n21505 , n21504 , n21458 );
xor ( n21506 , n21417 , n21419 );
xor ( n21507 , n21506 , n21455 );
xor ( n21508 , n21422 , n21423 );
xor ( n21509 , n21508 , n21452 );
xor ( n21510 , n21444 , n21446 );
xor ( n21511 , n21510 , n21449 );
and ( n21512 , n18255 , n18570 );
and ( n21513 , n18145 , n18568 );
nor ( n21514 , n21512 , n21513 );
xnor ( n21515 , n21514 , n18214 );
and ( n21516 , n18506 , n18077 );
and ( n21517 , n18203 , n18075 );
nor ( n21518 , n21516 , n21517 );
xnor ( n21519 , n21518 , n17919 );
and ( n21520 , n21515 , n21519 );
and ( n21521 , n18708 , n17797 );
and ( n21522 , n18654 , n17795 );
nor ( n21523 , n21521 , n21522 );
xnor ( n21524 , n21523 , n17726 );
and ( n21525 , n21519 , n21524 );
and ( n21526 , n21515 , n21524 );
or ( n21527 , n21520 , n21525 , n21526 );
xor ( n21528 , n21398 , n21402 );
xor ( n21529 , n21528 , n21381 );
and ( n21530 , n21527 , n21529 );
xor ( n21531 , n21432 , n21436 );
xor ( n21532 , n21531 , n21441 );
and ( n21533 , n21529 , n21532 );
and ( n21534 , n21527 , n21532 );
or ( n21535 , n21530 , n21533 , n21534 );
and ( n21536 , n21511 , n21535 );
xor ( n21537 , n21511 , n21535 );
xor ( n21538 , n21428 , n21431 );
and ( n21539 , n18145 , n18698 );
and ( n21540 , n17985 , n18695 );
nor ( n21541 , n21539 , n21540 );
xnor ( n21542 , n21541 , n18211 );
and ( n21543 , n18203 , n18570 );
and ( n21544 , n18255 , n18568 );
nor ( n21545 , n21543 , n21544 );
xnor ( n21546 , n21545 , n18214 );
and ( n21547 , n21542 , n21546 );
and ( n21548 , n21546 , n21429 );
and ( n21549 , n21542 , n21429 );
or ( n21550 , n21547 , n21548 , n21549 );
and ( n21551 , n21538 , n21550 );
xor ( n21552 , n21515 , n21519 );
xor ( n21553 , n21552 , n21524 );
and ( n21554 , n21550 , n21553 );
and ( n21555 , n21538 , n21553 );
or ( n21556 , n21551 , n21554 , n21555 );
xor ( n21557 , n21527 , n21529 );
xor ( n21558 , n21557 , n21532 );
and ( n21559 , n21556 , n21558 );
xor ( n21560 , n21556 , n21558 );
xor ( n21561 , n21538 , n21550 );
xor ( n21562 , n21561 , n21553 );
and ( n21563 , n18255 , n18698 );
and ( n21564 , n18145 , n18695 );
nor ( n21565 , n21563 , n21564 );
xnor ( n21566 , n21565 , n18211 );
and ( n21567 , n18708 , n18075 );
not ( n21568 , n21567 );
and ( n21569 , n21568 , n17919 );
and ( n21570 , n21566 , n21569 );
and ( n21571 , n18654 , n18077 );
and ( n21572 , n18506 , n18075 );
nor ( n21573 , n21571 , n21572 );
xnor ( n21574 , n21573 , n17919 );
and ( n21575 , n21570 , n21574 );
xor ( n21576 , n21542 , n21546 );
xor ( n21577 , n21576 , n21429 );
and ( n21578 , n21574 , n21577 );
and ( n21579 , n21570 , n21577 );
or ( n21580 , n21575 , n21578 , n21579 );
and ( n21581 , n21562 , n21580 );
xor ( n21582 , n21562 , n21580 );
xor ( n21583 , n21570 , n21574 );
xor ( n21584 , n21583 , n21577 );
xor ( n21585 , n21566 , n21569 );
and ( n21586 , n18506 , n18570 );
and ( n21587 , n18203 , n18568 );
nor ( n21588 , n21586 , n21587 );
xnor ( n21589 , n21588 , n18214 );
and ( n21590 , n21585 , n21589 );
and ( n21591 , n18708 , n18077 );
and ( n21592 , n18654 , n18075 );
nor ( n21593 , n21591 , n21592 );
xnor ( n21594 , n21593 , n17919 );
and ( n21595 , n21589 , n21594 );
and ( n21596 , n21585 , n21594 );
or ( n21597 , n21590 , n21595 , n21596 );
and ( n21598 , n21584 , n21597 );
xor ( n21599 , n21584 , n21597 );
and ( n21600 , n18203 , n18698 );
and ( n21601 , n18255 , n18695 );
nor ( n21602 , n21600 , n21601 );
xnor ( n21603 , n21602 , n18211 );
and ( n21604 , n18654 , n18570 );
and ( n21605 , n18506 , n18568 );
nor ( n21606 , n21604 , n21605 );
xnor ( n21607 , n21606 , n18214 );
and ( n21608 , n21603 , n21607 );
and ( n21609 , n21607 , n21567 );
and ( n21610 , n21603 , n21567 );
or ( n21611 , n21608 , n21609 , n21610 );
xor ( n21612 , n21585 , n21589 );
xor ( n21613 , n21612 , n21594 );
and ( n21614 , n21611 , n21613 );
xor ( n21615 , n21611 , n21613 );
xor ( n21616 , n21603 , n21607 );
xor ( n21617 , n21616 , n21567 );
and ( n21618 , n18506 , n18698 );
and ( n21619 , n18203 , n18695 );
nor ( n21620 , n21618 , n21619 );
xnor ( n21621 , n21620 , n18211 );
and ( n21622 , n18708 , n18568 );
not ( n21623 , n21622 );
and ( n21624 , n21623 , n18214 );
and ( n21625 , n21621 , n21624 );
and ( n21626 , n21617 , n21625 );
xor ( n21627 , n21617 , n21625 );
and ( n21628 , n18708 , n18570 );
and ( n21629 , n18654 , n18568 );
nor ( n21630 , n21628 , n21629 );
xnor ( n21631 , n21630 , n18214 );
xor ( n21632 , n21621 , n21624 );
and ( n21633 , n21631 , n21632 );
xor ( n21634 , n21631 , n21632 );
and ( n21635 , n18654 , n18698 );
and ( n21636 , n18506 , n18695 );
nor ( n21637 , n21635 , n21636 );
xnor ( n21638 , n21637 , n18211 );
and ( n21639 , n21638 , n21622 );
xor ( n21640 , n21638 , n21622 );
and ( n21641 , n18708 , n18698 );
and ( n21642 , n18654 , n18695 );
nor ( n21643 , n21641 , n21642 );
xnor ( n21644 , n21643 , n18211 );
and ( n21645 , n18708 , n18695 );
not ( n21646 , n21645 );
and ( n21647 , n21646 , n18211 );
and ( n21648 , n21644 , n21647 );
and ( n21649 , n21640 , n21648 );
or ( n21650 , n21639 , n21649 );
and ( n21651 , n21634 , n21650 );
or ( n21652 , n21633 , n21651 );
and ( n21653 , n21627 , n21652 );
or ( n21654 , n21626 , n21653 );
and ( n21655 , n21615 , n21654 );
or ( n21656 , n21614 , n21655 );
and ( n21657 , n21599 , n21656 );
or ( n21658 , n21598 , n21657 );
and ( n21659 , n21582 , n21658 );
or ( n21660 , n21581 , n21659 );
and ( n21661 , n21560 , n21660 );
or ( n21662 , n21559 , n21661 );
and ( n21663 , n21537 , n21662 );
or ( n21664 , n21536 , n21663 );
and ( n21665 , n21509 , n21664 );
and ( n21666 , n21507 , n21665 );
and ( n21667 , n21505 , n21666 );
and ( n21668 , n21503 , n21667 );
and ( n21669 , n21501 , n21668 );
and ( n21670 , n21499 , n21669 );
and ( n21671 , n21497 , n21670 );
and ( n21672 , n21495 , n21671 );
and ( n21673 , n21493 , n21672 );
and ( n21674 , n21491 , n21673 );
and ( n21675 , n21489 , n21674 );
and ( n21676 , n21487 , n21675 );
or ( n21677 , n21486 , n21676 );
and ( n21678 , n20887 , n21677 );
and ( n21679 , n20885 , n21678 );
or ( n21680 , n20884 , n21679 );
and ( n21681 , n20691 , n21680 );
and ( n21682 , n20689 , n21681 );
or ( n21683 , n20688 , n21682 );
and ( n21684 , n20471 , n21683 );
or ( n21685 , n20470 , n21684 );
and ( n21686 , n20366 , n21685 );
and ( n21687 , n20364 , n21686 );
or ( n21688 , n20363 , n21687 );
and ( n21689 , n20185 , n21688 );
and ( n21690 , n20183 , n21689 );
and ( n21691 , n20181 , n21690 );
and ( n21692 , n20179 , n21691 );
or ( n21693 , n20178 , n21692 );
and ( n21694 , n19822 , n21693 );
or ( n21695 , n19821 , n21694 );
and ( n21696 , n19692 , n21695 );
or ( n21697 , n19691 , n21696 );
and ( n21698 , n19377 , n21697 );
and ( n21699 , n19375 , n21698 );
and ( n21700 , n19373 , n21699 );
or ( n21701 , n19372 , n21700 );
and ( n21702 , n19181 , n21701 );
and ( n21703 , n19179 , n21702 );
and ( n21704 , n19177 , n21703 );
and ( n21705 , n19175 , n21704 );
and ( n21706 , n19173 , n21705 );
and ( n21707 , n19171 , n21706 );
and ( n21708 , n19169 , n21707 );
and ( n21709 , n19167 , n21708 );
and ( n21710 , n19165 , n21709 );
and ( n21711 , n19163 , n21710 );
and ( n21712 , n19161 , n21711 );
and ( n21713 , n19159 , n21712 );
and ( n21714 , n19157 , n21713 );
and ( n21715 , n19155 , n21714 );
and ( n21716 , n19153 , n21715 );
and ( n21717 , n19151 , n21716 );
and ( n21718 , n19149 , n21717 );
and ( n21719 , n19147 , n21718 );
and ( n21720 , n19145 , n21719 );
and ( n21721 , n19143 , n21720 );
and ( n21722 , n19141 , n21721 );
and ( n21723 , n19139 , n21722 );
and ( n21724 , n19137 , n21723 );
xor ( n21725 , n19135 , n21724 );
buf ( n548986 , n21725 );
buf ( n548987 , n548986 );
buf ( n21728 , n548987 );
buf ( n548989 , n1184 );
buf ( n21730 , n548989 );
buf ( n548991 , n1185 );
buf ( n21732 , n548991 );
xor ( n21733 , n21730 , n21732 );
not ( n21734 , n21732 );
and ( n21735 , n21733 , n21734 );
and ( n21736 , n21728 , n21735 );
and ( n21737 , n16112 , n16116 );
and ( n21738 , n16116 , n16118 );
and ( n21739 , n16112 , n16118 );
or ( n21740 , n21737 , n21738 , n21739 );
and ( n21741 , n16066 , n16093 );
not ( n21742 , n21741 );
xnor ( n21743 , n21742 , n16101 );
xor ( n21744 , n21740 , n21743 );
and ( n21745 , n16096 , n16087 );
not ( n21746 , n21745 );
xor ( n21747 , n21744 , n21746 );
and ( n21748 , n16109 , n16110 );
and ( n21749 , n16110 , n16119 );
and ( n21750 , n16109 , n16119 );
or ( n21751 , n21748 , n21749 , n21750 );
xor ( n21752 , n21747 , n21751 );
and ( n21753 , n16120 , n16176 );
and ( n21754 , n16176 , n19134 );
and ( n21755 , n16120 , n19134 );
or ( n21756 , n21753 , n21754 , n21755 );
xor ( n21757 , n21752 , n21756 );
and ( n21758 , n19135 , n21724 );
xor ( n21759 , n21757 , n21758 );
buf ( n549020 , n21759 );
buf ( n549021 , n549020 );
buf ( n21762 , n549021 );
and ( n21763 , n21762 , n21732 );
nor ( n21764 , n21736 , n21763 );
xnor ( n21765 , n21764 , n21730 );
xor ( n21766 , n19155 , n21714 );
buf ( n549027 , n21766 );
buf ( n549028 , n549027 );
buf ( n21769 , n549028 );
buf ( n549030 , n1176 );
buf ( n21771 , n549030 );
buf ( n549032 , n1177 );
buf ( n21773 , n549032 );
xor ( n21774 , n21771 , n21773 );
buf ( n549035 , n1178 );
buf ( n21776 , n549035 );
xor ( n21777 , n21773 , n21776 );
not ( n21778 , n21777 );
and ( n21779 , n21774 , n21778 );
and ( n21780 , n21769 , n21779 );
xor ( n21781 , n19153 , n21715 );
buf ( n549042 , n21781 );
buf ( n549043 , n549042 );
buf ( n21784 , n549043 );
and ( n21785 , n21784 , n21777 );
nor ( n21786 , n21780 , n21785 );
and ( n21787 , n21773 , n21776 );
not ( n21788 , n21787 );
and ( n21789 , n21771 , n21788 );
xnor ( n21790 , n21786 , n21789 );
xor ( n21791 , n19171 , n21706 );
buf ( n549052 , n21791 );
buf ( n549053 , n549052 );
buf ( n21794 , n549053 );
buf ( n549055 , n1168 );
buf ( n21796 , n549055 );
buf ( n549057 , n1169 );
buf ( n21798 , n549057 );
xor ( n21799 , n21796 , n21798 );
buf ( n549060 , n1170 );
buf ( n21801 , n549060 );
xor ( n21802 , n21798 , n21801 );
not ( n21803 , n21802 );
and ( n21804 , n21799 , n21803 );
and ( n21805 , n21794 , n21804 );
xor ( n21806 , n19169 , n21707 );
buf ( n549067 , n21806 );
buf ( n549068 , n549067 );
buf ( n21809 , n549068 );
and ( n21810 , n21809 , n21802 );
nor ( n21811 , n21805 , n21810 );
and ( n21812 , n21798 , n21801 );
not ( n21813 , n21812 );
and ( n21814 , n21796 , n21813 );
xnor ( n21815 , n21811 , n21814 );
and ( n21816 , n21790 , n21815 );
xor ( n21817 , n19175 , n21704 );
buf ( n549078 , n21817 );
buf ( n549079 , n549078 );
buf ( n21820 , n549079 );
buf ( n549081 , n1166 );
buf ( n21822 , n549081 );
buf ( n549083 , n1167 );
buf ( n21824 , n549083 );
xor ( n21825 , n21822 , n21824 );
xor ( n21826 , n21824 , n21796 );
not ( n21827 , n21826 );
and ( n21828 , n21825 , n21827 );
and ( n21829 , n21820 , n21828 );
xor ( n21830 , n19173 , n21705 );
buf ( n549091 , n21830 );
buf ( n549092 , n549091 );
buf ( n21833 , n549092 );
and ( n21834 , n21833 , n21826 );
nor ( n21835 , n21829 , n21834 );
and ( n21836 , n21824 , n21796 );
not ( n21837 , n21836 );
and ( n21838 , n21822 , n21837 );
xnor ( n21839 , n21835 , n21838 );
and ( n21840 , n21815 , n21839 );
and ( n21841 , n21790 , n21839 );
or ( n21842 , n21816 , n21840 , n21841 );
xor ( n21843 , n19149 , n21717 );
buf ( n549104 , n21843 );
buf ( n549105 , n549104 );
buf ( n21846 , n549105 );
buf ( n549107 , n1179 );
buf ( n21848 , n549107 );
xor ( n21849 , n21776 , n21848 );
buf ( n549110 , n1180 );
buf ( n21851 , n549110 );
xor ( n21852 , n21848 , n21851 );
not ( n21853 , n21852 );
and ( n21854 , n21849 , n21853 );
and ( n21855 , n21846 , n21854 );
xor ( n21856 , n19147 , n21718 );
buf ( n549117 , n21856 );
buf ( n549118 , n549117 );
buf ( n21859 , n549118 );
and ( n21860 , n21859 , n21852 );
nor ( n21861 , n21855 , n21860 );
and ( n21862 , n21848 , n21851 );
not ( n21863 , n21862 );
and ( n21864 , n21776 , n21863 );
xnor ( n21865 , n21861 , n21864 );
and ( n21866 , n21842 , n21865 );
xor ( n21867 , n19181 , n21701 );
buf ( n549128 , n21867 );
buf ( n549129 , n549128 );
buf ( n21870 , n549129 );
buf ( n549131 , n1162 );
buf ( n21872 , n549131 );
buf ( n549133 , n1163 );
buf ( n21874 , n549133 );
xor ( n21875 , n21872 , n21874 );
buf ( n549136 , n1164 );
buf ( n21877 , n549136 );
xor ( n21878 , n21874 , n21877 );
not ( n21879 , n21878 );
and ( n21880 , n21875 , n21879 );
and ( n21881 , n21870 , n21880 );
xor ( n21882 , n19179 , n21702 );
buf ( n549143 , n21882 );
buf ( n549144 , n549143 );
buf ( n21885 , n549144 );
and ( n21886 , n21885 , n21878 );
nor ( n21887 , n21881 , n21886 );
and ( n21888 , n21874 , n21877 );
not ( n21889 , n21888 );
and ( n21890 , n21872 , n21889 );
xnor ( n21891 , n21887 , n21890 );
xor ( n21892 , n19375 , n21698 );
buf ( n549153 , n21892 );
buf ( n549154 , n549153 );
buf ( n21895 , n549154 );
buf ( n549156 , n1160 );
buf ( n21897 , n549156 );
buf ( n549158 , n1161 );
buf ( n21899 , n549158 );
xor ( n21900 , n21897 , n21899 );
xor ( n21901 , n21899 , n21872 );
not ( n21902 , n21901 );
and ( n21903 , n21900 , n21902 );
and ( n21904 , n21895 , n21903 );
xor ( n21905 , n19373 , n21699 );
buf ( n549166 , n21905 );
buf ( n549167 , n549166 );
buf ( n21908 , n549167 );
and ( n21909 , n21908 , n21901 );
nor ( n21910 , n21904 , n21909 );
and ( n21911 , n21899 , n21872 );
not ( n21912 , n21911 );
and ( n21913 , n21897 , n21912 );
xnor ( n21914 , n21910 , n21913 );
xor ( n21915 , n21891 , n21914 );
xor ( n21916 , n19692 , n21695 );
buf ( n549177 , n21916 );
buf ( n549178 , n549177 );
buf ( n21919 , n549178 );
buf ( n549180 , n1158 );
buf ( n21921 , n549180 );
buf ( n549182 , n1159 );
buf ( n21923 , n549182 );
xor ( n21924 , n21921 , n21923 );
xor ( n21925 , n21923 , n21897 );
not ( n21926 , n21925 );
and ( n21927 , n21924 , n21926 );
and ( n21928 , n21919 , n21927 );
xor ( n21929 , n19377 , n21697 );
buf ( n549190 , n21929 );
buf ( n549191 , n549190 );
buf ( n21932 , n549191 );
and ( n21933 , n21932 , n21925 );
nor ( n21934 , n21928 , n21933 );
and ( n21935 , n21923 , n21897 );
not ( n21936 , n21935 );
and ( n21937 , n21921 , n21936 );
xnor ( n21938 , n21934 , n21937 );
xor ( n21939 , n21915 , n21938 );
and ( n21940 , n21865 , n21939 );
and ( n21941 , n21842 , n21939 );
or ( n21942 , n21866 , n21940 , n21941 );
xor ( n21943 , n21765 , n21942 );
xor ( n21944 , n19161 , n21711 );
buf ( n549205 , n21944 );
buf ( n549206 , n549205 );
buf ( n21947 , n549206 );
buf ( n549208 , n1172 );
buf ( n21949 , n549208 );
buf ( n549210 , n1173 );
buf ( n21951 , n549210 );
xor ( n21952 , n21949 , n21951 );
buf ( n549213 , n1174 );
buf ( n21954 , n549213 );
xor ( n21955 , n21951 , n21954 );
not ( n21956 , n21955 );
and ( n21957 , n21952 , n21956 );
and ( n21958 , n21947 , n21957 );
xor ( n21959 , n19159 , n21712 );
buf ( n549220 , n21959 );
buf ( n549221 , n549220 );
buf ( n21962 , n549221 );
and ( n21963 , n21962 , n21955 );
nor ( n21964 , n21958 , n21963 );
and ( n21965 , n21951 , n21954 );
not ( n21966 , n21965 );
and ( n21967 , n21949 , n21966 );
xnor ( n21968 , n21964 , n21967 );
xor ( n21969 , n19165 , n21709 );
buf ( n549230 , n21969 );
buf ( n549231 , n549230 );
buf ( n21972 , n549231 );
buf ( n549233 , n1171 );
buf ( n21974 , n549233 );
xor ( n21975 , n21801 , n21974 );
xor ( n21976 , n21974 , n21949 );
not ( n21977 , n21976 );
and ( n21978 , n21975 , n21977 );
and ( n21979 , n21972 , n21978 );
xor ( n21980 , n19163 , n21710 );
buf ( n549241 , n21980 );
buf ( n549242 , n549241 );
buf ( n21983 , n549242 );
and ( n21984 , n21983 , n21976 );
nor ( n21985 , n21979 , n21984 );
and ( n21986 , n21974 , n21949 );
not ( n21987 , n21986 );
and ( n21988 , n21801 , n21987 );
xnor ( n21989 , n21985 , n21988 );
and ( n21990 , n21968 , n21989 );
and ( n21991 , n21809 , n21804 );
xor ( n21992 , n19167 , n21708 );
buf ( n549253 , n21992 );
buf ( n549254 , n549253 );
buf ( n21995 , n549254 );
and ( n21996 , n21995 , n21802 );
nor ( n21997 , n21991 , n21996 );
xnor ( n21998 , n21997 , n21814 );
and ( n21999 , n21989 , n21998 );
and ( n22000 , n21968 , n21998 );
or ( n22001 , n21990 , n21999 , n22000 );
and ( n22002 , n21859 , n21854 );
xor ( n22003 , n19145 , n21719 );
buf ( n549264 , n22003 );
buf ( n549265 , n549264 );
buf ( n22006 , n549265 );
and ( n22007 , n22006 , n21852 );
nor ( n22008 , n22002 , n22007 );
xnor ( n22009 , n22008 , n21864 );
xor ( n22010 , n22001 , n22009 );
xor ( n22011 , n19822 , n21693 );
buf ( n549272 , n22011 );
buf ( n549273 , n549272 );
buf ( n22014 , n549273 );
buf ( n549275 , n1156 );
buf ( n22016 , n549275 );
buf ( n549277 , n1157 );
buf ( n22018 , n549277 );
xor ( n22019 , n22016 , n22018 );
xor ( n22020 , n22018 , n21921 );
not ( n22021 , n22020 );
and ( n22022 , n22019 , n22021 );
and ( n22023 , n22014 , n22022 );
and ( n22024 , n21919 , n22020 );
nor ( n22025 , n22023 , n22024 );
and ( n22026 , n22018 , n21921 );
not ( n22027 , n22026 );
and ( n22028 , n22016 , n22027 );
xnor ( n22029 , n22025 , n22028 );
xor ( n22030 , n20183 , n21689 );
buf ( n549291 , n22030 );
buf ( n549292 , n549291 );
buf ( n22033 , n549292 );
buf ( n549294 , n1154 );
buf ( n22035 , n549294 );
and ( n22036 , n22033 , n22035 );
xor ( n22037 , n22029 , n22036 );
xor ( n22038 , n20179 , n21691 );
buf ( n549299 , n22038 );
buf ( n549300 , n549299 );
buf ( n22041 , n549300 );
and ( n22042 , n22041 , n22022 );
and ( n22043 , n22014 , n22020 );
nor ( n22044 , n22042 , n22043 );
xnor ( n22045 , n22044 , n22028 );
xor ( n22046 , n20185 , n21688 );
buf ( n549307 , n22046 );
buf ( n549308 , n549307 );
buf ( n22049 , n549308 );
and ( n22050 , n22049 , n22035 );
and ( n22051 , n22045 , n22050 );
xor ( n22052 , n22037 , n22051 );
xor ( n22053 , n20181 , n21690 );
buf ( n549314 , n22053 );
buf ( n549315 , n549314 );
buf ( n22056 , n549315 );
buf ( n549317 , n1155 );
buf ( n22058 , n549317 );
xor ( n22059 , n22035 , n22058 );
xor ( n22060 , n22058 , n22016 );
not ( n22061 , n22060 );
and ( n22062 , n22059 , n22061 );
and ( n22063 , n22056 , n22062 );
and ( n22064 , n22041 , n22060 );
nor ( n22065 , n22063 , n22064 );
and ( n22066 , n22058 , n22016 );
not ( n22067 , n22066 );
and ( n22068 , n22035 , n22067 );
xnor ( n22069 , n22065 , n22068 );
xor ( n22070 , n22052 , n22069 );
xor ( n22071 , n22010 , n22070 );
xor ( n22072 , n21943 , n22071 );
and ( n22073 , n22049 , n22022 );
and ( n22074 , n22033 , n22020 );
nor ( n22075 , n22073 , n22074 );
xnor ( n22076 , n22075 , n22028 );
xor ( n22077 , n20471 , n21683 );
buf ( n549338 , n22077 );
buf ( n549339 , n549338 );
buf ( n22080 , n549339 );
and ( n22081 , n22080 , n22035 );
xor ( n22082 , n22076 , n22081 );
xor ( n22083 , n20364 , n21686 );
buf ( n549344 , n22083 );
buf ( n549345 , n549344 );
buf ( n22086 , n549345 );
and ( n22087 , n22086 , n22022 );
and ( n22088 , n22049 , n22020 );
nor ( n22089 , n22087 , n22088 );
xnor ( n22090 , n22089 , n22028 );
xor ( n22091 , n20689 , n21681 );
buf ( n549352 , n22091 );
buf ( n549353 , n549352 );
buf ( n22094 , n549353 );
and ( n22095 , n22094 , n22035 );
and ( n22096 , n22090 , n22095 );
and ( n22097 , n22082 , n22096 );
xor ( n22098 , n20366 , n21685 );
buf ( n549359 , n22098 );
buf ( n549360 , n549359 );
buf ( n22101 , n549360 );
and ( n22102 , n22101 , n22062 );
and ( n22103 , n22086 , n22060 );
nor ( n22104 , n22102 , n22103 );
xnor ( n22105 , n22104 , n22068 );
and ( n22106 , n22096 , n22105 );
and ( n22107 , n22082 , n22105 );
or ( n22108 , n22097 , n22106 , n22107 );
and ( n22109 , n21809 , n21978 );
and ( n22110 , n21995 , n21976 );
nor ( n22111 , n22109 , n22110 );
xnor ( n22112 , n22111 , n21988 );
and ( n22113 , n22108 , n22112 );
and ( n22114 , n21895 , n21880 );
and ( n22115 , n21908 , n21878 );
nor ( n22116 , n22114 , n22115 );
xnor ( n22117 , n22116 , n21890 );
and ( n22118 , n22112 , n22117 );
and ( n22119 , n22108 , n22117 );
or ( n22120 , n22113 , n22118 , n22119 );
xor ( n22121 , n19139 , n21722 );
buf ( n549382 , n22121 );
buf ( n549383 , n549382 );
buf ( n22124 , n549383 );
and ( n22125 , n22124 , n21735 );
xor ( n22126 , n19137 , n21723 );
buf ( n549387 , n22126 );
buf ( n549388 , n549387 );
buf ( n22129 , n549388 );
and ( n22130 , n22129 , n21732 );
nor ( n22131 , n22125 , n22130 );
xnor ( n22132 , n22131 , n21730 );
and ( n22133 , n22120 , n22132 );
xor ( n22134 , n19151 , n21716 );
buf ( n549395 , n22134 );
buf ( n549396 , n549395 );
buf ( n22137 , n549396 );
and ( n22138 , n22137 , n21854 );
and ( n22139 , n21846 , n21852 );
nor ( n22140 , n22138 , n22139 );
xnor ( n22141 , n22140 , n21864 );
and ( n22142 , n22132 , n22141 );
and ( n22143 , n22120 , n22141 );
or ( n22144 , n22133 , n22142 , n22143 );
xor ( n22145 , n19157 , n21713 );
buf ( n549406 , n22145 );
buf ( n549407 , n549406 );
buf ( n22148 , n549407 );
and ( n22149 , n22148 , n21779 );
and ( n22150 , n21769 , n21777 );
nor ( n22151 , n22149 , n22150 );
xnor ( n22152 , n22151 , n21789 );
and ( n22153 , n21972 , n21957 );
and ( n22154 , n21983 , n21955 );
nor ( n22155 , n22153 , n22154 );
xnor ( n22156 , n22155 , n21967 );
and ( n22157 , n22152 , n22156 );
and ( n22158 , n22086 , n22062 );
and ( n22159 , n22049 , n22060 );
nor ( n22160 , n22158 , n22159 );
xnor ( n22161 , n22160 , n22068 );
and ( n22162 , n22101 , n22035 );
xor ( n22163 , n22161 , n22162 );
and ( n22164 , n22076 , n22081 );
xor ( n22165 , n22163 , n22164 );
and ( n22166 , n22041 , n21927 );
and ( n22167 , n22014 , n21925 );
nor ( n22168 , n22166 , n22167 );
xnor ( n22169 , n22168 , n21937 );
xor ( n22170 , n22165 , n22169 );
and ( n22171 , n22156 , n22170 );
and ( n22172 , n22152 , n22170 );
or ( n22173 , n22157 , n22171 , n22172 );
and ( n22174 , n22163 , n22164 );
and ( n22175 , n22164 , n22169 );
and ( n22176 , n22163 , n22169 );
or ( n22177 , n22174 , n22175 , n22176 );
and ( n22178 , n21995 , n21978 );
and ( n22179 , n21972 , n21976 );
nor ( n22180 , n22178 , n22179 );
xnor ( n22181 , n22180 , n21988 );
xor ( n22182 , n22177 , n22181 );
and ( n22183 , n21908 , n21880 );
and ( n22184 , n21870 , n21878 );
nor ( n22185 , n22183 , n22184 );
xnor ( n22186 , n22185 , n21890 );
xor ( n22187 , n22182 , n22186 );
and ( n22188 , n22173 , n22187 );
buf ( n549449 , n1165 );
buf ( n22190 , n549449 );
xor ( n22191 , n21877 , n22190 );
xor ( n22192 , n22190 , n21822 );
not ( n22193 , n22192 );
and ( n22194 , n22191 , n22193 );
and ( n22195 , n21870 , n22194 );
and ( n22196 , n21885 , n22192 );
nor ( n22197 , n22195 , n22196 );
and ( n22198 , n22190 , n21822 );
not ( n22199 , n22198 );
and ( n22200 , n21877 , n22199 );
xnor ( n22201 , n22197 , n22200 );
and ( n22202 , n21919 , n21903 );
and ( n22203 , n21932 , n21901 );
nor ( n22204 , n22202 , n22203 );
xnor ( n22205 , n22204 , n21913 );
and ( n22206 , n22201 , n22205 );
and ( n22207 , n22033 , n22022 );
and ( n22208 , n22056 , n22020 );
nor ( n22209 , n22207 , n22208 );
xnor ( n22210 , n22209 , n22028 );
and ( n22211 , n22205 , n22210 );
and ( n22212 , n22201 , n22210 );
or ( n22213 , n22206 , n22211 , n22212 );
and ( n22214 , n21983 , n21957 );
and ( n22215 , n21947 , n21955 );
nor ( n22216 , n22214 , n22215 );
xnor ( n22217 , n22216 , n21967 );
xor ( n22218 , n22213 , n22217 );
and ( n22219 , n22049 , n22062 );
and ( n22220 , n22033 , n22060 );
nor ( n22221 , n22219 , n22220 );
xnor ( n22222 , n22221 , n22068 );
and ( n22223 , n22086 , n22035 );
xor ( n22224 , n22222 , n22223 );
and ( n22225 , n22161 , n22162 );
xor ( n22226 , n22224 , n22225 );
and ( n22227 , n22014 , n21927 );
and ( n22228 , n21919 , n21925 );
nor ( n22229 , n22227 , n22228 );
xnor ( n22230 , n22229 , n21937 );
xor ( n22231 , n22226 , n22230 );
xor ( n22232 , n22218 , n22231 );
and ( n22233 , n22187 , n22232 );
and ( n22234 , n22173 , n22232 );
or ( n22235 , n22188 , n22233 , n22234 );
and ( n22236 , n22144 , n22235 );
and ( n22237 , n22129 , n21735 );
and ( n22238 , n21728 , n21732 );
nor ( n22239 , n22237 , n22238 );
xnor ( n22240 , n22239 , n21730 );
xor ( n22241 , n19141 , n21721 );
buf ( n549502 , n22241 );
buf ( n549503 , n549502 );
buf ( n22244 , n549503 );
buf ( n549505 , n1182 );
buf ( n22246 , n549505 );
buf ( n549507 , n1183 );
buf ( n22248 , n549507 );
xor ( n22249 , n22246 , n22248 );
xor ( n22250 , n22248 , n21730 );
not ( n22251 , n22250 );
and ( n22252 , n22249 , n22251 );
and ( n22253 , n22244 , n22252 );
and ( n22254 , n22124 , n22250 );
nor ( n22255 , n22253 , n22254 );
and ( n22256 , n22248 , n21730 );
not ( n22257 , n22256 );
and ( n22258 , n22246 , n22257 );
xnor ( n22259 , n22255 , n22258 );
xor ( n22260 , n22240 , n22259 );
and ( n22261 , n22224 , n22225 );
and ( n22262 , n22225 , n22230 );
and ( n22263 , n22224 , n22230 );
or ( n22264 , n22261 , n22262 , n22263 );
and ( n22265 , n21833 , n21828 );
and ( n22266 , n21794 , n21826 );
nor ( n22267 , n22265 , n22266 );
xnor ( n22268 , n22267 , n21838 );
xor ( n22269 , n22264 , n22268 );
xor ( n22270 , n19177 , n21703 );
buf ( n549531 , n22270 );
buf ( n549532 , n549531 );
buf ( n22273 , n549532 );
and ( n22274 , n22273 , n22194 );
and ( n22275 , n21820 , n22192 );
nor ( n22276 , n22274 , n22275 );
xnor ( n22277 , n22276 , n22200 );
xor ( n22278 , n22269 , n22277 );
xor ( n22279 , n22260 , n22278 );
and ( n22280 , n22235 , n22279 );
and ( n22281 , n22144 , n22279 );
or ( n22282 , n22236 , n22280 , n22281 );
xor ( n22283 , n22072 , n22282 );
and ( n22284 , n21885 , n22194 );
and ( n22285 , n22273 , n22192 );
nor ( n22286 , n22284 , n22285 );
xnor ( n22287 , n22286 , n22200 );
and ( n22288 , n21932 , n21903 );
and ( n22289 , n21895 , n21901 );
nor ( n22290 , n22288 , n22289 );
xnor ( n22291 , n22290 , n21913 );
and ( n22292 , n22287 , n22291 );
and ( n22293 , n22056 , n22022 );
and ( n22294 , n22041 , n22020 );
nor ( n22295 , n22293 , n22294 );
xnor ( n22296 , n22295 , n22028 );
and ( n22297 , n22291 , n22296 );
and ( n22298 , n22287 , n22296 );
or ( n22299 , n22292 , n22297 , n22298 );
buf ( n549560 , n1181 );
buf ( n22301 , n549560 );
xor ( n22302 , n21851 , n22301 );
xor ( n22303 , n22301 , n22246 );
not ( n22304 , n22303 );
and ( n22305 , n22302 , n22304 );
and ( n22306 , n22006 , n22305 );
xor ( n22307 , n19143 , n21720 );
buf ( n549568 , n22307 );
buf ( n549569 , n549568 );
buf ( n22310 , n549569 );
and ( n22311 , n22310 , n22303 );
nor ( n22312 , n22306 , n22311 );
and ( n22313 , n22301 , n22246 );
not ( n22314 , n22313 );
and ( n22315 , n21851 , n22314 );
xnor ( n22316 , n22312 , n22315 );
and ( n22317 , n22299 , n22316 );
buf ( n549578 , n1175 );
buf ( n22319 , n549578 );
xor ( n22320 , n21954 , n22319 );
xor ( n22321 , n22319 , n21771 );
not ( n22322 , n22321 );
and ( n22323 , n22320 , n22322 );
and ( n22324 , n22148 , n22323 );
and ( n22325 , n21769 , n22321 );
nor ( n22326 , n22324 , n22325 );
and ( n22327 , n22319 , n21771 );
not ( n22328 , n22327 );
and ( n22329 , n21954 , n22328 );
xnor ( n22330 , n22326 , n22329 );
and ( n22331 , n22316 , n22330 );
and ( n22332 , n22299 , n22330 );
or ( n22333 , n22317 , n22331 , n22332 );
and ( n22334 , n22124 , n22252 );
and ( n22335 , n22129 , n22250 );
nor ( n22336 , n22334 , n22335 );
xnor ( n22337 , n22336 , n22258 );
xor ( n22338 , n22333 , n22337 );
and ( n22339 , n21995 , n21804 );
and ( n22340 , n21972 , n21802 );
nor ( n22341 , n22339 , n22340 );
xnor ( n22342 , n22341 , n21814 );
and ( n22343 , n21794 , n21828 );
and ( n22344 , n21809 , n21826 );
nor ( n22345 , n22343 , n22344 );
xnor ( n22346 , n22345 , n21838 );
xor ( n22347 , n22342 , n22346 );
and ( n22348 , n21820 , n22194 );
and ( n22349 , n21833 , n22192 );
nor ( n22350 , n22348 , n22349 );
xnor ( n22351 , n22350 , n22200 );
xor ( n22352 , n22347 , n22351 );
xor ( n22353 , n22338 , n22352 );
and ( n22354 , n22264 , n22268 );
and ( n22355 , n22268 , n22277 );
and ( n22356 , n22264 , n22277 );
or ( n22357 , n22354 , n22355 , n22356 );
and ( n22358 , n22310 , n22305 );
and ( n22359 , n22244 , n22303 );
nor ( n22360 , n22358 , n22359 );
xnor ( n22361 , n22360 , n22315 );
xor ( n22362 , n22357 , n22361 );
and ( n22363 , n21885 , n21880 );
and ( n22364 , n22273 , n21878 );
nor ( n22365 , n22363 , n22364 );
xnor ( n22366 , n22365 , n21890 );
and ( n22367 , n21908 , n21903 );
and ( n22368 , n21870 , n21901 );
nor ( n22369 , n22367 , n22368 );
xnor ( n22370 , n22369 , n21913 );
xor ( n22371 , n22366 , n22370 );
and ( n22372 , n21932 , n21927 );
and ( n22373 , n21895 , n21925 );
nor ( n22374 , n22372 , n22373 );
xnor ( n22375 , n22374 , n21937 );
xor ( n22376 , n22371 , n22375 );
xor ( n22377 , n22362 , n22376 );
xor ( n22378 , n22353 , n22377 );
and ( n22379 , n22240 , n22259 );
and ( n22380 , n22259 , n22278 );
and ( n22381 , n22240 , n22278 );
or ( n22382 , n22379 , n22380 , n22381 );
xor ( n22383 , n22378 , n22382 );
xor ( n22384 , n22283 , n22383 );
and ( n22385 , n21820 , n21804 );
and ( n22386 , n21833 , n21802 );
nor ( n22387 , n22385 , n22386 );
xnor ( n22388 , n22387 , n21814 );
and ( n22389 , n21885 , n21828 );
and ( n22390 , n22273 , n21826 );
nor ( n22391 , n22389 , n22390 );
xnor ( n22392 , n22391 , n21838 );
and ( n22393 , n22388 , n22392 );
and ( n22394 , n21932 , n21880 );
and ( n22395 , n21895 , n21878 );
nor ( n22396 , n22394 , n22395 );
xnor ( n22397 , n22396 , n21890 );
and ( n22398 , n22392 , n22397 );
and ( n22399 , n22388 , n22397 );
or ( n22400 , n22393 , n22398 , n22399 );
xor ( n22401 , n22090 , n22095 );
and ( n22402 , n22094 , n22062 );
and ( n22403 , n22080 , n22060 );
nor ( n22404 , n22402 , n22403 );
xnor ( n22405 , n22404 , n22068 );
xor ( n22406 , n20691 , n21680 );
buf ( n549667 , n22406 );
buf ( n549668 , n549667 );
buf ( n22409 , n549668 );
and ( n22410 , n22409 , n22035 );
and ( n22411 , n22405 , n22410 );
and ( n22412 , n22401 , n22411 );
and ( n22413 , n22080 , n22062 );
and ( n22414 , n22101 , n22060 );
nor ( n22415 , n22413 , n22414 );
xnor ( n22416 , n22415 , n22068 );
and ( n22417 , n22411 , n22416 );
and ( n22418 , n22401 , n22416 );
or ( n22419 , n22412 , n22417 , n22418 );
and ( n22420 , n21995 , n21957 );
and ( n22421 , n21972 , n21955 );
nor ( n22422 , n22420 , n22421 );
xnor ( n22423 , n22422 , n21967 );
and ( n22424 , n22419 , n22423 );
and ( n22425 , n21794 , n21978 );
and ( n22426 , n21809 , n21976 );
nor ( n22427 , n22425 , n22426 );
xnor ( n22428 , n22427 , n21988 );
and ( n22429 , n22423 , n22428 );
and ( n22430 , n22419 , n22428 );
or ( n22431 , n22424 , n22429 , n22430 );
and ( n22432 , n22400 , n22431 );
and ( n22433 , n21784 , n21854 );
and ( n22434 , n22137 , n21852 );
nor ( n22435 , n22433 , n22434 );
xnor ( n22436 , n22435 , n21864 );
and ( n22437 , n22431 , n22436 );
and ( n22438 , n22400 , n22436 );
or ( n22439 , n22432 , n22437 , n22438 );
and ( n22440 , n21908 , n22194 );
and ( n22441 , n21870 , n22192 );
nor ( n22442 , n22440 , n22441 );
xnor ( n22443 , n22442 , n22200 );
and ( n22444 , n22014 , n21903 );
and ( n22445 , n21919 , n21901 );
nor ( n22446 , n22444 , n22445 );
xnor ( n22447 , n22446 , n21913 );
and ( n22448 , n22443 , n22447 );
and ( n22449 , n22056 , n21927 );
and ( n22450 , n22041 , n21925 );
nor ( n22451 , n22449 , n22450 );
xnor ( n22452 , n22451 , n21937 );
and ( n22453 , n22447 , n22452 );
and ( n22454 , n22443 , n22452 );
or ( n22455 , n22448 , n22453 , n22454 );
and ( n22456 , n22006 , n22252 );
and ( n22457 , n22310 , n22250 );
nor ( n22458 , n22456 , n22457 );
xnor ( n22459 , n22458 , n22258 );
and ( n22460 , n22455 , n22459 );
xor ( n22461 , n22201 , n22205 );
xor ( n22462 , n22461 , n22210 );
and ( n22463 , n22459 , n22462 );
and ( n22464 , n22455 , n22462 );
or ( n22465 , n22460 , n22463 , n22464 );
and ( n22466 , n22439 , n22465 );
and ( n22467 , n22310 , n22252 );
and ( n22468 , n22244 , n22250 );
nor ( n22469 , n22467 , n22468 );
xnor ( n22470 , n22469 , n22258 );
and ( n22471 , n21962 , n22323 );
and ( n22472 , n22148 , n22321 );
nor ( n22473 , n22471 , n22472 );
xnor ( n22474 , n22473 , n22329 );
xor ( n22475 , n22470 , n22474 );
xor ( n22476 , n22287 , n22291 );
xor ( n22477 , n22476 , n22296 );
xor ( n22478 , n22475 , n22477 );
and ( n22479 , n22465 , n22478 );
and ( n22480 , n22439 , n22478 );
or ( n22481 , n22466 , n22479 , n22480 );
xor ( n22482 , n21842 , n21865 );
xor ( n22483 , n22482 , n21939 );
and ( n22484 , n22481 , n22483 );
and ( n22485 , n22213 , n22217 );
and ( n22486 , n22217 , n22231 );
and ( n22487 , n22213 , n22231 );
or ( n22488 , n22485 , n22486 , n22487 );
xor ( n22489 , n21968 , n21989 );
xor ( n22490 , n22489 , n21998 );
xor ( n22491 , n22488 , n22490 );
xor ( n22492 , n22299 , n22316 );
xor ( n22493 , n22492 , n22330 );
xor ( n22494 , n22491 , n22493 );
and ( n22495 , n22483 , n22494 );
and ( n22496 , n22481 , n22494 );
or ( n22497 , n22484 , n22495 , n22496 );
and ( n22498 , n22488 , n22490 );
and ( n22499 , n22490 , n22493 );
and ( n22500 , n22488 , n22493 );
or ( n22501 , n22498 , n22499 , n22500 );
and ( n22502 , n22470 , n22474 );
and ( n22503 , n22474 , n22477 );
and ( n22504 , n22470 , n22477 );
or ( n22505 , n22502 , n22503 , n22504 );
and ( n22506 , n21947 , n22323 );
and ( n22507 , n21962 , n22321 );
nor ( n22508 , n22506 , n22507 );
xnor ( n22509 , n22508 , n22329 );
and ( n22510 , n21833 , n21804 );
and ( n22511 , n21794 , n21802 );
nor ( n22512 , n22510 , n22511 );
xnor ( n22513 , n22512 , n21814 );
and ( n22514 , n22509 , n22513 );
and ( n22515 , n22273 , n21828 );
and ( n22516 , n21820 , n21826 );
nor ( n22517 , n22515 , n22516 );
xnor ( n22518 , n22517 , n21838 );
and ( n22519 , n22513 , n22518 );
and ( n22520 , n22509 , n22518 );
or ( n22521 , n22514 , n22519 , n22520 );
and ( n22522 , n21859 , n22305 );
and ( n22523 , n22006 , n22303 );
nor ( n22524 , n22522 , n22523 );
xnor ( n22525 , n22524 , n22315 );
and ( n22526 , n22521 , n22525 );
xor ( n22527 , n21790 , n21815 );
xor ( n22528 , n22527 , n21839 );
and ( n22529 , n22525 , n22528 );
and ( n22530 , n22521 , n22528 );
or ( n22531 , n22526 , n22529 , n22530 );
and ( n22532 , n22505 , n22531 );
and ( n22533 , n22177 , n22181 );
and ( n22534 , n22181 , n22186 );
and ( n22535 , n22177 , n22186 );
or ( n22536 , n22533 , n22534 , n22535 );
and ( n22537 , n21784 , n21779 );
and ( n22538 , n22137 , n21777 );
nor ( n22539 , n22537 , n22538 );
xnor ( n22540 , n22539 , n21789 );
xor ( n22541 , n22536 , n22540 );
xor ( n22542 , n22045 , n22050 );
and ( n22543 , n22222 , n22223 );
xor ( n22544 , n22542 , n22543 );
and ( n22545 , n22033 , n22062 );
and ( n22546 , n22056 , n22060 );
nor ( n22547 , n22545 , n22546 );
xnor ( n22548 , n22547 , n22068 );
xor ( n22549 , n22544 , n22548 );
xor ( n22550 , n22541 , n22549 );
and ( n22551 , n22531 , n22550 );
and ( n22552 , n22505 , n22550 );
or ( n22553 , n22532 , n22551 , n22552 );
xor ( n22554 , n22501 , n22553 );
and ( n22555 , n22536 , n22540 );
and ( n22556 , n22540 , n22549 );
and ( n22557 , n22536 , n22549 );
or ( n22558 , n22555 , n22556 , n22557 );
and ( n22559 , n21891 , n21914 );
and ( n22560 , n21914 , n21938 );
and ( n22561 , n21891 , n21938 );
or ( n22562 , n22559 , n22560 , n22561 );
and ( n22563 , n22137 , n21779 );
and ( n22564 , n21846 , n21777 );
nor ( n22565 , n22563 , n22564 );
xnor ( n22566 , n22565 , n21789 );
xor ( n22567 , n22562 , n22566 );
and ( n22568 , n21962 , n21957 );
and ( n22569 , n22148 , n21955 );
nor ( n22570 , n22568 , n22569 );
xnor ( n22571 , n22570 , n21967 );
xor ( n22572 , n22567 , n22571 );
xor ( n22573 , n22558 , n22572 );
and ( n22574 , n22542 , n22543 );
and ( n22575 , n22543 , n22548 );
and ( n22576 , n22542 , n22548 );
or ( n22577 , n22574 , n22575 , n22576 );
and ( n22578 , n21769 , n22323 );
and ( n22579 , n21784 , n22321 );
nor ( n22580 , n22578 , n22579 );
xnor ( n22581 , n22580 , n22329 );
xor ( n22582 , n22577 , n22581 );
and ( n22583 , n21983 , n21978 );
and ( n22584 , n21947 , n21976 );
nor ( n22585 , n22583 , n22584 );
xnor ( n22586 , n22585 , n21988 );
xor ( n22587 , n22582 , n22586 );
xor ( n22588 , n22573 , n22587 );
xor ( n22589 , n22554 , n22588 );
xor ( n22590 , n22497 , n22589 );
and ( n22591 , n22384 , n22590 );
and ( n22592 , n21769 , n21854 );
and ( n22593 , n21784 , n21852 );
nor ( n22594 , n22592 , n22593 );
xnor ( n22595 , n22594 , n21864 );
and ( n22596 , n21983 , n22323 );
and ( n22597 , n21947 , n22321 );
nor ( n22598 , n22596 , n22597 );
xnor ( n22599 , n22598 , n22329 );
and ( n22600 , n22595 , n22599 );
xor ( n22601 , n22082 , n22096 );
xor ( n22602 , n22601 , n22105 );
and ( n22603 , n22599 , n22602 );
and ( n22604 , n22595 , n22602 );
or ( n22605 , n22600 , n22603 , n22604 );
and ( n22606 , n22244 , n21735 );
and ( n22607 , n22124 , n21732 );
nor ( n22608 , n22606 , n22607 );
xnor ( n22609 , n22608 , n21730 );
and ( n22610 , n22605 , n22609 );
and ( n22611 , n21846 , n22305 );
and ( n22612 , n21859 , n22303 );
nor ( n22613 , n22611 , n22612 );
xnor ( n22614 , n22613 , n22315 );
and ( n22615 , n22609 , n22614 );
and ( n22616 , n22605 , n22614 );
or ( n22617 , n22610 , n22615 , n22616 );
xor ( n22618 , n22120 , n22132 );
xor ( n22619 , n22618 , n22141 );
and ( n22620 , n22617 , n22619 );
xor ( n22621 , n22521 , n22525 );
xor ( n22622 , n22621 , n22528 );
and ( n22623 , n22619 , n22622 );
and ( n22624 , n22617 , n22622 );
or ( n22625 , n22620 , n22623 , n22624 );
xor ( n22626 , n22509 , n22513 );
xor ( n22627 , n22626 , n22518 );
xor ( n22628 , n22108 , n22112 );
xor ( n22629 , n22628 , n22117 );
and ( n22630 , n22627 , n22629 );
xor ( n22631 , n22152 , n22156 );
xor ( n22632 , n22631 , n22170 );
and ( n22633 , n22629 , n22632 );
and ( n22634 , n22627 , n22632 );
or ( n22635 , n22630 , n22633 , n22634 );
and ( n22636 , n21895 , n22194 );
and ( n22637 , n21908 , n22192 );
nor ( n22638 , n22636 , n22637 );
xnor ( n22639 , n22638 , n22200 );
and ( n22640 , n22041 , n21903 );
and ( n22641 , n22014 , n21901 );
nor ( n22642 , n22640 , n22641 );
xnor ( n22643 , n22642 , n21913 );
and ( n22644 , n22639 , n22643 );
and ( n22645 , n22033 , n21927 );
and ( n22646 , n22056 , n21925 );
nor ( n22647 , n22645 , n22646 );
xnor ( n22648 , n22647 , n21937 );
and ( n22649 , n22643 , n22648 );
and ( n22650 , n22639 , n22648 );
or ( n22651 , n22644 , n22649 , n22650 );
and ( n22652 , n22409 , n22062 );
and ( n22653 , n22094 , n22060 );
nor ( n22654 , n22652 , n22653 );
xnor ( n22655 , n22654 , n22068 );
xor ( n22656 , n20885 , n21678 );
buf ( n549917 , n22656 );
buf ( n549918 , n549917 );
buf ( n22659 , n549918 );
and ( n22660 , n22659 , n22035 );
and ( n22661 , n22655 , n22660 );
and ( n549922 , n22049 , n21927 );
and ( n22662 , n22033 , n21925 );
nor ( n22663 , n549922 , n22662 );
xnor ( n22664 , n22663 , n21937 );
and ( n22665 , n22661 , n22664 );
and ( n22666 , n22101 , n22022 );
and ( n22667 , n22086 , n22020 );
nor ( n22668 , n22666 , n22667 );
xnor ( n22669 , n22668 , n22028 );
and ( n22670 , n22664 , n22669 );
and ( n22671 , n22661 , n22669 );
or ( n22672 , n22665 , n22670 , n22671 );
and ( n22673 , n21870 , n21828 );
and ( n22674 , n21885 , n21826 );
nor ( n22675 , n22673 , n22674 );
xnor ( n22676 , n22675 , n21838 );
and ( n22677 , n22672 , n22676 );
and ( n22678 , n21919 , n21880 );
and ( n22679 , n21932 , n21878 );
nor ( n22680 , n22678 , n22679 );
xnor ( n22681 , n22680 , n21890 );
and ( n22682 , n22676 , n22681 );
and ( n22683 , n22672 , n22681 );
or ( n22684 , n22677 , n22682 , n22683 );
and ( n22685 , n22651 , n22684 );
and ( n22686 , n21962 , n21779 );
and ( n22687 , n22148 , n21777 );
nor ( n22688 , n22686 , n22687 );
xnor ( n22689 , n22688 , n21789 );
and ( n22690 , n22684 , n22689 );
and ( n22691 , n22651 , n22689 );
or ( n22692 , n22685 , n22690 , n22691 );
xor ( n22693 , n22405 , n22410 );
and ( n22694 , n22014 , n21880 );
and ( n22695 , n21919 , n21878 );
nor ( n22696 , n22694 , n22695 );
xnor ( n22697 , n22696 , n21890 );
and ( n22698 , n22693 , n22697 );
and ( n22699 , n22056 , n21903 );
and ( n22700 , n22041 , n21901 );
nor ( n22701 , n22699 , n22700 );
xnor ( n22702 , n22701 , n21913 );
and ( n22703 , n22697 , n22702 );
and ( n22704 , n22693 , n22702 );
or ( n22705 , n22698 , n22703 , n22704 );
and ( n22706 , n21809 , n21957 );
and ( n22707 , n21995 , n21955 );
nor ( n22708 , n22706 , n22707 );
xnor ( n22709 , n22708 , n21967 );
and ( n22710 , n22705 , n22709 );
and ( n22711 , n22273 , n21804 );
and ( n22712 , n21820 , n21802 );
nor ( n22713 , n22711 , n22712 );
xnor ( n22714 , n22713 , n21814 );
and ( n22715 , n22709 , n22714 );
and ( n22716 , n22705 , n22714 );
or ( n22717 , n22710 , n22715 , n22716 );
and ( n22718 , n22310 , n21735 );
and ( n22719 , n22244 , n21732 );
nor ( n22720 , n22718 , n22719 );
xnor ( n22721 , n22720 , n21730 );
and ( n22722 , n22717 , n22721 );
xor ( n22723 , n22443 , n22447 );
xor ( n22724 , n22723 , n22452 );
and ( n22725 , n22721 , n22724 );
and ( n22726 , n22717 , n22724 );
or ( n22727 , n22722 , n22725 , n22726 );
and ( n22728 , n22692 , n22727 );
xor ( n22729 , n22455 , n22459 );
xor ( n22730 , n22729 , n22462 );
and ( n22731 , n22727 , n22730 );
and ( n22732 , n22692 , n22730 );
or ( n22733 , n22728 , n22731 , n22732 );
and ( n22734 , n22635 , n22733 );
xor ( n22735 , n22173 , n22187 );
xor ( n22736 , n22735 , n22232 );
and ( n22737 , n22733 , n22736 );
and ( n22738 , n22635 , n22736 );
or ( n22739 , n22734 , n22737 , n22738 );
and ( n22740 , n22625 , n22739 );
xor ( n22741 , n22505 , n22531 );
xor ( n22742 , n22741 , n22550 );
and ( n22743 , n22739 , n22742 );
and ( n22744 , n22625 , n22742 );
or ( n22745 , n22740 , n22743 , n22744 );
and ( n22746 , n22590 , n22745 );
and ( n22747 , n22384 , n22745 );
or ( n22748 , n22591 , n22746 , n22747 );
and ( n22749 , n22497 , n22589 );
and ( n22750 , n22333 , n22337 );
and ( n22751 , n22337 , n22352 );
and ( n22752 , n22333 , n22352 );
or ( n22753 , n22750 , n22751 , n22752 );
and ( n22754 , n22001 , n22009 );
and ( n22755 , n22009 , n22070 );
and ( n22756 , n22001 , n22070 );
or ( n22757 , n22754 , n22755 , n22756 );
and ( n22758 , n21784 , n22323 );
and ( n22759 , n22137 , n22321 );
nor ( n22760 , n22758 , n22759 );
xnor ( n22761 , n22760 , n22329 );
and ( n22762 , n21833 , n22194 );
and ( n22763 , n21794 , n22192 );
nor ( n22764 , n22762 , n22763 );
xnor ( n22765 , n22764 , n22200 );
xor ( n22766 , n22761 , n22765 );
and ( n22767 , n21895 , n21927 );
and ( n22768 , n21908 , n21925 );
nor ( n22769 , n22767 , n22768 );
xnor ( n22770 , n22769 , n21937 );
xor ( n22771 , n22766 , n22770 );
and ( n22772 , n21919 , n22022 );
and ( n22773 , n21932 , n22020 );
nor ( n22774 , n22772 , n22773 );
xnor ( n22775 , n22774 , n22028 );
xor ( n22776 , n22771 , n22775 );
xor ( n22777 , n22757 , n22776 );
and ( n22778 , n22029 , n22036 );
and ( n22779 , n21870 , n21903 );
and ( n22780 , n21885 , n21901 );
nor ( n22781 , n22779 , n22780 );
xnor ( n22782 , n22781 , n21913 );
xor ( n22783 , n22778 , n22782 );
and ( n22784 , n22041 , n22062 );
and ( n22785 , n22014 , n22060 );
nor ( n22786 , n22784 , n22785 );
xnor ( n22787 , n22786 , n22068 );
xor ( n22788 , n22783 , n22787 );
and ( n22789 , n22056 , n22035 );
xor ( n22790 , n22788 , n22789 );
xor ( n22791 , n22777 , n22790 );
xor ( n22792 , n22753 , n22791 );
and ( n22793 , n22353 , n22377 );
and ( n22794 , n22377 , n22382 );
and ( n22795 , n22353 , n22382 );
or ( n22796 , n22793 , n22794 , n22795 );
xor ( n22797 , n22792 , n22796 );
and ( n22798 , n22558 , n22572 );
and ( n22799 , n22572 , n22587 );
and ( n22800 , n22558 , n22587 );
or ( n22801 , n22798 , n22799 , n22800 );
and ( n22802 , n21762 , n21735 );
and ( n22803 , n21740 , n21743 );
and ( n22804 , n21743 , n21746 );
and ( n22805 , n21740 , n21746 );
or ( n22806 , n22803 , n22804 , n22805 );
buf ( n22807 , n21745 );
not ( n22808 , n16101 );
xor ( n22809 , n22807 , n22808 );
and ( n22810 , n16066 , n16087 );
xor ( n22811 , n22809 , n22810 );
xor ( n22812 , n22806 , n22811 );
and ( n22813 , n21747 , n21751 );
and ( n22814 , n21751 , n21756 );
and ( n22815 , n21747 , n21756 );
or ( n22816 , n22813 , n22814 , n22815 );
xor ( n22817 , n22812 , n22816 );
and ( n22818 , n21757 , n21758 );
xor ( n22819 , n22817 , n22818 );
buf ( n550081 , n22819 );
buf ( n550082 , n550081 );
buf ( n22822 , n550082 );
and ( n22823 , n22822 , n21732 );
nor ( n22824 , n22802 , n22823 );
xnor ( n22825 , n22824 , n21730 );
xor ( n22826 , n22801 , n22825 );
and ( n22827 , n22244 , n22305 );
and ( n22828 , n22124 , n22303 );
nor ( n22829 , n22827 , n22828 );
xnor ( n22830 , n22829 , n22315 );
and ( n22831 , n21846 , n21779 );
and ( n22832 , n21859 , n21777 );
nor ( n22833 , n22831 , n22832 );
xnor ( n22834 , n22833 , n21789 );
xor ( n22835 , n22830 , n22834 );
and ( n22836 , n21947 , n21978 );
and ( n22837 , n21962 , n21976 );
nor ( n22838 , n22836 , n22837 );
xnor ( n22839 , n22838 , n21988 );
and ( n22840 , n21809 , n21828 );
and ( n22841 , n21995 , n21826 );
nor ( n22842 , n22840 , n22841 );
xnor ( n22843 , n22842 , n21838 );
xor ( n22844 , n22839 , n22843 );
and ( n22845 , n22273 , n21880 );
and ( n22846 , n21820 , n21878 );
nor ( n22847 , n22845 , n22846 );
xnor ( n22848 , n22847 , n21890 );
xor ( n22849 , n22844 , n22848 );
xor ( n22850 , n22835 , n22849 );
xor ( n22851 , n22826 , n22850 );
xor ( n22852 , n22797 , n22851 );
xor ( n22853 , n22749 , n22852 );
and ( n22854 , n22501 , n22553 );
and ( n22855 , n22553 , n22588 );
and ( n22856 , n22501 , n22588 );
or ( n22857 , n22854 , n22855 , n22856 );
and ( n22858 , n22072 , n22282 );
and ( n22859 , n22282 , n22383 );
and ( n22860 , n22072 , n22383 );
or ( n22861 , n22858 , n22859 , n22860 );
xor ( n22862 , n22857 , n22861 );
and ( n22863 , n21765 , n21942 );
and ( n22864 , n21942 , n22071 );
and ( n22865 , n21765 , n22071 );
or ( n22866 , n22863 , n22864 , n22865 );
and ( n22867 , n22129 , n22252 );
and ( n22868 , n21728 , n22250 );
nor ( n22869 , n22867 , n22868 );
xnor ( n22870 , n22869 , n22258 );
and ( n22871 , n22562 , n22566 );
and ( n22872 , n22566 , n22571 );
and ( n22873 , n22562 , n22571 );
or ( n22874 , n22871 , n22872 , n22873 );
xor ( n22875 , n22870 , n22874 );
and ( n22876 , n22577 , n22581 );
and ( n22877 , n22581 , n22586 );
and ( n22878 , n22577 , n22586 );
or ( n22879 , n22876 , n22877 , n22878 );
xor ( n22880 , n22875 , n22879 );
xor ( n22881 , n22866 , n22880 );
and ( n22882 , n22357 , n22361 );
and ( n22883 , n22361 , n22376 );
and ( n22884 , n22357 , n22376 );
or ( n22885 , n22882 , n22883 , n22884 );
and ( n22886 , n22366 , n22370 );
and ( n22887 , n22370 , n22375 );
and ( n22888 , n22366 , n22375 );
or ( n22889 , n22886 , n22887 , n22888 );
and ( n22890 , n22342 , n22346 );
and ( n22891 , n22346 , n22351 );
and ( n22892 , n22342 , n22351 );
or ( n22893 , n22890 , n22891 , n22892 );
xor ( n22894 , n22889 , n22893 );
and ( n22895 , n22148 , n21957 );
and ( n22896 , n21769 , n21955 );
nor ( n22897 , n22895 , n22896 );
xnor ( n22898 , n22897 , n21967 );
xor ( n22899 , n22894 , n22898 );
xor ( n22900 , n22885 , n22899 );
and ( n22901 , n22037 , n22051 );
and ( n22902 , n22051 , n22069 );
and ( n22903 , n22037 , n22069 );
or ( n22904 , n22901 , n22902 , n22903 );
and ( n22905 , n22006 , n21854 );
and ( n22906 , n22310 , n21852 );
nor ( n22907 , n22905 , n22906 );
xnor ( n22908 , n22907 , n21864 );
xor ( n22909 , n22904 , n22908 );
and ( n22910 , n21972 , n21804 );
and ( n22911 , n21983 , n21802 );
nor ( n22912 , n22910 , n22911 );
xnor ( n22913 , n22912 , n21814 );
xor ( n22914 , n22909 , n22913 );
xor ( n22915 , n22900 , n22914 );
xor ( n22916 , n22881 , n22915 );
xor ( n22917 , n22862 , n22916 );
xor ( n22918 , n22853 , n22917 );
xor ( n22919 , n22748 , n22918 );
xor ( n22920 , n22144 , n22235 );
xor ( n22921 , n22920 , n22279 );
xor ( n22922 , n22481 , n22483 );
xor ( n22923 , n22922 , n22494 );
and ( n22924 , n22921 , n22923 );
and ( n22925 , n21859 , n22252 );
and ( n22926 , n22006 , n22250 );
nor ( n22927 , n22925 , n22926 );
xnor ( n22928 , n22927 , n22258 );
and ( n22929 , n22137 , n22305 );
and ( n22930 , n21846 , n22303 );
nor ( n22931 , n22929 , n22930 );
xnor ( n22932 , n22931 , n22315 );
and ( n22933 , n22928 , n22932 );
xor ( n22934 , n22388 , n22392 );
xor ( n22935 , n22934 , n22397 );
and ( n22936 , n22932 , n22935 );
and ( n22937 , n22928 , n22935 );
or ( n22938 , n22933 , n22936 , n22937 );
and ( n22939 , n21947 , n21779 );
and ( n22940 , n21962 , n21777 );
nor ( n22941 , n22939 , n22940 );
xnor ( n22942 , n22941 , n21789 );
and ( n22943 , n21833 , n21978 );
and ( n22944 , n21794 , n21976 );
nor ( n22945 , n22943 , n22944 );
xnor ( n22946 , n22945 , n21988 );
and ( n22947 , n22942 , n22946 );
xor ( n22948 , n22401 , n22411 );
xor ( n22949 , n22948 , n22416 );
and ( n22950 , n22946 , n22949 );
and ( n22951 , n22942 , n22949 );
or ( n22952 , n22947 , n22950 , n22951 );
xor ( n22953 , n22419 , n22423 );
xor ( n22954 , n22953 , n22428 );
and ( n22955 , n22952 , n22954 );
xor ( n22956 , n22595 , n22599 );
xor ( n22957 , n22956 , n22602 );
and ( n22958 , n22954 , n22957 );
and ( n22959 , n22952 , n22957 );
or ( n22960 , n22955 , n22958 , n22959 );
and ( n22961 , n22938 , n22960 );
xor ( n22962 , n22400 , n22431 );
xor ( n22963 , n22962 , n22436 );
and ( n22964 , n22960 , n22963 );
and ( n22965 , n22938 , n22963 );
or ( n22966 , n22961 , n22964 , n22965 );
xor ( n22967 , n22439 , n22465 );
xor ( n22968 , n22967 , n22478 );
and ( n22969 , n22966 , n22968 );
xor ( n22970 , n22617 , n22619 );
xor ( n22971 , n22970 , n22622 );
and ( n22972 , n22968 , n22971 );
and ( n22973 , n22966 , n22971 );
or ( n22974 , n22969 , n22972 , n22973 );
and ( n22975 , n22923 , n22974 );
and ( n22976 , n22921 , n22974 );
or ( n22977 , n22924 , n22975 , n22976 );
xor ( n22978 , n22655 , n22660 );
and ( n22979 , n22041 , n21880 );
and ( n22980 , n22014 , n21878 );
nor ( n22981 , n22979 , n22980 );
xnor ( n22982 , n22981 , n21890 );
and ( n22983 , n22978 , n22982 );
and ( n22984 , n22033 , n21903 );
and ( n22985 , n22056 , n21901 );
nor ( n22986 , n22984 , n22985 );
xnor ( n22987 , n22986 , n21913 );
and ( n22988 , n22982 , n22987 );
and ( n22989 , n22978 , n22987 );
or ( n22990 , n22983 , n22988 , n22989 );
and ( n22991 , n21995 , n22323 );
and ( n22992 , n21972 , n22321 );
nor ( n22993 , n22991 , n22992 );
xnor ( n22994 , n22993 , n22329 );
and ( n22995 , n22990 , n22994 );
and ( n22996 , n21794 , n21957 );
and ( n22997 , n21809 , n21955 );
nor ( n22998 , n22996 , n22997 );
xnor ( n22999 , n22998 , n21967 );
and ( n23000 , n22994 , n22999 );
and ( n23001 , n22990 , n22999 );
or ( n23002 , n22995 , n23000 , n23001 );
and ( n23003 , n21784 , n22305 );
and ( n23004 , n22137 , n22303 );
nor ( n23005 , n23003 , n23004 );
xnor ( n23006 , n23005 , n22315 );
and ( n23007 , n23002 , n23006 );
xor ( n23008 , n22672 , n22676 );
xor ( n23009 , n23008 , n22681 );
and ( n23010 , n23006 , n23009 );
and ( n23011 , n23002 , n23009 );
or ( n23012 , n23007 , n23010 , n23011 );
and ( n23013 , n21769 , n22305 );
and ( n23014 , n21784 , n22303 );
nor ( n23015 , n23013 , n23014 );
xnor ( n23016 , n23015 , n22315 );
and ( n23017 , n21983 , n21779 );
and ( n23018 , n21947 , n21777 );
nor ( n23019 , n23017 , n23018 );
xnor ( n23020 , n23019 , n21789 );
and ( n23021 , n23016 , n23020 );
xor ( n23022 , n22693 , n22697 );
xor ( n23023 , n23022 , n22702 );
and ( n23024 , n23020 , n23023 );
and ( n23025 , n23016 , n23023 );
or ( n23026 , n23021 , n23024 , n23025 );
and ( n23027 , n21846 , n22252 );
and ( n23028 , n21859 , n22250 );
nor ( n23029 , n23027 , n23028 );
xnor ( n23030 , n23029 , n22258 );
and ( n23031 , n23026 , n23030 );
xor ( n23032 , n22942 , n22946 );
xor ( n23033 , n23032 , n22949 );
and ( n23034 , n23030 , n23033 );
and ( n23035 , n23026 , n23033 );
or ( n23036 , n23031 , n23034 , n23035 );
and ( n23037 , n23012 , n23036 );
xor ( n23038 , n22928 , n22932 );
xor ( n23039 , n23038 , n22935 );
and ( n23040 , n23036 , n23039 );
and ( n23041 , n23012 , n23039 );
or ( n23042 , n23037 , n23040 , n23041 );
xor ( n23043 , n22938 , n22960 );
xor ( n23044 , n23043 , n22963 );
and ( n23045 , n23042 , n23044 );
xor ( n23046 , n22692 , n22727 );
xor ( n23047 , n23046 , n22730 );
and ( n23048 , n23044 , n23047 );
and ( n23049 , n23042 , n23047 );
or ( n23050 , n23045 , n23048 , n23049 );
and ( n23051 , n22006 , n21735 );
and ( n23052 , n22310 , n21732 );
nor ( n23053 , n23051 , n23052 );
xnor ( n23054 , n23053 , n21730 );
and ( n23055 , n22148 , n21854 );
and ( n23056 , n21769 , n21852 );
nor ( n23057 , n23055 , n23056 );
xnor ( n23058 , n23057 , n21864 );
and ( n23059 , n23054 , n23058 );
and ( n23060 , n21972 , n22323 );
and ( n23061 , n21983 , n22321 );
nor ( n23062 , n23060 , n23061 );
xnor ( n23063 , n23062 , n22329 );
and ( n23064 , n23058 , n23063 );
and ( n23065 , n23054 , n23063 );
or ( n23066 , n23059 , n23064 , n23065 );
and ( n23067 , n22659 , n22062 );
and ( n23068 , n22409 , n22060 );
nor ( n23069 , n23067 , n23068 );
xnor ( n23070 , n23069 , n22068 );
xor ( n23071 , n20887 , n21677 );
buf ( n550333 , n23071 );
buf ( n550334 , n550333 );
buf ( n23074 , n550334 );
and ( n23075 , n23074 , n22035 );
and ( n23076 , n23070 , n23075 );
and ( n23077 , n22086 , n21927 );
and ( n23078 , n22049 , n21925 );
nor ( n23079 , n23077 , n23078 );
xnor ( n23080 , n23079 , n21937 );
and ( n23081 , n23076 , n23080 );
and ( n23082 , n22080 , n22022 );
and ( n23083 , n22101 , n22020 );
nor ( n23084 , n23082 , n23083 );
xnor ( n23085 , n23084 , n22028 );
and ( n23086 , n23080 , n23085 );
and ( n23087 , n23076 , n23085 );
or ( n23088 , n23081 , n23086 , n23087 );
and ( n23089 , n21908 , n21828 );
and ( n23090 , n21870 , n21826 );
nor ( n23091 , n23089 , n23090 );
xnor ( n23092 , n23091 , n21838 );
and ( n23093 , n23088 , n23092 );
and ( n23094 , n21932 , n22194 );
and ( n23095 , n21895 , n22192 );
nor ( n23096 , n23094 , n23095 );
xnor ( n23097 , n23096 , n22200 );
and ( n23098 , n23092 , n23097 );
and ( n23099 , n23088 , n23097 );
or ( n23100 , n23093 , n23098 , n23099 );
and ( n23101 , n21820 , n21978 );
and ( n23102 , n21833 , n21976 );
nor ( n23103 , n23101 , n23102 );
xnor ( n23104 , n23103 , n21988 );
and ( n23105 , n21885 , n21804 );
and ( n23106 , n22273 , n21802 );
nor ( n23107 , n23105 , n23106 );
xnor ( n23108 , n23107 , n21814 );
and ( n23109 , n23104 , n23108 );
xor ( n23110 , n22661 , n22664 );
xor ( n23111 , n23110 , n22669 );
and ( n23112 , n23108 , n23111 );
and ( n23113 , n23104 , n23111 );
or ( n23114 , n23109 , n23112 , n23113 );
and ( n23115 , n23100 , n23114 );
xor ( n23116 , n22639 , n22643 );
xor ( n23117 , n23116 , n22648 );
and ( n23118 , n23114 , n23117 );
and ( n23119 , n23100 , n23117 );
or ( n23120 , n23115 , n23118 , n23119 );
and ( n23121 , n23066 , n23120 );
xor ( n23122 , n22651 , n22684 );
xor ( n23123 , n23122 , n22689 );
and ( n23124 , n23120 , n23123 );
and ( n23125 , n23066 , n23123 );
or ( n23126 , n23121 , n23124 , n23125 );
xor ( n23127 , n22605 , n22609 );
xor ( n23128 , n23127 , n22614 );
and ( n23129 , n23126 , n23128 );
xor ( n23130 , n22627 , n22629 );
xor ( n23131 , n23130 , n22632 );
and ( n23132 , n23128 , n23131 );
and ( n23133 , n23126 , n23131 );
or ( n23134 , n23129 , n23132 , n23133 );
and ( n23135 , n23050 , n23134 );
xor ( n23136 , n22635 , n22733 );
xor ( n23137 , n23136 , n22736 );
and ( n23138 , n23134 , n23137 );
and ( n23139 , n23050 , n23137 );
or ( n23140 , n23135 , n23138 , n23139 );
xor ( n23141 , n22625 , n22739 );
xor ( n23142 , n23141 , n22742 );
and ( n23143 , n23140 , n23142 );
and ( n23144 , n22977 , n23143 );
xor ( n23145 , n22384 , n22590 );
xor ( n23146 , n23145 , n22745 );
and ( n23147 , n23143 , n23146 );
and ( n23148 , n22977 , n23146 );
or ( n23149 , n23144 , n23147 , n23148 );
xor ( n23150 , n22919 , n23149 );
xor ( n23151 , n22977 , n23143 );
xor ( n23152 , n23151 , n23146 );
xor ( n23153 , n22921 , n22923 );
xor ( n23154 , n23153 , n22974 );
xor ( n23155 , n23140 , n23142 );
and ( n23156 , n23154 , n23155 );
xor ( n23157 , n23070 , n23075 );
and ( n23158 , n23074 , n22062 );
and ( n23159 , n22659 , n22060 );
nor ( n23160 , n23158 , n23159 );
xnor ( n23161 , n23160 , n22068 );
xor ( n23162 , n21487 , n21675 );
buf ( n550424 , n23162 );
buf ( n550425 , n550424 );
buf ( n23165 , n550425 );
and ( n23166 , n23165 , n22035 );
and ( n23167 , n23161 , n23166 );
and ( n23168 , n23157 , n23167 );
and ( n23169 , n22094 , n22022 );
and ( n23170 , n22080 , n22020 );
nor ( n23171 , n23169 , n23170 );
xnor ( n23172 , n23171 , n22028 );
and ( n23173 , n23167 , n23172 );
and ( n23174 , n23157 , n23172 );
or ( n23175 , n23168 , n23173 , n23174 );
and ( n23176 , n21895 , n21828 );
and ( n23177 , n21908 , n21826 );
nor ( n23178 , n23176 , n23177 );
xnor ( n23179 , n23178 , n21838 );
and ( n23180 , n23175 , n23179 );
and ( n23181 , n21919 , n22194 );
and ( n23182 , n21932 , n22192 );
nor ( n23183 , n23181 , n23182 );
xnor ( n23184 , n23183 , n22200 );
and ( n23185 , n23179 , n23184 );
and ( n23186 , n23175 , n23184 );
or ( n23187 , n23180 , n23185 , n23186 );
and ( n23188 , n22273 , n21978 );
and ( n23189 , n21820 , n21976 );
nor ( n23190 , n23188 , n23189 );
xnor ( n23191 , n23190 , n21988 );
and ( n23192 , n21870 , n21804 );
and ( n23193 , n21885 , n21802 );
nor ( n23194 , n23192 , n23193 );
xnor ( n23195 , n23194 , n21814 );
and ( n23196 , n23191 , n23195 );
xor ( n23197 , n23076 , n23080 );
xor ( n23198 , n23197 , n23085 );
and ( n23199 , n23195 , n23198 );
and ( n23200 , n23191 , n23198 );
or ( n23201 , n23196 , n23199 , n23200 );
and ( n23202 , n23187 , n23201 );
and ( n23203 , n21962 , n21854 );
and ( n23204 , n22148 , n21852 );
nor ( n23205 , n23203 , n23204 );
xnor ( n23206 , n23205 , n21864 );
and ( n23207 , n23201 , n23206 );
and ( n23208 , n23187 , n23206 );
or ( n23209 , n23202 , n23207 , n23208 );
and ( n23210 , n22137 , n22252 );
and ( n23211 , n21846 , n22250 );
nor ( n23212 , n23210 , n23211 );
xnor ( n23213 , n23212 , n22258 );
xor ( n23214 , n23088 , n23092 );
xor ( n23215 , n23214 , n23097 );
and ( n23216 , n23213 , n23215 );
xor ( n23217 , n23104 , n23108 );
xor ( n23218 , n23217 , n23111 );
and ( n23219 , n23215 , n23218 );
and ( n23220 , n23213 , n23218 );
or ( n23221 , n23216 , n23219 , n23220 );
and ( n23222 , n23209 , n23221 );
xor ( n23223 , n23002 , n23006 );
xor ( n23224 , n23223 , n23009 );
and ( n23225 , n23221 , n23224 );
and ( n23226 , n23209 , n23224 );
or ( n23227 , n23222 , n23225 , n23226 );
and ( n23228 , n22056 , n21880 );
and ( n23229 , n22041 , n21878 );
nor ( n23230 , n23228 , n23229 );
xnor ( n23231 , n23230 , n21890 );
and ( n23232 , n22049 , n21903 );
and ( n23233 , n22033 , n21901 );
nor ( n23234 , n23232 , n23233 );
xnor ( n23235 , n23234 , n21913 );
and ( n23236 , n23231 , n23235 );
and ( n23237 , n22101 , n21927 );
and ( n23238 , n22086 , n21925 );
nor ( n23239 , n23237 , n23238 );
xnor ( n23240 , n23239 , n21937 );
and ( n23241 , n23235 , n23240 );
and ( n23242 , n23231 , n23240 );
or ( n23243 , n23236 , n23241 , n23242 );
and ( n23244 , n21809 , n22323 );
and ( n23245 , n21995 , n22321 );
nor ( n23246 , n23244 , n23245 );
xnor ( n23247 , n23246 , n22329 );
and ( n23248 , n23243 , n23247 );
and ( n23249 , n21833 , n21957 );
and ( n23250 , n21794 , n21955 );
nor ( n23251 , n23249 , n23250 );
xnor ( n23252 , n23251 , n21967 );
and ( n23253 , n23247 , n23252 );
and ( n23254 , n23243 , n23252 );
or ( n23255 , n23248 , n23253 , n23254 );
and ( n23256 , n21947 , n21854 );
and ( n23257 , n21962 , n21852 );
nor ( n23258 , n23256 , n23257 );
xnor ( n23259 , n23258 , n21864 );
and ( n550521 , n21972 , n21779 );
and ( n23261 , n21983 , n21777 );
nor ( n550523 , n550521 , n23261 );
xnor ( n23263 , n550523 , n21789 );
and ( n23264 , n23259 , n23263 );
xor ( n23265 , n22978 , n22982 );
xor ( n23266 , n23265 , n22987 );
and ( n23267 , n23263 , n23266 );
and ( n23268 , n23259 , n23266 );
or ( n23269 , n23264 , n23267 , n23268 );
and ( n23270 , n23255 , n23269 );
xor ( n23271 , n22990 , n22994 );
xor ( n23272 , n23271 , n22999 );
and ( n23273 , n23269 , n23272 );
and ( n23274 , n23255 , n23272 );
or ( n23275 , n23270 , n23273 , n23274 );
xor ( n23276 , n23161 , n23166 );
and ( n23277 , n23165 , n22062 );
and ( n23278 , n23074 , n22060 );
nor ( n23279 , n23277 , n23278 );
xnor ( n23280 , n23279 , n22068 );
xor ( n23281 , n21489 , n21674 );
buf ( n550543 , n23281 );
buf ( n550544 , n550543 );
buf ( n23284 , n550544 );
and ( n23285 , n23284 , n22035 );
and ( n23286 , n23280 , n23285 );
and ( n23287 , n23276 , n23286 );
and ( n23288 , n22409 , n22022 );
and ( n23289 , n22094 , n22020 );
nor ( n23290 , n23288 , n23289 );
xnor ( n23291 , n23290 , n22028 );
and ( n23292 , n23286 , n23291 );
and ( n23293 , n23276 , n23291 );
or ( n23294 , n23287 , n23292 , n23293 );
and ( n23295 , n21885 , n21978 );
and ( n23296 , n22273 , n21976 );
nor ( n23297 , n23295 , n23296 );
xnor ( n23298 , n23297 , n21988 );
and ( n23299 , n23294 , n23298 );
and ( n23300 , n22014 , n22194 );
and ( n23301 , n21919 , n22192 );
nor ( n23302 , n23300 , n23301 );
xnor ( n23303 , n23302 , n22200 );
and ( n23304 , n23298 , n23303 );
and ( n23305 , n23294 , n23303 );
or ( n23306 , n23299 , n23304 , n23305 );
and ( n23307 , n21908 , n21804 );
and ( n23308 , n21870 , n21802 );
nor ( n23309 , n23307 , n23308 );
xnor ( n23310 , n23309 , n21814 );
and ( n23311 , n21932 , n21828 );
and ( n23312 , n21895 , n21826 );
nor ( n23313 , n23311 , n23312 );
xnor ( n23314 , n23313 , n21838 );
and ( n23315 , n23310 , n23314 );
xor ( n23316 , n23157 , n23167 );
xor ( n23317 , n23316 , n23172 );
and ( n23318 , n23314 , n23317 );
and ( n23319 , n23310 , n23317 );
or ( n23320 , n23315 , n23318 , n23319 );
and ( n23321 , n23306 , n23320 );
and ( n23322 , n22148 , n22305 );
and ( n550584 , n21769 , n22303 );
nor ( n23323 , n23322 , n550584 );
xnor ( n23324 , n23323 , n22315 );
and ( n23325 , n23320 , n23324 );
and ( n23326 , n23306 , n23324 );
or ( n23327 , n23321 , n23325 , n23326 );
and ( n23328 , n21859 , n21735 );
and ( n23329 , n22006 , n21732 );
nor ( n23330 , n23328 , n23329 );
xnor ( n23331 , n23330 , n21730 );
and ( n23332 , n23327 , n23331 );
xor ( n23333 , n23016 , n23020 );
xor ( n23334 , n23333 , n23023 );
and ( n23335 , n23331 , n23334 );
and ( n23336 , n23327 , n23334 );
or ( n23337 , n23332 , n23335 , n23336 );
and ( n23338 , n23275 , n23337 );
xor ( n23339 , n23026 , n23030 );
xor ( n23340 , n23339 , n23033 );
and ( n23341 , n23337 , n23340 );
and ( n23342 , n23275 , n23340 );
or ( n23343 , n23338 , n23341 , n23342 );
and ( n23344 , n23227 , n23343 );
xor ( n23345 , n23066 , n23120 );
xor ( n23346 , n23345 , n23123 );
and ( n23347 , n23343 , n23346 );
and ( n23348 , n23227 , n23346 );
or ( n23349 , n23344 , n23347 , n23348 );
xor ( n23350 , n23054 , n23058 );
xor ( n23351 , n23350 , n23063 );
xor ( n23352 , n22705 , n22709 );
xor ( n23353 , n23352 , n22714 );
and ( n23354 , n23351 , n23353 );
xor ( n23355 , n23100 , n23114 );
xor ( n23356 , n23355 , n23117 );
and ( n23357 , n23353 , n23356 );
and ( n23358 , n23351 , n23356 );
or ( n23359 , n23354 , n23357 , n23358 );
xor ( n23360 , n22717 , n22721 );
xor ( n23361 , n23360 , n22724 );
and ( n23362 , n23359 , n23361 );
xor ( n23363 , n22952 , n22954 );
xor ( n23364 , n23363 , n22957 );
and ( n23365 , n23361 , n23364 );
and ( n23366 , n23359 , n23364 );
or ( n23367 , n23362 , n23365 , n23366 );
and ( n23368 , n23349 , n23367 );
xor ( n23369 , n23126 , n23128 );
xor ( n23370 , n23369 , n23131 );
and ( n23371 , n23367 , n23370 );
and ( n23372 , n23349 , n23370 );
or ( n23373 , n23368 , n23371 , n23372 );
xor ( n23374 , n22966 , n22968 );
xor ( n23375 , n23374 , n22971 );
and ( n23376 , n23373 , n23375 );
xor ( n23377 , n23050 , n23134 );
xor ( n23378 , n23377 , n23137 );
and ( n23379 , n23375 , n23378 );
and ( n23380 , n23373 , n23378 );
or ( n23381 , n23376 , n23379 , n23380 );
and ( n23382 , n23155 , n23381 );
and ( n23383 , n23154 , n23381 );
or ( n23384 , n23156 , n23382 , n23383 );
and ( n23385 , n23152 , n23384 );
xor ( n23386 , n23152 , n23384 );
xor ( n23387 , n23154 , n23155 );
xor ( n23388 , n23387 , n23381 );
xor ( n23389 , n23373 , n23375 );
xor ( n23390 , n23389 , n23378 );
and ( n23391 , n21784 , n22252 );
and ( n23392 , n22137 , n22250 );
nor ( n23393 , n23391 , n23392 );
xnor ( n23394 , n23393 , n22258 );
xor ( n23395 , n23175 , n23179 );
xor ( n23396 , n23395 , n23184 );
and ( n23397 , n23394 , n23396 );
xor ( n23398 , n23191 , n23195 );
xor ( n23399 , n23398 , n23198 );
and ( n23400 , n23396 , n23399 );
and ( n23401 , n23394 , n23399 );
or ( n23402 , n23397 , n23400 , n23401 );
xor ( n23403 , n23187 , n23201 );
xor ( n23404 , n23403 , n23206 );
and ( n23405 , n23402 , n23404 );
xor ( n23406 , n23213 , n23215 );
xor ( n23407 , n23406 , n23218 );
and ( n23408 , n23404 , n23407 );
and ( n23409 , n23402 , n23407 );
or ( n23410 , n23405 , n23408 , n23409 );
xor ( n23411 , n23209 , n23221 );
xor ( n23412 , n23411 , n23224 );
and ( n23413 , n23410 , n23412 );
xor ( n23414 , n23351 , n23353 );
xor ( n23415 , n23414 , n23356 );
and ( n23416 , n23412 , n23415 );
and ( n23417 , n23410 , n23415 );
or ( n23418 , n23413 , n23416 , n23417 );
xor ( n23419 , n23012 , n23036 );
xor ( n23420 , n23419 , n23039 );
and ( n23421 , n23418 , n23420 );
xor ( n23422 , n23359 , n23361 );
xor ( n23423 , n23422 , n23364 );
and ( n23424 , n23420 , n23423 );
and ( n23425 , n23418 , n23423 );
or ( n23426 , n23421 , n23424 , n23425 );
xor ( n23427 , n23042 , n23044 );
xor ( n23428 , n23427 , n23047 );
and ( n23429 , n23426 , n23428 );
xor ( n23430 , n23349 , n23367 );
xor ( n23431 , n23430 , n23370 );
and ( n23432 , n23428 , n23431 );
and ( n23433 , n23426 , n23431 );
or ( n23434 , n23429 , n23432 , n23433 );
and ( n23435 , n23390 , n23434 );
xor ( n23436 , n23426 , n23428 );
xor ( n23437 , n23436 , n23431 );
xor ( n23438 , n23280 , n23285 );
and ( n23439 , n23284 , n22062 );
and ( n23440 , n23165 , n22060 );
nor ( n23441 , n23439 , n23440 );
xnor ( n23442 , n23441 , n22068 );
xor ( n23443 , n21491 , n21673 );
buf ( n550706 , n23443 );
buf ( n550707 , n550706 );
buf ( n23446 , n550707 );
and ( n23447 , n23446 , n22035 );
and ( n23448 , n23442 , n23447 );
and ( n23449 , n23438 , n23448 );
and ( n23450 , n22659 , n22022 );
and ( n23451 , n22409 , n22020 );
nor ( n23452 , n23450 , n23451 );
xnor ( n23453 , n23452 , n22028 );
and ( n23454 , n23448 , n23453 );
and ( n23455 , n23438 , n23453 );
or ( n23456 , n23449 , n23454 , n23455 );
and ( n23457 , n22086 , n21903 );
and ( n23458 , n22049 , n21901 );
nor ( n23459 , n23457 , n23458 );
xnor ( n23460 , n23459 , n21913 );
and ( n23461 , n23456 , n23460 );
and ( n23462 , n22080 , n21927 );
and ( n23463 , n22101 , n21925 );
nor ( n23464 , n23462 , n23463 );
xnor ( n23465 , n23464 , n21937 );
and ( n23466 , n23460 , n23465 );
and ( n23467 , n23456 , n23465 );
or ( n23468 , n23461 , n23466 , n23467 );
and ( n23469 , n21995 , n21779 );
and ( n23470 , n21972 , n21777 );
nor ( n23471 , n23469 , n23470 );
xnor ( n23472 , n23471 , n21789 );
and ( n23473 , n23468 , n23472 );
and ( n23474 , n21794 , n22323 );
and ( n23475 , n21809 , n22321 );
nor ( n23476 , n23474 , n23475 );
xnor ( n23477 , n23476 , n22329 );
and ( n23478 , n23472 , n23477 );
and ( n23479 , n23468 , n23477 );
or ( n23480 , n23473 , n23478 , n23479 );
and ( n23481 , n21769 , n22252 );
and ( n23482 , n21784 , n22250 );
nor ( n23483 , n23481 , n23482 );
xnor ( n23484 , n23483 , n22258 );
and ( n23485 , n21820 , n21957 );
and ( n23486 , n21833 , n21955 );
nor ( n23487 , n23485 , n23486 );
xnor ( n23488 , n23487 , n21967 );
and ( n23489 , n23484 , n23488 );
xor ( n23490 , n23231 , n23235 );
xor ( n23491 , n23490 , n23240 );
and ( n23492 , n23488 , n23491 );
and ( n23493 , n23484 , n23491 );
or ( n23494 , n23489 , n23492 , n23493 );
and ( n23495 , n23480 , n23494 );
and ( n23496 , n21846 , n21735 );
and ( n23497 , n21859 , n21732 );
nor ( n23498 , n23496 , n23497 );
xnor ( n23499 , n23498 , n21730 );
and ( n23500 , n23494 , n23499 );
and ( n23501 , n23480 , n23499 );
or ( n23502 , n23495 , n23500 , n23501 );
and ( n23503 , n22049 , n21880 );
and ( n23504 , n22033 , n21878 );
nor ( n23505 , n23503 , n23504 );
xnor ( n23506 , n23505 , n21890 );
and ( n23507 , n22101 , n21903 );
and ( n23508 , n22086 , n21901 );
nor ( n23509 , n23507 , n23508 );
xnor ( n23510 , n23509 , n21913 );
and ( n23511 , n23506 , n23510 );
and ( n23512 , n22094 , n21927 );
and ( n23513 , n22080 , n21925 );
nor ( n23514 , n23512 , n23513 );
xnor ( n23515 , n23514 , n21937 );
and ( n23516 , n23510 , n23515 );
and ( n23517 , n23506 , n23515 );
or ( n23518 , n23511 , n23516 , n23517 );
and ( n23519 , n22041 , n22194 );
and ( n23520 , n22014 , n22192 );
nor ( n23521 , n23519 , n23520 );
xnor ( n23522 , n23521 , n22200 );
and ( n23523 , n23518 , n23522 );
and ( n23524 , n22033 , n21880 );
and ( n23525 , n22056 , n21878 );
nor ( n23526 , n23524 , n23525 );
xnor ( n23527 , n23526 , n21890 );
and ( n23528 , n23522 , n23527 );
and ( n23529 , n23518 , n23527 );
or ( n23530 , n23523 , n23528 , n23529 );
and ( n23531 , n21870 , n21978 );
and ( n23532 , n21885 , n21976 );
nor ( n23533 , n23531 , n23532 );
xnor ( n23534 , n23533 , n21988 );
and ( n23535 , n21895 , n21804 );
and ( n23536 , n21908 , n21802 );
nor ( n23537 , n23535 , n23536 );
xnor ( n23538 , n23537 , n21814 );
and ( n23539 , n23534 , n23538 );
xor ( n23540 , n23276 , n23286 );
xor ( n23541 , n23540 , n23291 );
and ( n23542 , n23538 , n23541 );
and ( n23543 , n23534 , n23541 );
or ( n23544 , n23539 , n23542 , n23543 );
and ( n23545 , n23530 , n23544 );
and ( n23546 , n21983 , n21854 );
and ( n23547 , n21947 , n21852 );
nor ( n23548 , n23546 , n23547 );
xnor ( n23549 , n23548 , n21864 );
and ( n23550 , n23544 , n23549 );
and ( n23551 , n23530 , n23549 );
or ( n23552 , n23545 , n23550 , n23551 );
xor ( n23553 , n23243 , n23247 );
xor ( n23554 , n23553 , n23252 );
and ( n23555 , n23552 , n23554 );
xor ( n23556 , n23259 , n23263 );
xor ( n23557 , n23556 , n23266 );
and ( n23558 , n23554 , n23557 );
and ( n23559 , n23552 , n23557 );
or ( n23560 , n23555 , n23558 , n23559 );
and ( n23561 , n23502 , n23560 );
xor ( n23562 , n23255 , n23269 );
xor ( n23563 , n23562 , n23272 );
and ( n23564 , n23560 , n23563 );
and ( n23565 , n23502 , n23563 );
or ( n23566 , n23561 , n23564 , n23565 );
xor ( n23567 , n23442 , n23447 );
and ( n23568 , n23165 , n22022 );
and ( n23569 , n23074 , n22020 );
nor ( n23570 , n23568 , n23569 );
xnor ( n23571 , n23570 , n22028 );
xor ( n23572 , n21493 , n21672 );
buf ( n550835 , n23572 );
buf ( n550836 , n550835 );
buf ( n23575 , n550836 );
and ( n23576 , n23575 , n22035 );
and ( n23577 , n23571 , n23576 );
and ( n23578 , n23567 , n23577 );
and ( n23579 , n23074 , n22022 );
and ( n23580 , n22659 , n22020 );
nor ( n23581 , n23579 , n23580 );
xnor ( n23582 , n23581 , n22028 );
and ( n23583 , n23577 , n23582 );
and ( n23584 , n23567 , n23582 );
or ( n23585 , n23578 , n23583 , n23584 );
and ( n23586 , n22014 , n21828 );
and ( n23587 , n21919 , n21826 );
nor ( n23588 , n23586 , n23587 );
xnor ( n23589 , n23588 , n21838 );
and ( n23590 , n23585 , n23589 );
and ( n23591 , n22056 , n22194 );
and ( n23592 , n22041 , n22192 );
nor ( n23593 , n23591 , n23592 );
xnor ( n23594 , n23593 , n22200 );
and ( n23595 , n23589 , n23594 );
and ( n23596 , n23585 , n23594 );
or ( n23597 , n23590 , n23595 , n23596 );
and ( n23598 , n21809 , n21779 );
and ( n23599 , n21995 , n21777 );
nor ( n23600 , n23598 , n23599 );
xnor ( n23601 , n23600 , n21789 );
and ( n23602 , n23597 , n23601 );
and ( n23603 , n21919 , n21828 );
and ( n23604 , n21932 , n21826 );
nor ( n23605 , n23603 , n23604 );
xnor ( n23606 , n23605 , n21838 );
and ( n23607 , n23601 , n23606 );
and ( n23608 , n23597 , n23606 );
or ( n23609 , n23602 , n23607 , n23608 );
and ( n23610 , n21833 , n22323 );
and ( n23611 , n21794 , n22321 );
nor ( n23612 , n23610 , n23611 );
xnor ( n23613 , n23612 , n22329 );
and ( n23614 , n22273 , n21957 );
and ( n23615 , n21820 , n21955 );
nor ( n23616 , n23614 , n23615 );
xnor ( n23617 , n23616 , n21967 );
and ( n23618 , n23613 , n23617 );
xor ( n23619 , n23456 , n23460 );
xor ( n23620 , n23619 , n23465 );
and ( n23621 , n23617 , n23620 );
and ( n23622 , n23613 , n23620 );
or ( n23623 , n23618 , n23621 , n23622 );
and ( n23624 , n23609 , n23623 );
and ( n23625 , n22137 , n21735 );
and ( n23626 , n21846 , n21732 );
nor ( n23627 , n23625 , n23626 );
xnor ( n23628 , n23627 , n21730 );
and ( n23629 , n23623 , n23628 );
and ( n23630 , n23609 , n23628 );
or ( n23631 , n23624 , n23629 , n23630 );
and ( n23632 , n21962 , n22305 );
and ( n23633 , n22148 , n22303 );
nor ( n23634 , n23632 , n23633 );
xnor ( n23635 , n23634 , n22315 );
xor ( n23636 , n23294 , n23298 );
xor ( n23637 , n23636 , n23303 );
and ( n23638 , n23635 , n23637 );
xor ( n23639 , n23310 , n23314 );
xor ( n23640 , n23639 , n23317 );
and ( n23641 , n23637 , n23640 );
and ( n23642 , n23635 , n23640 );
or ( n23643 , n23638 , n23641 , n23642 );
and ( n23644 , n23631 , n23643 );
xor ( n23645 , n23306 , n23320 );
xor ( n23646 , n23645 , n23324 );
and ( n23647 , n23643 , n23646 );
and ( n23648 , n23631 , n23646 );
or ( n23649 , n23644 , n23647 , n23648 );
xor ( n23650 , n23327 , n23331 );
xor ( n23651 , n23650 , n23334 );
and ( n23652 , n23649 , n23651 );
xor ( n23653 , n23402 , n23404 );
xor ( n23654 , n23653 , n23407 );
and ( n23655 , n23651 , n23654 );
and ( n23656 , n23649 , n23654 );
or ( n23657 , n23652 , n23655 , n23656 );
and ( n23658 , n23566 , n23657 );
xor ( n23659 , n23275 , n23337 );
xor ( n23660 , n23659 , n23340 );
and ( n23661 , n23657 , n23660 );
and ( n23662 , n23566 , n23660 );
or ( n23663 , n23658 , n23661 , n23662 );
xor ( n23664 , n23227 , n23343 );
xor ( n23665 , n23664 , n23346 );
and ( n23666 , n23663 , n23665 );
xor ( n23667 , n23418 , n23420 );
xor ( n23668 , n23667 , n23423 );
and ( n23669 , n23665 , n23668 );
and ( n23670 , n23663 , n23668 );
or ( n23671 , n23666 , n23669 , n23670 );
and ( n23672 , n23437 , n23671 );
xor ( n23673 , n23663 , n23665 );
xor ( n23674 , n23673 , n23668 );
xor ( n23675 , n23410 , n23412 );
xor ( n23676 , n23675 , n23415 );
xor ( n23677 , n23566 , n23657 );
xor ( n23678 , n23677 , n23660 );
and ( n23679 , n23676 , n23678 );
xor ( n23680 , n23502 , n23560 );
xor ( n23681 , n23680 , n23563 );
and ( n23682 , n21947 , n22305 );
and ( n23683 , n21962 , n22303 );
nor ( n23684 , n23682 , n23683 );
xnor ( n23685 , n23684 , n22315 );
and ( n23686 , n21972 , n21854 );
and ( n23687 , n21983 , n21852 );
nor ( n23688 , n23686 , n23687 );
xnor ( n23689 , n23688 , n21864 );
and ( n23690 , n23685 , n23689 );
xor ( n23691 , n23518 , n23522 );
xor ( n23692 , n23691 , n23527 );
and ( n23693 , n23689 , n23692 );
and ( n23694 , n23685 , n23692 );
or ( n23695 , n23690 , n23693 , n23694 );
xor ( n23696 , n23468 , n23472 );
xor ( n23697 , n23696 , n23477 );
and ( n23698 , n23695 , n23697 );
xor ( n23699 , n23484 , n23488 );
xor ( n23700 , n23699 , n23491 );
and ( n23701 , n23697 , n23700 );
and ( n23702 , n23695 , n23700 );
or ( n23703 , n23698 , n23701 , n23702 );
xor ( n23704 , n23480 , n23494 );
xor ( n23705 , n23704 , n23499 );
and ( n23706 , n23703 , n23705 );
xor ( n23707 , n23394 , n23396 );
xor ( n23708 , n23707 , n23399 );
and ( n23709 , n23705 , n23708 );
and ( n23710 , n23703 , n23708 );
or ( n23711 , n23706 , n23709 , n23710 );
and ( n23712 , n23681 , n23711 );
xor ( n23713 , n23649 , n23651 );
xor ( n23714 , n23713 , n23654 );
and ( n23715 , n23711 , n23714 );
and ( n23716 , n23681 , n23714 );
or ( n23717 , n23712 , n23715 , n23716 );
and ( n23718 , n23678 , n23717 );
and ( n23719 , n23676 , n23717 );
or ( n23720 , n23679 , n23718 , n23719 );
and ( n23721 , n23674 , n23720 );
and ( n23722 , n21885 , n21957 );
and ( n23723 , n22273 , n21955 );
nor ( n23724 , n23722 , n23723 );
xnor ( n23725 , n23724 , n21967 );
and ( n23726 , n21908 , n21978 );
and ( n23727 , n21870 , n21976 );
nor ( n23728 , n23726 , n23727 );
xnor ( n23729 , n23728 , n21988 );
and ( n23730 , n23725 , n23729 );
xor ( n23731 , n23506 , n23510 );
xor ( n23732 , n23731 , n23515 );
and ( n23733 , n23729 , n23732 );
and ( n23734 , n23725 , n23732 );
or ( n23735 , n23730 , n23733 , n23734 );
and ( n23736 , n22086 , n21880 );
and ( n23737 , n22049 , n21878 );
nor ( n23738 , n23736 , n23737 );
xnor ( n23739 , n23738 , n21890 );
and ( n23740 , n22080 , n21903 );
and ( n23741 , n22101 , n21901 );
nor ( n23742 , n23740 , n23741 );
xnor ( n23743 , n23742 , n21913 );
and ( n23744 , n23739 , n23743 );
and ( n23745 , n22409 , n21927 );
and ( n23746 , n22094 , n21925 );
nor ( n23747 , n23745 , n23746 );
xnor ( n23748 , n23747 , n21937 );
and ( n23749 , n23743 , n23748 );
and ( n23750 , n23739 , n23748 );
or ( n23751 , n23744 , n23749 , n23750 );
and ( n23752 , n21932 , n21804 );
and ( n23753 , n21895 , n21802 );
nor ( n23754 , n23752 , n23753 );
xnor ( n23755 , n23754 , n21814 );
and ( n23756 , n23751 , n23755 );
xor ( n23757 , n23438 , n23448 );
xor ( n23758 , n23757 , n23453 );
and ( n23759 , n23755 , n23758 );
and ( n23760 , n23751 , n23758 );
or ( n23761 , n23756 , n23759 , n23760 );
and ( n23762 , n23735 , n23761 );
and ( n23763 , n22148 , n22252 );
and ( n23764 , n21769 , n22250 );
nor ( n23765 , n23763 , n23764 );
xnor ( n23766 , n23765 , n22258 );
and ( n23767 , n23761 , n23766 );
and ( n23768 , n23735 , n23766 );
or ( n23769 , n23762 , n23767 , n23768 );
xor ( n23770 , n23530 , n23544 );
xor ( n23771 , n23770 , n23549 );
and ( n23772 , n23769 , n23771 );
xor ( n23773 , n23635 , n23637 );
xor ( n23774 , n23773 , n23640 );
and ( n23775 , n23771 , n23774 );
and ( n23776 , n23769 , n23774 );
or ( n23777 , n23772 , n23775 , n23776 );
xor ( n23778 , n23631 , n23643 );
xor ( n23779 , n23778 , n23646 );
and ( n23780 , n23777 , n23779 );
xor ( n23781 , n23552 , n23554 );
xor ( n23782 , n23781 , n23557 );
and ( n23783 , n23779 , n23782 );
and ( n23784 , n23777 , n23782 );
or ( n23785 , n23780 , n23783 , n23784 );
xor ( n23786 , n23703 , n23705 );
xor ( n23787 , n23786 , n23708 );
and ( n23788 , n21962 , n22252 );
and ( n23789 , n22148 , n22250 );
nor ( n23790 , n23788 , n23789 );
xnor ( n23791 , n23790 , n22258 );
xor ( n23792 , n23585 , n23589 );
xor ( n23793 , n23792 , n23594 );
and ( n23794 , n23791 , n23793 );
xor ( n23795 , n23751 , n23755 );
xor ( n23796 , n23795 , n23758 );
and ( n23797 , n23793 , n23796 );
and ( n23798 , n23791 , n23796 );
or ( n23799 , n23794 , n23797 , n23798 );
and ( n23800 , n21870 , n21957 );
and ( n23801 , n21885 , n21955 );
nor ( n23802 , n23800 , n23801 );
xnor ( n23803 , n23802 , n21967 );
and ( n23804 , n21895 , n21978 );
and ( n23805 , n21908 , n21976 );
nor ( n23806 , n23804 , n23805 );
xnor ( n23807 , n23806 , n21988 );
and ( n23808 , n23803 , n23807 );
xor ( n23809 , n23739 , n23743 );
xor ( n23810 , n23809 , n23748 );
and ( n23811 , n23807 , n23810 );
and ( n23812 , n23803 , n23810 );
or ( n23813 , n23808 , n23811 , n23812 );
xor ( n23814 , n23571 , n23576 );
and ( n23815 , n22101 , n21880 );
and ( n23816 , n22086 , n21878 );
nor ( n23817 , n23815 , n23816 );
xnor ( n23818 , n23817 , n21890 );
and ( n23819 , n23814 , n23818 );
and ( n23820 , n22094 , n21903 );
and ( n23821 , n22080 , n21901 );
nor ( n23822 , n23820 , n23821 );
xnor ( n23823 , n23822 , n21913 );
and ( n23824 , n23818 , n23823 );
and ( n23825 , n23814 , n23823 );
or ( n23826 , n23819 , n23824 , n23825 );
and ( n23827 , n21919 , n21804 );
and ( n23828 , n21932 , n21802 );
nor ( n23829 , n23827 , n23828 );
xnor ( n23830 , n23829 , n21814 );
and ( n23831 , n23826 , n23830 );
xor ( n23832 , n23567 , n23577 );
xor ( n23833 , n23832 , n23582 );
and ( n23834 , n23830 , n23833 );
and ( n23835 , n23826 , n23833 );
or ( n23836 , n23831 , n23834 , n23835 );
and ( n23837 , n23813 , n23836 );
xor ( n23838 , n23725 , n23729 );
xor ( n23839 , n23838 , n23732 );
and ( n23840 , n23836 , n23839 );
and ( n23841 , n23813 , n23839 );
or ( n23842 , n23837 , n23840 , n23841 );
and ( n23843 , n23799 , n23842 );
xor ( n23844 , n23685 , n23689 );
xor ( n23845 , n23844 , n23692 );
and ( n23846 , n23842 , n23845 );
and ( n23847 , n23799 , n23845 );
or ( n23848 , n23843 , n23846 , n23847 );
xor ( n23849 , n23695 , n23697 );
xor ( n23850 , n23849 , n23700 );
and ( n23851 , n23848 , n23850 );
xor ( n23852 , n23769 , n23771 );
xor ( n23853 , n23852 , n23774 );
and ( n23854 , n23850 , n23853 );
and ( n23855 , n23848 , n23853 );
or ( n23856 , n23851 , n23854 , n23855 );
and ( n23857 , n23787 , n23856 );
and ( n23858 , n21784 , n21735 );
and ( n23859 , n22137 , n21732 );
nor ( n23860 , n23858 , n23859 );
xnor ( n23861 , n23860 , n21730 );
and ( n23862 , n21769 , n21735 );
and ( n23863 , n21784 , n21732 );
nor ( n23864 , n23862 , n23863 );
xnor ( n23865 , n23864 , n21730 );
and ( n23866 , n21983 , n22305 );
and ( n23867 , n21947 , n22303 );
nor ( n23868 , n23866 , n23867 );
xnor ( n23869 , n23868 , n22315 );
and ( n23870 , n23865 , n23869 );
and ( n23871 , n21995 , n21854 );
and ( n23872 , n21972 , n21852 );
nor ( n23873 , n23871 , n23872 );
xnor ( n23874 , n23873 , n21864 );
and ( n23875 , n23869 , n23874 );
and ( n23876 , n23865 , n23874 );
or ( n23877 , n23870 , n23875 , n23876 );
and ( n23878 , n23861 , n23877 );
xor ( n23879 , n23534 , n23538 );
xor ( n23880 , n23879 , n23541 );
and ( n23881 , n23877 , n23880 );
and ( n23882 , n23861 , n23880 );
or ( n23883 , n23878 , n23881 , n23882 );
xor ( n23884 , n23609 , n23623 );
xor ( n23885 , n23884 , n23628 );
and ( n23886 , n23883 , n23885 );
and ( n23887 , n22148 , n21735 );
and ( n23888 , n21769 , n21732 );
nor ( n23889 , n23887 , n23888 );
xnor ( n23890 , n23889 , n21730 );
and ( n23891 , n21947 , n22252 );
and ( n23892 , n21962 , n22250 );
nor ( n23893 , n23891 , n23892 );
xnor ( n23894 , n23893 , n22258 );
and ( n23895 , n23890 , n23894 );
and ( n23896 , n21972 , n22305 );
and ( n23897 , n21983 , n22303 );
nor ( n23898 , n23896 , n23897 );
xnor ( n23899 , n23898 , n22315 );
and ( n23900 , n23894 , n23899 );
and ( n23901 , n23890 , n23899 );
or ( n23902 , n23895 , n23900 , n23901 );
xor ( n23903 , n23865 , n23869 );
xor ( n23904 , n23903 , n23874 );
and ( n23905 , n23902 , n23904 );
and ( n23906 , n21809 , n21854 );
and ( n23907 , n21995 , n21852 );
nor ( n23908 , n23906 , n23907 );
xnor ( n23909 , n23908 , n21864 );
and ( n23910 , n21983 , n22252 );
and ( n23911 , n21947 , n22250 );
nor ( n23912 , n23910 , n23911 );
xnor ( n23913 , n23912 , n22258 );
and ( n23914 , n21995 , n22305 );
and ( n23915 , n21972 , n22303 );
nor ( n23916 , n23914 , n23915 );
xnor ( n23917 , n23916 , n22315 );
and ( n23918 , n23913 , n23917 );
and ( n23919 , n23909 , n23918 );
xor ( n23920 , n23890 , n23894 );
xor ( n23921 , n23920 , n23899 );
and ( n23922 , n23918 , n23921 );
and ( n23923 , n23909 , n23921 );
or ( n23924 , n23919 , n23922 , n23923 );
and ( n23925 , n23904 , n23924 );
and ( n23926 , n23902 , n23924 );
or ( n23927 , n23905 , n23925 , n23926 );
xor ( n23928 , n23597 , n23601 );
xor ( n23929 , n23928 , n23606 );
and ( n23930 , n23927 , n23929 );
xor ( n23931 , n23735 , n23761 );
xor ( n23932 , n23931 , n23766 );
and ( n23933 , n23929 , n23932 );
and ( n23934 , n23927 , n23932 );
or ( n23935 , n23930 , n23933 , n23934 );
and ( n23936 , n23885 , n23935 );
and ( n23937 , n23883 , n23935 );
or ( n23938 , n23886 , n23936 , n23937 );
and ( n23939 , n23856 , n23938 );
and ( n23940 , n23787 , n23938 );
or ( n23941 , n23857 , n23939 , n23940 );
and ( n23942 , n23785 , n23941 );
xor ( n23943 , n23777 , n23779 );
xor ( n23944 , n23943 , n23782 );
xor ( n23945 , n23613 , n23617 );
xor ( n23946 , n23945 , n23620 );
and ( n23947 , n23284 , n22022 );
and ( n23948 , n23165 , n22020 );
nor ( n23949 , n23947 , n23948 );
xnor ( n23950 , n23949 , n22028 );
xor ( n23951 , n21495 , n21671 );
buf ( n551214 , n23951 );
buf ( n551215 , n551214 );
buf ( n23954 , n551215 );
and ( n23955 , n23954 , n22035 );
and ( n23956 , n23950 , n23955 );
and ( n23957 , n22659 , n21927 );
and ( n23958 , n22409 , n21925 );
nor ( n23959 , n23957 , n23958 );
xnor ( n23960 , n23959 , n21937 );
and ( n23961 , n23956 , n23960 );
and ( n23962 , n23446 , n22062 );
and ( n23963 , n23284 , n22060 );
nor ( n23964 , n23962 , n23963 );
xnor ( n23965 , n23964 , n22068 );
and ( n23966 , n23960 , n23965 );
and ( n23967 , n23956 , n23965 );
or ( n23968 , n23961 , n23966 , n23967 );
and ( n23969 , n22041 , n21828 );
and ( n23970 , n22014 , n21826 );
nor ( n23971 , n23969 , n23970 );
xnor ( n23972 , n23971 , n21838 );
and ( n23973 , n23968 , n23972 );
and ( n23974 , n22033 , n22194 );
and ( n23975 , n22056 , n22192 );
nor ( n23976 , n23974 , n23975 );
xnor ( n23977 , n23976 , n22200 );
and ( n23978 , n23972 , n23977 );
and ( n23979 , n23968 , n23977 );
or ( n23980 , n23973 , n23978 , n23979 );
and ( n23981 , n21794 , n21779 );
and ( n23982 , n21809 , n21777 );
nor ( n23983 , n23981 , n23982 );
xnor ( n23984 , n23983 , n21789 );
and ( n23985 , n23980 , n23984 );
and ( n23986 , n21820 , n22323 );
and ( n23987 , n21833 , n22321 );
nor ( n23988 , n23986 , n23987 );
xnor ( n23989 , n23988 , n22329 );
and ( n23990 , n23984 , n23989 );
and ( n23991 , n23980 , n23989 );
or ( n23992 , n23985 , n23990 , n23991 );
and ( n23993 , n23946 , n23992 );
xor ( n23994 , n23861 , n23877 );
xor ( n23995 , n23994 , n23880 );
and ( n23996 , n23992 , n23995 );
and ( n23997 , n23946 , n23995 );
or ( n23998 , n23993 , n23996 , n23997 );
xor ( n23999 , n23848 , n23850 );
xor ( n24000 , n23999 , n23853 );
and ( n24001 , n23998 , n24000 );
xor ( n24002 , n23799 , n23842 );
xor ( n24003 , n24002 , n23845 );
and ( n24004 , n23954 , n22062 );
and ( n24005 , n23575 , n22060 );
nor ( n24006 , n24004 , n24005 );
xnor ( n24007 , n24006 , n22068 );
xor ( n24008 , n21497 , n21670 );
buf ( n551271 , n24008 );
buf ( n551272 , n551271 );
buf ( n24011 , n551272 );
and ( n24012 , n24011 , n22035 );
and ( n24013 , n24007 , n24012 );
and ( n24014 , n23074 , n21927 );
and ( n24015 , n22659 , n21925 );
nor ( n24016 , n24014 , n24015 );
xnor ( n24017 , n24016 , n21937 );
and ( n24018 , n24013 , n24017 );
and ( n24019 , n23575 , n22062 );
and ( n24020 , n23446 , n22060 );
nor ( n24021 , n24019 , n24020 );
xnor ( n24022 , n24021 , n22068 );
and ( n24023 , n24017 , n24022 );
and ( n24024 , n24013 , n24022 );
or ( n24025 , n24018 , n24023 , n24024 );
and ( n24026 , n22014 , n21804 );
and ( n24027 , n21919 , n21802 );
nor ( n24028 , n24026 , n24027 );
xnor ( n24029 , n24028 , n21814 );
and ( n24030 , n24025 , n24029 );
and ( n24031 , n22049 , n22194 );
and ( n24032 , n22033 , n22192 );
nor ( n24033 , n24031 , n24032 );
xnor ( n24034 , n24033 , n22200 );
and ( n24035 , n24029 , n24034 );
and ( n24036 , n24025 , n24034 );
or ( n24037 , n24030 , n24035 , n24036 );
and ( n24038 , n21833 , n21779 );
and ( n24039 , n21794 , n21777 );
nor ( n24040 , n24038 , n24039 );
xnor ( n24041 , n24040 , n21789 );
and ( n24042 , n24037 , n24041 );
and ( n24043 , n22273 , n22323 );
and ( n24044 , n21820 , n22321 );
nor ( n24045 , n24043 , n24044 );
xnor ( n24046 , n24045 , n22329 );
and ( n24047 , n24041 , n24046 );
and ( n24048 , n24037 , n24046 );
or ( n24049 , n24042 , n24047 , n24048 );
xor ( n24050 , n23980 , n23984 );
xor ( n24051 , n24050 , n23989 );
and ( n24052 , n24049 , n24051 );
and ( n24053 , n24003 , n24052 );
xor ( n24054 , n23803 , n23807 );
xor ( n24055 , n24054 , n23810 );
and ( n24056 , n21962 , n21735 );
and ( n24057 , n22148 , n21732 );
nor ( n24058 , n24056 , n24057 );
xnor ( n24059 , n24058 , n21730 );
and ( n24060 , n22056 , n21828 );
and ( n24061 , n22041 , n21826 );
nor ( n24062 , n24060 , n24061 );
xnor ( n24063 , n24062 , n21838 );
and ( n24064 , n24059 , n24063 );
and ( n24065 , n21794 , n21854 );
and ( n24066 , n21809 , n21852 );
nor ( n24067 , n24065 , n24066 );
xnor ( n24068 , n24067 , n21864 );
and ( n24069 , n21885 , n22323 );
and ( n24070 , n22273 , n22321 );
nor ( n24071 , n24069 , n24070 );
xnor ( n24072 , n24071 , n22329 );
xor ( n24073 , n24068 , n24072 );
and ( n24074 , n21908 , n21957 );
and ( n24075 , n21870 , n21955 );
nor ( n24076 , n24074 , n24075 );
xnor ( n24077 , n24076 , n21967 );
xor ( n24078 , n24073 , n24077 );
and ( n24079 , n24063 , n24078 );
and ( n24080 , n24059 , n24078 );
or ( n24081 , n24064 , n24079 , n24080 );
and ( n24082 , n24055 , n24081 );
xor ( n24083 , n23909 , n23918 );
xor ( n24084 , n24083 , n23921 );
and ( n24085 , n24081 , n24084 );
and ( n24086 , n24055 , n24084 );
or ( n24087 , n24082 , n24085 , n24086 );
xor ( n24088 , n23902 , n23904 );
xor ( n24089 , n24088 , n23924 );
and ( n24090 , n24087 , n24089 );
xor ( n24091 , n23791 , n23793 );
xor ( n24092 , n24091 , n23796 );
and ( n24093 , n24089 , n24092 );
and ( n24094 , n24087 , n24092 );
or ( n24095 , n24090 , n24093 , n24094 );
and ( n24096 , n24052 , n24095 );
and ( n24097 , n24003 , n24095 );
or ( n24098 , n24053 , n24096 , n24097 );
and ( n24099 , n24000 , n24098 );
and ( n24100 , n23998 , n24098 );
or ( n24101 , n24001 , n24099 , n24100 );
and ( n24102 , n23944 , n24101 );
xor ( n24103 , n23787 , n23856 );
xor ( n24104 , n24103 , n23938 );
and ( n24105 , n24101 , n24104 );
and ( n24106 , n23944 , n24104 );
or ( n24107 , n24102 , n24105 , n24106 );
and ( n24108 , n23941 , n24107 );
and ( n24109 , n23785 , n24107 );
or ( n24110 , n23942 , n24108 , n24109 );
xor ( n24111 , n23676 , n23678 );
xor ( n24112 , n24111 , n23717 );
and ( n24113 , n24110 , n24112 );
xor ( n24114 , n23681 , n23711 );
xor ( n24115 , n24114 , n23714 );
xor ( n24116 , n23785 , n23941 );
xor ( n24117 , n24116 , n24107 );
and ( n24118 , n24115 , n24117 );
xor ( n24119 , n23883 , n23885 );
xor ( n24120 , n24119 , n23935 );
xor ( n24121 , n23927 , n23929 );
xor ( n24122 , n24121 , n23932 );
xor ( n24123 , n23946 , n23992 );
xor ( n24124 , n24123 , n23995 );
and ( n24125 , n24122 , n24124 );
xor ( n24126 , n23813 , n23836 );
xor ( n24127 , n24126 , n23839 );
xor ( n24128 , n23968 , n23972 );
xor ( n24129 , n24128 , n23977 );
xor ( n24130 , n23826 , n23830 );
xor ( n24131 , n24130 , n23833 );
and ( n24132 , n24129 , n24131 );
xor ( n24133 , n23913 , n23917 );
and ( n24134 , n21833 , n21854 );
and ( n24135 , n21794 , n21852 );
nor ( n24136 , n24134 , n24135 );
xnor ( n24137 , n24136 , n21864 );
and ( n24138 , n22273 , n21779 );
and ( n24139 , n21820 , n21777 );
nor ( n24140 , n24138 , n24139 );
xnor ( n24141 , n24140 , n21789 );
and ( n24142 , n24137 , n24141 );
and ( n24143 , n24133 , n24142 );
xor ( n24144 , n23956 , n23960 );
xor ( n24145 , n24144 , n23965 );
and ( n24146 , n24142 , n24145 );
and ( n24147 , n24133 , n24145 );
or ( n24148 , n24143 , n24146 , n24147 );
and ( n24149 , n24131 , n24148 );
and ( n24150 , n24129 , n24148 );
or ( n24151 , n24132 , n24149 , n24150 );
and ( n24152 , n24127 , n24151 );
xor ( n24153 , n24049 , n24051 );
and ( n24154 , n24151 , n24153 );
and ( n24155 , n24127 , n24153 );
or ( n24156 , n24152 , n24154 , n24155 );
and ( n24157 , n24124 , n24156 );
and ( n24158 , n24122 , n24156 );
or ( n24159 , n24125 , n24157 , n24158 );
and ( n24160 , n24120 , n24159 );
xor ( n24161 , n23998 , n24000 );
xor ( n24162 , n24161 , n24098 );
and ( n24163 , n24159 , n24162 );
and ( n24164 , n24120 , n24162 );
or ( n24165 , n24160 , n24163 , n24164 );
xor ( n24166 , n23944 , n24101 );
xor ( n24167 , n24166 , n24104 );
and ( n24168 , n24165 , n24167 );
and ( n24169 , n24068 , n24072 );
and ( n24170 , n24072 , n24077 );
and ( n24171 , n24068 , n24077 );
or ( n24172 , n24169 , n24170 , n24171 );
and ( n24173 , n22094 , n21880 );
and ( n24174 , n22080 , n21878 );
nor ( n24175 , n24173 , n24174 );
xnor ( n24176 , n24175 , n21890 );
and ( n24177 , n22659 , n21903 );
and ( n24178 , n22409 , n21901 );
nor ( n24179 , n24177 , n24178 );
xnor ( n24180 , n24179 , n21913 );
and ( n24181 , n24176 , n24180 );
and ( n24182 , n23446 , n22022 );
and ( n24183 , n23284 , n22020 );
nor ( n24184 , n24182 , n24183 );
xnor ( n24185 , n24184 , n22028 );
and ( n24186 , n24180 , n24185 );
and ( n24187 , n24176 , n24185 );
or ( n24188 , n24181 , n24186 , n24187 );
and ( n24189 , n22041 , n21804 );
and ( n24190 , n22014 , n21802 );
nor ( n24191 , n24189 , n24190 );
xnor ( n24192 , n24191 , n21814 );
and ( n24193 , n24188 , n24192 );
and ( n24194 , n22033 , n21828 );
and ( n24195 , n22056 , n21826 );
nor ( n24196 , n24194 , n24195 );
xnor ( n24197 , n24196 , n21838 );
and ( n24198 , n24192 , n24197 );
and ( n24199 , n24188 , n24197 );
or ( n24200 , n24193 , n24198 , n24199 );
and ( n24201 , n21820 , n21779 );
and ( n24202 , n21833 , n21777 );
nor ( n24203 , n24201 , n24202 );
xnor ( n24204 , n24203 , n21789 );
and ( n24205 , n24200 , n24204 );
xor ( n24206 , n24025 , n24029 );
xor ( n24207 , n24206 , n24034 );
and ( n24208 , n24204 , n24207 );
and ( n24209 , n24200 , n24207 );
or ( n24210 , n24205 , n24208 , n24209 );
and ( n24211 , n24172 , n24210 );
xor ( n24212 , n24037 , n24041 );
xor ( n24213 , n24212 , n24046 );
and ( n24214 , n24210 , n24213 );
and ( n24215 , n24172 , n24213 );
or ( n24216 , n24211 , n24214 , n24215 );
and ( n24217 , n22409 , n21903 );
and ( n24218 , n22094 , n21901 );
nor ( n24219 , n24217 , n24218 );
xnor ( n24220 , n24219 , n21913 );
xor ( n24221 , n23950 , n23955 );
and ( n24222 , n24220 , n24221 );
and ( n24223 , n21919 , n21978 );
and ( n24224 , n21932 , n21976 );
nor ( n24225 , n24223 , n24224 );
xnor ( n24226 , n24225 , n21988 );
xor ( n24227 , n24137 , n24141 );
and ( n24228 , n24226 , n24227 );
and ( n24229 , n21983 , n21735 );
and ( n24230 , n21947 , n21732 );
nor ( n24231 , n24229 , n24230 );
xnor ( n24232 , n24231 , n21730 );
and ( n24233 , n21995 , n22252 );
and ( n24234 , n21972 , n22250 );
nor ( n24235 , n24233 , n24234 );
xnor ( n24236 , n24235 , n22258 );
and ( n24237 , n24232 , n24236 );
and ( n24238 , n21794 , n22305 );
and ( n24239 , n21809 , n22303 );
nor ( n24240 , n24238 , n24239 );
xnor ( n24241 , n24240 , n22315 );
and ( n24242 , n24236 , n24241 );
and ( n24243 , n24232 , n24241 );
or ( n24244 , n24237 , n24242 , n24243 );
and ( n24245 , n24227 , n24244 );
and ( n24246 , n24226 , n24244 );
or ( n24247 , n24228 , n24245 , n24246 );
and ( n24248 , n24222 , n24247 );
xor ( n24249 , n24059 , n24063 );
xor ( n24250 , n24249 , n24078 );
and ( n24251 , n24247 , n24250 );
and ( n24252 , n24222 , n24250 );
or ( n24253 , n24248 , n24251 , n24252 );
xor ( n24254 , n24055 , n24081 );
xor ( n24255 , n24254 , n24084 );
and ( n24256 , n24253 , n24255 );
and ( n24257 , n22086 , n22194 );
and ( n24258 , n22049 , n22192 );
nor ( n24259 , n24257 , n24258 );
xnor ( n24260 , n24259 , n22200 );
and ( n24261 , n22080 , n21880 );
and ( n24262 , n22101 , n21878 );
nor ( n24263 , n24261 , n24262 );
xnor ( n24264 , n24263 , n21890 );
and ( n24265 , n24260 , n24264 );
xor ( n24266 , n24013 , n24017 );
xor ( n24267 , n24266 , n24022 );
and ( n24268 , n24264 , n24267 );
and ( n24269 , n24260 , n24267 );
or ( n24270 , n24265 , n24268 , n24269 );
and ( n24271 , n21932 , n21978 );
and ( n24272 , n21895 , n21976 );
nor ( n24273 , n24271 , n24272 );
xnor ( n24274 , n24273 , n21988 );
and ( n24275 , n24270 , n24274 );
xor ( n24276 , n23814 , n23818 );
xor ( n24277 , n24276 , n23823 );
and ( n24278 , n24274 , n24277 );
and ( n24279 , n24270 , n24277 );
or ( n24280 , n24275 , n24278 , n24279 );
and ( n24281 , n24255 , n24280 );
and ( n24282 , n24253 , n24280 );
or ( n24283 , n24256 , n24281 , n24282 );
and ( n24284 , n24216 , n24283 );
and ( n24285 , n22086 , n21828 );
and ( n24286 , n22049 , n21826 );
nor ( n24287 , n24285 , n24286 );
xnor ( n24288 , n24287 , n21838 );
and ( n24289 , n22080 , n22194 );
and ( n24290 , n22101 , n22192 );
nor ( n24291 , n24289 , n24290 );
xnor ( n24292 , n24291 , n22200 );
and ( n24293 , n24288 , n24292 );
and ( n24294 , n22409 , n21880 );
and ( n24295 , n22094 , n21878 );
nor ( n24296 , n24294 , n24295 );
xnor ( n24297 , n24296 , n21890 );
and ( n24298 , n24292 , n24297 );
and ( n24299 , n24288 , n24297 );
or ( n24300 , n24293 , n24298 , n24299 );
and ( n24301 , n22056 , n21804 );
and ( n24302 , n22041 , n21802 );
nor ( n24303 , n24301 , n24302 );
xnor ( n24304 , n24303 , n21814 );
and ( n24305 , n24300 , n24304 );
xor ( n24306 , n24176 , n24180 );
xor ( n24307 , n24306 , n24185 );
and ( n24308 , n24304 , n24307 );
and ( n24309 , n24300 , n24307 );
or ( n24310 , n24305 , n24308 , n24309 );
and ( n24311 , n21972 , n22252 );
and ( n24312 , n21983 , n22250 );
nor ( n24313 , n24311 , n24312 );
xnor ( n24314 , n24313 , n22258 );
and ( n24315 , n24310 , n24314 );
and ( n24316 , n21809 , n22305 );
and ( n24317 , n21995 , n22303 );
nor ( n24318 , n24316 , n24317 );
xnor ( n24319 , n24318 , n22315 );
and ( n24320 , n24314 , n24319 );
and ( n24321 , n24310 , n24319 );
or ( n24322 , n24315 , n24320 , n24321 );
and ( n24323 , n21885 , n21779 );
and ( n24324 , n22273 , n21777 );
nor ( n24325 , n24323 , n24324 );
xnor ( n24326 , n24325 , n21789 );
and ( n24327 , n21908 , n22323 );
and ( n24328 , n21870 , n22321 );
nor ( n24329 , n24327 , n24328 );
xnor ( n24330 , n24329 , n22329 );
and ( n24331 , n24326 , n24330 );
and ( n24332 , n21932 , n21957 );
and ( n24333 , n21895 , n21955 );
nor ( n24334 , n24332 , n24333 );
xnor ( n24335 , n24334 , n21967 );
and ( n24336 , n24330 , n24335 );
and ( n24337 , n24326 , n24335 );
or ( n24338 , n24331 , n24336 , n24337 );
and ( n24339 , n21947 , n21735 );
and ( n24340 , n21962 , n21732 );
nor ( n24341 , n24339 , n24340 );
xnor ( n24342 , n24341 , n21730 );
and ( n24343 , n24338 , n24342 );
xor ( n24344 , n24188 , n24192 );
xor ( n24345 , n24344 , n24197 );
and ( n24346 , n24342 , n24345 );
and ( n24347 , n24338 , n24345 );
or ( n24348 , n24343 , n24346 , n24347 );
and ( n24349 , n24322 , n24348 );
and ( n24350 , n21820 , n21854 );
and ( n24351 , n21833 , n21852 );
nor ( n24352 , n24350 , n24351 );
xnor ( n24353 , n24352 , n21864 );
and ( n24354 , n22014 , n21978 );
and ( n24355 , n21919 , n21976 );
nor ( n24356 , n24354 , n24355 );
xnor ( n24357 , n24356 , n21988 );
and ( n24358 , n24353 , n24357 );
and ( n24359 , n22049 , n21828 );
and ( n24360 , n22033 , n21826 );
nor ( n24361 , n24359 , n24360 );
xnor ( n24362 , n24361 , n21838 );
and ( n24363 , n24357 , n24362 );
and ( n24364 , n24353 , n24362 );
or ( n24365 , n24358 , n24363 , n24364 );
xor ( n24366 , n24220 , n24221 );
and ( n24367 , n24365 , n24366 );
and ( n24368 , n22101 , n22194 );
and ( n24369 , n22086 , n22192 );
nor ( n24370 , n24368 , n24369 );
xnor ( n24371 , n24370 , n22200 );
and ( n24372 , n23165 , n21927 );
and ( n24373 , n23074 , n21925 );
nor ( n24374 , n24372 , n24373 );
xnor ( n24375 , n24374 , n21937 );
and ( n24376 , n24371 , n24375 );
xor ( n24377 , n24326 , n24330 );
xor ( n24378 , n24377 , n24335 );
and ( n24379 , n24375 , n24378 );
and ( n24380 , n24371 , n24378 );
or ( n24381 , n24376 , n24379 , n24380 );
and ( n24382 , n24366 , n24381 );
and ( n24383 , n24365 , n24381 );
or ( n24384 , n24367 , n24382 , n24383 );
and ( n24385 , n24348 , n24384 );
and ( n24386 , n24322 , n24384 );
or ( n24387 , n24349 , n24385 , n24386 );
xor ( n24388 , n24007 , n24012 );
and ( n24389 , n23074 , n21903 );
and ( n24390 , n22659 , n21901 );
nor ( n24391 , n24389 , n24390 );
xnor ( n24392 , n24391 , n21913 );
and ( n24393 , n23575 , n22022 );
and ( n24394 , n23446 , n22020 );
nor ( n24395 , n24393 , n24394 );
xnor ( n24396 , n24395 , n22028 );
and ( n24397 , n24392 , n24396 );
and ( n24398 , n24388 , n24397 );
and ( n24399 , n21972 , n21735 );
and ( n24400 , n21983 , n21732 );
nor ( n24401 , n24399 , n24400 );
xnor ( n24402 , n24401 , n21730 );
and ( n24403 , n21833 , n22305 );
and ( n24404 , n21794 , n22303 );
nor ( n24405 , n24403 , n24404 );
xnor ( n24406 , n24405 , n22315 );
and ( n24407 , n24402 , n24406 );
and ( n24408 , n22273 , n21854 );
and ( n24409 , n21820 , n21852 );
nor ( n24410 , n24408 , n24409 );
xnor ( n24411 , n24410 , n21864 );
and ( n24412 , n24406 , n24411 );
and ( n24413 , n24402 , n24411 );
or ( n24414 , n24407 , n24412 , n24413 );
and ( n24415 , n24397 , n24414 );
and ( n24416 , n24388 , n24414 );
or ( n24417 , n24398 , n24415 , n24416 );
and ( n24418 , n21870 , n21779 );
and ( n24419 , n21885 , n21777 );
nor ( n24420 , n24418 , n24419 );
xnor ( n24421 , n24420 , n21789 );
and ( n24422 , n21919 , n21957 );
and ( n24423 , n21932 , n21955 );
nor ( n24424 , n24422 , n24423 );
xnor ( n24425 , n24424 , n21967 );
and ( n24426 , n24421 , n24425 );
and ( n24427 , n22041 , n21978 );
and ( n24428 , n22014 , n21976 );
nor ( n24429 , n24427 , n24428 );
xnor ( n24430 , n24429 , n21988 );
and ( n24431 , n24425 , n24430 );
and ( n24432 , n24421 , n24430 );
or ( n24433 , n24426 , n24431 , n24432 );
and ( n24434 , n22033 , n21804 );
and ( n24435 , n22056 , n21802 );
nor ( n24436 , n24434 , n24435 );
xnor ( n24437 , n24436 , n21814 );
and ( n24438 , n24011 , n22062 );
and ( n24439 , n23954 , n22060 );
nor ( n24440 , n24438 , n24439 );
xnor ( n24441 , n24440 , n22068 );
and ( n24442 , n24437 , n24441 );
xor ( n24443 , n21499 , n21669 );
buf ( n551706 , n24443 );
buf ( n551707 , n551706 );
buf ( n24446 , n551707 );
and ( n24447 , n24446 , n22035 );
and ( n24448 , n24441 , n24447 );
and ( n24449 , n24437 , n24447 );
or ( n24450 , n24442 , n24448 , n24449 );
and ( n24451 , n24433 , n24450 );
xor ( n24452 , n24232 , n24236 );
xor ( n24453 , n24452 , n24241 );
and ( n24454 , n24450 , n24453 );
and ( n24455 , n24433 , n24453 );
or ( n24456 , n24451 , n24454 , n24455 );
and ( n24457 , n24417 , n24456 );
xor ( n24458 , n24226 , n24227 );
xor ( n24459 , n24458 , n24244 );
and ( n24460 , n24456 , n24459 );
and ( n24461 , n24417 , n24459 );
or ( n24462 , n24457 , n24460 , n24461 );
xor ( n24463 , n24133 , n24142 );
xor ( n24464 , n24463 , n24145 );
and ( n24465 , n24462 , n24464 );
xor ( n24466 , n24222 , n24247 );
xor ( n24467 , n24466 , n24250 );
and ( n24468 , n24464 , n24467 );
and ( n24469 , n24462 , n24467 );
or ( n24470 , n24465 , n24468 , n24469 );
and ( n24471 , n24387 , n24470 );
xor ( n24472 , n24129 , n24131 );
xor ( n24473 , n24472 , n24148 );
and ( n24474 , n24470 , n24473 );
and ( n24475 , n24387 , n24473 );
or ( n24476 , n24471 , n24474 , n24475 );
and ( n24477 , n24283 , n24476 );
and ( n24478 , n24216 , n24476 );
or ( n24479 , n24284 , n24477 , n24478 );
xor ( n24480 , n24003 , n24052 );
xor ( n24481 , n24480 , n24095 );
and ( n24482 , n24479 , n24481 );
xor ( n24483 , n24087 , n24089 );
xor ( n24484 , n24483 , n24092 );
xor ( n24485 , n24172 , n24210 );
xor ( n24486 , n24485 , n24213 );
xor ( n24487 , n24270 , n24274 );
xor ( n24488 , n24487 , n24277 );
xor ( n24489 , n24200 , n24204 );
xor ( n24490 , n24489 , n24207 );
and ( n24491 , n24488 , n24490 );
and ( n24492 , n21870 , n22323 );
and ( n24493 , n21885 , n22321 );
nor ( n24494 , n24492 , n24493 );
xnor ( n24495 , n24494 , n22329 );
and ( n24496 , n21895 , n21957 );
and ( n24497 , n21908 , n21955 );
nor ( n24498 , n24496 , n24497 );
xnor ( n24499 , n24498 , n21967 );
and ( n24500 , n24495 , n24499 );
xor ( n24501 , n24260 , n24264 );
xor ( n24502 , n24501 , n24267 );
and ( n24503 , n24499 , n24502 );
and ( n24504 , n24495 , n24502 );
or ( n24505 , n24500 , n24503 , n24504 );
and ( n24506 , n24490 , n24505 );
and ( n24507 , n24488 , n24505 );
or ( n24508 , n24491 , n24506 , n24507 );
and ( n24509 , n24486 , n24508 );
xor ( n24510 , n24310 , n24314 );
xor ( n24511 , n24510 , n24319 );
xor ( n24512 , n24338 , n24342 );
xor ( n24513 , n24512 , n24345 );
and ( n24514 , n24511 , n24513 );
xor ( n24515 , n24353 , n24357 );
xor ( n24516 , n24515 , n24362 );
xor ( n24517 , n24300 , n24304 );
xor ( n24518 , n24517 , n24307 );
and ( n24519 , n24516 , n24518 );
and ( n24520 , n21809 , n22252 );
and ( n24521 , n21995 , n22250 );
nor ( n24522 , n24520 , n24521 );
xnor ( n24523 , n24522 , n22258 );
and ( n24524 , n21895 , n22323 );
and ( n24525 , n21908 , n22321 );
nor ( n24526 , n24524 , n24525 );
xnor ( n24527 , n24526 , n22329 );
and ( n24528 , n24523 , n24527 );
xor ( n24529 , n24288 , n24292 );
xor ( n24530 , n24529 , n24297 );
and ( n24531 , n24527 , n24530 );
and ( n24532 , n24523 , n24530 );
or ( n24533 , n24528 , n24531 , n24532 );
and ( n24534 , n24518 , n24533 );
and ( n24535 , n24516 , n24533 );
or ( n24536 , n24519 , n24534 , n24535 );
and ( n24537 , n24446 , n22062 );
and ( n24538 , n24011 , n22060 );
nor ( n24539 , n24537 , n24538 );
xnor ( n24540 , n24539 , n22068 );
xor ( n24541 , n21501 , n21668 );
buf ( n551804 , n24541 );
buf ( n551805 , n551804 );
buf ( n24544 , n551805 );
and ( n24545 , n24544 , n22035 );
and ( n24546 , n24540 , n24545 );
and ( n24547 , n23284 , n21927 );
and ( n24548 , n23165 , n21925 );
nor ( n24549 , n24547 , n24548 );
xnor ( n24550 , n24549 , n21937 );
and ( n24551 , n24546 , n24550 );
xor ( n24552 , n24392 , n24396 );
and ( n24553 , n22659 , n21880 );
and ( n24554 , n22409 , n21878 );
nor ( n24555 , n24553 , n24554 );
xnor ( n24556 , n24555 , n21890 );
and ( n24557 , n23165 , n21903 );
and ( n24558 , n23074 , n21901 );
nor ( n24559 , n24557 , n24558 );
xnor ( n24560 , n24559 , n21913 );
and ( n24561 , n24556 , n24560 );
and ( n24562 , n23446 , n21927 );
and ( n24563 , n23284 , n21925 );
nor ( n24564 , n24562 , n24563 );
xnor ( n24565 , n24564 , n21937 );
and ( n24566 , n24560 , n24565 );
and ( n24567 , n24556 , n24565 );
or ( n24568 , n24561 , n24566 , n24567 );
and ( n24569 , n24552 , n24568 );
and ( n24570 , n21794 , n22252 );
and ( n24571 , n21809 , n22250 );
nor ( n24572 , n24570 , n24571 );
xnor ( n24573 , n24572 , n22258 );
and ( n24574 , n21820 , n22305 );
and ( n24575 , n21833 , n22303 );
nor ( n24576 , n24574 , n24575 );
xnor ( n24577 , n24576 , n22315 );
and ( n24578 , n24573 , n24577 );
and ( n24579 , n21932 , n22323 );
and ( n24580 , n21895 , n22321 );
nor ( n24581 , n24579 , n24580 );
xnor ( n24582 , n24581 , n22329 );
and ( n24583 , n24577 , n24582 );
and ( n24584 , n24573 , n24582 );
or ( n24585 , n24578 , n24583 , n24584 );
and ( n24586 , n24568 , n24585 );
and ( n24587 , n24552 , n24585 );
or ( n24588 , n24569 , n24586 , n24587 );
and ( n24589 , n24551 , n24588 );
and ( n24590 , n21995 , n21735 );
and ( n24591 , n21972 , n21732 );
nor ( n24592 , n24590 , n24591 );
xnor ( n24593 , n24592 , n21730 );
and ( n24594 , n21885 , n21854 );
and ( n24595 , n22273 , n21852 );
nor ( n24596 , n24594 , n24595 );
xnor ( n24597 , n24596 , n21864 );
and ( n24598 , n24593 , n24597 );
and ( n24599 , n21908 , n21779 );
and ( n24600 , n21870 , n21777 );
nor ( n24601 , n24599 , n24600 );
xnor ( n24602 , n24601 , n21789 );
and ( n24603 , n24597 , n24602 );
and ( n24604 , n24593 , n24602 );
or ( n24605 , n24598 , n24603 , n24604 );
and ( n24606 , n22014 , n21957 );
and ( n24607 , n21919 , n21955 );
nor ( n24608 , n24606 , n24607 );
xnor ( n24609 , n24608 , n21967 );
and ( n24610 , n22056 , n21978 );
and ( n24611 , n22041 , n21976 );
nor ( n24612 , n24610 , n24611 );
xnor ( n24613 , n24612 , n21988 );
and ( n24614 , n24609 , n24613 );
and ( n24615 , n22049 , n21804 );
and ( n24616 , n22033 , n21802 );
nor ( n24617 , n24615 , n24616 );
xnor ( n24618 , n24617 , n21814 );
and ( n24619 , n24613 , n24618 );
and ( n24620 , n24609 , n24618 );
or ( n24621 , n24614 , n24619 , n24620 );
and ( n24622 , n24605 , n24621 );
and ( n24623 , n22101 , n21828 );
and ( n24624 , n22086 , n21826 );
nor ( n24625 , n24623 , n24624 );
xnor ( n24626 , n24625 , n21838 );
and ( n24627 , n22094 , n22194 );
and ( n24628 , n22080 , n22192 );
nor ( n24629 , n24627 , n24628 );
xnor ( n24630 , n24629 , n22200 );
and ( n24631 , n24626 , n24630 );
and ( n24632 , n23954 , n22022 );
and ( n24633 , n23575 , n22020 );
nor ( n24634 , n24632 , n24633 );
xnor ( n24635 , n24634 , n22028 );
and ( n24636 , n24630 , n24635 );
and ( n24637 , n24626 , n24635 );
or ( n24638 , n24631 , n24636 , n24637 );
and ( n24639 , n24621 , n24638 );
and ( n24640 , n24605 , n24638 );
or ( n24641 , n24622 , n24639 , n24640 );
and ( n24642 , n24588 , n24641 );
and ( n24643 , n24551 , n24641 );
or ( n24644 , n24589 , n24642 , n24643 );
and ( n24645 , n24536 , n24644 );
xor ( n24646 , n24402 , n24406 );
xor ( n24647 , n24646 , n24411 );
xor ( n24648 , n24421 , n24425 );
xor ( n24649 , n24648 , n24430 );
and ( n24650 , n24647 , n24649 );
xor ( n24651 , n24437 , n24441 );
xor ( n24652 , n24651 , n24447 );
and ( n24653 , n24649 , n24652 );
and ( n24654 , n24647 , n24652 );
or ( n24655 , n24650 , n24653 , n24654 );
xor ( n24656 , n24371 , n24375 );
xor ( n24657 , n24656 , n24378 );
and ( n24658 , n24655 , n24657 );
xor ( n24659 , n24388 , n24397 );
xor ( n24660 , n24659 , n24414 );
and ( n24661 , n24657 , n24660 );
and ( n24662 , n24655 , n24660 );
or ( n24663 , n24658 , n24661 , n24662 );
and ( n24664 , n24644 , n24663 );
and ( n24665 , n24536 , n24663 );
or ( n24666 , n24645 , n24664 , n24665 );
and ( n24667 , n24514 , n24666 );
xor ( n24668 , n24322 , n24348 );
xor ( n24669 , n24668 , n24384 );
and ( n24670 , n24666 , n24669 );
and ( n24671 , n24514 , n24669 );
or ( n24672 , n24667 , n24670 , n24671 );
and ( n24673 , n24508 , n24672 );
and ( n24674 , n24486 , n24672 );
or ( n24675 , n24509 , n24673 , n24674 );
and ( n24676 , n24484 , n24675 );
xor ( n24677 , n24127 , n24151 );
xor ( n24678 , n24677 , n24153 );
and ( n24679 , n24675 , n24678 );
and ( n24680 , n24484 , n24678 );
or ( n24681 , n24676 , n24679 , n24680 );
and ( n24682 , n24481 , n24681 );
and ( n24683 , n24479 , n24681 );
or ( n24684 , n24482 , n24682 , n24683 );
xor ( n24685 , n24120 , n24159 );
xor ( n24686 , n24685 , n24162 );
and ( n24687 , n24684 , n24686 );
xor ( n24688 , n24122 , n24124 );
xor ( n24689 , n24688 , n24156 );
xor ( n24690 , n24216 , n24283 );
xor ( n24691 , n24690 , n24476 );
xor ( n24692 , n24253 , n24255 );
xor ( n24693 , n24692 , n24280 );
xor ( n24694 , n24387 , n24470 );
xor ( n24695 , n24694 , n24473 );
and ( n24696 , n24693 , n24695 );
xor ( n24697 , n24462 , n24464 );
xor ( n24698 , n24697 , n24467 );
xor ( n24699 , n24365 , n24366 );
xor ( n24700 , n24699 , n24381 );
xor ( n24701 , n24417 , n24456 );
xor ( n24702 , n24701 , n24459 );
and ( n24703 , n24700 , n24702 );
xor ( n24704 , n24495 , n24499 );
xor ( n24705 , n24704 , n24502 );
and ( n24706 , n24702 , n24705 );
and ( n24707 , n24700 , n24705 );
or ( n24708 , n24703 , n24706 , n24707 );
and ( n24709 , n24698 , n24708 );
xor ( n24710 , n24511 , n24513 );
xor ( n24711 , n24433 , n24450 );
xor ( n24712 , n24711 , n24453 );
xor ( n24713 , n24523 , n24527 );
xor ( n24714 , n24713 , n24530 );
xor ( n24715 , n24546 , n24550 );
and ( n24716 , n24714 , n24715 );
xor ( n24717 , n24556 , n24560 );
xor ( n24718 , n24717 , n24565 );
xor ( n24719 , n24573 , n24577 );
xor ( n24720 , n24719 , n24582 );
and ( n24721 , n24718 , n24720 );
xor ( n24722 , n24540 , n24545 );
and ( n24723 , n24720 , n24722 );
and ( n24724 , n24718 , n24722 );
or ( n24725 , n24721 , n24723 , n24724 );
and ( n24726 , n24715 , n24725 );
and ( n24727 , n24714 , n24725 );
or ( n24728 , n24716 , n24726 , n24727 );
and ( n24729 , n24712 , n24728 );
and ( n24730 , n21833 , n22252 );
and ( n24731 , n21794 , n22250 );
nor ( n24732 , n24730 , n24731 );
xnor ( n24733 , n24732 , n22258 );
and ( n24734 , n21870 , n21854 );
and ( n24735 , n21885 , n21852 );
nor ( n24736 , n24734 , n24735 );
xnor ( n24737 , n24736 , n21864 );
and ( n24738 , n24733 , n24737 );
and ( n24739 , n21919 , n22323 );
and ( n24740 , n21932 , n22321 );
nor ( n24741 , n24739 , n24740 );
xnor ( n24742 , n24741 , n22329 );
and ( n24743 , n24737 , n24742 );
and ( n24744 , n24733 , n24742 );
or ( n24745 , n24738 , n24743 , n24744 );
and ( n24746 , n24544 , n22062 );
and ( n24747 , n24446 , n22060 );
nor ( n24748 , n24746 , n24747 );
xnor ( n24749 , n24748 , n22068 );
xor ( n24750 , n21503 , n21667 );
buf ( n552013 , n24750 );
buf ( n552014 , n552013 );
buf ( n24753 , n552014 );
and ( n24754 , n24753 , n22035 );
and ( n24755 , n24749 , n24754 );
and ( n24756 , n24745 , n24755 );
and ( n24757 , n22409 , n22194 );
and ( n24758 , n22094 , n22192 );
nor ( n24759 , n24757 , n24758 );
xnor ( n24760 , n24759 , n22200 );
and ( n24761 , n23074 , n21880 );
and ( n24762 , n22659 , n21878 );
nor ( n24763 , n24761 , n24762 );
xnor ( n24764 , n24763 , n21890 );
and ( n24765 , n24760 , n24764 );
and ( n24766 , n24755 , n24765 );
and ( n24767 , n24745 , n24765 );
or ( n24768 , n24756 , n24766 , n24767 );
and ( n24769 , n22273 , n22305 );
and ( n24770 , n21820 , n22303 );
nor ( n24771 , n24769 , n24770 );
xnor ( n24772 , n24771 , n22315 );
and ( n24773 , n21895 , n21779 );
and ( n24774 , n21908 , n21777 );
nor ( n24775 , n24773 , n24774 );
xnor ( n24776 , n24775 , n21789 );
and ( n24777 , n24772 , n24776 );
and ( n24778 , n22041 , n21957 );
and ( n24779 , n22014 , n21955 );
nor ( n24780 , n24778 , n24779 );
xnor ( n24781 , n24780 , n21967 );
and ( n24782 , n24776 , n24781 );
and ( n24783 , n24772 , n24781 );
or ( n24784 , n24777 , n24782 , n24783 );
xor ( n24785 , n24593 , n24597 );
xor ( n24786 , n24785 , n24602 );
and ( n24787 , n24784 , n24786 );
xor ( n24788 , n24609 , n24613 );
xor ( n24789 , n24788 , n24618 );
and ( n24790 , n24786 , n24789 );
and ( n24791 , n24784 , n24789 );
or ( n24792 , n24787 , n24790 , n24791 );
and ( n24793 , n24768 , n24792 );
xor ( n24794 , n24552 , n24568 );
xor ( n24795 , n24794 , n24585 );
and ( n24796 , n24792 , n24795 );
and ( n24797 , n24768 , n24795 );
or ( n24798 , n24793 , n24796 , n24797 );
and ( n24799 , n24728 , n24798 );
and ( n24800 , n24712 , n24798 );
or ( n24801 , n24729 , n24799 , n24800 );
and ( n24802 , n24710 , n24801 );
xor ( n24803 , n24516 , n24518 );
xor ( n24804 , n24803 , n24533 );
xor ( n24805 , n24551 , n24588 );
xor ( n24806 , n24805 , n24641 );
and ( n24807 , n24804 , n24806 );
xor ( n24808 , n24655 , n24657 );
xor ( n24809 , n24808 , n24660 );
and ( n24810 , n24806 , n24809 );
and ( n24811 , n24804 , n24809 );
or ( n24812 , n24807 , n24810 , n24811 );
and ( n24813 , n24801 , n24812 );
and ( n24814 , n24710 , n24812 );
or ( n24815 , n24802 , n24813 , n24814 );
and ( n24816 , n24708 , n24815 );
and ( n24817 , n24698 , n24815 );
or ( n24818 , n24709 , n24816 , n24817 );
and ( n24819 , n24695 , n24818 );
and ( n24820 , n24693 , n24818 );
or ( n24821 , n24696 , n24819 , n24820 );
and ( n24822 , n24691 , n24821 );
xor ( n24823 , n24484 , n24675 );
xor ( n24824 , n24823 , n24678 );
and ( n24825 , n24821 , n24824 );
and ( n24826 , n24691 , n24824 );
or ( n24827 , n24822 , n24825 , n24826 );
and ( n24828 , n24689 , n24827 );
xor ( n24829 , n24479 , n24481 );
xor ( n24830 , n24829 , n24681 );
and ( n24831 , n24827 , n24830 );
and ( n24832 , n24689 , n24830 );
or ( n24833 , n24828 , n24831 , n24832 );
and ( n24834 , n24686 , n24833 );
and ( n24835 , n24684 , n24833 );
or ( n24836 , n24687 , n24834 , n24835 );
and ( n24837 , n24167 , n24836 );
and ( n24838 , n24165 , n24836 );
or ( n24839 , n24168 , n24837 , n24838 );
and ( n24840 , n24117 , n24839 );
and ( n24841 , n24115 , n24839 );
or ( n24842 , n24118 , n24840 , n24841 );
and ( n24843 , n24112 , n24842 );
and ( n24844 , n24110 , n24842 );
or ( n24845 , n24113 , n24843 , n24844 );
and ( n24846 , n23720 , n24845 );
and ( n24847 , n23674 , n24845 );
or ( n24848 , n23721 , n24846 , n24847 );
and ( n24849 , n23671 , n24848 );
and ( n24850 , n23437 , n24848 );
or ( n24851 , n23672 , n24849 , n24850 );
and ( n24852 , n23434 , n24851 );
and ( n24853 , n23390 , n24851 );
or ( n24854 , n23435 , n24852 , n24853 );
and ( n24855 , n23388 , n24854 );
xor ( n24856 , n23388 , n24854 );
xor ( n24857 , n23390 , n23434 );
xor ( n24858 , n24857 , n24851 );
xor ( n24859 , n23437 , n23671 );
xor ( n24860 , n24859 , n24848 );
xor ( n24861 , n23674 , n23720 );
xor ( n24862 , n24861 , n24845 );
xor ( n24863 , n24110 , n24112 );
xor ( n24864 , n24863 , n24842 );
xor ( n24865 , n24115 , n24117 );
xor ( n24866 , n24865 , n24839 );
xor ( n24867 , n24165 , n24167 );
xor ( n24868 , n24867 , n24836 );
xor ( n24869 , n24684 , n24686 );
xor ( n24870 , n24869 , n24833 );
xor ( n24871 , n24689 , n24827 );
xor ( n24872 , n24871 , n24830 );
xor ( n24873 , n24486 , n24508 );
xor ( n24874 , n24873 , n24672 );
xor ( n24875 , n24488 , n24490 );
xor ( n24876 , n24875 , n24505 );
xor ( n24877 , n24514 , n24666 );
xor ( n24878 , n24877 , n24669 );
and ( n24879 , n24876 , n24878 );
xor ( n24880 , n24536 , n24644 );
xor ( n24881 , n24880 , n24663 );
xor ( n24882 , n24605 , n24621 );
xor ( n24883 , n24882 , n24638 );
xor ( n24884 , n24647 , n24649 );
xor ( n24885 , n24884 , n24652 );
and ( n24886 , n24883 , n24885 );
xor ( n24887 , n24626 , n24630 );
xor ( n24888 , n24887 , n24635 );
and ( n24889 , n24753 , n22062 );
and ( n24890 , n24544 , n22060 );
nor ( n24891 , n24889 , n24890 );
xnor ( n24892 , n24891 , n22068 );
xor ( n24893 , n21505 , n21666 );
buf ( n552156 , n24893 );
buf ( n552157 , n552156 );
buf ( n24896 , n552157 );
and ( n24897 , n24896 , n22035 );
and ( n24898 , n24892 , n24897 );
and ( n24899 , n24011 , n22022 );
and ( n24900 , n23954 , n22020 );
nor ( n24901 , n24899 , n24900 );
xnor ( n24902 , n24901 , n22028 );
and ( n24903 , n24898 , n24902 );
and ( n24904 , n24888 , n24903 );
and ( n24905 , n22086 , n21804 );
and ( n24906 , n22049 , n21802 );
nor ( n24907 , n24905 , n24906 );
xnor ( n24908 , n24907 , n21814 );
and ( n24909 , n22080 , n21828 );
and ( n24910 , n22101 , n21826 );
nor ( n24911 , n24909 , n24910 );
xnor ( n24912 , n24911 , n21838 );
and ( n24913 , n24908 , n24912 );
xor ( n24914 , n24733 , n24737 );
xor ( n24915 , n24914 , n24742 );
and ( n24916 , n24912 , n24915 );
and ( n24917 , n24908 , n24915 );
or ( n24918 , n24913 , n24916 , n24917 );
and ( n24919 , n24903 , n24918 );
and ( n24920 , n24888 , n24918 );
or ( n24921 , n24904 , n24919 , n24920 );
and ( n24922 , n24885 , n24921 );
and ( n24923 , n24883 , n24921 );
or ( n24924 , n24886 , n24922 , n24923 );
xor ( n24925 , n24749 , n24754 );
xor ( n24926 , n24760 , n24764 );
and ( n24927 , n24925 , n24926 );
and ( n24928 , n21794 , n21735 );
and ( n24929 , n21809 , n21732 );
nor ( n24930 , n24928 , n24929 );
xnor ( n24931 , n24930 , n21730 );
and ( n24932 , n21820 , n22252 );
and ( n24933 , n21833 , n22250 );
nor ( n24934 , n24932 , n24933 );
xnor ( n24935 , n24934 , n22258 );
and ( n24936 , n24931 , n24935 );
and ( n24937 , n21885 , n22305 );
and ( n24938 , n22273 , n22303 );
nor ( n24939 , n24937 , n24938 );
xnor ( n24940 , n24939 , n22315 );
and ( n24941 , n24935 , n24940 );
and ( n24942 , n24931 , n24940 );
or ( n24943 , n24936 , n24941 , n24942 );
and ( n24944 , n24926 , n24943 );
and ( n24945 , n24925 , n24943 );
or ( n24946 , n24927 , n24944 , n24945 );
xor ( n24947 , n24718 , n24720 );
xor ( n24948 , n24947 , n24722 );
and ( n24949 , n24946 , n24948 );
xor ( n24950 , n24745 , n24755 );
xor ( n24951 , n24950 , n24765 );
and ( n24952 , n24948 , n24951 );
and ( n24953 , n24946 , n24951 );
or ( n24954 , n24949 , n24952 , n24953 );
xor ( n24955 , n24714 , n24715 );
xor ( n24956 , n24955 , n24725 );
and ( n24957 , n24954 , n24956 );
xor ( n24958 , n24768 , n24792 );
xor ( n24959 , n24958 , n24795 );
and ( n24960 , n24956 , n24959 );
and ( n24961 , n24954 , n24959 );
or ( n24962 , n24957 , n24960 , n24961 );
and ( n24963 , n24924 , n24962 );
xor ( n24964 , n24712 , n24728 );
xor ( n24965 , n24964 , n24798 );
and ( n24966 , n24962 , n24965 );
and ( n24967 , n24924 , n24965 );
or ( n24968 , n24963 , n24966 , n24967 );
and ( n24969 , n24881 , n24968 );
xor ( n24970 , n24700 , n24702 );
xor ( n24971 , n24970 , n24705 );
and ( n24972 , n24968 , n24971 );
and ( n24973 , n24881 , n24971 );
or ( n24974 , n24969 , n24972 , n24973 );
and ( n24975 , n24878 , n24974 );
and ( n24976 , n24876 , n24974 );
or ( n24977 , n24879 , n24975 , n24976 );
and ( n24978 , n24874 , n24977 );
xor ( n24979 , n24693 , n24695 );
xor ( n24980 , n24979 , n24818 );
and ( n24981 , n24977 , n24980 );
and ( n24982 , n24874 , n24980 );
or ( n24983 , n24978 , n24981 , n24982 );
xor ( n24984 , n24691 , n24821 );
xor ( n24985 , n24984 , n24824 );
and ( n24986 , n24983 , n24985 );
xor ( n24987 , n24983 , n24985 );
xor ( n24988 , n24698 , n24708 );
xor ( n24989 , n24988 , n24815 );
xor ( n24990 , n24710 , n24801 );
xor ( n24991 , n24990 , n24812 );
xor ( n24992 , n24804 , n24806 );
xor ( n24993 , n24992 , n24809 );
xor ( n24994 , n24784 , n24786 );
xor ( n24995 , n24994 , n24789 );
xor ( n24996 , n24892 , n24897 );
and ( n24997 , n24896 , n22062 );
and ( n24998 , n24753 , n22060 );
nor ( n24999 , n24997 , n24998 );
xnor ( n25000 , n24999 , n22068 );
xor ( n25001 , n21507 , n21665 );
buf ( n552264 , n25001 );
buf ( n552265 , n552264 );
buf ( n25004 , n552265 );
and ( n25005 , n25004 , n22035 );
and ( n25006 , n25000 , n25005 );
and ( n25007 , n24996 , n25006 );
and ( n25008 , n24446 , n22022 );
and ( n25009 , n24011 , n22020 );
nor ( n25010 , n25008 , n25009 );
xnor ( n25011 , n25010 , n22028 );
and ( n25012 , n25006 , n25011 );
and ( n25013 , n24996 , n25011 );
or ( n25014 , n25007 , n25012 , n25013 );
and ( n25015 , n23284 , n21903 );
and ( n25016 , n23165 , n21901 );
nor ( n25017 , n25015 , n25016 );
xnor ( n25018 , n25017 , n21913 );
and ( n25019 , n25014 , n25018 );
and ( n25020 , n23575 , n21927 );
and ( n25021 , n23446 , n21925 );
nor ( n25022 , n25020 , n25021 );
xnor ( n25023 , n25022 , n21937 );
and ( n25024 , n25018 , n25023 );
and ( n25025 , n25014 , n25023 );
or ( n25026 , n25019 , n25024 , n25025 );
and ( n25027 , n24995 , n25026 );
and ( n25028 , n22049 , n21978 );
and ( n25029 , n22033 , n21976 );
nor ( n25030 , n25028 , n25029 );
xnor ( n25031 , n25030 , n21988 );
and ( n25032 , n22101 , n21804 );
and ( n25033 , n22086 , n21802 );
nor ( n25034 , n25032 , n25033 );
xnor ( n25035 , n25034 , n21814 );
and ( n25036 , n25031 , n25035 );
and ( n25037 , n22094 , n21828 );
and ( n25038 , n22080 , n21826 );
nor ( n25039 , n25037 , n25038 );
xnor ( n25040 , n25039 , n21838 );
and ( n25041 , n25035 , n25040 );
and ( n25042 , n25031 , n25040 );
or ( n25043 , n25036 , n25041 , n25042 );
xor ( n25044 , n24772 , n24776 );
xor ( n25045 , n25044 , n24781 );
and ( n25046 , n25043 , n25045 );
xor ( n25047 , n24898 , n24902 );
and ( n25048 , n25045 , n25047 );
and ( n25049 , n25043 , n25047 );
or ( n25050 , n25046 , n25048 , n25049 );
and ( n25051 , n25026 , n25050 );
and ( n25052 , n24995 , n25050 );
or ( n25053 , n25027 , n25051 , n25052 );
and ( n25054 , n23165 , n21880 );
and ( n25055 , n23074 , n21878 );
nor ( n25056 , n25054 , n25055 );
xnor ( n25057 , n25056 , n21890 );
and ( n25058 , n23954 , n21927 );
and ( n25059 , n23575 , n21925 );
nor ( n25060 , n25058 , n25059 );
xnor ( n25061 , n25060 , n21937 );
and ( n25062 , n25057 , n25061 );
and ( n25063 , n23284 , n21880 );
and ( n25064 , n23165 , n21878 );
nor ( n25065 , n25063 , n25064 );
xnor ( n25066 , n25065 , n21890 );
and ( n25067 , n24011 , n21927 );
and ( n25068 , n23954 , n21925 );
nor ( n25069 , n25067 , n25068 );
xnor ( n25070 , n25069 , n21937 );
and ( n25071 , n25066 , n25070 );
and ( n25072 , n25061 , n25071 );
and ( n25073 , n25057 , n25071 );
or ( n25074 , n25062 , n25072 , n25073 );
and ( n25075 , n21833 , n21735 );
and ( n25076 , n21794 , n21732 );
nor ( n25077 , n25075 , n25076 );
xnor ( n25078 , n25077 , n21730 );
and ( n552341 , n22273 , n22252 );
and ( n552342 , n21820 , n22250 );
nor ( n25079 , n552341 , n552342 );
xnor ( n25080 , n25079 , n22258 );
and ( n25081 , n25078 , n25080 );
and ( n25082 , n21895 , n21854 );
and ( n25083 , n21908 , n21852 );
nor ( n25084 , n25082 , n25083 );
xnor ( n25085 , n25084 , n21864 );
and ( n25086 , n22041 , n22323 );
and ( n25087 , n22014 , n22321 );
nor ( n25088 , n25086 , n25087 );
xnor ( n25089 , n25088 , n22329 );
and ( n25090 , n25085 , n25089 );
and ( n25091 , n22033 , n21957 );
and ( n25092 , n22056 , n21955 );
nor ( n25093 , n25091 , n25092 );
xnor ( n25094 , n25093 , n21967 );
and ( n25095 , n25089 , n25094 );
and ( n25096 , n25085 , n25094 );
or ( n25097 , n25090 , n25095 , n25096 );
and ( n25098 , n25081 , n25097 );
and ( n25099 , n22080 , n21804 );
and ( n25100 , n22101 , n21802 );
nor ( n25101 , n25099 , n25100 );
xnor ( n25102 , n25101 , n21814 );
and ( n25103 , n23074 , n22194 );
and ( n25104 , n22659 , n22192 );
nor ( n25105 , n25103 , n25104 );
xnor ( n25106 , n25105 , n22200 );
and ( n25107 , n25102 , n25106 );
and ( n25108 , n23575 , n21903 );
and ( n25109 , n23446 , n21901 );
nor ( n25110 , n25108 , n25109 );
xnor ( n25111 , n25110 , n21913 );
and ( n25112 , n25106 , n25111 );
and ( n25113 , n25102 , n25111 );
or ( n25114 , n25107 , n25112 , n25113 );
and ( n25115 , n25097 , n25114 );
and ( n25116 , n25081 , n25114 );
or ( n25117 , n25098 , n25115 , n25116 );
and ( n25118 , n25074 , n25117 );
xor ( n25119 , n24908 , n24912 );
xor ( n25120 , n25119 , n24915 );
and ( n25121 , n25117 , n25120 );
and ( n25122 , n25074 , n25120 );
or ( n25123 , n25118 , n25121 , n25122 );
xor ( n25124 , n24888 , n24903 );
xor ( n25125 , n25124 , n24918 );
and ( n25126 , n25123 , n25125 );
xor ( n25127 , n24946 , n24948 );
xor ( n25128 , n25127 , n24951 );
and ( n25129 , n25125 , n25128 );
and ( n25130 , n25123 , n25128 );
or ( n25131 , n25126 , n25129 , n25130 );
and ( n25132 , n25053 , n25131 );
xor ( n25133 , n24883 , n24885 );
xor ( n25134 , n25133 , n24921 );
and ( n25135 , n25131 , n25134 );
and ( n25136 , n25053 , n25134 );
or ( n25137 , n25132 , n25135 , n25136 );
and ( n25138 , n24993 , n25137 );
xor ( n25139 , n24924 , n24962 );
xor ( n25140 , n25139 , n24965 );
and ( n25141 , n25137 , n25140 );
and ( n25142 , n24993 , n25140 );
or ( n25143 , n25138 , n25141 , n25142 );
and ( n25144 , n24991 , n25143 );
xor ( n25145 , n24881 , n24968 );
xor ( n25146 , n25145 , n24971 );
and ( n25147 , n25143 , n25146 );
and ( n25148 , n24991 , n25146 );
or ( n25149 , n25144 , n25147 , n25148 );
and ( n25150 , n24989 , n25149 );
xor ( n25151 , n24876 , n24878 );
xor ( n25152 , n25151 , n24974 );
and ( n25153 , n25149 , n25152 );
and ( n25154 , n24989 , n25152 );
or ( n25155 , n25150 , n25153 , n25154 );
xor ( n25156 , n24874 , n24977 );
xor ( n25157 , n25156 , n24980 );
and ( n25158 , n25155 , n25157 );
xor ( n25159 , n25155 , n25157 );
xor ( n25160 , n24989 , n25149 );
xor ( n25161 , n25160 , n25152 );
xor ( n25162 , n24991 , n25143 );
xor ( n25163 , n25162 , n25146 );
xor ( n25164 , n24954 , n24956 );
xor ( n25165 , n25164 , n24959 );
and ( n25166 , n22659 , n22194 );
and ( n25167 , n22409 , n22192 );
nor ( n25168 , n25166 , n25167 );
xnor ( n25169 , n25168 , n22200 );
and ( n25170 , n23446 , n21903 );
and ( n25171 , n23284 , n21901 );
nor ( n25172 , n25170 , n25171 );
xnor ( n25173 , n25172 , n21913 );
and ( n25174 , n25169 , n25173 );
xor ( n25175 , n24996 , n25006 );
xor ( n25176 , n25175 , n25011 );
and ( n25177 , n25173 , n25176 );
and ( n25178 , n25169 , n25176 );
or ( n25179 , n25174 , n25177 , n25178 );
and ( n25180 , n22033 , n21978 );
and ( n25181 , n22056 , n21976 );
nor ( n25182 , n25180 , n25181 );
xnor ( n25183 , n25182 , n21988 );
and ( n25184 , n25179 , n25183 );
xor ( n25185 , n25014 , n25018 );
xor ( n25186 , n25185 , n25023 );
and ( n25187 , n25183 , n25186 );
and ( n25188 , n25179 , n25186 );
or ( n25189 , n25184 , n25187 , n25188 );
xor ( n25190 , n24925 , n24926 );
xor ( n25191 , n25190 , n24943 );
xor ( n25192 , n24931 , n24935 );
xor ( n25193 , n25192 , n24940 );
xor ( n25194 , n25031 , n25035 );
xor ( n25195 , n25194 , n25040 );
and ( n25196 , n25193 , n25195 );
and ( n25197 , n24544 , n22022 );
and ( n25198 , n24446 , n22020 );
nor ( n25199 , n25197 , n25198 );
xnor ( n25200 , n25199 , n22028 );
xor ( n25201 , n25000 , n25005 );
and ( n25202 , n25200 , n25201 );
xor ( n25203 , n25066 , n25070 );
and ( n25204 , n25201 , n25203 );
and ( n25205 , n25200 , n25203 );
or ( n25206 , n25202 , n25204 , n25205 );
and ( n25207 , n25195 , n25206 );
and ( n25208 , n25193 , n25206 );
or ( n25209 , n25196 , n25207 , n25208 );
and ( n25210 , n25191 , n25209 );
xor ( n25211 , n25078 , n25080 );
and ( n25212 , n22659 , n21828 );
and ( n25213 , n22409 , n21826 );
nor ( n25214 , n25212 , n25213 );
xnor ( n25215 , n25214 , n21838 );
and ( n25216 , n23165 , n22194 );
and ( n25217 , n23074 , n22192 );
nor ( n25218 , n25216 , n25217 );
xnor ( n25219 , n25218 , n22200 );
and ( n25220 , n25215 , n25219 );
and ( n25221 , n23446 , n21880 );
and ( n25222 , n23284 , n21878 );
nor ( n25223 , n25221 , n25222 );
xnor ( n25224 , n25223 , n21890 );
and ( n25225 , n25219 , n25224 );
and ( n25226 , n25215 , n25224 );
or ( n25227 , n25220 , n25225 , n25226 );
and ( n25228 , n25211 , n25227 );
and ( n25229 , n21885 , n22252 );
and ( n25230 , n22273 , n22250 );
nor ( n25231 , n25229 , n25230 );
xnor ( n25232 , n25231 , n22258 );
and ( n25233 , n21932 , n21854 );
and ( n25234 , n21895 , n21852 );
nor ( n25235 , n25233 , n25234 );
xnor ( n25236 , n25235 , n21864 );
and ( n25237 , n25232 , n25236 );
and ( n25238 , n22014 , n21779 );
and ( n25239 , n21919 , n21777 );
nor ( n25240 , n25238 , n25239 );
xnor ( n25241 , n25240 , n21789 );
and ( n25242 , n25236 , n25241 );
and ( n25243 , n25232 , n25241 );
or ( n25244 , n25237 , n25242 , n25243 );
and ( n25245 , n25227 , n25244 );
and ( n25246 , n25211 , n25244 );
or ( n25247 , n25228 , n25245 , n25246 );
and ( n25248 , n22056 , n22323 );
and ( n25249 , n22041 , n22321 );
nor ( n25250 , n25248 , n25249 );
xnor ( n25251 , n25250 , n22329 );
and ( n25252 , n22094 , n21804 );
and ( n25253 , n22080 , n21802 );
nor ( n25254 , n25252 , n25253 );
xnor ( n25255 , n25254 , n21814 );
and ( n25256 , n25251 , n25255 );
and ( n25257 , n24753 , n22022 );
and ( n25258 , n24544 , n22020 );
nor ( n25259 , n25257 , n25258 );
xnor ( n25260 , n25259 , n22028 );
and ( n25261 , n25255 , n25260 );
and ( n25262 , n25251 , n25260 );
or ( n25263 , n25256 , n25261 , n25262 );
xor ( n25264 , n25085 , n25089 );
xor ( n25265 , n25264 , n25094 );
and ( n25266 , n25263 , n25265 );
xor ( n25267 , n25102 , n25106 );
xor ( n25268 , n25267 , n25111 );
and ( n25269 , n25265 , n25268 );
and ( n25270 , n25263 , n25268 );
or ( n25271 , n25266 , n25269 , n25270 );
and ( n25272 , n25247 , n25271 );
xor ( n25273 , n25057 , n25061 );
xor ( n25274 , n25273 , n25071 );
and ( n25275 , n25271 , n25274 );
and ( n25276 , n25247 , n25274 );
or ( n25277 , n25272 , n25275 , n25276 );
and ( n25278 , n25209 , n25277 );
and ( n25279 , n25191 , n25277 );
or ( n25280 , n25210 , n25278 , n25279 );
and ( n25281 , n25189 , n25280 );
xor ( n25282 , n24995 , n25026 );
xor ( n25283 , n25282 , n25050 );
and ( n25284 , n25280 , n25283 );
and ( n25285 , n25189 , n25283 );
or ( n25286 , n25281 , n25284 , n25285 );
and ( n25287 , n25165 , n25286 );
xor ( n25288 , n25053 , n25131 );
xor ( n25289 , n25288 , n25134 );
and ( n25290 , n25286 , n25289 );
and ( n25291 , n25165 , n25289 );
or ( n25292 , n25287 , n25290 , n25291 );
xor ( n25293 , n24993 , n25137 );
xor ( n25294 , n25293 , n25140 );
and ( n25295 , n25292 , n25294 );
xor ( n25296 , n25123 , n25125 );
xor ( n25297 , n25296 , n25128 );
and ( n25298 , n22014 , n22323 );
and ( n25299 , n21919 , n22321 );
nor ( n25300 , n25298 , n25299 );
xnor ( n25301 , n25300 , n22329 );
and ( n25302 , n22056 , n21957 );
and ( n25303 , n22041 , n21955 );
nor ( n25304 , n25302 , n25303 );
xnor ( n25305 , n25304 , n21967 );
and ( n25306 , n25301 , n25305 );
xor ( n25307 , n25169 , n25173 );
xor ( n25308 , n25307 , n25176 );
and ( n25309 , n25305 , n25308 );
and ( n25310 , n25301 , n25308 );
or ( n25311 , n25306 , n25309 , n25310 );
and ( n25312 , n21809 , n21735 );
and ( n25313 , n21995 , n21732 );
nor ( n25314 , n25312 , n25313 );
xnor ( n25315 , n25314 , n21730 );
and ( n25316 , n25311 , n25315 );
xor ( n25317 , n25179 , n25183 );
xor ( n25318 , n25317 , n25186 );
and ( n25319 , n25315 , n25318 );
and ( n25320 , n25311 , n25318 );
or ( n25321 , n25316 , n25319 , n25320 );
and ( n25322 , n25297 , n25321 );
xor ( n25323 , n25043 , n25045 );
xor ( n25324 , n25323 , n25047 );
xor ( n25325 , n25074 , n25117 );
xor ( n25326 , n25325 , n25120 );
and ( n25327 , n25324 , n25326 );
xor ( n25328 , n25081 , n25097 );
xor ( n25329 , n25328 , n25114 );
and ( n25330 , n25004 , n22062 );
and ( n25331 , n24896 , n22060 );
nor ( n25332 , n25330 , n25331 );
xnor ( n25333 , n25332 , n22068 );
xor ( n25334 , n21509 , n21664 );
buf ( n552599 , n25334 );
buf ( n552600 , n552599 );
buf ( n25337 , n552600 );
and ( n25338 , n25337 , n22035 );
and ( n25339 , n25333 , n25338 );
and ( n25340 , n24896 , n22022 );
and ( n25341 , n24753 , n22020 );
nor ( n25342 , n25340 , n25341 );
xnor ( n25343 , n25342 , n22028 );
xor ( n25344 , n21537 , n21662 );
buf ( n552609 , n25344 );
buf ( n552610 , n552609 );
buf ( n25347 , n552610 );
and ( n25348 , n25347 , n22035 );
and ( n25349 , n25343 , n25348 );
and ( n25350 , n25338 , n25349 );
and ( n25351 , n25333 , n25349 );
or ( n25352 , n25339 , n25350 , n25351 );
and ( n25353 , n22273 , n21735 );
and ( n25354 , n21820 , n21732 );
nor ( n25355 , n25353 , n25354 );
xnor ( n25356 , n25355 , n21730 );
and ( n25357 , n21870 , n22252 );
and ( n25358 , n21885 , n22250 );
nor ( n25359 , n25357 , n25358 );
xnor ( n25360 , n25359 , n22258 );
and ( n25361 , n25356 , n25360 );
and ( n25362 , n21895 , n22305 );
and ( n25363 , n21908 , n22303 );
nor ( n25364 , n25362 , n25363 );
xnor ( n25365 , n25364 , n22315 );
and ( n25366 , n25360 , n25365 );
and ( n25367 , n25356 , n25365 );
or ( n25368 , n25361 , n25366 , n25367 );
and ( n25369 , n21919 , n21854 );
and ( n25370 , n21932 , n21852 );
nor ( n25371 , n25369 , n25370 );
xnor ( n25372 , n25371 , n21864 );
and ( n25373 , n22033 , n22323 );
and ( n25374 , n22056 , n22321 );
nor ( n25375 , n25373 , n25374 );
xnor ( n25376 , n25375 , n22329 );
and ( n25377 , n25372 , n25376 );
and ( n25378 , n22080 , n21978 );
and ( n25379 , n22101 , n21976 );
nor ( n25380 , n25378 , n25379 );
xnor ( n25381 , n25380 , n21988 );
and ( n25382 , n25376 , n25381 );
and ( n25383 , n25372 , n25381 );
or ( n25384 , n25377 , n25382 , n25383 );
and ( n25385 , n25368 , n25384 );
xor ( n25386 , n25232 , n25236 );
xor ( n25387 , n25386 , n25241 );
and ( n25388 , n25384 , n25387 );
and ( n25389 , n25368 , n25387 );
or ( n25390 , n25385 , n25388 , n25389 );
and ( n25391 , n25352 , n25390 );
xor ( n25392 , n25200 , n25201 );
xor ( n25393 , n25392 , n25203 );
and ( n25394 , n25390 , n25393 );
and ( n25395 , n25352 , n25393 );
or ( n25396 , n25391 , n25394 , n25395 );
and ( n25397 , n25329 , n25396 );
xor ( n25398 , n25193 , n25195 );
xor ( n25399 , n25398 , n25206 );
and ( n25400 , n25396 , n25399 );
and ( n25401 , n25329 , n25399 );
or ( n25402 , n25397 , n25400 , n25401 );
and ( n25403 , n25326 , n25402 );
and ( n25404 , n25324 , n25402 );
or ( n25405 , n25327 , n25403 , n25404 );
and ( n25406 , n25321 , n25405 );
and ( n25407 , n25297 , n25405 );
or ( n25408 , n25322 , n25406 , n25407 );
xor ( n25409 , n25165 , n25286 );
xor ( n25410 , n25409 , n25289 );
and ( n25411 , n25408 , n25410 );
xor ( n25412 , n25189 , n25280 );
xor ( n25413 , n25412 , n25283 );
xor ( n25414 , n25191 , n25209 );
xor ( n25415 , n25414 , n25277 );
xor ( n25416 , n25311 , n25315 );
xor ( n25417 , n25416 , n25318 );
and ( n25418 , n25415 , n25417 );
xor ( n25419 , n25343 , n25348 );
and ( n25420 , n25347 , n22062 );
and ( n25421 , n25337 , n22060 );
nor ( n25422 , n25420 , n25421 );
xnor ( n25423 , n25422 , n22068 );
xor ( n25424 , n21560 , n21660 );
buf ( n552689 , n25424 );
buf ( n552690 , n552689 );
buf ( n25427 , n552690 );
and ( n25428 , n25427 , n22035 );
and ( n25429 , n25423 , n25428 );
and ( n25430 , n25419 , n25429 );
and ( n25431 , n25337 , n22062 );
and ( n25432 , n25004 , n22060 );
nor ( n25433 , n25431 , n25432 );
xnor ( n25434 , n25433 , n22068 );
and ( n25435 , n25429 , n25434 );
and ( n25436 , n25419 , n25434 );
or ( n25437 , n25430 , n25435 , n25436 );
and ( n25438 , n23954 , n21903 );
and ( n25439 , n23575 , n21901 );
nor ( n25440 , n25438 , n25439 );
xnor ( n25441 , n25440 , n21913 );
and ( n25442 , n25437 , n25441 );
and ( n25443 , n24446 , n21927 );
and ( n25444 , n24011 , n21925 );
nor ( n25445 , n25443 , n25444 );
xnor ( n25446 , n25445 , n21937 );
and ( n25447 , n25441 , n25446 );
and ( n25448 , n25437 , n25446 );
or ( n25449 , n25442 , n25447 , n25448 );
and ( n25450 , n22086 , n21978 );
and ( n25451 , n22049 , n21976 );
nor ( n25452 , n25450 , n25451 );
xnor ( n25453 , n25452 , n21988 );
and ( n25454 , n25449 , n25453 );
and ( n25455 , n22409 , n21828 );
and ( n25456 , n22094 , n21826 );
nor ( n25457 , n25455 , n25456 );
xnor ( n25458 , n25457 , n21838 );
and ( n25459 , n25453 , n25458 );
and ( n25460 , n25449 , n25458 );
or ( n25461 , n25454 , n25459 , n25460 );
and ( n25462 , n21908 , n21854 );
and ( n25463 , n21870 , n21852 );
nor ( n25464 , n25462 , n25463 );
xnor ( n25465 , n25464 , n21864 );
and ( n25466 , n25461 , n25465 );
and ( n25467 , n21932 , n21779 );
and ( n25468 , n21895 , n21777 );
nor ( n25469 , n25467 , n25468 );
xnor ( n25470 , n25469 , n21789 );
and ( n25471 , n25465 , n25470 );
and ( n25472 , n25461 , n25470 );
or ( n25473 , n25466 , n25471 , n25472 );
and ( n25474 , n25417 , n25473 );
and ( n25475 , n25415 , n25473 );
or ( n25476 , n25418 , n25474 , n25475 );
and ( n25477 , n25413 , n25476 );
xor ( n25478 , n25297 , n25321 );
xor ( n25479 , n25478 , n25405 );
and ( n25480 , n25476 , n25479 );
and ( n25481 , n25413 , n25479 );
or ( n25482 , n25477 , n25480 , n25481 );
and ( n25483 , n25410 , n25482 );
and ( n25484 , n25408 , n25482 );
or ( n25485 , n25411 , n25483 , n25484 );
and ( n25486 , n25294 , n25485 );
and ( n25487 , n25292 , n25485 );
or ( n25488 , n25295 , n25486 , n25487 );
and ( n25489 , n25163 , n25488 );
xor ( n25490 , n25163 , n25488 );
xor ( n25491 , n25292 , n25294 );
xor ( n25492 , n25491 , n25485 );
xor ( n25493 , n25408 , n25410 );
xor ( n25494 , n25493 , n25482 );
xor ( n25495 , n25247 , n25271 );
xor ( n25496 , n25495 , n25274 );
xor ( n25497 , n25301 , n25305 );
xor ( n25498 , n25497 , n25308 );
and ( n25499 , n25496 , n25498 );
xor ( n25500 , n25211 , n25227 );
xor ( n25501 , n25500 , n25244 );
xor ( n25502 , n25263 , n25265 );
xor ( n25503 , n25502 , n25268 );
and ( n25504 , n25501 , n25503 );
xor ( n25505 , n25251 , n25255 );
xor ( n25506 , n25505 , n25260 );
and ( n25507 , n21885 , n21735 );
and ( n25508 , n22273 , n21732 );
nor ( n25509 , n25507 , n25508 );
xnor ( n25510 , n25509 , n21730 );
and ( n25511 , n21932 , n22305 );
and ( n25512 , n21895 , n22303 );
nor ( n25513 , n25511 , n25512 );
xnor ( n25514 , n25513 , n22315 );
and ( n25515 , n25510 , n25514 );
and ( n25516 , n21908 , n22252 );
and ( n25517 , n21870 , n22250 );
nor ( n25518 , n25516 , n25517 );
xnor ( n25519 , n25518 , n22258 );
and ( n25520 , n22056 , n21779 );
and ( n25521 , n22041 , n21777 );
nor ( n25522 , n25520 , n25521 );
xnor ( n25523 , n25522 , n21789 );
and ( n25524 , n25519 , n25523 );
and ( n25525 , n22049 , n22323 );
and ( n25526 , n22033 , n22321 );
nor ( n25527 , n25525 , n25526 );
xnor ( n25528 , n25527 , n22329 );
and ( n25529 , n25523 , n25528 );
and ( n25530 , n25519 , n25528 );
or ( n25531 , n25524 , n25529 , n25530 );
and ( n25532 , n25515 , n25531 );
and ( n25533 , n22101 , n21957 );
and ( n25534 , n22086 , n21955 );
nor ( n25535 , n25533 , n25534 );
xnor ( n25536 , n25535 , n21967 );
and ( n25537 , n23446 , n22194 );
and ( n25538 , n23284 , n22192 );
nor ( n25539 , n25537 , n25538 );
xnor ( n25540 , n25539 , n22200 );
and ( n25541 , n25536 , n25540 );
and ( n25542 , n23954 , n21880 );
and ( n25543 , n23575 , n21878 );
nor ( n25544 , n25542 , n25543 );
xnor ( n25545 , n25544 , n21890 );
and ( n25546 , n25540 , n25545 );
and ( n25547 , n25536 , n25545 );
or ( n25548 , n25541 , n25546 , n25547 );
and ( n25549 , n25531 , n25548 );
and ( n25550 , n25515 , n25548 );
or ( n25551 , n25532 , n25549 , n25550 );
and ( n25552 , n25506 , n25551 );
xor ( n25553 , n25333 , n25338 );
xor ( n25554 , n25553 , n25349 );
and ( n25555 , n25551 , n25554 );
and ( n25556 , n25506 , n25554 );
or ( n25557 , n25552 , n25555 , n25556 );
and ( n25558 , n25503 , n25557 );
and ( n25559 , n25501 , n25557 );
or ( n25560 , n25504 , n25558 , n25559 );
and ( n25561 , n25498 , n25560 );
and ( n25562 , n25496 , n25560 );
or ( n25563 , n25499 , n25561 , n25562 );
xor ( n25564 , n25324 , n25326 );
xor ( n25565 , n25564 , n25402 );
and ( n25566 , n25563 , n25565 );
and ( n25567 , n21870 , n22305 );
and ( n25568 , n21885 , n22303 );
nor ( n25569 , n25567 , n25568 );
xnor ( n25570 , n25569 , n22315 );
and ( n25571 , n21919 , n21779 );
and ( n25572 , n21932 , n21777 );
nor ( n25573 , n25571 , n25572 );
xnor ( n25574 , n25573 , n21789 );
and ( n25575 , n25570 , n25574 );
xor ( n25576 , n25449 , n25453 );
xor ( n25577 , n25576 , n25458 );
and ( n25578 , n25574 , n25577 );
and ( n25579 , n25570 , n25577 );
or ( n25580 , n25575 , n25578 , n25579 );
xor ( n25581 , n25461 , n25465 );
xor ( n25582 , n25581 , n25470 );
and ( n25583 , n25580 , n25582 );
and ( n25584 , n25565 , n25583 );
and ( n25585 , n25563 , n25583 );
or ( n25586 , n25566 , n25584 , n25585 );
xor ( n25587 , n25413 , n25476 );
xor ( n25588 , n25587 , n25479 );
and ( n25589 , n25586 , n25588 );
xor ( n25590 , n25329 , n25396 );
xor ( n25591 , n25590 , n25399 );
xor ( n25592 , n25352 , n25390 );
xor ( n25593 , n25592 , n25393 );
and ( n25594 , n23284 , n22194 );
and ( n25595 , n23165 , n22192 );
nor ( n25596 , n25594 , n25595 );
xnor ( n25597 , n25596 , n22200 );
and ( n25598 , n23575 , n21880 );
and ( n25599 , n23446 , n21878 );
nor ( n25600 , n25598 , n25599 );
xnor ( n25601 , n25600 , n21890 );
and ( n25602 , n25597 , n25601 );
xor ( n25603 , n25419 , n25429 );
xor ( n25604 , n25603 , n25434 );
and ( n25605 , n25601 , n25604 );
and ( n25606 , n25597 , n25604 );
or ( n25607 , n25602 , n25605 , n25606 );
and ( n25608 , n22049 , n21957 );
and ( n25609 , n22033 , n21955 );
nor ( n25610 , n25608 , n25609 );
xnor ( n25611 , n25610 , n21967 );
and ( n25612 , n25607 , n25611 );
and ( n25613 , n22101 , n21978 );
and ( n25614 , n22086 , n21976 );
nor ( n25615 , n25613 , n25614 );
xnor ( n25616 , n25615 , n21988 );
and ( n25617 , n25611 , n25616 );
and ( n25618 , n25607 , n25616 );
or ( n25619 , n25612 , n25617 , n25618 );
and ( n25620 , n25593 , n25619 );
and ( n25621 , n24896 , n21927 );
and ( n25622 , n24753 , n21925 );
nor ( n25623 , n25621 , n25622 );
xnor ( n25624 , n25623 , n21937 );
and ( n25625 , n25427 , n22062 );
and ( n25626 , n25347 , n22060 );
nor ( n25627 , n25625 , n25626 );
xnor ( n25628 , n25627 , n22068 );
and ( n25629 , n25624 , n25628 );
xor ( n25630 , n21582 , n21658 );
buf ( n552895 , n25630 );
buf ( n552896 , n552895 );
buf ( n25633 , n552896 );
and ( n25634 , n25633 , n22035 );
and ( n25635 , n25628 , n25634 );
and ( n25636 , n25624 , n25634 );
or ( n25637 , n25629 , n25635 , n25636 );
and ( n25638 , n24446 , n21903 );
and ( n25639 , n24011 , n21901 );
nor ( n25640 , n25638 , n25639 );
xnor ( n25641 , n25640 , n21913 );
and ( n25642 , n25637 , n25641 );
and ( n25643 , n25004 , n22022 );
and ( n25644 , n24896 , n22020 );
nor ( n25645 , n25643 , n25644 );
xnor ( n25646 , n25645 , n22028 );
and ( n25647 , n25641 , n25646 );
and ( n25648 , n25637 , n25646 );
or ( n25649 , n25642 , n25647 , n25648 );
and ( n25650 , n22409 , n21804 );
and ( n25651 , n22094 , n21802 );
nor ( n25652 , n25650 , n25651 );
xnor ( n25653 , n25652 , n21814 );
and ( n25654 , n25649 , n25653 );
and ( n25655 , n23074 , n21828 );
and ( n25656 , n22659 , n21826 );
nor ( n25657 , n25655 , n25656 );
xnor ( n25658 , n25657 , n21838 );
and ( n25659 , n25653 , n25658 );
and ( n25660 , n25649 , n25658 );
or ( n25661 , n25654 , n25659 , n25660 );
xor ( n25662 , n25215 , n25219 );
xor ( n25663 , n25662 , n25224 );
and ( n25664 , n25661 , n25663 );
xor ( n25665 , n25437 , n25441 );
xor ( n25666 , n25665 , n25446 );
and ( n25667 , n25663 , n25666 );
and ( n25668 , n25661 , n25666 );
or ( n25669 , n25664 , n25667 , n25668 );
and ( n25670 , n25619 , n25669 );
and ( n25671 , n25593 , n25669 );
or ( n25672 , n25620 , n25670 , n25671 );
and ( n25673 , n25591 , n25672 );
xor ( n25674 , n25496 , n25498 );
xor ( n25675 , n25674 , n25560 );
and ( n25676 , n25672 , n25675 );
and ( n25677 , n25591 , n25675 );
or ( n25678 , n25673 , n25676 , n25677 );
xor ( n25679 , n25415 , n25417 );
xor ( n25680 , n25679 , n25473 );
and ( n25681 , n25678 , n25680 );
xor ( n25682 , n25580 , n25582 );
xor ( n25683 , n25368 , n25384 );
xor ( n25684 , n25683 , n25387 );
and ( n25685 , n24753 , n21927 );
and ( n25686 , n24544 , n21925 );
nor ( n25687 , n25685 , n25686 );
xnor ( n25688 , n25687 , n21937 );
xor ( n25689 , n25423 , n25428 );
and ( n25690 , n25688 , n25689 );
and ( n25691 , n24011 , n21903 );
and ( n25692 , n23954 , n21901 );
nor ( n25693 , n25691 , n25692 );
xnor ( n25694 , n25693 , n21913 );
and ( n25695 , n25690 , n25694 );
and ( n25696 , n24544 , n21927 );
and ( n25697 , n24446 , n21925 );
nor ( n25698 , n25696 , n25697 );
xnor ( n25699 , n25698 , n21937 );
and ( n25700 , n25694 , n25699 );
and ( n25701 , n25690 , n25699 );
or ( n25702 , n25695 , n25700 , n25701 );
and ( n25703 , n25684 , n25702 );
xor ( n25704 , n25356 , n25360 );
xor ( n25705 , n25704 , n25365 );
xor ( n25706 , n25372 , n25376 );
xor ( n25707 , n25706 , n25381 );
and ( n25708 , n25705 , n25707 );
xor ( n25709 , n25510 , n25514 );
and ( n25710 , n22080 , n21957 );
and ( n25711 , n22101 , n21955 );
nor ( n25712 , n25710 , n25711 );
xnor ( n25713 , n25712 , n21967 );
and ( n25714 , n23284 , n21828 );
and ( n25715 , n23165 , n21826 );
nor ( n25716 , n25714 , n25715 );
xnor ( n25717 , n25716 , n21838 );
and ( n25718 , n25713 , n25717 );
and ( n25719 , n23575 , n22194 );
and ( n25720 , n23446 , n22192 );
nor ( n25721 , n25719 , n25720 );
xnor ( n25722 , n25721 , n22200 );
and ( n25723 , n25717 , n25722 );
and ( n25724 , n25713 , n25722 );
or ( n25725 , n25718 , n25723 , n25724 );
and ( n25726 , n25709 , n25725 );
xor ( n25727 , n25519 , n25523 );
xor ( n25728 , n25727 , n25528 );
and ( n25729 , n25725 , n25728 );
and ( n25730 , n25709 , n25728 );
or ( n25731 , n25726 , n25729 , n25730 );
and ( n25732 , n25707 , n25731 );
and ( n25733 , n25705 , n25731 );
or ( n25734 , n25708 , n25732 , n25733 );
and ( n25735 , n25702 , n25734 );
and ( n25736 , n25684 , n25734 );
or ( n25737 , n25703 , n25735 , n25736 );
xor ( n25738 , n25501 , n25503 );
xor ( n25739 , n25738 , n25557 );
and ( n25740 , n25737 , n25739 );
and ( n25741 , n25347 , n22022 );
and ( n25742 , n25337 , n22020 );
nor ( n25743 , n25741 , n25742 );
xnor ( n25744 , n25743 , n22028 );
and ( n25745 , n25633 , n22062 );
and ( n25746 , n25427 , n22060 );
nor ( n25747 , n25745 , n25746 );
xnor ( n25748 , n25747 , n22068 );
and ( n25749 , n25744 , n25748 );
xor ( n25750 , n21599 , n21656 );
buf ( n553015 , n25750 );
buf ( n553016 , n553015 );
buf ( n25753 , n553016 );
and ( n25754 , n25753 , n22035 );
and ( n25755 , n25748 , n25754 );
and ( n25756 , n25744 , n25754 );
or ( n25757 , n25749 , n25755 , n25756 );
and ( n25758 , n24544 , n21903 );
and ( n25759 , n24446 , n21901 );
nor ( n25760 , n25758 , n25759 );
xnor ( n25761 , n25760 , n21913 );
and ( n25762 , n25757 , n25761 );
and ( n25763 , n25337 , n22022 );
and ( n25764 , n25004 , n22020 );
nor ( n25765 , n25763 , n25764 );
xnor ( n25766 , n25765 , n22028 );
and ( n25767 , n25761 , n25766 );
and ( n25768 , n25757 , n25766 );
or ( n25769 , n25762 , n25767 , n25768 );
and ( n25770 , n22659 , n21804 );
and ( n25771 , n22409 , n21802 );
nor ( n25772 , n25770 , n25771 );
xnor ( n25773 , n25772 , n21814 );
and ( n25774 , n25769 , n25773 );
and ( n25775 , n23165 , n21828 );
and ( n25776 , n23074 , n21826 );
nor ( n25777 , n25775 , n25776 );
xnor ( n25778 , n25777 , n21838 );
and ( n25779 , n25773 , n25778 );
and ( n25780 , n25769 , n25778 );
or ( n25781 , n25774 , n25779 , n25780 );
and ( n25782 , n22086 , n21957 );
and ( n25783 , n22049 , n21955 );
nor ( n25784 , n25782 , n25783 );
xnor ( n25785 , n25784 , n21967 );
and ( n25786 , n25781 , n25785 );
xor ( n25787 , n25597 , n25601 );
xor ( n25788 , n25787 , n25604 );
and ( n25789 , n25785 , n25788 );
and ( n25790 , n25781 , n25788 );
or ( n25791 , n25786 , n25789 , n25790 );
and ( n25792 , n21908 , n22305 );
and ( n25793 , n21870 , n22303 );
nor ( n25794 , n25792 , n25793 );
xnor ( n25795 , n25794 , n22315 );
and ( n25796 , n25791 , n25795 );
xor ( n25797 , n25607 , n25611 );
xor ( n25798 , n25797 , n25616 );
and ( n25799 , n25795 , n25798 );
and ( n25800 , n25791 , n25798 );
or ( n25801 , n25796 , n25799 , n25800 );
and ( n25802 , n25739 , n25801 );
and ( n25803 , n25737 , n25801 );
or ( n25804 , n25740 , n25802 , n25803 );
and ( n25805 , n25682 , n25804 );
xor ( n25806 , n25591 , n25672 );
xor ( n25807 , n25806 , n25675 );
and ( n25808 , n25804 , n25807 );
and ( n25809 , n25682 , n25807 );
or ( n25810 , n25805 , n25808 , n25809 );
and ( n25811 , n25680 , n25810 );
and ( n25812 , n25678 , n25810 );
or ( n25813 , n25681 , n25811 , n25812 );
and ( n25814 , n25588 , n25813 );
and ( n25815 , n25586 , n25813 );
or ( n25816 , n25589 , n25814 , n25815 );
and ( n25817 , n25494 , n25816 );
xor ( n25818 , n25494 , n25816 );
xor ( n25819 , n25563 , n25565 );
xor ( n25820 , n25819 , n25583 );
and ( n25821 , n25427 , n22022 );
and ( n25822 , n25347 , n22020 );
nor ( n25823 , n25821 , n25822 );
xnor ( n25824 , n25823 , n22028 );
and ( n25825 , n25753 , n22062 );
and ( n25826 , n25633 , n22060 );
nor ( n25827 , n25825 , n25826 );
xnor ( n25828 , n25827 , n22068 );
and ( n25829 , n25824 , n25828 );
xor ( n25830 , n21615 , n21654 );
buf ( n553095 , n25830 );
buf ( n553096 , n553095 );
buf ( n25833 , n553096 );
and ( n25834 , n25833 , n22035 );
and ( n25835 , n25828 , n25834 );
and ( n25836 , n25824 , n25834 );
or ( n25837 , n25829 , n25835 , n25836 );
and ( n25838 , n24753 , n21903 );
and ( n25839 , n24544 , n21901 );
nor ( n25840 , n25838 , n25839 );
xnor ( n25841 , n25840 , n21913 );
and ( n25842 , n25837 , n25841 );
and ( n25843 , n25004 , n21927 );
and ( n25844 , n24896 , n21925 );
nor ( n25845 , n25843 , n25844 );
xnor ( n25846 , n25845 , n21937 );
and ( n25847 , n25841 , n25846 );
and ( n25848 , n25837 , n25846 );
or ( n25849 , n25842 , n25847 , n25848 );
and ( n25850 , n24011 , n21880 );
and ( n25851 , n23954 , n21878 );
nor ( n25852 , n25850 , n25851 );
xnor ( n25853 , n25852 , n21890 );
and ( n25854 , n25849 , n25853 );
xor ( n25855 , n25624 , n25628 );
xor ( n25856 , n25855 , n25634 );
and ( n25857 , n25853 , n25856 );
and ( n25858 , n25849 , n25856 );
or ( n25859 , n25854 , n25857 , n25858 );
and ( n25860 , n22094 , n21978 );
and ( n25861 , n22080 , n21976 );
nor ( n25862 , n25860 , n25861 );
xnor ( n25863 , n25862 , n21988 );
and ( n25864 , n25859 , n25863 );
xor ( n25865 , n25637 , n25641 );
xor ( n25866 , n25865 , n25646 );
and ( n25867 , n25863 , n25866 );
and ( n25868 , n25859 , n25866 );
or ( n25869 , n25864 , n25867 , n25868 );
and ( n25870 , n22041 , n21779 );
and ( n25871 , n22014 , n21777 );
nor ( n25872 , n25870 , n25871 );
xnor ( n25873 , n25872 , n21789 );
and ( n25874 , n25869 , n25873 );
xor ( n25875 , n25649 , n25653 );
xor ( n25876 , n25875 , n25658 );
and ( n25877 , n25873 , n25876 );
and ( n25878 , n25869 , n25876 );
or ( n25879 , n25874 , n25877 , n25878 );
and ( n25880 , n21820 , n21735 );
and ( n25881 , n21833 , n21732 );
nor ( n25882 , n25880 , n25881 );
xnor ( n25883 , n25882 , n21730 );
and ( n25884 , n25879 , n25883 );
xor ( n25885 , n25661 , n25663 );
xor ( n25886 , n25885 , n25666 );
and ( n25887 , n25883 , n25886 );
and ( n25888 , n25879 , n25886 );
or ( n25889 , n25884 , n25887 , n25888 );
xor ( n25890 , n25570 , n25574 );
xor ( n25891 , n25890 , n25577 );
and ( n25892 , n25889 , n25891 );
xor ( n25893 , n25506 , n25551 );
xor ( n25894 , n25893 , n25554 );
xor ( n25895 , n25515 , n25531 );
xor ( n25896 , n25895 , n25548 );
xor ( n25897 , n25690 , n25694 );
xor ( n25898 , n25897 , n25699 );
and ( n25899 , n25896 , n25898 );
xor ( n25900 , n25536 , n25540 );
xor ( n25901 , n25900 , n25545 );
xor ( n25902 , n25688 , n25689 );
and ( n25903 , n25901 , n25902 );
xor ( n25904 , n25709 , n25725 );
xor ( n25905 , n25904 , n25728 );
and ( n25906 , n25902 , n25905 );
and ( n25907 , n25901 , n25905 );
or ( n25908 , n25903 , n25906 , n25907 );
and ( n25909 , n25898 , n25908 );
and ( n25910 , n25896 , n25908 );
or ( n25911 , n25899 , n25909 , n25910 );
and ( n25912 , n25894 , n25911 );
xor ( n25913 , n25684 , n25702 );
xor ( n25914 , n25913 , n25734 );
and ( n25915 , n25911 , n25914 );
and ( n25916 , n25894 , n25914 );
or ( n25917 , n25912 , n25915 , n25916 );
xor ( n25918 , n25593 , n25619 );
xor ( n25919 , n25918 , n25669 );
and ( n25920 , n25917 , n25919 );
xor ( n25921 , n25737 , n25739 );
xor ( n25922 , n25921 , n25801 );
and ( n25923 , n25919 , n25922 );
and ( n25924 , n25917 , n25922 );
or ( n25925 , n25920 , n25923 , n25924 );
and ( n25926 , n25892 , n25925 );
xor ( n25927 , n25682 , n25804 );
xor ( n25928 , n25927 , n25807 );
and ( n25929 , n25925 , n25928 );
and ( n25930 , n25892 , n25928 );
or ( n25931 , n25926 , n25929 , n25930 );
and ( n25932 , n25820 , n25931 );
xor ( n25933 , n25678 , n25680 );
xor ( n25934 , n25933 , n25810 );
and ( n25935 , n25931 , n25934 );
and ( n25936 , n25820 , n25934 );
or ( n25937 , n25932 , n25935 , n25936 );
xor ( n25938 , n25586 , n25588 );
xor ( n25939 , n25938 , n25813 );
and ( n25940 , n25937 , n25939 );
xor ( n25941 , n25937 , n25939 );
xor ( n25942 , n25820 , n25931 );
xor ( n25943 , n25942 , n25934 );
xor ( n25944 , n25889 , n25891 );
xor ( n25945 , n25791 , n25795 );
xor ( n25946 , n25945 , n25798 );
xor ( n25947 , n25894 , n25911 );
xor ( n25948 , n25947 , n25914 );
and ( n25949 , n25946 , n25948 );
xor ( n25950 , n25879 , n25883 );
xor ( n25951 , n25950 , n25886 );
and ( n25952 , n25948 , n25951 );
and ( n25953 , n25946 , n25951 );
or ( n25954 , n25949 , n25952 , n25953 );
and ( n25955 , n25944 , n25954 );
xor ( n25956 , n25917 , n25919 );
xor ( n25957 , n25956 , n25922 );
and ( n25958 , n25954 , n25957 );
and ( n25959 , n25944 , n25957 );
or ( n25960 , n25955 , n25958 , n25959 );
xor ( n25961 , n25892 , n25925 );
xor ( n25962 , n25961 , n25928 );
and ( n25963 , n25960 , n25962 );
xor ( n25964 , n25869 , n25873 );
xor ( n25965 , n25964 , n25876 );
xor ( n25966 , n25781 , n25785 );
xor ( n25967 , n25966 , n25788 );
and ( n25968 , n25965 , n25967 );
xor ( n25969 , n25705 , n25707 );
xor ( n25970 , n25969 , n25731 );
xor ( n25971 , n25896 , n25898 );
xor ( n25972 , n25971 , n25908 );
and ( n25973 , n25970 , n25972 );
and ( n25974 , n25633 , n22022 );
and ( n25975 , n25427 , n22020 );
nor ( n25976 , n25974 , n25975 );
xnor ( n25977 , n25976 , n22028 );
and ( n25978 , n25833 , n22062 );
and ( n25979 , n25753 , n22060 );
nor ( n25980 , n25978 , n25979 );
xnor ( n25981 , n25980 , n22068 );
and ( n25982 , n25977 , n25981 );
xor ( n25983 , n21627 , n21652 );
buf ( n553248 , n25983 );
buf ( n553249 , n553248 );
buf ( n25986 , n553249 );
and ( n25987 , n25986 , n22035 );
and ( n25988 , n25981 , n25987 );
and ( n25989 , n25977 , n25987 );
or ( n25990 , n25982 , n25988 , n25989 );
and ( n25991 , n24896 , n21903 );
and ( n25992 , n24753 , n21901 );
nor ( n25993 , n25991 , n25992 );
xnor ( n25994 , n25993 , n21913 );
and ( n25995 , n25990 , n25994 );
and ( n25996 , n25337 , n21927 );
and ( n25997 , n25004 , n21925 );
nor ( n25998 , n25996 , n25997 );
xnor ( n25999 , n25998 , n21937 );
and ( n26000 , n25994 , n25999 );
and ( n26001 , n25990 , n25999 );
or ( n26002 , n25995 , n26000 , n26001 );
and ( n26003 , n24446 , n21880 );
and ( n26004 , n24011 , n21878 );
nor ( n26005 , n26003 , n26004 );
xnor ( n26006 , n26005 , n21890 );
and ( n26007 , n26002 , n26006 );
xor ( n26008 , n25744 , n25748 );
xor ( n26009 , n26008 , n25754 );
and ( n26010 , n26006 , n26009 );
and ( n26011 , n26002 , n26009 );
or ( n26012 , n26007 , n26010 , n26011 );
and ( n26013 , n22409 , n21978 );
and ( n26014 , n22094 , n21976 );
nor ( n26015 , n26013 , n26014 );
xnor ( n26016 , n26015 , n21988 );
and ( n26017 , n26012 , n26016 );
and ( n26018 , n23074 , n21804 );
and ( n26019 , n22659 , n21802 );
nor ( n26020 , n26018 , n26019 );
xnor ( n26021 , n26020 , n21814 );
and ( n26022 , n26016 , n26021 );
and ( n26023 , n26012 , n26021 );
or ( n26024 , n26017 , n26022 , n26023 );
and ( n26025 , n22014 , n21854 );
and ( n26026 , n21919 , n21852 );
nor ( n26027 , n26025 , n26026 );
xnor ( n26028 , n26027 , n21864 );
and ( n26029 , n26024 , n26028 );
xor ( n26030 , n25859 , n25863 );
xor ( n26031 , n26030 , n25866 );
and ( n26032 , n26028 , n26031 );
and ( n26033 , n26024 , n26031 );
or ( n26034 , n26029 , n26032 , n26033 );
and ( n26035 , n25972 , n26034 );
and ( n26036 , n25970 , n26034 );
or ( n26037 , n25973 , n26035 , n26036 );
and ( n26038 , n25968 , n26037 );
xor ( n26039 , n25769 , n25773 );
xor ( n26040 , n26039 , n25778 );
xor ( n26041 , n25901 , n25902 );
xor ( n26042 , n26041 , n25905 );
and ( n26043 , n26040 , n26042 );
and ( n26044 , n23165 , n21804 );
and ( n26045 , n23074 , n21802 );
nor ( n26046 , n26044 , n26045 );
xnor ( n26047 , n26046 , n21814 );
and ( n26048 , n23954 , n22194 );
and ( n26049 , n23575 , n22192 );
nor ( n26050 , n26048 , n26049 );
xnor ( n26051 , n26050 , n22200 );
and ( n26052 , n26047 , n26051 );
xor ( n26053 , n25837 , n25841 );
xor ( n26054 , n26053 , n25846 );
and ( n26055 , n26051 , n26054 );
and ( n26056 , n26047 , n26054 );
or ( n26057 , n26052 , n26055 , n26056 );
and ( n26058 , n22086 , n22323 );
and ( n26059 , n22049 , n22321 );
nor ( n26060 , n26058 , n26059 );
xnor ( n26061 , n26060 , n22329 );
and ( n26062 , n26057 , n26061 );
xor ( n26063 , n25849 , n25853 );
xor ( n26064 , n26063 , n25856 );
and ( n26065 , n26061 , n26064 );
and ( n26066 , n26057 , n26064 );
or ( n26067 , n26062 , n26065 , n26066 );
and ( n26068 , n26042 , n26067 );
and ( n26069 , n26040 , n26067 );
or ( n26070 , n26043 , n26068 , n26069 );
xor ( n26071 , n25965 , n25967 );
and ( n26072 , n26070 , n26071 );
xor ( n26073 , n26024 , n26028 );
xor ( n26074 , n26073 , n26031 );
and ( n26075 , n21870 , n21735 );
and ( n26076 , n21885 , n21732 );
nor ( n26077 , n26075 , n26076 );
xnor ( n26078 , n26077 , n21730 );
and ( n26079 , n21919 , n22305 );
and ( n26080 , n21932 , n22303 );
nor ( n26081 , n26079 , n26080 );
xnor ( n26082 , n26081 , n22315 );
and ( n26083 , n26078 , n26082 );
xor ( n26084 , n26057 , n26061 );
xor ( n26085 , n26084 , n26064 );
and ( n26086 , n26082 , n26085 );
and ( n26087 , n26078 , n26085 );
or ( n26088 , n26083 , n26086 , n26087 );
and ( n26089 , n26074 , n26088 );
xor ( n26090 , n25713 , n25717 );
xor ( n26091 , n26090 , n25722 );
xor ( n26092 , n25757 , n25761 );
xor ( n26093 , n26092 , n25766 );
and ( n26094 , n26091 , n26093 );
and ( n26095 , n25753 , n22022 );
and ( n26096 , n25633 , n22020 );
nor ( n26097 , n26095 , n26096 );
xnor ( n26098 , n26097 , n22028 );
and ( n26099 , n25986 , n22062 );
and ( n26100 , n25833 , n22060 );
nor ( n26101 , n26099 , n26100 );
xnor ( n26102 , n26101 , n22068 );
and ( n26103 , n26098 , n26102 );
xor ( n26104 , n21634 , n21650 );
buf ( n553369 , n26104 );
buf ( n553370 , n553369 );
buf ( n26107 , n553370 );
and ( n26108 , n26107 , n22035 );
and ( n26109 , n26102 , n26108 );
and ( n26110 , n26098 , n26108 );
or ( n26111 , n26103 , n26109 , n26110 );
and ( n26112 , n25347 , n21927 );
and ( n26113 , n25337 , n21925 );
nor ( n26114 , n26112 , n26113 );
xnor ( n26115 , n26114 , n21937 );
and ( n26116 , n26111 , n26115 );
xor ( n26117 , n25977 , n25981 );
xor ( n26118 , n26117 , n25987 );
and ( n26119 , n26115 , n26118 );
and ( n26120 , n26111 , n26118 );
or ( n26121 , n26116 , n26119 , n26120 );
and ( n26122 , n24544 , n21880 );
and ( n26123 , n24446 , n21878 );
nor ( n26124 , n26122 , n26123 );
xnor ( n26125 , n26124 , n21890 );
and ( n26126 , n26121 , n26125 );
xor ( n26127 , n25824 , n25828 );
xor ( n26128 , n26127 , n25834 );
and ( n26129 , n26125 , n26128 );
and ( n26130 , n26121 , n26128 );
or ( n26131 , n26126 , n26129 , n26130 );
and ( n26132 , n22659 , n21978 );
and ( n26133 , n22409 , n21976 );
nor ( n26134 , n26132 , n26133 );
xnor ( n26135 , n26134 , n21988 );
and ( n26136 , n26131 , n26135 );
and ( n26137 , n23446 , n21828 );
and ( n26138 , n23284 , n21826 );
nor ( n26139 , n26137 , n26138 );
xnor ( n26140 , n26139 , n21838 );
and ( n26141 , n26135 , n26140 );
and ( n26142 , n26131 , n26140 );
or ( n26143 , n26136 , n26141 , n26142 );
and ( n26144 , n26093 , n26143 );
and ( n26145 , n26091 , n26143 );
or ( n26146 , n26094 , n26144 , n26145 );
and ( n26147 , n26088 , n26146 );
and ( n26148 , n26074 , n26146 );
or ( n26149 , n26089 , n26147 , n26148 );
and ( n26150 , n26071 , n26149 );
and ( n26151 , n26070 , n26149 );
or ( n26152 , n26072 , n26150 , n26151 );
and ( n26153 , n26037 , n26152 );
and ( n26154 , n25968 , n26152 );
or ( n26155 , n26038 , n26153 , n26154 );
xor ( n26156 , n25944 , n25954 );
xor ( n26157 , n26156 , n25957 );
and ( n26158 , n26155 , n26157 );
xor ( n26159 , n25946 , n25948 );
xor ( n26160 , n26159 , n25951 );
xor ( n26161 , n25970 , n25972 );
xor ( n26162 , n26161 , n26034 );
xor ( n26163 , n26040 , n26042 );
xor ( n26164 , n26163 , n26067 );
and ( n26165 , n23284 , n21804 );
and ( n26166 , n23165 , n21802 );
nor ( n26167 , n26165 , n26166 );
xnor ( n26168 , n26167 , n21814 );
and ( n26169 , n23575 , n21828 );
and ( n26170 , n23446 , n21826 );
nor ( n26171 , n26169 , n26170 );
xnor ( n26172 , n26171 , n21838 );
and ( n26173 , n26168 , n26172 );
xor ( n26174 , n26121 , n26125 );
xor ( n26175 , n26174 , n26128 );
and ( n26176 , n26172 , n26175 );
and ( n26177 , n26168 , n26175 );
or ( n26178 , n26173 , n26176 , n26177 );
and ( n26179 , n22049 , n21779 );
and ( n26180 , n22033 , n21777 );
nor ( n26181 , n26179 , n26180 );
xnor ( n26182 , n26181 , n21789 );
and ( n26183 , n26178 , n26182 );
xor ( n26184 , n26047 , n26051 );
xor ( n26185 , n26184 , n26054 );
and ( n26186 , n26182 , n26185 );
and ( n26187 , n26178 , n26185 );
or ( n26188 , n26183 , n26186 , n26187 );
and ( n26189 , n21895 , n22252 );
and ( n26190 , n21908 , n22250 );
nor ( n26191 , n26189 , n26190 );
xnor ( n26192 , n26191 , n22258 );
and ( n26193 , n26188 , n26192 );
and ( n26194 , n22041 , n21854 );
and ( n26195 , n22014 , n21852 );
nor ( n26196 , n26194 , n26195 );
xnor ( n26197 , n26196 , n21864 );
and ( n26198 , n26192 , n26197 );
and ( n26199 , n26188 , n26197 );
or ( n26200 , n26193 , n26198 , n26199 );
and ( n26201 , n26164 , n26200 );
and ( n26202 , n25833 , n22022 );
and ( n26203 , n25753 , n22020 );
nor ( n26204 , n26202 , n26203 );
xnor ( n26205 , n26204 , n22028 );
and ( n26206 , n26107 , n22062 );
and ( n26207 , n25986 , n22060 );
nor ( n26208 , n26206 , n26207 );
xnor ( n26209 , n26208 , n22068 );
and ( n26210 , n26205 , n26209 );
xor ( n26211 , n21640 , n21648 );
buf ( n553476 , n26211 );
buf ( n553477 , n553476 );
buf ( n26214 , n553477 );
and ( n26215 , n26214 , n22035 );
and ( n26216 , n26209 , n26215 );
and ( n26217 , n26205 , n26215 );
or ( n26218 , n26210 , n26216 , n26217 );
and ( n26219 , n25427 , n21927 );
and ( n26220 , n25347 , n21925 );
nor ( n26221 , n26219 , n26220 );
xnor ( n26222 , n26221 , n21937 );
and ( n26223 , n26218 , n26222 );
xor ( n26224 , n26098 , n26102 );
xor ( n26225 , n26224 , n26108 );
and ( n26226 , n26222 , n26225 );
and ( n26227 , n26218 , n26225 );
or ( n26228 , n26223 , n26226 , n26227 );
and ( n26229 , n24753 , n21880 );
and ( n26230 , n24544 , n21878 );
nor ( n26231 , n26229 , n26230 );
xnor ( n26232 , n26231 , n21890 );
and ( n26233 , n26228 , n26232 );
and ( n26234 , n25004 , n21903 );
and ( n26235 , n24896 , n21901 );
nor ( n26236 , n26234 , n26235 );
xnor ( n26237 , n26236 , n21913 );
and ( n26238 , n26232 , n26237 );
and ( n26239 , n26228 , n26237 );
or ( n26240 , n26233 , n26238 , n26239 );
and ( n26241 , n24011 , n22194 );
and ( n26242 , n23954 , n22192 );
nor ( n26243 , n26241 , n26242 );
xnor ( n26244 , n26243 , n22200 );
and ( n26245 , n26240 , n26244 );
xor ( n26246 , n25990 , n25994 );
xor ( n26247 , n26246 , n25999 );
and ( n26248 , n26244 , n26247 );
and ( n26249 , n26240 , n26247 );
or ( n26250 , n26245 , n26248 , n26249 );
and ( n26251 , n22094 , n21957 );
and ( n26252 , n22080 , n21955 );
nor ( n26253 , n26251 , n26252 );
xnor ( n26254 , n26253 , n21967 );
and ( n26255 , n26250 , n26254 );
xor ( n26256 , n26002 , n26006 );
xor ( n26257 , n26256 , n26009 );
and ( n26258 , n26254 , n26257 );
and ( n26259 , n26250 , n26257 );
or ( n26260 , n26255 , n26258 , n26259 );
and ( n26261 , n22033 , n21779 );
and ( n26262 , n22056 , n21777 );
nor ( n26263 , n26261 , n26262 );
xnor ( n26264 , n26263 , n21789 );
and ( n26265 , n26260 , n26264 );
xor ( n26266 , n26012 , n26016 );
xor ( n26267 , n26266 , n26021 );
and ( n26268 , n26264 , n26267 );
and ( n26269 , n26260 , n26267 );
or ( n26270 , n26265 , n26268 , n26269 );
and ( n26271 , n26200 , n26270 );
and ( n26272 , n26164 , n26270 );
or ( n26273 , n26201 , n26271 , n26272 );
and ( n26274 , n26162 , n26273 );
xor ( n26275 , n26070 , n26071 );
xor ( n26276 , n26275 , n26149 );
and ( n26277 , n26273 , n26276 );
and ( n26278 , n26162 , n26276 );
or ( n26279 , n26274 , n26277 , n26278 );
and ( n26280 , n26160 , n26279 );
xor ( n26281 , n25968 , n26037 );
xor ( n26282 , n26281 , n26152 );
and ( n26283 , n26279 , n26282 );
and ( n26284 , n26160 , n26282 );
or ( n26285 , n26280 , n26283 , n26284 );
and ( n26286 , n26157 , n26285 );
and ( n26287 , n26155 , n26285 );
or ( n26288 , n26158 , n26286 , n26287 );
and ( n26289 , n25962 , n26288 );
and ( n26290 , n25960 , n26288 );
or ( n26291 , n25963 , n26289 , n26290 );
and ( n26292 , n25943 , n26291 );
xor ( n26293 , n25943 , n26291 );
xor ( n26294 , n25960 , n25962 );
xor ( n26295 , n26294 , n26288 );
xor ( n26296 , n26155 , n26157 );
xor ( n26297 , n26296 , n26285 );
xor ( n26298 , n26160 , n26279 );
xor ( n26299 , n26298 , n26282 );
xor ( n26300 , n26078 , n26082 );
xor ( n26301 , n26300 , n26085 );
and ( n26302 , n23954 , n21828 );
and ( n26303 , n23575 , n21826 );
nor ( n26304 , n26302 , n26303 );
xnor ( n26305 , n26304 , n21838 );
and ( n26306 , n24446 , n22194 );
and ( n26307 , n24011 , n22192 );
nor ( n26308 , n26306 , n26307 );
xnor ( n26309 , n26308 , n22200 );
and ( n26310 , n26305 , n26309 );
xor ( n26311 , n26111 , n26115 );
xor ( n26312 , n26311 , n26118 );
and ( n26313 , n26309 , n26312 );
and ( n26314 , n26305 , n26312 );
or ( n26315 , n26310 , n26313 , n26314 );
and ( n26316 , n22409 , n21957 );
and ( n26317 , n22094 , n21955 );
nor ( n26318 , n26316 , n26317 );
xnor ( n26319 , n26318 , n21967 );
and ( n26320 , n26315 , n26319 );
and ( n26321 , n23074 , n21978 );
and ( n26322 , n22659 , n21976 );
nor ( n26323 , n26321 , n26322 );
xnor ( n26324 , n26323 , n21988 );
and ( n26325 , n26319 , n26324 );
and ( n26326 , n26315 , n26324 );
or ( n26327 , n26320 , n26325 , n26326 );
and ( n26328 , n22101 , n22323 );
and ( n26329 , n22086 , n22321 );
nor ( n26330 , n26328 , n26329 );
xnor ( n26331 , n26330 , n22329 );
and ( n26332 , n26327 , n26331 );
xor ( n26333 , n26131 , n26135 );
xor ( n26334 , n26333 , n26140 );
and ( n26335 , n26331 , n26334 );
and ( n26336 , n26327 , n26334 );
or ( n26337 , n26332 , n26335 , n26336 );
and ( n26338 , n26301 , n26337 );
xor ( n26339 , n26091 , n26093 );
xor ( n26340 , n26339 , n26143 );
and ( n26341 , n26337 , n26340 );
and ( n26342 , n26301 , n26340 );
or ( n26343 , n26338 , n26341 , n26342 );
xor ( n26344 , n26074 , n26088 );
xor ( n26345 , n26344 , n26146 );
and ( n26346 , n26343 , n26345 );
xor ( n26347 , n26164 , n26200 );
xor ( n26348 , n26347 , n26270 );
and ( n26349 , n26345 , n26348 );
and ( n26350 , n26343 , n26348 );
or ( n26351 , n26346 , n26349 , n26350 );
xor ( n26352 , n26162 , n26273 );
xor ( n26353 , n26352 , n26276 );
and ( n26354 , n26351 , n26353 );
xor ( n26355 , n26343 , n26345 );
xor ( n26356 , n26355 , n26348 );
buf ( n26357 , n21645 );
buf ( n553622 , n26357 );
buf ( n553623 , n553622 );
buf ( n26360 , n553623 );
and ( n26361 , n26360 , n22060 );
not ( n26362 , n26361 );
and ( n26363 , n26362 , n22068 );
and ( n26364 , n26360 , n22062 );
xor ( n26365 , n21644 , n21647 );
buf ( n553630 , n26365 );
buf ( n553631 , n553630 );
buf ( n26368 , n553631 );
and ( n26369 , n26368 , n22060 );
nor ( n26370 , n26364 , n26369 );
xnor ( n26371 , n26370 , n22068 );
and ( n26372 , n26363 , n26371 );
and ( n26373 , n26368 , n22062 );
and ( n26374 , n26214 , n22060 );
nor ( n26375 , n26373 , n26374 );
xnor ( n26376 , n26375 , n22068 );
and ( n26377 , n26372 , n26376 );
and ( n26378 , n26360 , n22035 );
and ( n26379 , n26376 , n26378 );
and ( n26380 , n26372 , n26378 );
or ( n26381 , n26377 , n26379 , n26380 );
and ( n26382 , n26214 , n22062 );
and ( n26383 , n26107 , n22060 );
nor ( n26384 , n26382 , n26383 );
xnor ( n26385 , n26384 , n22068 );
and ( n26386 , n26381 , n26385 );
and ( n26387 , n26368 , n22035 );
and ( n26388 , n26385 , n26387 );
and ( n26389 , n26381 , n26387 );
or ( n26390 , n26386 , n26388 , n26389 );
and ( n26391 , n25633 , n21927 );
and ( n26392 , n25427 , n21925 );
nor ( n26393 , n26391 , n26392 );
xnor ( n26394 , n26393 , n21937 );
and ( n26395 , n26390 , n26394 );
xor ( n26396 , n26205 , n26209 );
xor ( n26397 , n26396 , n26215 );
and ( n26398 , n26394 , n26397 );
and ( n26399 , n26390 , n26397 );
or ( n26400 , n26395 , n26398 , n26399 );
and ( n26401 , n24896 , n21880 );
and ( n26402 , n24753 , n21878 );
nor ( n26403 , n26401 , n26402 );
xnor ( n26404 , n26403 , n21890 );
and ( n26405 , n26400 , n26404 );
and ( n26406 , n25337 , n21903 );
and ( n26407 , n25004 , n21901 );
nor ( n26408 , n26406 , n26407 );
xnor ( n26409 , n26408 , n21913 );
and ( n26410 , n26404 , n26409 );
and ( n26411 , n26400 , n26409 );
or ( n26412 , n26405 , n26410 , n26411 );
and ( n26413 , n23165 , n21978 );
and ( n26414 , n23074 , n21976 );
nor ( n26415 , n26413 , n26414 );
xnor ( n26416 , n26415 , n21988 );
and ( n26417 , n26412 , n26416 );
xor ( n26418 , n26228 , n26232 );
xor ( n26419 , n26418 , n26237 );
and ( n26420 , n26416 , n26419 );
and ( n26421 , n26412 , n26419 );
or ( n26422 , n26417 , n26420 , n26421 );
and ( n26423 , n22086 , n21779 );
and ( n26424 , n22049 , n21777 );
nor ( n26425 , n26423 , n26424 );
xnor ( n26426 , n26425 , n21789 );
and ( n26427 , n26422 , n26426 );
xor ( n26428 , n26240 , n26244 );
xor ( n26429 , n26428 , n26247 );
and ( n26430 , n26426 , n26429 );
and ( n26431 , n26422 , n26429 );
or ( n26432 , n26427 , n26430 , n26431 );
and ( n26433 , n22014 , n22305 );
and ( n26434 , n21919 , n22303 );
nor ( n26435 , n26433 , n26434 );
xnor ( n26436 , n26435 , n22315 );
and ( n26437 , n26432 , n26436 );
and ( n26438 , n22056 , n21854 );
and ( n26439 , n22041 , n21852 );
nor ( n26440 , n26438 , n26439 );
xnor ( n26441 , n26440 , n21864 );
and ( n26442 , n26436 , n26441 );
and ( n26443 , n26432 , n26441 );
or ( n26444 , n26437 , n26442 , n26443 );
and ( n26445 , n21932 , n22252 );
and ( n26446 , n21895 , n22250 );
nor ( n26447 , n26445 , n26446 );
xnor ( n26448 , n26447 , n22258 );
xor ( n26449 , n26250 , n26254 );
xor ( n26450 , n26449 , n26257 );
and ( n26451 , n26448 , n26450 );
xor ( n26452 , n26178 , n26182 );
xor ( n26453 , n26452 , n26185 );
and ( n26454 , n26450 , n26453 );
and ( n26455 , n26448 , n26453 );
or ( n26456 , n26451 , n26454 , n26455 );
and ( n26457 , n26444 , n26456 );
xor ( n26458 , n26188 , n26192 );
xor ( n26459 , n26458 , n26197 );
and ( n26460 , n26456 , n26459 );
and ( n26461 , n26444 , n26459 );
or ( n26462 , n26457 , n26460 , n26461 );
and ( n26463 , n26356 , n26462 );
xor ( n26464 , n26260 , n26264 );
xor ( n26465 , n26464 , n26267 );
xor ( n26466 , n26301 , n26337 );
xor ( n26467 , n26466 , n26340 );
and ( n26468 , n26465 , n26467 );
and ( n26469 , n22041 , n22305 );
and ( n26470 , n22014 , n22303 );
nor ( n26471 , n26469 , n26470 );
xnor ( n26472 , n26471 , n22315 );
and ( n26473 , n22033 , n21854 );
and ( n26474 , n22056 , n21852 );
nor ( n26475 , n26473 , n26474 );
xnor ( n26476 , n26475 , n21864 );
and ( n26477 , n26472 , n26476 );
xor ( n26478 , n26315 , n26319 );
xor ( n26479 , n26478 , n26324 );
and ( n26480 , n26476 , n26479 );
and ( n26481 , n26472 , n26479 );
or ( n26482 , n26477 , n26480 , n26481 );
and ( n26483 , n25753 , n21927 );
and ( n26484 , n25633 , n21925 );
nor ( n26485 , n26483 , n26484 );
xnor ( n26486 , n26485 , n21937 );
and ( n26487 , n25986 , n22022 );
and ( n26488 , n25833 , n22020 );
nor ( n26489 , n26487 , n26488 );
xnor ( n26490 , n26489 , n22028 );
and ( n26491 , n26486 , n26490 );
xor ( n26492 , n26381 , n26385 );
xor ( n26493 , n26492 , n26387 );
and ( n26494 , n26490 , n26493 );
and ( n26495 , n26486 , n26493 );
or ( n26496 , n26491 , n26494 , n26495 );
and ( n26497 , n25347 , n21903 );
and ( n26498 , n25337 , n21901 );
nor ( n26499 , n26497 , n26498 );
xnor ( n26500 , n26499 , n21913 );
and ( n26501 , n26496 , n26500 );
xor ( n26502 , n26390 , n26394 );
xor ( n26503 , n26502 , n26397 );
and ( n26504 , n26500 , n26503 );
and ( n26505 , n26496 , n26503 );
or ( n26506 , n26501 , n26504 , n26505 );
and ( n26507 , n24544 , n22194 );
and ( n26508 , n24446 , n22192 );
nor ( n26509 , n26507 , n26508 );
xnor ( n26510 , n26509 , n22200 );
and ( n26511 , n26506 , n26510 );
xor ( n26512 , n26218 , n26222 );
xor ( n26513 , n26512 , n26225 );
and ( n26514 , n26510 , n26513 );
and ( n26515 , n26506 , n26513 );
or ( n26516 , n26511 , n26514 , n26515 );
and ( n26517 , n22659 , n21957 );
and ( n26518 , n22409 , n21955 );
nor ( n26519 , n26517 , n26518 );
xnor ( n26520 , n26519 , n21967 );
and ( n26521 , n26516 , n26520 );
and ( n26522 , n23446 , n21804 );
and ( n26523 , n23284 , n21802 );
nor ( n26524 , n26522 , n26523 );
xnor ( n26525 , n26524 , n21814 );
and ( n26526 , n26520 , n26525 );
and ( n26527 , n26516 , n26525 );
or ( n26528 , n26521 , n26526 , n26527 );
and ( n26529 , n22080 , n22323 );
and ( n26530 , n22101 , n22321 );
nor ( n26531 , n26529 , n26530 );
xnor ( n26532 , n26531 , n22329 );
and ( n26533 , n26528 , n26532 );
xor ( n26534 , n26168 , n26172 );
xor ( n26535 , n26534 , n26175 );
and ( n26536 , n26532 , n26535 );
and ( n26537 , n26528 , n26535 );
or ( n26538 , n26533 , n26536 , n26537 );
and ( n26539 , n26482 , n26538 );
and ( n26540 , n21908 , n21735 );
and ( n26541 , n21870 , n21732 );
nor ( n26542 , n26540 , n26541 );
xnor ( n26543 , n26542 , n21730 );
and ( n26544 , n26538 , n26543 );
and ( n26545 , n26482 , n26543 );
or ( n26546 , n26539 , n26544 , n26545 );
and ( n26547 , n26467 , n26546 );
and ( n26548 , n26465 , n26546 );
or ( n26549 , n26468 , n26547 , n26548 );
and ( n26550 , n26462 , n26549 );
and ( n26551 , n26356 , n26549 );
or ( n26552 , n26463 , n26550 , n26551 );
and ( n26553 , n26353 , n26552 );
and ( n26554 , n26351 , n26552 );
or ( n26555 , n26354 , n26553 , n26554 );
and ( n26556 , n26299 , n26555 );
xor ( n26557 , n26299 , n26555 );
xor ( n26558 , n26351 , n26353 );
xor ( n26559 , n26558 , n26552 );
and ( n26560 , n22049 , n21854 );
and ( n26561 , n22033 , n21852 );
nor ( n26562 , n26560 , n26561 );
xnor ( n26563 , n26562 , n21864 );
and ( n26564 , n22101 , n21779 );
and ( n26565 , n22086 , n21777 );
nor ( n26566 , n26564 , n26565 );
xnor ( n26567 , n26566 , n21789 );
and ( n26568 , n26563 , n26567 );
xor ( n26569 , n26412 , n26416 );
xor ( n26570 , n26569 , n26419 );
and ( n26571 , n26567 , n26570 );
and ( n26572 , n26563 , n26570 );
or ( n26573 , n26568 , n26571 , n26572 );
xor ( n26574 , n26363 , n26371 );
and ( n26575 , n26360 , n22020 );
not ( n26576 , n26575 );
and ( n26577 , n26576 , n22028 );
and ( n26578 , n26360 , n22022 );
and ( n26579 , n26368 , n22020 );
nor ( n26580 , n26578 , n26579 );
xnor ( n26581 , n26580 , n22028 );
and ( n26582 , n26577 , n26581 );
and ( n26583 , n26368 , n22022 );
and ( n26584 , n26214 , n22020 );
nor ( n26585 , n26583 , n26584 );
xnor ( n26586 , n26585 , n22028 );
and ( n26587 , n26582 , n26586 );
and ( n26588 , n26586 , n26361 );
and ( n26589 , n26582 , n26361 );
or ( n26590 , n26587 , n26588 , n26589 );
and ( n26591 , n26574 , n26590 );
and ( n26592 , n26214 , n22022 );
and ( n26593 , n26107 , n22020 );
nor ( n26594 , n26592 , n26593 );
xnor ( n26595 , n26594 , n22028 );
and ( n26596 , n26590 , n26595 );
and ( n26597 , n26574 , n26595 );
or ( n26598 , n26591 , n26596 , n26597 );
and ( n26599 , n26107 , n22022 );
and ( n26600 , n25986 , n22020 );
nor ( n26601 , n26599 , n26600 );
xnor ( n26602 , n26601 , n22028 );
and ( n26603 , n26598 , n26602 );
xor ( n26604 , n26372 , n26376 );
xor ( n26605 , n26604 , n26378 );
and ( n26606 , n26602 , n26605 );
and ( n26607 , n26598 , n26605 );
or ( n26608 , n26603 , n26606 , n26607 );
and ( n26609 , n25427 , n21903 );
and ( n26610 , n25347 , n21901 );
nor ( n26611 , n26609 , n26610 );
xnor ( n26612 , n26611 , n21913 );
and ( n26613 , n26608 , n26612 );
xor ( n26614 , n26486 , n26490 );
xor ( n26615 , n26614 , n26493 );
and ( n26616 , n26612 , n26615 );
and ( n26617 , n26608 , n26615 );
or ( n26618 , n26613 , n26616 , n26617 );
and ( n26619 , n24753 , n22194 );
and ( n26620 , n24544 , n22192 );
nor ( n26621 , n26619 , n26620 );
xnor ( n26622 , n26621 , n22200 );
and ( n26623 , n26618 , n26622 );
and ( n26624 , n25004 , n21880 );
and ( n26625 , n24896 , n21878 );
nor ( n26626 , n26624 , n26625 );
xnor ( n26627 , n26626 , n21890 );
and ( n26628 , n26622 , n26627 );
and ( n26629 , n26618 , n26627 );
or ( n26630 , n26623 , n26628 , n26629 );
and ( n26631 , n24011 , n21828 );
and ( n26632 , n23954 , n21826 );
nor ( n26633 , n26631 , n26632 );
xnor ( n26634 , n26633 , n21838 );
and ( n26635 , n26630 , n26634 );
xor ( n26636 , n26400 , n26404 );
xor ( n26637 , n26636 , n26409 );
and ( n26638 , n26634 , n26637 );
and ( n26639 , n26630 , n26637 );
or ( n26640 , n26635 , n26638 , n26639 );
and ( n26641 , n22094 , n22323 );
and ( n26642 , n22080 , n22321 );
nor ( n26643 , n26641 , n26642 );
xnor ( n26644 , n26643 , n22329 );
and ( n26645 , n26640 , n26644 );
xor ( n26646 , n26305 , n26309 );
xor ( n26647 , n26646 , n26312 );
and ( n26648 , n26644 , n26647 );
and ( n26649 , n26640 , n26647 );
or ( n26650 , n26645 , n26648 , n26649 );
and ( n26651 , n26573 , n26650 );
xor ( n26652 , n26422 , n26426 );
xor ( n26653 , n26652 , n26429 );
and ( n26654 , n26650 , n26653 );
and ( n26655 , n26573 , n26653 );
or ( n26656 , n26651 , n26654 , n26655 );
xor ( n26657 , n26432 , n26436 );
xor ( n26658 , n26657 , n26441 );
and ( n26659 , n26656 , n26658 );
xor ( n26660 , n26327 , n26331 );
xor ( n26661 , n26660 , n26334 );
and ( n26662 , n26658 , n26661 );
and ( n26663 , n26656 , n26661 );
or ( n26664 , n26659 , n26662 , n26663 );
and ( n26665 , n21895 , n21735 );
and ( n26666 , n21908 , n21732 );
nor ( n26667 , n26665 , n26666 );
xnor ( n26668 , n26667 , n21730 );
and ( n26669 , n21919 , n22252 );
and ( n26670 , n21932 , n22250 );
nor ( n26671 , n26669 , n26670 );
xnor ( n26672 , n26671 , n22258 );
and ( n26673 , n26668 , n26672 );
xor ( n26674 , n26528 , n26532 );
xor ( n26675 , n26674 , n26535 );
and ( n26676 , n26672 , n26675 );
and ( n26677 , n26668 , n26675 );
or ( n26678 , n26673 , n26676 , n26677 );
xor ( n26679 , n26482 , n26538 );
xor ( n26680 , n26679 , n26543 );
and ( n26681 , n26678 , n26680 );
xor ( n26682 , n26448 , n26450 );
xor ( n26683 , n26682 , n26453 );
and ( n26684 , n26680 , n26683 );
and ( n26685 , n26678 , n26683 );
or ( n26686 , n26681 , n26684 , n26685 );
and ( n26687 , n26664 , n26686 );
xor ( n26688 , n26444 , n26456 );
xor ( n26689 , n26688 , n26459 );
and ( n26690 , n26686 , n26689 );
and ( n26691 , n26664 , n26689 );
or ( n26692 , n26687 , n26690 , n26691 );
xor ( n26693 , n26356 , n26462 );
xor ( n26694 , n26693 , n26549 );
and ( n26695 , n26692 , n26694 );
xor ( n26696 , n26465 , n26467 );
xor ( n26697 , n26696 , n26546 );
xor ( n26698 , n26664 , n26686 );
xor ( n26699 , n26698 , n26689 );
and ( n26700 , n26697 , n26699 );
and ( n26701 , n23074 , n21957 );
and ( n26702 , n22659 , n21955 );
nor ( n26703 , n26701 , n26702 );
xnor ( n26704 , n26703 , n21967 );
and ( n26705 , n23284 , n21978 );
and ( n26706 , n23165 , n21976 );
nor ( n26707 , n26705 , n26706 );
xnor ( n26708 , n26707 , n21988 );
and ( n26709 , n26704 , n26708 );
and ( n26710 , n23575 , n21804 );
and ( n26711 , n23446 , n21802 );
nor ( n26712 , n26710 , n26711 );
xnor ( n26713 , n26712 , n21814 );
and ( n26714 , n26708 , n26713 );
and ( n26715 , n26704 , n26713 );
or ( n26716 , n26709 , n26714 , n26715 );
and ( n26717 , n23954 , n21804 );
and ( n26718 , n23575 , n21802 );
nor ( n26719 , n26717 , n26718 );
xnor ( n26720 , n26719 , n21814 );
and ( n26721 , n24446 , n21828 );
and ( n26722 , n24011 , n21826 );
nor ( n26723 , n26721 , n26722 );
xnor ( n26724 , n26723 , n21838 );
and ( n26725 , n26720 , n26724 );
xor ( n26726 , n26496 , n26500 );
xor ( n26727 , n26726 , n26503 );
and ( n26728 , n26724 , n26727 );
and ( n26729 , n26720 , n26727 );
or ( n26730 , n26725 , n26728 , n26729 );
xor ( n26731 , n26630 , n26634 );
xor ( n26732 , n26731 , n26637 );
and ( n26733 , n26730 , n26732 );
xor ( n26734 , n26506 , n26510 );
xor ( n26735 , n26734 , n26513 );
and ( n26736 , n26732 , n26735 );
and ( n26737 , n26730 , n26735 );
or ( n26738 , n26733 , n26736 , n26737 );
and ( n26739 , n26716 , n26738 );
xor ( n26740 , n26516 , n26520 );
xor ( n26741 , n26740 , n26525 );
and ( n26742 , n26738 , n26741 );
and ( n26743 , n26716 , n26741 );
or ( n26744 , n26739 , n26742 , n26743 );
and ( n26745 , n22014 , n22252 );
and ( n26746 , n21919 , n22250 );
nor ( n26747 , n26745 , n26746 );
xnor ( n26748 , n26747 , n22258 );
and ( n26749 , n22056 , n22305 );
and ( n26750 , n22041 , n22303 );
nor ( n26751 , n26749 , n26750 );
xnor ( n26752 , n26751 , n22315 );
and ( n26753 , n26748 , n26752 );
xor ( n26754 , n26640 , n26644 );
xor ( n26755 , n26754 , n26647 );
and ( n26756 , n26752 , n26755 );
and ( n26757 , n26748 , n26755 );
or ( n26758 , n26753 , n26756 , n26757 );
and ( n26759 , n26744 , n26758 );
xor ( n26760 , n26472 , n26476 );
xor ( n26761 , n26760 , n26479 );
and ( n26762 , n26758 , n26761 );
and ( n26763 , n26744 , n26761 );
or ( n26764 , n26759 , n26762 , n26763 );
and ( n26765 , n25753 , n21903 );
and ( n26766 , n25633 , n21901 );
nor ( n26767 , n26765 , n26766 );
xnor ( n26768 , n26767 , n21913 );
and ( n26769 , n25986 , n21927 );
and ( n26770 , n25833 , n21925 );
nor ( n26771 , n26769 , n26770 );
xnor ( n26772 , n26771 , n21937 );
and ( n26773 , n26768 , n26772 );
xor ( n26774 , n26574 , n26590 );
xor ( n26775 , n26774 , n26595 );
and ( n26776 , n26772 , n26775 );
and ( n26777 , n26768 , n26775 );
or ( n26778 , n26773 , n26776 , n26777 );
and ( n26779 , n25347 , n21880 );
and ( n26780 , n25337 , n21878 );
nor ( n26781 , n26779 , n26780 );
xnor ( n26782 , n26781 , n21890 );
and ( n26783 , n26778 , n26782 );
and ( n26784 , n25633 , n21903 );
and ( n26785 , n25427 , n21901 );
nor ( n26786 , n26784 , n26785 );
xnor ( n26787 , n26786 , n21913 );
and ( n26788 , n25833 , n21927 );
and ( n26789 , n25753 , n21925 );
nor ( n26790 , n26788 , n26789 );
xnor ( n26791 , n26790 , n21937 );
xor ( n26792 , n26787 , n26791 );
xor ( n26793 , n26598 , n26602 );
xor ( n26794 , n26793 , n26605 );
xor ( n26795 , n26792 , n26794 );
and ( n26796 , n26782 , n26795 );
and ( n26797 , n26778 , n26795 );
or ( n26798 , n26783 , n26796 , n26797 );
and ( n26799 , n24544 , n21828 );
and ( n26800 , n24446 , n21826 );
nor ( n26801 , n26799 , n26800 );
xnor ( n26802 , n26801 , n21838 );
and ( n26803 , n26798 , n26802 );
and ( n26804 , n24896 , n22194 );
and ( n26805 , n24753 , n22192 );
nor ( n26806 , n26804 , n26805 );
xnor ( n26807 , n26806 , n22200 );
and ( n26808 , n26802 , n26807 );
and ( n26809 , n26798 , n26807 );
or ( n26810 , n26803 , n26808 , n26809 );
and ( n26811 , n23165 , n21957 );
and ( n26812 , n23074 , n21955 );
nor ( n26813 , n26811 , n26812 );
xnor ( n26814 , n26813 , n21967 );
and ( n26815 , n26810 , n26814 );
xor ( n26816 , n26720 , n26724 );
xor ( n26817 , n26816 , n26727 );
and ( n26818 , n26814 , n26817 );
and ( n26819 , n26810 , n26817 );
or ( n26820 , n26815 , n26818 , n26819 );
and ( n26821 , n22086 , n21854 );
and ( n26822 , n22049 , n21852 );
nor ( n26823 , n26821 , n26822 );
xnor ( n26824 , n26823 , n21864 );
and ( n26825 , n26820 , n26824 );
xor ( n26826 , n26704 , n26708 );
xor ( n26827 , n26826 , n26713 );
and ( n26828 , n26824 , n26827 );
and ( n26829 , n26820 , n26827 );
or ( n26830 , n26825 , n26828 , n26829 );
xor ( n26831 , n26577 , n26581 );
and ( n26832 , n26360 , n21925 );
not ( n26833 , n26832 );
and ( n26834 , n26833 , n21937 );
and ( n26835 , n26360 , n21927 );
and ( n26836 , n26368 , n21925 );
nor ( n26837 , n26835 , n26836 );
xnor ( n26838 , n26837 , n21937 );
and ( n26839 , n26834 , n26838 );
and ( n26840 , n26368 , n21927 );
and ( n26841 , n26214 , n21925 );
nor ( n26842 , n26840 , n26841 );
xnor ( n26843 , n26842 , n21937 );
and ( n26844 , n26839 , n26843 );
and ( n26845 , n26843 , n26575 );
and ( n26846 , n26839 , n26575 );
or ( n26847 , n26844 , n26845 , n26846 );
and ( n26848 , n26831 , n26847 );
and ( n26849 , n26214 , n21927 );
and ( n26850 , n26107 , n21925 );
nor ( n26851 , n26849 , n26850 );
xnor ( n26852 , n26851 , n21937 );
and ( n26853 , n26847 , n26852 );
and ( n26854 , n26831 , n26852 );
or ( n26855 , n26848 , n26853 , n26854 );
and ( n26856 , n26107 , n21927 );
and ( n26857 , n25986 , n21925 );
nor ( n26858 , n26856 , n26857 );
xnor ( n26859 , n26858 , n21937 );
and ( n26860 , n26855 , n26859 );
xor ( n26861 , n26582 , n26586 );
xor ( n26862 , n26861 , n26361 );
and ( n26863 , n26859 , n26862 );
and ( n26864 , n26855 , n26862 );
or ( n26865 , n26860 , n26863 , n26864 );
and ( n26866 , n25427 , n21880 );
and ( n26867 , n25347 , n21878 );
nor ( n26868 , n26866 , n26867 );
xnor ( n26869 , n26868 , n21890 );
and ( n26870 , n26865 , n26869 );
xor ( n26871 , n26768 , n26772 );
xor ( n26872 , n26871 , n26775 );
and ( n26873 , n26869 , n26872 );
and ( n26874 , n26865 , n26872 );
or ( n26875 , n26870 , n26873 , n26874 );
and ( n26876 , n24753 , n21828 );
and ( n26877 , n24544 , n21826 );
nor ( n26878 , n26876 , n26877 );
xnor ( n26879 , n26878 , n21838 );
and ( n26880 , n26875 , n26879 );
and ( n26881 , n25004 , n22194 );
and ( n26882 , n24896 , n22192 );
nor ( n26883 , n26881 , n26882 );
xnor ( n26884 , n26883 , n22200 );
and ( n26885 , n26879 , n26884 );
and ( n26886 , n26875 , n26884 );
or ( n26887 , n26880 , n26885 , n26886 );
and ( n26888 , n24011 , n21804 );
and ( n26889 , n23954 , n21802 );
nor ( n26890 , n26888 , n26889 );
xnor ( n26891 , n26890 , n21814 );
and ( n26892 , n26887 , n26891 );
and ( n26893 , n26787 , n26791 );
and ( n26894 , n26791 , n26794 );
and ( n26895 , n26787 , n26794 );
or ( n26896 , n26893 , n26894 , n26895 );
and ( n26897 , n25337 , n21880 );
and ( n26898 , n25004 , n21878 );
nor ( n26899 , n26897 , n26898 );
xnor ( n26900 , n26899 , n21890 );
xor ( n26901 , n26896 , n26900 );
xor ( n26902 , n26608 , n26612 );
xor ( n26903 , n26902 , n26615 );
xor ( n26904 , n26901 , n26903 );
and ( n26905 , n26891 , n26904 );
and ( n26906 , n26887 , n26904 );
or ( n26907 , n26892 , n26905 , n26906 );
and ( n26908 , n22094 , n21779 );
and ( n26909 , n22080 , n21777 );
nor ( n26910 , n26908 , n26909 );
xnor ( n26911 , n26910 , n21789 );
and ( n26912 , n26907 , n26911 );
and ( n26913 , n22659 , n22323 );
and ( n26914 , n22409 , n22321 );
nor ( n26915 , n26913 , n26914 );
xnor ( n26916 , n26915 , n22329 );
and ( n26917 , n26911 , n26916 );
and ( n26918 , n26907 , n26916 );
or ( n26919 , n26912 , n26917 , n26918 );
and ( n26920 , n22041 , n22252 );
and ( n26921 , n22014 , n22250 );
nor ( n26922 , n26920 , n26921 );
xnor ( n26923 , n26922 , n22258 );
and ( n26924 , n26919 , n26923 );
xor ( n26925 , n26730 , n26732 );
xor ( n26926 , n26925 , n26735 );
and ( n26927 , n26923 , n26926 );
and ( n26928 , n26919 , n26926 );
or ( n26929 , n26924 , n26927 , n26928 );
and ( n26930 , n26830 , n26929 );
xor ( n26931 , n26716 , n26738 );
xor ( n26932 , n26931 , n26741 );
and ( n26933 , n26929 , n26932 );
and ( n26934 , n26830 , n26932 );
or ( n26935 , n26930 , n26933 , n26934 );
and ( n26936 , n26896 , n26900 );
and ( n26937 , n26900 , n26903 );
and ( n26938 , n26896 , n26903 );
or ( n26939 , n26936 , n26937 , n26938 );
and ( n26940 , n23446 , n21978 );
and ( n26941 , n23284 , n21976 );
nor ( n26942 , n26940 , n26941 );
xnor ( n26943 , n26942 , n21988 );
and ( n26944 , n26939 , n26943 );
xor ( n26945 , n26618 , n26622 );
xor ( n26946 , n26945 , n26627 );
and ( n26947 , n26943 , n26946 );
and ( n26948 , n26939 , n26946 );
or ( n26949 , n26944 , n26947 , n26948 );
and ( n26950 , n22080 , n21779 );
and ( n26951 , n22101 , n21777 );
nor ( n26952 , n26950 , n26951 );
xnor ( n26953 , n26952 , n21789 );
and ( n26954 , n26949 , n26953 );
and ( n26955 , n22409 , n22323 );
and ( n26956 , n22094 , n22321 );
nor ( n26957 , n26955 , n26956 );
xnor ( n26958 , n26957 , n22329 );
and ( n26959 , n26953 , n26958 );
and ( n26960 , n26949 , n26958 );
or ( n26961 , n26954 , n26959 , n26960 );
and ( n26962 , n21932 , n21735 );
and ( n26963 , n21895 , n21732 );
nor ( n26964 , n26962 , n26963 );
xnor ( n26965 , n26964 , n21730 );
and ( n26966 , n26961 , n26965 );
xor ( n26967 , n26563 , n26567 );
xor ( n26968 , n26967 , n26570 );
and ( n26969 , n26965 , n26968 );
and ( n26970 , n26961 , n26968 );
or ( n26971 , n26966 , n26969 , n26970 );
and ( n26972 , n26935 , n26971 );
xor ( n26973 , n26573 , n26650 );
xor ( n26974 , n26973 , n26653 );
and ( n26975 , n26971 , n26974 );
and ( n26976 , n26935 , n26974 );
or ( n26977 , n26972 , n26975 , n26976 );
and ( n26978 , n26764 , n26977 );
xor ( n26979 , n26656 , n26658 );
xor ( n26980 , n26979 , n26661 );
and ( n26981 , n26977 , n26980 );
and ( n26982 , n26764 , n26980 );
or ( n26983 , n26978 , n26981 , n26982 );
and ( n26984 , n26699 , n26983 );
and ( n26985 , n26697 , n26983 );
or ( n26986 , n26700 , n26984 , n26985 );
and ( n26987 , n26694 , n26986 );
and ( n26988 , n26692 , n26986 );
or ( n26989 , n26695 , n26987 , n26988 );
and ( n26990 , n26559 , n26989 );
xor ( n26991 , n26559 , n26989 );
xor ( n26992 , n26692 , n26694 );
xor ( n26993 , n26992 , n26986 );
and ( n26994 , n22049 , n22305 );
and ( n26995 , n22033 , n22303 );
nor ( n26996 , n26994 , n26995 );
xnor ( n26997 , n26996 , n22315 );
and ( n26998 , n22101 , n21854 );
and ( n26999 , n22086 , n21852 );
nor ( n27000 , n26998 , n26999 );
xnor ( n27001 , n27000 , n21864 );
and ( n27002 , n26997 , n27001 );
xor ( n27003 , n26939 , n26943 );
xor ( n27004 , n27003 , n26946 );
and ( n27005 , n27001 , n27004 );
and ( n27006 , n26997 , n27004 );
or ( n27007 , n27002 , n27005 , n27006 );
and ( n27008 , n21919 , n21735 );
and ( n27009 , n21932 , n21732 );
nor ( n27010 , n27008 , n27009 );
xnor ( n27011 , n27010 , n21730 );
and ( n27012 , n27007 , n27011 );
and ( n27013 , n22033 , n22305 );
and ( n27014 , n22056 , n22303 );
nor ( n27015 , n27013 , n27014 );
xnor ( n27016 , n27015 , n22315 );
and ( n27017 , n27011 , n27016 );
and ( n27018 , n27007 , n27016 );
or ( n27019 , n27012 , n27017 , n27018 );
xor ( n27020 , n26961 , n26965 );
xor ( n27021 , n27020 , n26968 );
and ( n27022 , n27019 , n27021 );
xor ( n27023 , n26748 , n26752 );
xor ( n27024 , n27023 , n26755 );
and ( n27025 , n27021 , n27024 );
and ( n27026 , n27019 , n27024 );
or ( n27027 , n27022 , n27025 , n27026 );
xor ( n27028 , n26744 , n26758 );
xor ( n27029 , n27028 , n26761 );
and ( n27030 , n27027 , n27029 );
xor ( n27031 , n26668 , n26672 );
xor ( n27032 , n27031 , n26675 );
and ( n27033 , n27029 , n27032 );
and ( n27034 , n27027 , n27032 );
or ( n27035 , n27030 , n27033 , n27034 );
xor ( n27036 , n26764 , n26977 );
xor ( n27037 , n27036 , n26980 );
and ( n27038 , n27035 , n27037 );
xor ( n27039 , n26678 , n26680 );
xor ( n27040 , n27039 , n26683 );
and ( n27041 , n27037 , n27040 );
and ( n27042 , n27035 , n27040 );
or ( n27043 , n27038 , n27041 , n27042 );
xor ( n27044 , n26697 , n26699 );
xor ( n27045 , n27044 , n26983 );
and ( n27046 , n27043 , n27045 );
xor ( n27047 , n27043 , n27045 );
xor ( n27048 , n27035 , n27037 );
xor ( n27049 , n27048 , n27040 );
and ( n27050 , n23284 , n21957 );
and ( n27051 , n23165 , n21955 );
nor ( n27052 , n27050 , n27051 );
xnor ( n27053 , n27052 , n21967 );
and ( n27054 , n23575 , n21978 );
and ( n27055 , n23446 , n21976 );
nor ( n27056 , n27054 , n27055 );
xnor ( n27057 , n27056 , n21988 );
and ( n27058 , n27053 , n27057 );
xor ( n27059 , n26798 , n26802 );
xor ( n27060 , n27059 , n26807 );
and ( n27061 , n27057 , n27060 );
and ( n27062 , n27053 , n27060 );
or ( n27063 , n27058 , n27061 , n27062 );
and ( n27064 , n23954 , n21978 );
and ( n27065 , n23575 , n21976 );
nor ( n27066 , n27064 , n27065 );
xnor ( n27067 , n27066 , n21988 );
and ( n27068 , n24446 , n21804 );
and ( n27069 , n24011 , n21802 );
nor ( n27070 , n27068 , n27069 );
xnor ( n27071 , n27070 , n21814 );
and ( n27072 , n27067 , n27071 );
xor ( n27073 , n26778 , n26782 );
xor ( n27074 , n27073 , n26795 );
and ( n27075 , n27071 , n27074 );
and ( n27076 , n27067 , n27074 );
or ( n27077 , n27072 , n27075 , n27076 );
and ( n27078 , n23074 , n22323 );
and ( n27079 , n22659 , n22321 );
nor ( n27080 , n27078 , n27079 );
xnor ( n27081 , n27080 , n22329 );
and ( n27082 , n27077 , n27081 );
xor ( n27083 , n26887 , n26891 );
xor ( n27084 , n27083 , n26904 );
and ( n27085 , n27081 , n27084 );
and ( n27086 , n27077 , n27084 );
or ( n27087 , n27082 , n27085 , n27086 );
and ( n27088 , n27063 , n27087 );
xor ( n27089 , n26810 , n26814 );
xor ( n27090 , n27089 , n26817 );
and ( n27091 , n27087 , n27090 );
and ( n27092 , n27063 , n27090 );
or ( n27093 , n27088 , n27091 , n27092 );
xor ( n27094 , n26949 , n26953 );
xor ( n27095 , n27094 , n26958 );
and ( n27096 , n27093 , n27095 );
xor ( n27097 , n26820 , n26824 );
xor ( n27098 , n27097 , n26827 );
and ( n27099 , n27095 , n27098 );
and ( n27100 , n27093 , n27098 );
or ( n27101 , n27096 , n27099 , n27100 );
and ( n27102 , n25633 , n21880 );
and ( n27103 , n25427 , n21878 );
nor ( n27104 , n27102 , n27103 );
xnor ( n27105 , n27104 , n21890 );
and ( n27106 , n25833 , n21903 );
and ( n27107 , n25753 , n21901 );
nor ( n27108 , n27106 , n27107 );
xnor ( n27109 , n27108 , n21913 );
and ( n27110 , n27105 , n27109 );
xor ( n27111 , n26855 , n26859 );
xor ( n27112 , n27111 , n26862 );
and ( n27113 , n27109 , n27112 );
and ( n27114 , n27105 , n27112 );
or ( n27115 , n27110 , n27113 , n27114 );
and ( n27116 , n24896 , n21828 );
and ( n27117 , n24753 , n21826 );
nor ( n27118 , n27116 , n27117 );
xnor ( n27119 , n27118 , n21838 );
and ( n27120 , n27115 , n27119 );
and ( n27121 , n25337 , n22194 );
and ( n27122 , n25004 , n22192 );
nor ( n27123 , n27121 , n27122 );
xnor ( n27124 , n27123 , n22200 );
and ( n27125 , n27119 , n27124 );
and ( n27126 , n27115 , n27124 );
or ( n27127 , n27120 , n27125 , n27126 );
and ( n27128 , n23165 , n22323 );
and ( n27129 , n23074 , n22321 );
nor ( n27130 , n27128 , n27129 );
xnor ( n27131 , n27130 , n22329 );
and ( n27132 , n27127 , n27131 );
xor ( n27133 , n26875 , n26879 );
xor ( n27134 , n27133 , n26884 );
and ( n27135 , n27131 , n27134 );
and ( n27136 , n27127 , n27134 );
or ( n27137 , n27132 , n27135 , n27136 );
and ( n27138 , n22086 , n22305 );
and ( n27139 , n22049 , n22303 );
nor ( n27140 , n27138 , n27139 );
xnor ( n27141 , n27140 , n22315 );
and ( n27142 , n27137 , n27141 );
and ( n27143 , n22409 , n21779 );
and ( n27144 , n22094 , n21777 );
nor ( n27145 , n27143 , n27144 );
xnor ( n27146 , n27145 , n21789 );
and ( n27147 , n27141 , n27146 );
and ( n27148 , n27137 , n27146 );
or ( n27149 , n27142 , n27147 , n27148 );
and ( n27150 , n22014 , n21735 );
and ( n27151 , n21919 , n21732 );
nor ( n27152 , n27150 , n27151 );
xnor ( n27153 , n27152 , n21730 );
and ( n27154 , n27149 , n27153 );
and ( n27155 , n22056 , n22252 );
and ( n27156 , n22041 , n22250 );
nor ( n27157 , n27155 , n27156 );
xnor ( n27158 , n27157 , n22258 );
and ( n27159 , n27153 , n27158 );
and ( n27160 , n27149 , n27158 );
or ( n27161 , n27154 , n27159 , n27160 );
and ( n27162 , n25753 , n21880 );
and ( n27163 , n25633 , n21878 );
nor ( n27164 , n27162 , n27163 );
xnor ( n27165 , n27164 , n21890 );
and ( n27166 , n25986 , n21903 );
and ( n27167 , n25833 , n21901 );
nor ( n27168 , n27166 , n27167 );
xnor ( n27169 , n27168 , n21913 );
and ( n27170 , n27165 , n27169 );
xor ( n27171 , n26831 , n26847 );
xor ( n27172 , n27171 , n26852 );
and ( n27173 , n27169 , n27172 );
and ( n27174 , n27165 , n27172 );
or ( n27175 , n27170 , n27173 , n27174 );
and ( n27176 , n25347 , n22194 );
and ( n27177 , n25337 , n22192 );
nor ( n27178 , n27176 , n27177 );
xnor ( n27179 , n27178 , n22200 );
and ( n27180 , n27175 , n27179 );
xor ( n27181 , n27105 , n27109 );
xor ( n27182 , n27181 , n27112 );
and ( n27183 , n27179 , n27182 );
and ( n27184 , n27175 , n27182 );
or ( n27185 , n27180 , n27183 , n27184 );
and ( n27186 , n24544 , n21804 );
and ( n27187 , n24446 , n21802 );
nor ( n27188 , n27186 , n27187 );
xnor ( n27189 , n27188 , n21814 );
and ( n27190 , n27185 , n27189 );
xor ( n27191 , n26865 , n26869 );
xor ( n27192 , n27191 , n26872 );
and ( n27193 , n27189 , n27192 );
and ( n27194 , n27185 , n27192 );
or ( n27195 , n27190 , n27193 , n27194 );
and ( n27196 , n23446 , n21957 );
and ( n27197 , n23284 , n21955 );
nor ( n27198 , n27196 , n27197 );
xnor ( n27199 , n27198 , n21967 );
and ( n27200 , n27195 , n27199 );
xor ( n27201 , n27067 , n27071 );
xor ( n27202 , n27201 , n27074 );
and ( n27203 , n27199 , n27202 );
and ( n27204 , n27195 , n27202 );
or ( n27205 , n27200 , n27203 , n27204 );
and ( n27206 , n22080 , n21854 );
and ( n27207 , n22101 , n21852 );
nor ( n27208 , n27206 , n27207 );
xnor ( n27209 , n27208 , n21864 );
and ( n27210 , n27205 , n27209 );
xor ( n27211 , n27053 , n27057 );
xor ( n27212 , n27211 , n27060 );
and ( n27213 , n27209 , n27212 );
and ( n27214 , n27205 , n27212 );
or ( n27215 , n27210 , n27213 , n27214 );
xor ( n27216 , n26907 , n26911 );
xor ( n27217 , n27216 , n26916 );
and ( n27218 , n27215 , n27217 );
xor ( n27219 , n26997 , n27001 );
xor ( n27220 , n27219 , n27004 );
and ( n27221 , n27217 , n27220 );
and ( n27222 , n27215 , n27220 );
or ( n27223 , n27218 , n27221 , n27222 );
and ( n27224 , n27161 , n27223 );
xor ( n27225 , n26919 , n26923 );
xor ( n27226 , n27225 , n26926 );
and ( n27227 , n27223 , n27226 );
and ( n27228 , n27161 , n27226 );
or ( n27229 , n27224 , n27227 , n27228 );
and ( n27230 , n27101 , n27229 );
xor ( n27231 , n26830 , n26929 );
xor ( n27232 , n27231 , n26932 );
and ( n27233 , n27229 , n27232 );
and ( n27234 , n27101 , n27232 );
or ( n27235 , n27230 , n27233 , n27234 );
xor ( n27236 , n26935 , n26971 );
xor ( n27237 , n27236 , n26974 );
and ( n27238 , n27235 , n27237 );
xor ( n27239 , n27027 , n27029 );
xor ( n27240 , n27239 , n27032 );
and ( n27241 , n27237 , n27240 );
and ( n27242 , n27235 , n27240 );
or ( n27243 , n27238 , n27241 , n27242 );
and ( n27244 , n27049 , n27243 );
xor ( n27245 , n27049 , n27243 );
xor ( n27246 , n27235 , n27237 );
xor ( n27247 , n27246 , n27240 );
and ( n27248 , n22041 , n21735 );
and ( n27249 , n22014 , n21732 );
nor ( n27250 , n27248 , n27249 );
xnor ( n27251 , n27250 , n21730 );
and ( n27252 , n22033 , n22252 );
and ( n27253 , n22056 , n22250 );
nor ( n27254 , n27252 , n27253 );
xnor ( n27255 , n27254 , n22258 );
and ( n27256 , n27251 , n27255 );
xor ( n27257 , n27077 , n27081 );
xor ( n27258 , n27257 , n27084 );
and ( n27259 , n27255 , n27258 );
and ( n27260 , n27251 , n27258 );
or ( n27261 , n27256 , n27259 , n27260 );
xor ( n27262 , n27149 , n27153 );
xor ( n27263 , n27262 , n27158 );
and ( n27264 , n27261 , n27263 );
xor ( n27265 , n27063 , n27087 );
xor ( n27266 , n27265 , n27090 );
and ( n27267 , n27263 , n27266 );
and ( n27268 , n27261 , n27266 );
or ( n27269 , n27264 , n27267 , n27268 );
xor ( n27270 , n27007 , n27011 );
xor ( n27271 , n27270 , n27016 );
and ( n27272 , n27269 , n27271 );
xor ( n27273 , n27093 , n27095 );
xor ( n27274 , n27273 , n27098 );
and ( n27275 , n27271 , n27274 );
and ( n27276 , n27269 , n27274 );
or ( n27277 , n27272 , n27275 , n27276 );
xor ( n27278 , n27101 , n27229 );
xor ( n27279 , n27278 , n27232 );
and ( n27280 , n27277 , n27279 );
xor ( n27281 , n27019 , n27021 );
xor ( n27282 , n27281 , n27024 );
and ( n27283 , n27279 , n27282 );
and ( n27284 , n27277 , n27282 );
or ( n27285 , n27280 , n27283 , n27284 );
and ( n27286 , n27247 , n27285 );
xor ( n27287 , n27247 , n27285 );
xor ( n27288 , n27277 , n27279 );
xor ( n27289 , n27288 , n27282 );
xor ( n27290 , n26834 , n26838 );
and ( n27291 , n26360 , n21901 );
not ( n27292 , n27291 );
and ( n27293 , n27292 , n21913 );
and ( n27294 , n26360 , n21903 );
and ( n27295 , n26368 , n21901 );
nor ( n27296 , n27294 , n27295 );
xnor ( n27297 , n27296 , n21913 );
and ( n27298 , n27293 , n27297 );
and ( n27299 , n26368 , n21903 );
and ( n27300 , n26214 , n21901 );
nor ( n27301 , n27299 , n27300 );
xnor ( n27302 , n27301 , n21913 );
and ( n27303 , n27298 , n27302 );
and ( n27304 , n27302 , n26832 );
and ( n27305 , n27298 , n26832 );
or ( n27306 , n27303 , n27304 , n27305 );
and ( n27307 , n27290 , n27306 );
and ( n27308 , n26214 , n21903 );
and ( n27309 , n26107 , n21901 );
nor ( n27310 , n27308 , n27309 );
xnor ( n27311 , n27310 , n21913 );
and ( n27312 , n27306 , n27311 );
and ( n27313 , n27290 , n27311 );
or ( n27314 , n27307 , n27312 , n27313 );
and ( n27315 , n26107 , n21903 );
and ( n27316 , n25986 , n21901 );
nor ( n27317 , n27315 , n27316 );
xnor ( n27318 , n27317 , n21913 );
and ( n27319 , n27314 , n27318 );
xor ( n27320 , n26839 , n26843 );
xor ( n27321 , n27320 , n26575 );
and ( n27322 , n27318 , n27321 );
and ( n27323 , n27314 , n27321 );
or ( n27324 , n27319 , n27322 , n27323 );
and ( n27325 , n25427 , n22194 );
and ( n27326 , n25347 , n22192 );
nor ( n27327 , n27325 , n27326 );
xnor ( n27328 , n27327 , n22200 );
and ( n27329 , n27324 , n27328 );
xor ( n27330 , n27165 , n27169 );
xor ( n27331 , n27330 , n27172 );
and ( n27332 , n27328 , n27331 );
and ( n27333 , n27324 , n27331 );
or ( n27334 , n27329 , n27332 , n27333 );
and ( n27335 , n24753 , n21804 );
and ( n27336 , n24544 , n21802 );
nor ( n27337 , n27335 , n27336 );
xnor ( n27338 , n27337 , n21814 );
and ( n27339 , n27334 , n27338 );
and ( n27340 , n25004 , n21828 );
and ( n27341 , n24896 , n21826 );
nor ( n27342 , n27340 , n27341 );
xnor ( n27343 , n27342 , n21838 );
and ( n27344 , n27338 , n27343 );
and ( n27345 , n27334 , n27343 );
or ( n27346 , n27339 , n27344 , n27345 );
and ( n27347 , n24011 , n21978 );
and ( n27348 , n23954 , n21976 );
nor ( n27349 , n27347 , n27348 );
xnor ( n27350 , n27349 , n21988 );
and ( n27351 , n27346 , n27350 );
xor ( n27352 , n27115 , n27119 );
xor ( n27353 , n27352 , n27124 );
and ( n27354 , n27350 , n27353 );
and ( n27355 , n27346 , n27353 );
or ( n27356 , n27351 , n27354 , n27355 );
and ( n27357 , n22094 , n21854 );
and ( n27358 , n22080 , n21852 );
nor ( n27359 , n27357 , n27358 );
xnor ( n27360 , n27359 , n21864 );
and ( n27361 , n27356 , n27360 );
and ( n27362 , n22659 , n21779 );
and ( n27363 , n22409 , n21777 );
nor ( n27364 , n27362 , n27363 );
xnor ( n27365 , n27364 , n21789 );
and ( n27366 , n27360 , n27365 );
and ( n27367 , n27356 , n27365 );
or ( n27368 , n27361 , n27366 , n27367 );
and ( n27369 , n22049 , n22252 );
and ( n27370 , n22033 , n22250 );
nor ( n27371 , n27369 , n27370 );
xnor ( n27372 , n27371 , n22258 );
and ( n27373 , n22101 , n22305 );
and ( n27374 , n22086 , n22303 );
nor ( n27375 , n27373 , n27374 );
xnor ( n27376 , n27375 , n22315 );
and ( n27377 , n27372 , n27376 );
xor ( n27378 , n27127 , n27131 );
xor ( n27379 , n27378 , n27134 );
and ( n27380 , n27376 , n27379 );
and ( n27381 , n27372 , n27379 );
or ( n27382 , n27377 , n27380 , n27381 );
and ( n27383 , n27368 , n27382 );
xor ( n27384 , n27137 , n27141 );
xor ( n27385 , n27384 , n27146 );
and ( n27386 , n27382 , n27385 );
and ( n27387 , n27368 , n27385 );
or ( n27388 , n27383 , n27386 , n27387 );
and ( n27389 , n25633 , n22194 );
and ( n27390 , n25427 , n22192 );
nor ( n27391 , n27389 , n27390 );
xnor ( n27392 , n27391 , n22200 );
and ( n27393 , n25833 , n21880 );
and ( n27394 , n25753 , n21878 );
nor ( n27395 , n27393 , n27394 );
xnor ( n27396 , n27395 , n21890 );
and ( n27397 , n27392 , n27396 );
xor ( n27398 , n27314 , n27318 );
xor ( n27399 , n27398 , n27321 );
and ( n27400 , n27396 , n27399 );
and ( n27401 , n27392 , n27399 );
or ( n27402 , n27397 , n27400 , n27401 );
and ( n27403 , n24896 , n21804 );
and ( n27404 , n24753 , n21802 );
nor ( n27405 , n27403 , n27404 );
xnor ( n27406 , n27405 , n21814 );
and ( n27407 , n27402 , n27406 );
and ( n27408 , n25337 , n21828 );
and ( n27409 , n25004 , n21826 );
nor ( n27410 , n27408 , n27409 );
xnor ( n27411 , n27410 , n21838 );
and ( n27412 , n27406 , n27411 );
and ( n27413 , n27402 , n27411 );
or ( n27414 , n27407 , n27412 , n27413 );
and ( n27415 , n25753 , n22194 );
and ( n27416 , n25633 , n22192 );
nor ( n27417 , n27415 , n27416 );
xnor ( n27418 , n27417 , n22200 );
and ( n27419 , n25986 , n21880 );
and ( n27420 , n25833 , n21878 );
nor ( n27421 , n27419 , n27420 );
xnor ( n27422 , n27421 , n21890 );
and ( n27423 , n27418 , n27422 );
xor ( n27424 , n27290 , n27306 );
xor ( n27425 , n27424 , n27311 );
and ( n27426 , n27422 , n27425 );
and ( n27427 , n27418 , n27425 );
or ( n27428 , n27423 , n27426 , n27427 );
and ( n27429 , n25347 , n21828 );
and ( n27430 , n25337 , n21826 );
nor ( n27431 , n27429 , n27430 );
xnor ( n27432 , n27431 , n21838 );
and ( n27433 , n27428 , n27432 );
xor ( n27434 , n27392 , n27396 );
xor ( n27435 , n27434 , n27399 );
and ( n27436 , n27432 , n27435 );
and ( n27437 , n27428 , n27435 );
or ( n27438 , n27433 , n27436 , n27437 );
and ( n27439 , n24544 , n21978 );
and ( n27440 , n24446 , n21976 );
nor ( n27441 , n27439 , n27440 );
xnor ( n27442 , n27441 , n21988 );
and ( n27443 , n27438 , n27442 );
xor ( n27444 , n27324 , n27328 );
xor ( n27445 , n27444 , n27331 );
and ( n27446 , n27442 , n27445 );
and ( n27447 , n27438 , n27445 );
or ( n27448 , n27443 , n27446 , n27447 );
and ( n27449 , n27414 , n27448 );
xor ( n27450 , n27334 , n27338 );
xor ( n27451 , n27450 , n27343 );
and ( n27452 , n27448 , n27451 );
and ( n27453 , n27414 , n27451 );
or ( n27454 , n27449 , n27452 , n27453 );
and ( n27455 , n22086 , n22252 );
and ( n27456 , n22049 , n22250 );
nor ( n27457 , n27455 , n27456 );
xnor ( n27458 , n27457 , n22258 );
and ( n27459 , n27454 , n27458 );
xor ( n27460 , n27346 , n27350 );
xor ( n27461 , n27460 , n27353 );
and ( n27462 , n27458 , n27461 );
and ( n27463 , n27454 , n27461 );
or ( n27464 , n27459 , n27462 , n27463 );
and ( n27465 , n22056 , n21735 );
and ( n27466 , n22041 , n21732 );
nor ( n27467 , n27465 , n27466 );
xnor ( n27468 , n27467 , n21730 );
and ( n27469 , n27464 , n27468 );
xor ( n27470 , n27356 , n27360 );
xor ( n27471 , n27470 , n27365 );
and ( n27472 , n27468 , n27471 );
and ( n27473 , n27464 , n27471 );
or ( n27474 , n27469 , n27472 , n27473 );
and ( n27475 , n23954 , n21957 );
and ( n27476 , n23575 , n21955 );
nor ( n27477 , n27475 , n27476 );
xnor ( n27478 , n27477 , n21967 );
and ( n27479 , n24446 , n21978 );
and ( n27480 , n24011 , n21976 );
nor ( n27481 , n27479 , n27480 );
xnor ( n27482 , n27481 , n21988 );
and ( n27483 , n27478 , n27482 );
xor ( n27484 , n27175 , n27179 );
xor ( n27485 , n27484 , n27182 );
and ( n27486 , n27482 , n27485 );
and ( n27487 , n27478 , n27485 );
or ( n27488 , n27483 , n27486 , n27487 );
and ( n27489 , n22409 , n21854 );
and ( n27490 , n22094 , n21852 );
nor ( n27491 , n27489 , n27490 );
xnor ( n27492 , n27491 , n21864 );
and ( n27493 , n27488 , n27492 );
and ( n27494 , n23074 , n21779 );
and ( n27495 , n22659 , n21777 );
nor ( n27496 , n27494 , n27495 );
xnor ( n27497 , n27496 , n21789 );
and ( n27498 , n27492 , n27497 );
and ( n27499 , n27488 , n27497 );
or ( n27500 , n27493 , n27498 , n27499 );
and ( n27501 , n23284 , n22323 );
and ( n27502 , n23165 , n22321 );
nor ( n27503 , n27501 , n27502 );
xnor ( n27504 , n27503 , n22329 );
and ( n27505 , n23575 , n21957 );
and ( n27506 , n23446 , n21955 );
nor ( n27507 , n27505 , n27506 );
xnor ( n27508 , n27507 , n21967 );
and ( n27509 , n27504 , n27508 );
xor ( n27510 , n27185 , n27189 );
xor ( n27511 , n27510 , n27192 );
and ( n27512 , n27508 , n27511 );
and ( n27513 , n27504 , n27511 );
or ( n27514 , n27509 , n27512 , n27513 );
and ( n27515 , n27500 , n27514 );
xor ( n27516 , n27195 , n27199 );
xor ( n27517 , n27516 , n27202 );
and ( n27518 , n27514 , n27517 );
and ( n27519 , n27500 , n27517 );
or ( n27520 , n27515 , n27518 , n27519 );
and ( n27521 , n27474 , n27520 );
xor ( n27522 , n27205 , n27209 );
xor ( n27523 , n27522 , n27212 );
and ( n27524 , n27520 , n27523 );
and ( n27525 , n27474 , n27523 );
or ( n27526 , n27521 , n27524 , n27525 );
and ( n27527 , n27388 , n27526 );
xor ( n27528 , n27215 , n27217 );
xor ( n27529 , n27528 , n27220 );
and ( n27530 , n27526 , n27529 );
and ( n27531 , n27388 , n27529 );
or ( n27532 , n27527 , n27530 , n27531 );
xor ( n27533 , n27269 , n27271 );
xor ( n27534 , n27533 , n27274 );
and ( n27535 , n27532 , n27534 );
xor ( n27536 , n27161 , n27223 );
xor ( n27537 , n27536 , n27226 );
and ( n27538 , n27534 , n27537 );
and ( n27539 , n27532 , n27537 );
or ( n27540 , n27535 , n27538 , n27539 );
and ( n27541 , n27289 , n27540 );
xor ( n27542 , n27289 , n27540 );
xor ( n27543 , n27532 , n27534 );
xor ( n27544 , n27543 , n27537 );
xor ( n27545 , n27293 , n27297 );
and ( n27546 , n26360 , n21878 );
not ( n27547 , n27546 );
and ( n27548 , n27547 , n21890 );
and ( n27549 , n26360 , n21880 );
and ( n27550 , n26368 , n21878 );
nor ( n27551 , n27549 , n27550 );
xnor ( n27552 , n27551 , n21890 );
and ( n27553 , n27548 , n27552 );
and ( n27554 , n26368 , n21880 );
and ( n27555 , n26214 , n21878 );
nor ( n27556 , n27554 , n27555 );
xnor ( n27557 , n27556 , n21890 );
and ( n27558 , n27553 , n27557 );
and ( n27559 , n27557 , n27291 );
and ( n27560 , n27553 , n27291 );
or ( n27561 , n27558 , n27559 , n27560 );
and ( n27562 , n27545 , n27561 );
and ( n27563 , n26214 , n21880 );
and ( n27564 , n26107 , n21878 );
nor ( n27565 , n27563 , n27564 );
xnor ( n27566 , n27565 , n21890 );
and ( n27567 , n27561 , n27566 );
and ( n27568 , n27545 , n27566 );
or ( n27569 , n27562 , n27567 , n27568 );
and ( n27570 , n26107 , n21880 );
and ( n27571 , n25986 , n21878 );
nor ( n27572 , n27570 , n27571 );
xnor ( n27573 , n27572 , n21890 );
and ( n27574 , n27569 , n27573 );
xor ( n27575 , n27298 , n27302 );
xor ( n27576 , n27575 , n26832 );
and ( n27577 , n27573 , n27576 );
and ( n27578 , n27569 , n27576 );
or ( n27579 , n27574 , n27577 , n27578 );
and ( n27580 , n25427 , n21828 );
and ( n27581 , n25347 , n21826 );
nor ( n27582 , n27580 , n27581 );
xnor ( n27583 , n27582 , n21838 );
and ( n27584 , n27579 , n27583 );
xor ( n27585 , n27418 , n27422 );
xor ( n27586 , n27585 , n27425 );
and ( n27587 , n27583 , n27586 );
and ( n27588 , n27579 , n27586 );
or ( n27589 , n27584 , n27587 , n27588 );
and ( n27590 , n24753 , n21978 );
and ( n27591 , n24544 , n21976 );
nor ( n27592 , n27590 , n27591 );
xnor ( n27593 , n27592 , n21988 );
and ( n27594 , n27589 , n27593 );
and ( n27595 , n25004 , n21804 );
and ( n27596 , n24896 , n21802 );
nor ( n27597 , n27595 , n27596 );
xnor ( n27598 , n27597 , n21814 );
and ( n27599 , n27593 , n27598 );
and ( n27600 , n27589 , n27598 );
or ( n27601 , n27594 , n27599 , n27600 );
and ( n27602 , n24011 , n21957 );
and ( n27603 , n23954 , n21955 );
nor ( n27604 , n27602 , n27603 );
xnor ( n27605 , n27604 , n21967 );
and ( n27606 , n27601 , n27605 );
xor ( n27607 , n27402 , n27406 );
xor ( n27608 , n27607 , n27411 );
and ( n27609 , n27605 , n27608 );
and ( n27610 , n27601 , n27608 );
or ( n27611 , n27606 , n27609 , n27610 );
and ( n27612 , n22094 , n22305 );
and ( n27613 , n22080 , n22303 );
nor ( n27614 , n27612 , n27613 );
xnor ( n27615 , n27614 , n22315 );
and ( n27616 , n27611 , n27615 );
xor ( n27617 , n27478 , n27482 );
xor ( n27618 , n27617 , n27485 );
and ( n27619 , n27615 , n27618 );
and ( n27620 , n27611 , n27618 );
or ( n27621 , n27616 , n27619 , n27620 );
and ( n27622 , n22033 , n21735 );
and ( n27623 , n22056 , n21732 );
nor ( n27624 , n27622 , n27623 );
xnor ( n27625 , n27624 , n21730 );
and ( n27626 , n27621 , n27625 );
xor ( n27627 , n27488 , n27492 );
xor ( n27628 , n27627 , n27497 );
and ( n27629 , n27625 , n27628 );
and ( n27630 , n27621 , n27628 );
or ( n27631 , n27626 , n27629 , n27630 );
and ( n27632 , n22659 , n21854 );
and ( n27633 , n22409 , n21852 );
nor ( n27634 , n27632 , n27633 );
xnor ( n27635 , n27634 , n21864 );
and ( n27636 , n23165 , n21779 );
and ( n27637 , n23074 , n21777 );
nor ( n27638 , n27636 , n27637 );
xnor ( n27639 , n27638 , n21789 );
and ( n27640 , n27635 , n27639 );
and ( n27641 , n23446 , n22323 );
and ( n27642 , n23284 , n22321 );
nor ( n27643 , n27641 , n27642 );
xnor ( n27644 , n27643 , n22329 );
and ( n27645 , n27639 , n27644 );
and ( n27646 , n27635 , n27644 );
or ( n27647 , n27640 , n27645 , n27646 );
and ( n27648 , n22080 , n22305 );
and ( n27649 , n22101 , n22303 );
nor ( n27650 , n27648 , n27649 );
xnor ( n27651 , n27650 , n22315 );
and ( n27652 , n27647 , n27651 );
xor ( n27653 , n27504 , n27508 );
xor ( n27654 , n27653 , n27511 );
and ( n27655 , n27651 , n27654 );
and ( n27656 , n27647 , n27654 );
or ( n27657 , n27652 , n27655 , n27656 );
and ( n27658 , n27631 , n27657 );
xor ( n27659 , n27372 , n27376 );
xor ( n27660 , n27659 , n27379 );
and ( n27661 , n27657 , n27660 );
and ( n27662 , n27631 , n27660 );
or ( n27663 , n27658 , n27661 , n27662 );
xor ( n27664 , n27368 , n27382 );
xor ( n27665 , n27664 , n27385 );
and ( n27666 , n27663 , n27665 );
xor ( n27667 , n27251 , n27255 );
xor ( n27668 , n27667 , n27258 );
and ( n27669 , n27665 , n27668 );
and ( n27670 , n27663 , n27668 );
or ( n27671 , n27666 , n27669 , n27670 );
xor ( n27672 , n27388 , n27526 );
xor ( n27673 , n27672 , n27529 );
and ( n27674 , n27671 , n27673 );
xor ( n27675 , n27261 , n27263 );
xor ( n27676 , n27675 , n27266 );
and ( n27677 , n27673 , n27676 );
and ( n27678 , n27671 , n27676 );
or ( n27679 , n27674 , n27677 , n27678 );
and ( n27680 , n27544 , n27679 );
xor ( n27681 , n27544 , n27679 );
xor ( n27682 , n27464 , n27468 );
xor ( n27683 , n27682 , n27471 );
xor ( n27684 , n27631 , n27657 );
xor ( n27685 , n27684 , n27660 );
and ( n27686 , n27683 , n27685 );
xor ( n27687 , n27500 , n27514 );
xor ( n27688 , n27687 , n27517 );
and ( n27689 , n27685 , n27688 );
and ( n27690 , n27683 , n27688 );
or ( n27691 , n27686 , n27689 , n27690 );
xor ( n27692 , n27474 , n27520 );
xor ( n27693 , n27692 , n27523 );
and ( n27694 , n27691 , n27693 );
xor ( n27695 , n27663 , n27665 );
xor ( n27696 , n27695 , n27668 );
and ( n27697 , n27693 , n27696 );
and ( n27698 , n27691 , n27696 );
or ( n27699 , n27694 , n27697 , n27698 );
xor ( n27700 , n27671 , n27673 );
xor ( n27701 , n27700 , n27676 );
and ( n27702 , n27699 , n27701 );
xor ( n27703 , n27699 , n27701 );
xor ( n27704 , n27691 , n27693 );
xor ( n27705 , n27704 , n27696 );
and ( n27706 , n25633 , n21828 );
and ( n27707 , n25427 , n21826 );
nor ( n27708 , n27706 , n27707 );
xnor ( n27709 , n27708 , n21838 );
and ( n27710 , n25833 , n22194 );
and ( n27711 , n25753 , n22192 );
nor ( n27712 , n27710 , n27711 );
xnor ( n27713 , n27712 , n22200 );
and ( n27714 , n27709 , n27713 );
xor ( n27715 , n27569 , n27573 );
xor ( n27716 , n27715 , n27576 );
and ( n27717 , n27713 , n27716 );
and ( n27718 , n27709 , n27716 );
or ( n27719 , n27714 , n27717 , n27718 );
and ( n27720 , n24896 , n21978 );
and ( n27721 , n24753 , n21976 );
nor ( n27722 , n27720 , n27721 );
xnor ( n27723 , n27722 , n21988 );
and ( n27724 , n27719 , n27723 );
and ( n27725 , n25337 , n21804 );
and ( n27726 , n25004 , n21802 );
nor ( n27727 , n27725 , n27726 );
xnor ( n27728 , n27727 , n21814 );
and ( n27729 , n27723 , n27728 );
and ( n27730 , n27719 , n27728 );
or ( n27731 , n27724 , n27729 , n27730 );
and ( n27732 , n24446 , n21957 );
and ( n27733 , n24011 , n21955 );
nor ( n27734 , n27732 , n27733 );
xnor ( n27735 , n27734 , n21967 );
and ( n27736 , n27731 , n27735 );
xor ( n27737 , n27428 , n27432 );
xor ( n27738 , n27737 , n27435 );
and ( n27739 , n27735 , n27738 );
and ( n27740 , n27731 , n27738 );
or ( n27741 , n27736 , n27739 , n27740 );
and ( n27742 , n23284 , n21779 );
and ( n27743 , n23165 , n21777 );
nor ( n27744 , n27742 , n27743 );
xnor ( n27745 , n27744 , n21789 );
and ( n27746 , n27741 , n27745 );
and ( n27747 , n23575 , n22323 );
and ( n27748 , n23446 , n22321 );
nor ( n27749 , n27747 , n27748 );
xnor ( n27750 , n27749 , n22329 );
and ( n27751 , n27745 , n27750 );
and ( n27752 , n27741 , n27750 );
or ( n27753 , n27746 , n27751 , n27752 );
and ( n27754 , n23074 , n21854 );
and ( n27755 , n22659 , n21852 );
nor ( n27756 , n27754 , n27755 );
xnor ( n27757 , n27756 , n21864 );
xor ( n27758 , n27601 , n27605 );
xor ( n27759 , n27758 , n27608 );
and ( n27760 , n27757 , n27759 );
xor ( n27761 , n27438 , n27442 );
xor ( n27762 , n27761 , n27445 );
and ( n27763 , n27759 , n27762 );
and ( n27764 , n27757 , n27762 );
or ( n27765 , n27760 , n27763 , n27764 );
and ( n27766 , n27753 , n27765 );
xor ( n27767 , n27635 , n27639 );
xor ( n27768 , n27767 , n27644 );
and ( n27769 , n27765 , n27768 );
and ( n27770 , n27753 , n27768 );
or ( n27771 , n27766 , n27769 , n27770 );
and ( n27772 , n22049 , n21735 );
and ( n27773 , n22033 , n21732 );
nor ( n27774 , n27772 , n27773 );
xnor ( n27775 , n27774 , n21730 );
and ( n27776 , n22101 , n22252 );
and ( n27777 , n22086 , n22250 );
nor ( n27778 , n27776 , n27777 );
xnor ( n27779 , n27778 , n22258 );
and ( n27780 , n27775 , n27779 );
xor ( n27781 , n27414 , n27448 );
xor ( n27782 , n27781 , n27451 );
and ( n27783 , n27779 , n27782 );
and ( n27784 , n27775 , n27782 );
or ( n27785 , n27780 , n27783 , n27784 );
and ( n27786 , n27771 , n27785 );
xor ( n27787 , n27454 , n27458 );
xor ( n27788 , n27787 , n27461 );
and ( n27789 , n27785 , n27788 );
and ( n27790 , n27771 , n27788 );
or ( n27791 , n27786 , n27789 , n27790 );
and ( n27792 , n22086 , n21735 );
and ( n27793 , n22049 , n21732 );
nor ( n27794 , n27792 , n27793 );
xnor ( n27795 , n27794 , n21730 );
and ( n27796 , n22080 , n22252 );
and ( n27797 , n22101 , n22250 );
nor ( n27798 , n27796 , n27797 );
xnor ( n27799 , n27798 , n22258 );
and ( n27800 , n27795 , n27799 );
and ( n27801 , n22409 , n22305 );
and ( n27802 , n22094 , n22303 );
nor ( n27803 , n27801 , n27802 );
xnor ( n27804 , n27803 , n22315 );
and ( n27805 , n27799 , n27804 );
and ( n27806 , n27795 , n27804 );
or ( n27807 , n27800 , n27805 , n27806 );
and ( n27808 , n25753 , n21828 );
and ( n27809 , n25633 , n21826 );
nor ( n27810 , n27808 , n27809 );
xnor ( n27811 , n27810 , n21838 );
and ( n27812 , n25986 , n22194 );
and ( n27813 , n25833 , n22192 );
nor ( n27814 , n27812 , n27813 );
xnor ( n27815 , n27814 , n22200 );
and ( n27816 , n27811 , n27815 );
xor ( n27817 , n27545 , n27561 );
xor ( n27818 , n27817 , n27566 );
and ( n27819 , n27815 , n27818 );
and ( n27820 , n27811 , n27818 );
or ( n27821 , n27816 , n27819 , n27820 );
and ( n27822 , n25347 , n21804 );
and ( n27823 , n25337 , n21802 );
nor ( n27824 , n27822 , n27823 );
xnor ( n27825 , n27824 , n21814 );
and ( n27826 , n27821 , n27825 );
xor ( n27827 , n27709 , n27713 );
xor ( n27828 , n27827 , n27716 );
and ( n27829 , n27825 , n27828 );
and ( n27830 , n27821 , n27828 );
or ( n27831 , n27826 , n27829 , n27830 );
and ( n27832 , n24544 , n21957 );
and ( n27833 , n24446 , n21955 );
nor ( n27834 , n27832 , n27833 );
xnor ( n27835 , n27834 , n21967 );
and ( n27836 , n27831 , n27835 );
xor ( n27837 , n27579 , n27583 );
xor ( n27838 , n27837 , n27586 );
and ( n27839 , n27835 , n27838 );
and ( n27840 , n27831 , n27838 );
or ( n27841 , n27836 , n27839 , n27840 );
and ( n27842 , n23954 , n22323 );
and ( n27843 , n23575 , n22321 );
nor ( n27844 , n27842 , n27843 );
xnor ( n27845 , n27844 , n22329 );
and ( n27846 , n27841 , n27845 );
xor ( n27847 , n27589 , n27593 );
xor ( n27848 , n27847 , n27598 );
and ( n27849 , n27845 , n27848 );
and ( n27850 , n27841 , n27848 );
or ( n27851 , n27846 , n27849 , n27850 );
and ( n27852 , n23165 , n21854 );
and ( n27853 , n23074 , n21852 );
nor ( n27854 , n27852 , n27853 );
xnor ( n27855 , n27854 , n21864 );
and ( n27856 , n23446 , n21779 );
and ( n27857 , n23284 , n21777 );
nor ( n27858 , n27856 , n27857 );
xnor ( n27859 , n27858 , n21789 );
and ( n27860 , n27855 , n27859 );
xor ( n27861 , n27731 , n27735 );
xor ( n27862 , n27861 , n27738 );
and ( n27863 , n27859 , n27862 );
and ( n27864 , n27855 , n27862 );
or ( n27865 , n27860 , n27863 , n27864 );
and ( n27866 , n27851 , n27865 );
xor ( n27867 , n27741 , n27745 );
xor ( n27868 , n27867 , n27750 );
and ( n27869 , n27865 , n27868 );
and ( n27870 , n27851 , n27868 );
or ( n27871 , n27866 , n27869 , n27870 );
and ( n27872 , n27807 , n27871 );
xor ( n27873 , n27611 , n27615 );
xor ( n27874 , n27873 , n27618 );
and ( n27875 , n27871 , n27874 );
and ( n27876 , n27807 , n27874 );
or ( n27877 , n27872 , n27875 , n27876 );
xor ( n27878 , n27621 , n27625 );
xor ( n27879 , n27878 , n27628 );
and ( n27880 , n27877 , n27879 );
xor ( n27881 , n27647 , n27651 );
xor ( n27882 , n27881 , n27654 );
and ( n27883 , n27879 , n27882 );
and ( n27884 , n27877 , n27882 );
or ( n27885 , n27880 , n27883 , n27884 );
and ( n27886 , n27791 , n27885 );
xor ( n27887 , n27683 , n27685 );
xor ( n27888 , n27887 , n27688 );
and ( n27889 , n27885 , n27888 );
and ( n27890 , n27791 , n27888 );
or ( n27891 , n27886 , n27889 , n27890 );
and ( n27892 , n27705 , n27891 );
xor ( n27893 , n27705 , n27891 );
xor ( n27894 , n27791 , n27885 );
xor ( n27895 , n27894 , n27888 );
xor ( n27896 , n27753 , n27765 );
xor ( n27897 , n27896 , n27768 );
xor ( n27898 , n27775 , n27779 );
xor ( n27899 , n27898 , n27782 );
and ( n27900 , n27897 , n27899 );
xor ( n27901 , n27807 , n27871 );
xor ( n27902 , n27901 , n27874 );
and ( n27903 , n27899 , n27902 );
and ( n27904 , n27897 , n27902 );
or ( n27905 , n27900 , n27903 , n27904 );
xor ( n27906 , n27771 , n27785 );
xor ( n27907 , n27906 , n27788 );
and ( n27908 , n27905 , n27907 );
xor ( n27909 , n27877 , n27879 );
xor ( n27910 , n27909 , n27882 );
and ( n27911 , n27907 , n27910 );
and ( n27912 , n27905 , n27910 );
or ( n27913 , n27908 , n27911 , n27912 );
and ( n27914 , n27895 , n27913 );
xor ( n27915 , n27895 , n27913 );
xor ( n27916 , n27905 , n27907 );
xor ( n27917 , n27916 , n27910 );
xor ( n27918 , n27548 , n27552 );
and ( n27919 , n26360 , n22192 );
not ( n27920 , n27919 );
and ( n27921 , n27920 , n22200 );
and ( n27922 , n26360 , n22194 );
and ( n27923 , n26368 , n22192 );
nor ( n27924 , n27922 , n27923 );
xnor ( n27925 , n27924 , n22200 );
and ( n27926 , n27921 , n27925 );
and ( n27927 , n26368 , n22194 );
and ( n27928 , n26214 , n22192 );
nor ( n27929 , n27927 , n27928 );
xnor ( n27930 , n27929 , n22200 );
and ( n27931 , n27926 , n27930 );
and ( n27932 , n27930 , n27546 );
and ( n27933 , n27926 , n27546 );
or ( n27934 , n27931 , n27932 , n27933 );
and ( n27935 , n27918 , n27934 );
and ( n27936 , n26214 , n22194 );
and ( n27937 , n26107 , n22192 );
nor ( n27938 , n27936 , n27937 );
xnor ( n27939 , n27938 , n22200 );
and ( n27940 , n27934 , n27939 );
and ( n27941 , n27918 , n27939 );
or ( n27942 , n27935 , n27940 , n27941 );
and ( n27943 , n25633 , n21804 );
and ( n27944 , n25427 , n21802 );
nor ( n27945 , n27943 , n27944 );
xnor ( n27946 , n27945 , n21814 );
and ( n27947 , n27942 , n27946 );
and ( n27948 , n25833 , n21828 );
and ( n27949 , n25753 , n21826 );
nor ( n27950 , n27948 , n27949 );
xnor ( n27951 , n27950 , n21838 );
and ( n27952 , n26107 , n22194 );
and ( n27953 , n25986 , n22192 );
nor ( n27954 , n27952 , n27953 );
xnor ( n27955 , n27954 , n22200 );
xor ( n27956 , n27951 , n27955 );
xor ( n27957 , n27553 , n27557 );
xor ( n27958 , n27957 , n27291 );
xor ( n27959 , n27956 , n27958 );
and ( n27960 , n27946 , n27959 );
and ( n27961 , n27942 , n27959 );
or ( n27962 , n27947 , n27960 , n27961 );
and ( n27963 , n25337 , n21978 );
and ( n27964 , n25004 , n21976 );
nor ( n27965 , n27963 , n27964 );
xnor ( n27966 , n27965 , n21988 );
and ( n27967 , n27962 , n27966 );
and ( n27968 , n27951 , n27955 );
and ( n27969 , n27955 , n27958 );
and ( n27970 , n27951 , n27958 );
or ( n27971 , n27968 , n27969 , n27970 );
and ( n27972 , n25427 , n21804 );
and ( n27973 , n25347 , n21802 );
nor ( n27974 , n27972 , n27973 );
xnor ( n27975 , n27974 , n21814 );
xor ( n27976 , n27971 , n27975 );
xor ( n27977 , n27811 , n27815 );
xor ( n27978 , n27977 , n27818 );
xor ( n27979 , n27976 , n27978 );
and ( n27980 , n27966 , n27979 );
and ( n27981 , n27962 , n27979 );
or ( n27982 , n27967 , n27980 , n27981 );
and ( n27983 , n24446 , n22323 );
and ( n27984 , n24011 , n22321 );
nor ( n27985 , n27983 , n27984 );
xnor ( n27986 , n27985 , n22329 );
and ( n27987 , n27982 , n27986 );
xor ( n27988 , n27821 , n27825 );
xor ( n27989 , n27988 , n27828 );
and ( n27990 , n27986 , n27989 );
and ( n27991 , n27982 , n27989 );
or ( n27992 , n27987 , n27990 , n27991 );
and ( n27993 , n23284 , n21854 );
and ( n27994 , n23165 , n21852 );
nor ( n27995 , n27993 , n27994 );
xnor ( n27996 , n27995 , n21864 );
and ( n27997 , n27992 , n27996 );
and ( n27998 , n23575 , n21779 );
and ( n27999 , n23446 , n21777 );
nor ( n28000 , n27998 , n27999 );
xnor ( n28001 , n28000 , n21789 );
and ( n28002 , n27996 , n28001 );
and ( n28003 , n27992 , n28001 );
or ( n28004 , n27997 , n28002 , n28003 );
and ( n28005 , n23165 , n22305 );
and ( n28006 , n23074 , n22303 );
nor ( n28007 , n28005 , n28006 );
xnor ( n28008 , n28007 , n22315 );
and ( n28009 , n23954 , n21779 );
and ( n28010 , n23575 , n21777 );
nor ( n28011 , n28009 , n28010 );
xnor ( n28012 , n28011 , n21789 );
and ( n28013 , n28008 , n28012 );
and ( n28014 , n27971 , n27975 );
and ( n28015 , n27975 , n27978 );
and ( n28016 , n27971 , n27978 );
or ( n28017 , n28014 , n28015 , n28016 );
and ( n28018 , n24753 , n21957 );
and ( n28019 , n24544 , n21955 );
nor ( n28020 , n28018 , n28019 );
xnor ( n28021 , n28020 , n21967 );
xor ( n28022 , n28017 , n28021 );
and ( n28023 , n25004 , n21978 );
and ( n28024 , n24896 , n21976 );
nor ( n28025 , n28023 , n28024 );
xnor ( n28026 , n28025 , n21988 );
xor ( n28027 , n28022 , n28026 );
and ( n28028 , n28012 , n28027 );
and ( n28029 , n28008 , n28027 );
or ( n28030 , n28013 , n28028 , n28029 );
and ( n28031 , n22080 , n21735 );
and ( n28032 , n22101 , n21732 );
nor ( n28033 , n28031 , n28032 );
xnor ( n28034 , n28033 , n21730 );
and ( n28035 , n28030 , n28034 );
and ( n28036 , n28017 , n28021 );
and ( n28037 , n28021 , n28026 );
and ( n28038 , n28017 , n28026 );
or ( n28039 , n28036 , n28037 , n28038 );
and ( n28040 , n24011 , n22323 );
and ( n28041 , n23954 , n22321 );
nor ( n28042 , n28040 , n28041 );
xnor ( n28043 , n28042 , n22329 );
xor ( n28044 , n28039 , n28043 );
xor ( n28045 , n27719 , n27723 );
xor ( n28046 , n28045 , n27728 );
xor ( n28047 , n28044 , n28046 );
and ( n28048 , n28034 , n28047 );
and ( n28049 , n28030 , n28047 );
or ( n28050 , n28035 , n28048 , n28049 );
and ( n28051 , n28004 , n28050 );
and ( n28052 , n22409 , n22252 );
and ( n28053 , n22094 , n22250 );
nor ( n28054 , n28052 , n28053 );
xnor ( n28055 , n28054 , n22258 );
and ( n28056 , n23074 , n22305 );
and ( n28057 , n22659 , n22303 );
nor ( n28058 , n28056 , n28057 );
xnor ( n28059 , n28058 , n22315 );
and ( n28060 , n28055 , n28059 );
xor ( n28061 , n27831 , n27835 );
xor ( n28062 , n28061 , n27838 );
and ( n28063 , n28059 , n28062 );
and ( n28064 , n28055 , n28062 );
or ( n28065 , n28060 , n28063 , n28064 );
and ( n28066 , n28050 , n28065 );
and ( n28067 , n28004 , n28065 );
or ( n28068 , n28051 , n28066 , n28067 );
and ( n28069 , n22101 , n21735 );
and ( n28070 , n22086 , n21732 );
nor ( n28071 , n28069 , n28070 );
xnor ( n28072 , n28071 , n21730 );
xor ( n28073 , n27841 , n27845 );
xor ( n28074 , n28073 , n27848 );
and ( n28075 , n28072 , n28074 );
xor ( n28076 , n27855 , n27859 );
xor ( n28077 , n28076 , n27862 );
and ( n28078 , n28074 , n28077 );
and ( n28079 , n28072 , n28077 );
or ( n28080 , n28075 , n28078 , n28079 );
and ( n28081 , n28068 , n28080 );
xor ( n28082 , n27851 , n27865 );
xor ( n28083 , n28082 , n27868 );
and ( n28084 , n28080 , n28083 );
and ( n28085 , n28068 , n28083 );
or ( n28086 , n28081 , n28084 , n28085 );
and ( n28087 , n28039 , n28043 );
and ( n28088 , n28043 , n28046 );
and ( n28089 , n28039 , n28046 );
or ( n28090 , n28087 , n28088 , n28089 );
and ( n28091 , n22094 , n22252 );
and ( n28092 , n22080 , n22250 );
nor ( n28093 , n28091 , n28092 );
xnor ( n28094 , n28093 , n22258 );
and ( n28095 , n28090 , n28094 );
and ( n28096 , n22659 , n22305 );
and ( n28097 , n22409 , n22303 );
nor ( n28098 , n28096 , n28097 );
xnor ( n28099 , n28098 , n22315 );
and ( n28100 , n28094 , n28099 );
and ( n28101 , n28090 , n28099 );
or ( n28102 , n28095 , n28100 , n28101 );
xor ( n28103 , n27795 , n27799 );
xor ( n28104 , n28103 , n27804 );
and ( n28105 , n28102 , n28104 );
xor ( n28106 , n27757 , n27759 );
xor ( n28107 , n28106 , n27762 );
and ( n28108 , n28104 , n28107 );
and ( n28109 , n28102 , n28107 );
or ( n28110 , n28105 , n28108 , n28109 );
and ( n28111 , n28086 , n28110 );
xor ( n28112 , n27897 , n27899 );
xor ( n28113 , n28112 , n27902 );
and ( n28114 , n28110 , n28113 );
and ( n28115 , n28086 , n28113 );
or ( n28116 , n28111 , n28114 , n28115 );
and ( n28117 , n27917 , n28116 );
xor ( n28118 , n27917 , n28116 );
and ( n28119 , n25753 , n21804 );
and ( n28120 , n25633 , n21802 );
nor ( n28121 , n28119 , n28120 );
xnor ( n28122 , n28121 , n21814 );
and ( n28123 , n25986 , n21828 );
and ( n28124 , n25833 , n21826 );
nor ( n28125 , n28123 , n28124 );
xnor ( n28126 , n28125 , n21838 );
and ( n28127 , n28122 , n28126 );
xor ( n28128 , n27918 , n27934 );
xor ( n28129 , n28128 , n27939 );
and ( n28130 , n28126 , n28129 );
and ( n28131 , n28122 , n28129 );
or ( n28132 , n28127 , n28130 , n28131 );
and ( n28133 , n25347 , n21978 );
and ( n28134 , n25337 , n21976 );
nor ( n28135 , n28133 , n28134 );
xnor ( n28136 , n28135 , n21988 );
and ( n28137 , n28132 , n28136 );
xor ( n28138 , n27942 , n27946 );
xor ( n28139 , n28138 , n27959 );
and ( n28140 , n28136 , n28139 );
and ( n28141 , n28132 , n28139 );
or ( n28142 , n28137 , n28140 , n28141 );
and ( n28143 , n24544 , n22323 );
and ( n28144 , n24446 , n22321 );
nor ( n28145 , n28143 , n28144 );
xnor ( n28146 , n28145 , n22329 );
and ( n28147 , n28142 , n28146 );
and ( n28148 , n24896 , n21957 );
and ( n28149 , n24753 , n21955 );
nor ( n28150 , n28148 , n28149 );
xnor ( n28151 , n28150 , n21967 );
and ( n28152 , n28146 , n28151 );
and ( n28153 , n28142 , n28151 );
or ( n28154 , n28147 , n28152 , n28153 );
and ( n28155 , n22659 , n22252 );
and ( n28156 , n22409 , n22250 );
nor ( n28157 , n28155 , n28156 );
xnor ( n28158 , n28157 , n22258 );
and ( n28159 , n28154 , n28158 );
and ( n28160 , n23446 , n21854 );
and ( n28161 , n23284 , n21852 );
nor ( n28162 , n28160 , n28161 );
xnor ( n28163 , n28162 , n21864 );
and ( n28164 , n28158 , n28163 );
and ( n28165 , n28154 , n28163 );
or ( n28166 , n28159 , n28164 , n28165 );
xor ( n28167 , n27992 , n27996 );
xor ( n28168 , n28167 , n28001 );
and ( n28169 , n28166 , n28168 );
xor ( n28170 , n28055 , n28059 );
xor ( n28171 , n28170 , n28062 );
and ( n28172 , n28168 , n28171 );
and ( n28173 , n28166 , n28171 );
or ( n28174 , n28169 , n28172 , n28173 );
xor ( n28175 , n28090 , n28094 );
xor ( n28176 , n28175 , n28099 );
and ( n28177 , n28174 , n28176 );
xor ( n28178 , n28072 , n28074 );
xor ( n28179 , n28178 , n28077 );
and ( n28180 , n28176 , n28179 );
and ( n28181 , n28174 , n28179 );
or ( n28182 , n28177 , n28180 , n28181 );
xor ( n28183 , n28068 , n28080 );
xor ( n28184 , n28183 , n28083 );
and ( n28185 , n28182 , n28184 );
xor ( n28186 , n28102 , n28104 );
xor ( n28187 , n28186 , n28107 );
and ( n28188 , n28184 , n28187 );
and ( n28189 , n28182 , n28187 );
or ( n28190 , n28185 , n28188 , n28189 );
xor ( n28191 , n28086 , n28110 );
xor ( n28192 , n28191 , n28113 );
and ( n28193 , n28190 , n28192 );
xor ( n28194 , n28190 , n28192 );
xor ( n28195 , n28182 , n28184 );
xor ( n28196 , n28195 , n28187 );
and ( n28197 , n23954 , n21854 );
and ( n28198 , n23575 , n21852 );
nor ( n28199 , n28197 , n28198 );
xnor ( n28200 , n28199 , n21864 );
and ( n28201 , n24446 , n21779 );
and ( n28202 , n24011 , n21777 );
nor ( n28203 , n28201 , n28202 );
xnor ( n28204 , n28203 , n21789 );
and ( n28205 , n28200 , n28204 );
xor ( n28206 , n28132 , n28136 );
xor ( n28207 , n28206 , n28139 );
and ( n28208 , n28204 , n28207 );
and ( n28209 , n28200 , n28207 );
or ( n28210 , n28205 , n28208 , n28209 );
and ( n28211 , n23284 , n22305 );
and ( n28212 , n23165 , n22303 );
nor ( n28213 , n28211 , n28212 );
xnor ( n28214 , n28213 , n22315 );
and ( n28215 , n28210 , n28214 );
and ( n28216 , n23575 , n21854 );
and ( n28217 , n23446 , n21852 );
nor ( n28218 , n28216 , n28217 );
xnor ( n28219 , n28218 , n21864 );
and ( n28220 , n28214 , n28219 );
and ( n28221 , n28210 , n28219 );
or ( n28222 , n28215 , n28220 , n28221 );
xor ( n28223 , n28154 , n28158 );
xor ( n28224 , n28223 , n28163 );
and ( n28225 , n28222 , n28224 );
xor ( n28226 , n28008 , n28012 );
xor ( n28227 , n28226 , n28027 );
and ( n28228 , n28224 , n28227 );
and ( n28229 , n28222 , n28227 );
or ( n28230 , n28225 , n28228 , n28229 );
and ( n28231 , n25833 , n21804 );
and ( n28232 , n25753 , n21802 );
nor ( n28233 , n28231 , n28232 );
xnor ( n28234 , n28233 , n21814 );
and ( n28235 , n26107 , n21828 );
and ( n28236 , n25986 , n21826 );
nor ( n28237 , n28235 , n28236 );
xnor ( n28238 , n28237 , n21838 );
and ( n28239 , n28234 , n28238 );
xor ( n28240 , n27926 , n27930 );
xor ( n28241 , n28240 , n27546 );
and ( n28242 , n28238 , n28241 );
and ( n28243 , n28234 , n28241 );
or ( n28244 , n28239 , n28242 , n28243 );
and ( n28245 , n25427 , n21978 );
and ( n28246 , n25347 , n21976 );
nor ( n28247 , n28245 , n28246 );
xnor ( n28248 , n28247 , n21988 );
and ( n28249 , n28244 , n28248 );
xor ( n28250 , n28122 , n28126 );
xor ( n28251 , n28250 , n28129 );
and ( n28252 , n28248 , n28251 );
and ( n28253 , n28244 , n28251 );
or ( n28254 , n28249 , n28252 , n28253 );
and ( n28255 , n24753 , n22323 );
and ( n28256 , n24544 , n22321 );
nor ( n28257 , n28255 , n28256 );
xnor ( n28258 , n28257 , n22329 );
and ( n28259 , n28254 , n28258 );
and ( n28260 , n25004 , n21957 );
and ( n28261 , n24896 , n21955 );
nor ( n28262 , n28260 , n28261 );
xnor ( n28263 , n28262 , n21967 );
and ( n28264 , n28258 , n28263 );
and ( n28265 , n28254 , n28263 );
or ( n28266 , n28259 , n28264 , n28265 );
and ( n28267 , n24011 , n21779 );
and ( n28268 , n23954 , n21777 );
nor ( n28269 , n28267 , n28268 );
xnor ( n28270 , n28269 , n21789 );
and ( n28271 , n28266 , n28270 );
xor ( n28272 , n27962 , n27966 );
xor ( n28273 , n28272 , n27979 );
and ( n28274 , n28270 , n28273 );
and ( n28275 , n28266 , n28273 );
or ( n28276 , n28271 , n28274 , n28275 );
and ( n28277 , n22094 , n21735 );
and ( n28278 , n22080 , n21732 );
nor ( n28279 , n28277 , n28278 );
xnor ( n28280 , n28279 , n21730 );
and ( n28281 , n28276 , n28280 );
xor ( n28282 , n27982 , n27986 );
xor ( n28283 , n28282 , n27989 );
and ( n28284 , n28280 , n28283 );
and ( n28285 , n28276 , n28283 );
or ( n28286 , n28281 , n28284 , n28285 );
and ( n28287 , n28230 , n28286 );
xor ( n28288 , n28030 , n28034 );
xor ( n28289 , n28288 , n28047 );
and ( n28290 , n28286 , n28289 );
and ( n28291 , n28230 , n28289 );
or ( n28292 , n28287 , n28290 , n28291 );
xor ( n28293 , n28004 , n28050 );
xor ( n28294 , n28293 , n28065 );
and ( n28295 , n28292 , n28294 );
xor ( n28296 , n28174 , n28176 );
xor ( n28297 , n28296 , n28179 );
and ( n28298 , n28294 , n28297 );
and ( n28299 , n28292 , n28297 );
or ( n28300 , n28295 , n28298 , n28299 );
and ( n28301 , n28196 , n28300 );
xor ( n28302 , n28196 , n28300 );
and ( n28303 , n22409 , n21735 );
and ( n28304 , n22094 , n21732 );
nor ( n28305 , n28303 , n28304 );
xnor ( n28306 , n28305 , n21730 );
and ( n28307 , n23074 , n22252 );
and ( n28308 , n22659 , n22250 );
nor ( n28309 , n28307 , n28308 );
xnor ( n28310 , n28309 , n22258 );
and ( n28311 , n28306 , n28310 );
xor ( n28312 , n28142 , n28146 );
xor ( n28313 , n28312 , n28151 );
and ( n28314 , n28310 , n28313 );
and ( n28315 , n28306 , n28313 );
or ( n28316 , n28311 , n28314 , n28315 );
and ( n28317 , n22659 , n21735 );
and ( n28318 , n22409 , n21732 );
nor ( n28319 , n28317 , n28318 );
xnor ( n28320 , n28319 , n21730 );
and ( n28321 , n23165 , n22252 );
and ( n28322 , n23074 , n22250 );
nor ( n28323 , n28321 , n28322 );
xnor ( n28324 , n28323 , n22258 );
and ( n28325 , n28320 , n28324 );
and ( n28326 , n23446 , n22305 );
and ( n28327 , n23284 , n22303 );
nor ( n28328 , n28326 , n28327 );
xnor ( n28329 , n28328 , n22315 );
and ( n28330 , n28324 , n28329 );
and ( n28331 , n28320 , n28329 );
or ( n28332 , n28325 , n28330 , n28331 );
and ( n28333 , n25753 , n21978 );
and ( n28334 , n25633 , n21976 );
nor ( n28335 , n28333 , n28334 );
xnor ( n28336 , n28335 , n21988 );
and ( n28337 , n25986 , n21804 );
and ( n28338 , n25833 , n21802 );
nor ( n28339 , n28337 , n28338 );
xnor ( n28340 , n28339 , n21814 );
and ( n28341 , n28336 , n28340 );
xor ( n28342 , n27921 , n27925 );
and ( n28343 , n26360 , n21826 );
not ( n28344 , n28343 );
and ( n28345 , n28344 , n21838 );
and ( n28346 , n26360 , n21828 );
and ( n28347 , n26368 , n21826 );
nor ( n28348 , n28346 , n28347 );
xnor ( n28349 , n28348 , n21838 );
and ( n28350 , n28345 , n28349 );
and ( n28351 , n26368 , n21828 );
and ( n28352 , n26214 , n21826 );
nor ( n28353 , n28351 , n28352 );
xnor ( n28354 , n28353 , n21838 );
and ( n28355 , n28350 , n28354 );
and ( n28356 , n28354 , n27919 );
and ( n28357 , n28350 , n27919 );
or ( n28358 , n28355 , n28356 , n28357 );
xor ( n28359 , n28342 , n28358 );
and ( n28360 , n26214 , n21828 );
and ( n28361 , n26107 , n21826 );
nor ( n28362 , n28360 , n28361 );
xnor ( n28363 , n28362 , n21838 );
xor ( n28364 , n28359 , n28363 );
and ( n28365 , n28340 , n28364 );
and ( n28366 , n28336 , n28364 );
or ( n28367 , n28341 , n28365 , n28366 );
and ( n28368 , n25347 , n21957 );
and ( n28369 , n25337 , n21955 );
nor ( n28370 , n28368 , n28369 );
xnor ( n28371 , n28370 , n21967 );
and ( n28372 , n28367 , n28371 );
and ( n28373 , n28342 , n28358 );
and ( n28374 , n28358 , n28363 );
and ( n28375 , n28342 , n28363 );
or ( n28376 , n28373 , n28374 , n28375 );
and ( n28377 , n25633 , n21978 );
and ( n28378 , n25427 , n21976 );
nor ( n28379 , n28377 , n28378 );
xnor ( n28380 , n28379 , n21988 );
xor ( n28381 , n28376 , n28380 );
xor ( n28382 , n28234 , n28238 );
xor ( n28383 , n28382 , n28241 );
xor ( n28384 , n28381 , n28383 );
and ( n28385 , n28371 , n28384 );
and ( n28386 , n28367 , n28384 );
or ( n28387 , n28372 , n28385 , n28386 );
and ( n28388 , n24544 , n21779 );
and ( n28389 , n24446 , n21777 );
nor ( n28390 , n28388 , n28389 );
xnor ( n28391 , n28390 , n21789 );
and ( n28392 , n28387 , n28391 );
and ( n28393 , n25337 , n21957 );
and ( n28394 , n25004 , n21955 );
nor ( n28395 , n28393 , n28394 );
xnor ( n28396 , n28395 , n21967 );
and ( n28397 , n28391 , n28396 );
and ( n28398 , n28387 , n28396 );
or ( n28399 , n28392 , n28397 , n28398 );
and ( n28400 , n28376 , n28380 );
and ( n28401 , n28380 , n28383 );
and ( n28402 , n28376 , n28383 );
or ( n28403 , n28400 , n28401 , n28402 );
and ( n28404 , n24896 , n22323 );
and ( n28405 , n24753 , n22321 );
nor ( n28406 , n28404 , n28405 );
xnor ( n28407 , n28406 , n22329 );
and ( n28408 , n28403 , n28407 );
xor ( n28409 , n28244 , n28248 );
xor ( n28410 , n28409 , n28251 );
and ( n28411 , n28407 , n28410 );
and ( n28412 , n28403 , n28410 );
or ( n28413 , n28408 , n28411 , n28412 );
and ( n28414 , n28399 , n28413 );
xor ( n28415 , n28254 , n28258 );
xor ( n28416 , n28415 , n28263 );
and ( n28417 , n28413 , n28416 );
and ( n28418 , n28399 , n28416 );
or ( n28419 , n28414 , n28417 , n28418 );
and ( n28420 , n28332 , n28419 );
xor ( n28421 , n28266 , n28270 );
xor ( n28422 , n28421 , n28273 );
and ( n28423 , n28419 , n28422 );
and ( n28424 , n28332 , n28422 );
or ( n28425 , n28420 , n28423 , n28424 );
and ( n28426 , n28316 , n28425 );
xor ( n28427 , n28276 , n28280 );
xor ( n28428 , n28427 , n28283 );
and ( n28429 , n28425 , n28428 );
and ( n28430 , n28316 , n28428 );
or ( n28431 , n28426 , n28429 , n28430 );
xor ( n28432 , n28230 , n28286 );
xor ( n28433 , n28432 , n28289 );
and ( n28434 , n28431 , n28433 );
xor ( n28435 , n28166 , n28168 );
xor ( n28436 , n28435 , n28171 );
and ( n28437 , n28433 , n28436 );
and ( n28438 , n28431 , n28436 );
or ( n28439 , n28434 , n28437 , n28438 );
xor ( n28440 , n28292 , n28294 );
xor ( n28441 , n28440 , n28297 );
and ( n28442 , n28439 , n28441 );
xor ( n28443 , n28439 , n28441 );
xor ( n28444 , n28431 , n28433 );
xor ( n28445 , n28444 , n28436 );
and ( n28446 , n25833 , n21978 );
and ( n28447 , n25753 , n21976 );
nor ( n28448 , n28446 , n28447 );
xnor ( n28449 , n28448 , n21988 );
and ( n28450 , n26107 , n21804 );
and ( n28451 , n25986 , n21802 );
nor ( n28452 , n28450 , n28451 );
xnor ( n28453 , n28452 , n21814 );
and ( n28454 , n28449 , n28453 );
xor ( n28455 , n28350 , n28354 );
xor ( n28456 , n28455 , n27919 );
and ( n28457 , n28453 , n28456 );
and ( n28458 , n28449 , n28456 );
or ( n28459 , n28454 , n28457 , n28458 );
and ( n28460 , n25427 , n21957 );
and ( n28461 , n25347 , n21955 );
nor ( n28462 , n28460 , n28461 );
xnor ( n28463 , n28462 , n21967 );
and ( n28464 , n28459 , n28463 );
xor ( n28465 , n28336 , n28340 );
xor ( n28466 , n28465 , n28364 );
and ( n28467 , n28463 , n28466 );
and ( n28468 , n28459 , n28466 );
or ( n28469 , n28464 , n28467 , n28468 );
and ( n28470 , n24753 , n21779 );
and ( n28471 , n24544 , n21777 );
nor ( n28472 , n28470 , n28471 );
xnor ( n28473 , n28472 , n21789 );
and ( n28474 , n28469 , n28473 );
and ( n28475 , n25004 , n22323 );
and ( n28476 , n24896 , n22321 );
nor ( n28477 , n28475 , n28476 );
xnor ( n28478 , n28477 , n22329 );
and ( n28479 , n28473 , n28478 );
and ( n28480 , n28469 , n28478 );
or ( n28481 , n28474 , n28479 , n28480 );
and ( n28482 , n24011 , n21854 );
and ( n28483 , n23954 , n21852 );
nor ( n28484 , n28482 , n28483 );
xnor ( n28485 , n28484 , n21864 );
and ( n28486 , n28481 , n28485 );
xor ( n28487 , n28403 , n28407 );
xor ( n28488 , n28487 , n28410 );
and ( n28489 , n28485 , n28488 );
and ( n28490 , n28481 , n28488 );
or ( n28491 , n28486 , n28489 , n28490 );
xor ( n28492 , n28399 , n28413 );
xor ( n28493 , n28492 , n28416 );
and ( n28494 , n28491 , n28493 );
xor ( n28495 , n28200 , n28204 );
xor ( n28496 , n28495 , n28207 );
and ( n28497 , n28493 , n28496 );
and ( n28498 , n28491 , n28496 );
or ( n28499 , n28494 , n28497 , n28498 );
xor ( n28500 , n28210 , n28214 );
xor ( n28501 , n28500 , n28219 );
and ( n28502 , n28499 , n28501 );
xor ( n28503 , n28306 , n28310 );
xor ( n28504 , n28503 , n28313 );
and ( n28505 , n28501 , n28504 );
and ( n28506 , n28499 , n28504 );
or ( n28507 , n28502 , n28505 , n28506 );
xor ( n28508 , n28222 , n28224 );
xor ( n28509 , n28508 , n28227 );
and ( n28510 , n28507 , n28509 );
xor ( n28511 , n28316 , n28425 );
xor ( n28512 , n28511 , n28428 );
and ( n28513 , n28509 , n28512 );
and ( n28514 , n28507 , n28512 );
or ( n28515 , n28510 , n28513 , n28514 );
and ( n28516 , n28445 , n28515 );
xor ( n28517 , n28445 , n28515 );
xor ( n28518 , n28507 , n28509 );
xor ( n28519 , n28518 , n28512 );
and ( n28520 , n23074 , n21735 );
and ( n28521 , n22659 , n21732 );
nor ( n28522 , n28520 , n28521 );
xnor ( n28523 , n28522 , n21730 );
and ( n28524 , n23284 , n22252 );
and ( n28525 , n23165 , n22250 );
nor ( n28526 , n28524 , n28525 );
xnor ( n28527 , n28526 , n22258 );
and ( n28528 , n28523 , n28527 );
and ( n28529 , n23575 , n22305 );
and ( n28530 , n23446 , n22303 );
nor ( n28531 , n28529 , n28530 );
xnor ( n28532 , n28531 , n22315 );
and ( n28533 , n28527 , n28532 );
and ( n28534 , n28523 , n28532 );
or ( n28535 , n28528 , n28533 , n28534 );
xor ( n28536 , n28345 , n28349 );
and ( n28537 , n26360 , n21802 );
not ( n28538 , n28537 );
and ( n28539 , n28538 , n21814 );
and ( n28540 , n26360 , n21804 );
and ( n28541 , n26368 , n21802 );
nor ( n28542 , n28540 , n28541 );
xnor ( n28543 , n28542 , n21814 );
and ( n28544 , n28539 , n28543 );
and ( n28545 , n26368 , n21804 );
and ( n28546 , n26214 , n21802 );
nor ( n28547 , n28545 , n28546 );
xnor ( n28548 , n28547 , n21814 );
and ( n28549 , n28544 , n28548 );
and ( n28550 , n28548 , n28343 );
and ( n28551 , n28544 , n28343 );
or ( n28552 , n28549 , n28550 , n28551 );
and ( n28553 , n28536 , n28552 );
and ( n28554 , n26214 , n21804 );
and ( n28555 , n26107 , n21802 );
nor ( n28556 , n28554 , n28555 );
xnor ( n28557 , n28556 , n21814 );
and ( n28558 , n28552 , n28557 );
and ( n28559 , n28536 , n28557 );
or ( n28560 , n28553 , n28558 , n28559 );
and ( n28561 , n25633 , n21957 );
and ( n28562 , n25427 , n21955 );
nor ( n28563 , n28561 , n28562 );
xnor ( n28564 , n28563 , n21967 );
and ( n28565 , n28560 , n28564 );
xor ( n28566 , n28449 , n28453 );
xor ( n28567 , n28566 , n28456 );
and ( n28568 , n28564 , n28567 );
and ( n28569 , n28560 , n28567 );
or ( n28570 , n28565 , n28568 , n28569 );
and ( n28571 , n24896 , n21779 );
and ( n28572 , n24753 , n21777 );
nor ( n28573 , n28571 , n28572 );
xnor ( n28574 , n28573 , n21789 );
and ( n28575 , n28570 , n28574 );
xor ( n28576 , n28459 , n28463 );
xor ( n28577 , n28576 , n28466 );
and ( n28578 , n28574 , n28577 );
and ( n28579 , n28570 , n28577 );
or ( n28580 , n28575 , n28578 , n28579 );
and ( n28581 , n24446 , n21854 );
and ( n28582 , n24011 , n21852 );
nor ( n28583 , n28581 , n28582 );
xnor ( n28584 , n28583 , n21864 );
and ( n28585 , n28580 , n28584 );
xor ( n28586 , n28367 , n28371 );
xor ( n28587 , n28586 , n28384 );
and ( n28588 , n28584 , n28587 );
and ( n28589 , n28580 , n28587 );
or ( n28590 , n28585 , n28588 , n28589 );
xor ( n28591 , n28387 , n28391 );
xor ( n28592 , n28591 , n28396 );
and ( n28593 , n28590 , n28592 );
xor ( n28594 , n28481 , n28485 );
xor ( n28595 , n28594 , n28488 );
and ( n28596 , n28592 , n28595 );
and ( n28597 , n28590 , n28595 );
or ( n28598 , n28593 , n28596 , n28597 );
and ( n28599 , n28535 , n28598 );
xor ( n28600 , n28320 , n28324 );
xor ( n28601 , n28600 , n28329 );
and ( n28602 , n28598 , n28601 );
and ( n28603 , n28535 , n28601 );
or ( n28604 , n28599 , n28602 , n28603 );
xor ( n28605 , n28499 , n28501 );
xor ( n28606 , n28605 , n28504 );
and ( n28607 , n28604 , n28606 );
xor ( n28608 , n28332 , n28419 );
xor ( n28609 , n28608 , n28422 );
and ( n28610 , n28606 , n28609 );
and ( n28611 , n28604 , n28609 );
or ( n28612 , n28607 , n28610 , n28611 );
and ( n28613 , n28519 , n28612 );
xor ( n28614 , n28519 , n28612 );
xor ( n28615 , n28604 , n28606 );
xor ( n28616 , n28615 , n28609 );
and ( n28617 , n23165 , n21735 );
and ( n28618 , n23074 , n21732 );
nor ( n28619 , n28617 , n28618 );
xnor ( n28620 , n28619 , n21730 );
and ( n28621 , n23954 , n22305 );
and ( n28622 , n23575 , n22303 );
nor ( n28623 , n28621 , n28622 );
xnor ( n28624 , n28623 , n22315 );
and ( n28625 , n28620 , n28624 );
xor ( n28626 , n28469 , n28473 );
xor ( n28627 , n28626 , n28478 );
and ( n28628 , n28624 , n28627 );
and ( n28629 , n28620 , n28627 );
or ( n28630 , n28625 , n28628 , n28629 );
and ( n28631 , n25753 , n21957 );
and ( n28632 , n25633 , n21955 );
nor ( n28633 , n28631 , n28632 );
xnor ( n28634 , n28633 , n21967 );
and ( n28635 , n25986 , n21978 );
and ( n28636 , n25833 , n21976 );
nor ( n28637 , n28635 , n28636 );
xnor ( n28638 , n28637 , n21988 );
and ( n28639 , n28634 , n28638 );
xor ( n28640 , n28536 , n28552 );
xor ( n28641 , n28640 , n28557 );
and ( n28642 , n28638 , n28641 );
and ( n28643 , n28634 , n28641 );
or ( n28644 , n28639 , n28642 , n28643 );
and ( n28645 , n25347 , n22323 );
and ( n28646 , n25337 , n22321 );
nor ( n28647 , n28645 , n28646 );
xnor ( n28648 , n28647 , n22329 );
and ( n28649 , n28644 , n28648 );
xor ( n28650 , n28560 , n28564 );
xor ( n28651 , n28650 , n28567 );
and ( n28652 , n28648 , n28651 );
and ( n28653 , n28644 , n28651 );
or ( n28654 , n28649 , n28652 , n28653 );
and ( n28655 , n24544 , n21854 );
and ( n28656 , n24446 , n21852 );
nor ( n28657 , n28655 , n28656 );
xnor ( n28658 , n28657 , n21864 );
and ( n28659 , n28654 , n28658 );
and ( n28660 , n25337 , n22323 );
and ( n28661 , n25004 , n22321 );
nor ( n28662 , n28660 , n28661 );
xnor ( n28663 , n28662 , n22329 );
and ( n28664 , n28658 , n28663 );
and ( n28665 , n28654 , n28663 );
or ( n28666 , n28659 , n28664 , n28665 );
and ( n28667 , n23446 , n22252 );
and ( n28668 , n23284 , n22250 );
nor ( n28669 , n28667 , n28668 );
xnor ( n28670 , n28669 , n22258 );
and ( n28671 , n28666 , n28670 );
xor ( n28672 , n28580 , n28584 );
xor ( n28673 , n28672 , n28587 );
and ( n28674 , n28670 , n28673 );
and ( n28675 , n28666 , n28673 );
or ( n28676 , n28671 , n28674 , n28675 );
and ( n28677 , n28630 , n28676 );
xor ( n28678 , n28523 , n28527 );
xor ( n28679 , n28678 , n28532 );
and ( n28680 , n28676 , n28679 );
and ( n28681 , n28630 , n28679 );
or ( n28682 , n28677 , n28680 , n28681 );
xor ( n28683 , n28535 , n28598 );
xor ( n28684 , n28683 , n28601 );
and ( n28685 , n28682 , n28684 );
xor ( n28686 , n28491 , n28493 );
xor ( n28687 , n28686 , n28496 );
and ( n28688 , n28684 , n28687 );
and ( n28689 , n28682 , n28687 );
or ( n28690 , n28685 , n28688 , n28689 );
and ( n28691 , n28616 , n28690 );
xor ( n28692 , n28616 , n28690 );
xor ( n28693 , n28682 , n28684 );
xor ( n28694 , n28693 , n28687 );
and ( n28695 , n25833 , n21957 );
and ( n28696 , n25753 , n21955 );
nor ( n28697 , n28695 , n28696 );
xnor ( n28698 , n28697 , n21967 );
and ( n28699 , n26107 , n21978 );
and ( n28700 , n25986 , n21976 );
nor ( n28701 , n28699 , n28700 );
xnor ( n28702 , n28701 , n21988 );
and ( n28703 , n28698 , n28702 );
xor ( n28704 , n28544 , n28548 );
xor ( n28705 , n28704 , n28343 );
and ( n28706 , n28702 , n28705 );
and ( n28707 , n28698 , n28705 );
or ( n28708 , n28703 , n28706 , n28707 );
and ( n28709 , n25427 , n22323 );
and ( n28710 , n25347 , n22321 );
nor ( n28711 , n28709 , n28710 );
xnor ( n28712 , n28711 , n22329 );
and ( n28713 , n28708 , n28712 );
xor ( n28714 , n28634 , n28638 );
xor ( n28715 , n28714 , n28641 );
and ( n28716 , n28712 , n28715 );
and ( n28717 , n28708 , n28715 );
or ( n28718 , n28713 , n28716 , n28717 );
and ( n28719 , n24753 , n21854 );
and ( n28720 , n24544 , n21852 );
nor ( n28721 , n28719 , n28720 );
xnor ( n28722 , n28721 , n21864 );
and ( n28723 , n28718 , n28722 );
and ( n28724 , n25004 , n21779 );
and ( n28725 , n24896 , n21777 );
nor ( n28726 , n28724 , n28725 );
xnor ( n28727 , n28726 , n21789 );
and ( n28728 , n28722 , n28727 );
and ( n28729 , n28718 , n28727 );
or ( n28730 , n28723 , n28728 , n28729 );
and ( n28731 , n24011 , n22305 );
and ( n28732 , n23954 , n22303 );
nor ( n28733 , n28731 , n28732 );
xnor ( n28734 , n28733 , n22315 );
and ( n28735 , n28730 , n28734 );
xor ( n28736 , n28570 , n28574 );
xor ( n28737 , n28736 , n28577 );
and ( n28738 , n28734 , n28737 );
and ( n28739 , n28730 , n28737 );
or ( n28740 , n28735 , n28738 , n28739 );
xor ( n28741 , n28620 , n28624 );
xor ( n28742 , n28741 , n28627 );
and ( n28743 , n28740 , n28742 );
xor ( n28744 , n28666 , n28670 );
xor ( n28745 , n28744 , n28673 );
and ( n28746 , n28742 , n28745 );
and ( n28747 , n28740 , n28745 );
or ( n28748 , n28743 , n28746 , n28747 );
xor ( n28749 , n28630 , n28676 );
xor ( n28750 , n28749 , n28679 );
and ( n28751 , n28748 , n28750 );
xor ( n28752 , n28590 , n28592 );
xor ( n28753 , n28752 , n28595 );
and ( n28754 , n28750 , n28753 );
and ( n28755 , n28748 , n28753 );
or ( n28756 , n28751 , n28754 , n28755 );
and ( n28757 , n28694 , n28756 );
xor ( n28758 , n28694 , n28756 );
xor ( n28759 , n28748 , n28750 );
xor ( n28760 , n28759 , n28753 );
and ( n28761 , n23284 , n21735 );
and ( n28762 , n23165 , n21732 );
nor ( n28763 , n28761 , n28762 );
xnor ( n28764 , n28763 , n21730 );
and ( n28765 , n23575 , n22252 );
and ( n28766 , n23446 , n22250 );
nor ( n28767 , n28765 , n28766 );
xnor ( n28768 , n28767 , n22258 );
and ( n28769 , n28764 , n28768 );
xor ( n28770 , n28654 , n28658 );
xor ( n28771 , n28770 , n28663 );
and ( n28772 , n28768 , n28771 );
and ( n28773 , n28764 , n28771 );
or ( n28774 , n28769 , n28772 , n28773 );
and ( n28775 , n23446 , n21735 );
and ( n28776 , n23284 , n21732 );
nor ( n28777 , n28775 , n28776 );
xnor ( n28778 , n28777 , n21730 );
and ( n28779 , n23954 , n22252 );
and ( n28780 , n23575 , n22250 );
nor ( n28781 , n28779 , n28780 );
xnor ( n28782 , n28781 , n22258 );
and ( n28783 , n28778 , n28782 );
xor ( n28784 , n28718 , n28722 );
xor ( n28785 , n28784 , n28727 );
and ( n28786 , n28782 , n28785 );
and ( n28787 , n28778 , n28785 );
or ( n28788 , n28783 , n28786 , n28787 );
xor ( n28789 , n28539 , n28543 );
and ( n28790 , n26360 , n21976 );
not ( n28791 , n28790 );
and ( n28792 , n28791 , n21988 );
and ( n28793 , n26360 , n21978 );
and ( n28794 , n26368 , n21976 );
nor ( n28795 , n28793 , n28794 );
xnor ( n28796 , n28795 , n21988 );
and ( n28797 , n28792 , n28796 );
and ( n28798 , n26368 , n21978 );
and ( n28799 , n26214 , n21976 );
nor ( n28800 , n28798 , n28799 );
xnor ( n28801 , n28800 , n21988 );
and ( n28802 , n28797 , n28801 );
and ( n28803 , n28801 , n28537 );
and ( n28804 , n28797 , n28537 );
or ( n28805 , n28802 , n28803 , n28804 );
and ( n28806 , n28789 , n28805 );
and ( n28807 , n26214 , n21978 );
and ( n28808 , n26107 , n21976 );
nor ( n28809 , n28807 , n28808 );
xnor ( n28810 , n28809 , n21988 );
and ( n28811 , n28805 , n28810 );
and ( n28812 , n28789 , n28810 );
or ( n28813 , n28806 , n28811 , n28812 );
and ( n28814 , n25633 , n22323 );
and ( n28815 , n25427 , n22321 );
nor ( n28816 , n28814 , n28815 );
xnor ( n28817 , n28816 , n22329 );
and ( n28818 , n28813 , n28817 );
xor ( n28819 , n28698 , n28702 );
xor ( n28820 , n28819 , n28705 );
and ( n28821 , n28817 , n28820 );
and ( n28822 , n28813 , n28820 );
or ( n28823 , n28818 , n28821 , n28822 );
and ( n28824 , n24896 , n21854 );
and ( n28825 , n24753 , n21852 );
nor ( n28826 , n28824 , n28825 );
xnor ( n28827 , n28826 , n21864 );
and ( n28828 , n28823 , n28827 );
and ( n28829 , n25337 , n21779 );
and ( n28830 , n25004 , n21777 );
nor ( n28831 , n28829 , n28830 );
xnor ( n28832 , n28831 , n21789 );
and ( n28833 , n28827 , n28832 );
and ( n28834 , n28823 , n28832 );
or ( n28835 , n28828 , n28833 , n28834 );
and ( n28836 , n24446 , n22305 );
and ( n28837 , n24011 , n22303 );
nor ( n28838 , n28836 , n28837 );
xnor ( n28839 , n28838 , n22315 );
and ( n28840 , n28835 , n28839 );
xor ( n28841 , n28644 , n28648 );
xor ( n28842 , n28841 , n28651 );
and ( n28843 , n28839 , n28842 );
and ( n28844 , n28835 , n28842 );
or ( n28845 , n28840 , n28843 , n28844 );
and ( n28846 , n28788 , n28845 );
xor ( n28847 , n28730 , n28734 );
xor ( n28848 , n28847 , n28737 );
and ( n28849 , n28845 , n28848 );
and ( n28850 , n28788 , n28848 );
or ( n28851 , n28846 , n28849 , n28850 );
and ( n28852 , n28774 , n28851 );
xor ( n28853 , n28740 , n28742 );
xor ( n28854 , n28853 , n28745 );
and ( n28855 , n28851 , n28854 );
and ( n28856 , n28774 , n28854 );
or ( n28857 , n28852 , n28855 , n28856 );
and ( n28858 , n28760 , n28857 );
xor ( n28859 , n28760 , n28857 );
xor ( n28860 , n28792 , n28796 );
and ( n28861 , n26360 , n21955 );
not ( n28862 , n28861 );
and ( n28863 , n28862 , n21967 );
and ( n28864 , n26360 , n21957 );
and ( n28865 , n26368 , n21955 );
nor ( n28866 , n28864 , n28865 );
xnor ( n28867 , n28866 , n21967 );
and ( n28868 , n28863 , n28867 );
and ( n28869 , n26368 , n21957 );
and ( n28870 , n26214 , n21955 );
nor ( n28871 , n28869 , n28870 );
xnor ( n28872 , n28871 , n21967 );
and ( n28873 , n28868 , n28872 );
and ( n28874 , n28872 , n28790 );
and ( n28875 , n28868 , n28790 );
or ( n28876 , n28873 , n28874 , n28875 );
and ( n28877 , n28860 , n28876 );
and ( n28878 , n26214 , n21957 );
and ( n28879 , n26107 , n21955 );
nor ( n28880 , n28878 , n28879 );
xnor ( n28881 , n28880 , n21967 );
and ( n28882 , n28876 , n28881 );
and ( n28883 , n28860 , n28881 );
or ( n28884 , n28877 , n28882 , n28883 );
and ( n28885 , n26107 , n21957 );
and ( n28886 , n25986 , n21955 );
nor ( n28887 , n28885 , n28886 );
xnor ( n28888 , n28887 , n21967 );
and ( n28889 , n28884 , n28888 );
xor ( n28890 , n28797 , n28801 );
xor ( n28891 , n28890 , n28537 );
and ( n28892 , n28888 , n28891 );
and ( n28893 , n28884 , n28891 );
or ( n28894 , n28889 , n28892 , n28893 );
and ( n28895 , n25427 , n21779 );
and ( n28896 , n25347 , n21777 );
nor ( n28897 , n28895 , n28896 );
xnor ( n28898 , n28897 , n21789 );
and ( n28899 , n28894 , n28898 );
and ( n28900 , n25753 , n22323 );
and ( n28901 , n25633 , n22321 );
nor ( n28902 , n28900 , n28901 );
xnor ( n28903 , n28902 , n22329 );
and ( n28904 , n25986 , n21957 );
and ( n28905 , n25833 , n21955 );
nor ( n28906 , n28904 , n28905 );
xnor ( n28907 , n28906 , n21967 );
xor ( n28908 , n28903 , n28907 );
xor ( n28909 , n28789 , n28805 );
xor ( n28910 , n28909 , n28810 );
xor ( n28911 , n28908 , n28910 );
and ( n28912 , n28898 , n28911 );
and ( n28913 , n28894 , n28911 );
or ( n28914 , n28899 , n28912 , n28913 );
and ( n28915 , n24753 , n22305 );
and ( n28916 , n24544 , n22303 );
nor ( n28917 , n28915 , n28916 );
xnor ( n28918 , n28917 , n22315 );
and ( n28919 , n28914 , n28918 );
and ( n28920 , n25004 , n21854 );
and ( n28921 , n24896 , n21852 );
nor ( n28922 , n28920 , n28921 );
xnor ( n28923 , n28922 , n21864 );
and ( n28924 , n28918 , n28923 );
and ( n28925 , n28914 , n28923 );
or ( n28926 , n28919 , n28924 , n28925 );
and ( n28927 , n24011 , n22252 );
and ( n28928 , n23954 , n22250 );
nor ( n28929 , n28927 , n28928 );
xnor ( n28930 , n28929 , n22258 );
and ( n28931 , n28926 , n28930 );
xor ( n28932 , n28823 , n28827 );
xor ( n28933 , n28932 , n28832 );
and ( n28934 , n28930 , n28933 );
and ( n28935 , n28926 , n28933 );
or ( n28936 , n28931 , n28934 , n28935 );
and ( n28937 , n28903 , n28907 );
and ( n28938 , n28907 , n28910 );
and ( n28939 , n28903 , n28910 );
or ( n28940 , n28937 , n28938 , n28939 );
and ( n28941 , n25347 , n21779 );
and ( n28942 , n25337 , n21777 );
nor ( n28943 , n28941 , n28942 );
xnor ( n28944 , n28943 , n21789 );
and ( n28945 , n28940 , n28944 );
xor ( n28946 , n28813 , n28817 );
xor ( n28947 , n28946 , n28820 );
and ( n28948 , n28944 , n28947 );
and ( n28949 , n28940 , n28947 );
or ( n28950 , n28945 , n28948 , n28949 );
and ( n28951 , n24544 , n22305 );
and ( n28952 , n24446 , n22303 );
nor ( n28953 , n28951 , n28952 );
xnor ( n28954 , n28953 , n22315 );
and ( n28955 , n28950 , n28954 );
xor ( n28956 , n28708 , n28712 );
xor ( n28957 , n28956 , n28715 );
and ( n28958 , n28954 , n28957 );
and ( n28959 , n28950 , n28957 );
or ( n28960 , n28955 , n28958 , n28959 );
and ( n28961 , n28936 , n28960 );
xor ( n28962 , n28835 , n28839 );
xor ( n28963 , n28962 , n28842 );
and ( n28964 , n28960 , n28963 );
and ( n28965 , n28936 , n28963 );
or ( n28966 , n28961 , n28964 , n28965 );
xor ( n28967 , n28764 , n28768 );
xor ( n28968 , n28967 , n28771 );
and ( n28969 , n28966 , n28968 );
xor ( n28970 , n28788 , n28845 );
xor ( n28971 , n28970 , n28848 );
and ( n28972 , n28968 , n28971 );
and ( n28973 , n28966 , n28971 );
or ( n28974 , n28969 , n28972 , n28973 );
xor ( n28975 , n28774 , n28851 );
xor ( n28976 , n28975 , n28854 );
and ( n28977 , n28974 , n28976 );
xor ( n28978 , n28974 , n28976 );
xor ( n28979 , n28966 , n28968 );
xor ( n28980 , n28979 , n28971 );
and ( n28981 , n23954 , n21735 );
and ( n28982 , n23575 , n21732 );
nor ( n28983 , n28981 , n28982 );
xnor ( n28984 , n28983 , n21730 );
and ( n28985 , n24446 , n22252 );
and ( n28986 , n24011 , n22250 );
nor ( n28987 , n28985 , n28986 );
xnor ( n28988 , n28987 , n22258 );
and ( n28989 , n28984 , n28988 );
xor ( n28990 , n28940 , n28944 );
xor ( n28991 , n28990 , n28947 );
and ( n28992 , n28988 , n28991 );
and ( n28993 , n28984 , n28991 );
or ( n28994 , n28989 , n28992 , n28993 );
and ( n28995 , n23575 , n21735 );
and ( n28996 , n23446 , n21732 );
nor ( n28997 , n28995 , n28996 );
xnor ( n28998 , n28997 , n21730 );
and ( n28999 , n28994 , n28998 );
xor ( n29000 , n28950 , n28954 );
xor ( n29001 , n29000 , n28957 );
and ( n29002 , n28998 , n29001 );
and ( n29003 , n28994 , n29001 );
or ( n29004 , n28999 , n29002 , n29003 );
xor ( n29005 , n28778 , n28782 );
xor ( n29006 , n29005 , n28785 );
and ( n29007 , n29004 , n29006 );
xor ( n29008 , n28936 , n28960 );
xor ( n29009 , n29008 , n28963 );
and ( n29010 , n29006 , n29009 );
and ( n29011 , n29004 , n29009 );
or ( n29012 , n29007 , n29010 , n29011 );
and ( n29013 , n28980 , n29012 );
xor ( n29014 , n28980 , n29012 );
xor ( n29015 , n29004 , n29006 );
xor ( n29016 , n29015 , n29009 );
xor ( n29017 , n28926 , n28930 );
xor ( n29018 , n29017 , n28933 );
xor ( n29019 , n28994 , n28998 );
xor ( n29020 , n29019 , n29001 );
and ( n29021 , n29018 , n29020 );
and ( n29022 , n25753 , n21779 );
and ( n29023 , n25633 , n21777 );
nor ( n29024 , n29022 , n29023 );
xnor ( n29025 , n29024 , n21789 );
and ( n29026 , n25986 , n22323 );
and ( n29027 , n25833 , n22321 );
nor ( n29028 , n29026 , n29027 );
xnor ( n29029 , n29028 , n22329 );
and ( n29030 , n29025 , n29029 );
xor ( n29031 , n28860 , n28876 );
xor ( n29032 , n29031 , n28881 );
and ( n29033 , n29029 , n29032 );
and ( n29034 , n29025 , n29032 );
or ( n29035 , n29030 , n29033 , n29034 );
and ( n29036 , n25347 , n21854 );
and ( n29037 , n25337 , n21852 );
nor ( n29038 , n29036 , n29037 );
xnor ( n29039 , n29038 , n21864 );
and ( n29040 , n29035 , n29039 );
and ( n29041 , n25633 , n21779 );
and ( n29042 , n25427 , n21777 );
nor ( n29043 , n29041 , n29042 );
xnor ( n29044 , n29043 , n21789 );
and ( n29045 , n25833 , n22323 );
and ( n29046 , n25753 , n22321 );
nor ( n29047 , n29045 , n29046 );
xnor ( n29048 , n29047 , n22329 );
xor ( n29049 , n29044 , n29048 );
xor ( n29050 , n28884 , n28888 );
xor ( n29051 , n29050 , n28891 );
xor ( n29052 , n29049 , n29051 );
and ( n29053 , n29039 , n29052 );
and ( n29054 , n29035 , n29052 );
or ( n29055 , n29040 , n29053 , n29054 );
and ( n29056 , n24544 , n22252 );
and ( n29057 , n24446 , n22250 );
nor ( n29058 , n29056 , n29057 );
xnor ( n29059 , n29058 , n22258 );
and ( n29060 , n29055 , n29059 );
and ( n29061 , n25337 , n21854 );
and ( n29062 , n25004 , n21852 );
nor ( n29063 , n29061 , n29062 );
xnor ( n29064 , n29063 , n21864 );
and ( n29065 , n29059 , n29064 );
and ( n29066 , n29055 , n29064 );
or ( n29067 , n29060 , n29065 , n29066 );
and ( n29068 , n29044 , n29048 );
and ( n29069 , n29048 , n29051 );
and ( n29070 , n29044 , n29051 );
or ( n29071 , n29068 , n29069 , n29070 );
and ( n29072 , n24896 , n22305 );
and ( n29073 , n24753 , n22303 );
nor ( n29074 , n29072 , n29073 );
xnor ( n29075 , n29074 , n22315 );
and ( n29076 , n29071 , n29075 );
xor ( n29077 , n28894 , n28898 );
xor ( n29078 , n29077 , n28911 );
and ( n29079 , n29075 , n29078 );
and ( n29080 , n29071 , n29078 );
or ( n29081 , n29076 , n29079 , n29080 );
and ( n29082 , n29067 , n29081 );
xor ( n29083 , n28914 , n28918 );
xor ( n29084 , n29083 , n28923 );
and ( n29085 , n29081 , n29084 );
and ( n29086 , n29067 , n29084 );
or ( n29087 , n29082 , n29085 , n29086 );
and ( n29088 , n29020 , n29087 );
and ( n29089 , n29018 , n29087 );
or ( n29090 , n29021 , n29088 , n29089 );
and ( n29091 , n29016 , n29090 );
xor ( n29092 , n29016 , n29090 );
xor ( n29093 , n28863 , n28867 );
and ( n29094 , n26360 , n22321 );
not ( n29095 , n29094 );
and ( n29096 , n29095 , n22329 );
and ( n29097 , n26360 , n22323 );
and ( n29098 , n26368 , n22321 );
nor ( n29099 , n29097 , n29098 );
xnor ( n29100 , n29099 , n22329 );
and ( n29101 , n29096 , n29100 );
and ( n29102 , n26368 , n22323 );
and ( n29103 , n26214 , n22321 );
nor ( n29104 , n29102 , n29103 );
xnor ( n29105 , n29104 , n22329 );
and ( n29106 , n29101 , n29105 );
and ( n29107 , n29105 , n28861 );
and ( n29108 , n29101 , n28861 );
or ( n29109 , n29106 , n29107 , n29108 );
and ( n29110 , n29093 , n29109 );
and ( n29111 , n26214 , n22323 );
and ( n29112 , n26107 , n22321 );
nor ( n29113 , n29111 , n29112 );
xnor ( n29114 , n29113 , n22329 );
and ( n29115 , n29109 , n29114 );
and ( n29116 , n29093 , n29114 );
or ( n29117 , n29110 , n29115 , n29116 );
and ( n29118 , n26107 , n22323 );
and ( n29119 , n25986 , n22321 );
nor ( n29120 , n29118 , n29119 );
xnor ( n29121 , n29120 , n22329 );
and ( n29122 , n29117 , n29121 );
xor ( n29123 , n28868 , n28872 );
xor ( n29124 , n29123 , n28790 );
and ( n29125 , n29121 , n29124 );
and ( n29126 , n29117 , n29124 );
or ( n29127 , n29122 , n29125 , n29126 );
and ( n29128 , n25427 , n21854 );
and ( n29129 , n25347 , n21852 );
nor ( n29130 , n29128 , n29129 );
xnor ( n29131 , n29130 , n21864 );
and ( n29132 , n29127 , n29131 );
xor ( n29133 , n29025 , n29029 );
xor ( n29134 , n29133 , n29032 );
and ( n29135 , n29131 , n29134 );
and ( n29136 , n29127 , n29134 );
or ( n29137 , n29132 , n29135 , n29136 );
and ( n29138 , n24753 , n22252 );
and ( n29139 , n24544 , n22250 );
nor ( n29140 , n29138 , n29139 );
xnor ( n29141 , n29140 , n22258 );
and ( n29142 , n29137 , n29141 );
and ( n29143 , n25004 , n22305 );
and ( n29144 , n24896 , n22303 );
nor ( n29145 , n29143 , n29144 );
xnor ( n29146 , n29145 , n22315 );
and ( n29147 , n29141 , n29146 );
and ( n29148 , n29137 , n29146 );
or ( n29149 , n29142 , n29147 , n29148 );
and ( n29150 , n24011 , n21735 );
and ( n29151 , n23954 , n21732 );
nor ( n29152 , n29150 , n29151 );
xnor ( n29153 , n29152 , n21730 );
and ( n29154 , n29149 , n29153 );
xor ( n29155 , n29071 , n29075 );
xor ( n29156 , n29155 , n29078 );
and ( n29157 , n29153 , n29156 );
and ( n29158 , n29149 , n29156 );
or ( n29159 , n29154 , n29157 , n29158 );
xor ( n29160 , n29067 , n29081 );
xor ( n29161 , n29160 , n29084 );
and ( n29162 , n29159 , n29161 );
xor ( n29163 , n28984 , n28988 );
xor ( n29164 , n29163 , n28991 );
and ( n29165 , n29161 , n29164 );
and ( n29166 , n29159 , n29164 );
or ( n29167 , n29162 , n29165 , n29166 );
xor ( n29168 , n29018 , n29020 );
xor ( n29169 , n29168 , n29087 );
and ( n29170 , n29167 , n29169 );
xor ( n29171 , n29167 , n29169 );
and ( n29172 , n25633 , n21854 );
and ( n29173 , n25427 , n21852 );
nor ( n29174 , n29172 , n29173 );
xnor ( n29175 , n29174 , n21864 );
and ( n29176 , n25833 , n21779 );
and ( n29177 , n25753 , n21777 );
nor ( n29178 , n29176 , n29177 );
xnor ( n29179 , n29178 , n21789 );
and ( n29180 , n29175 , n29179 );
xor ( n29181 , n29117 , n29121 );
xor ( n29182 , n29181 , n29124 );
and ( n29183 , n29179 , n29182 );
and ( n29184 , n29175 , n29182 );
or ( n29185 , n29180 , n29183 , n29184 );
and ( n29186 , n24896 , n22252 );
and ( n29187 , n24753 , n22250 );
nor ( n29188 , n29186 , n29187 );
xnor ( n29189 , n29188 , n22258 );
and ( n29190 , n29185 , n29189 );
xor ( n29191 , n29127 , n29131 );
xor ( n29192 , n29191 , n29134 );
and ( n29193 , n29189 , n29192 );
and ( n29194 , n29185 , n29192 );
or ( n29195 , n29190 , n29193 , n29194 );
and ( n29196 , n24446 , n21735 );
and ( n29197 , n24011 , n21732 );
nor ( n29198 , n29196 , n29197 );
xnor ( n29199 , n29198 , n21730 );
and ( n29200 , n29195 , n29199 );
xor ( n29201 , n29035 , n29039 );
xor ( n29202 , n29201 , n29052 );
and ( n29203 , n29199 , n29202 );
and ( n29204 , n29195 , n29202 );
or ( n29205 , n29200 , n29203 , n29204 );
xor ( n29206 , n29055 , n29059 );
xor ( n29207 , n29206 , n29064 );
and ( n29208 , n29205 , n29207 );
xor ( n29209 , n29149 , n29153 );
xor ( n29210 , n29209 , n29156 );
and ( n29211 , n29207 , n29210 );
and ( n29212 , n29205 , n29210 );
or ( n29213 , n29208 , n29211 , n29212 );
xor ( n29214 , n29159 , n29161 );
xor ( n29215 , n29214 , n29164 );
and ( n29216 , n29213 , n29215 );
xor ( n29217 , n29213 , n29215 );
xor ( n29218 , n29205 , n29207 );
xor ( n29219 , n29218 , n29210 );
and ( n29220 , n25753 , n21854 );
and ( n29221 , n25633 , n21852 );
nor ( n29222 , n29220 , n29221 );
xnor ( n29223 , n29222 , n21864 );
and ( n29224 , n25986 , n21779 );
and ( n29225 , n25833 , n21777 );
nor ( n29226 , n29224 , n29225 );
xnor ( n29227 , n29226 , n21789 );
and ( n29228 , n29223 , n29227 );
xor ( n29229 , n29093 , n29109 );
xor ( n29230 , n29229 , n29114 );
and ( n29231 , n29227 , n29230 );
and ( n29232 , n29223 , n29230 );
or ( n29233 , n29228 , n29231 , n29232 );
and ( n29234 , n25347 , n22305 );
and ( n29235 , n25337 , n22303 );
nor ( n29236 , n29234 , n29235 );
xnor ( n29237 , n29236 , n22315 );
and ( n29238 , n29233 , n29237 );
xor ( n29239 , n29175 , n29179 );
xor ( n29240 , n29239 , n29182 );
and ( n29241 , n29237 , n29240 );
and ( n29242 , n29233 , n29240 );
or ( n29243 , n29238 , n29241 , n29242 );
and ( n29244 , n24544 , n21735 );
and ( n29245 , n24446 , n21732 );
nor ( n29246 , n29244 , n29245 );
xnor ( n29247 , n29246 , n21730 );
and ( n29248 , n29243 , n29247 );
and ( n29249 , n25337 , n22305 );
and ( n29250 , n25004 , n22303 );
nor ( n29251 , n29249 , n29250 );
xnor ( n29252 , n29251 , n22315 );
and ( n29253 , n29247 , n29252 );
and ( n29254 , n29243 , n29252 );
or ( n29255 , n29248 , n29253 , n29254 );
xor ( n29256 , n29137 , n29141 );
xor ( n29257 , n29256 , n29146 );
and ( n29258 , n29255 , n29257 );
xor ( n29259 , n29195 , n29199 );
xor ( n29260 , n29259 , n29202 );
and ( n29261 , n29257 , n29260 );
and ( n29262 , n29255 , n29260 );
or ( n29263 , n29258 , n29261 , n29262 );
and ( n29264 , n29219 , n29263 );
xor ( n29265 , n29219 , n29263 );
xor ( n29266 , n29255 , n29257 );
xor ( n29267 , n29266 , n29260 );
xor ( n29268 , n29096 , n29100 );
and ( n29269 , n26360 , n21777 );
not ( n29270 , n29269 );
and ( n29271 , n29270 , n21789 );
and ( n29272 , n26360 , n21779 );
and ( n29273 , n26368 , n21777 );
nor ( n29274 , n29272 , n29273 );
xnor ( n29275 , n29274 , n21789 );
and ( n29276 , n29271 , n29275 );
and ( n29277 , n26368 , n21779 );
and ( n29278 , n26214 , n21777 );
nor ( n29279 , n29277 , n29278 );
xnor ( n29280 , n29279 , n21789 );
and ( n29281 , n29276 , n29280 );
and ( n29282 , n29280 , n29094 );
and ( n29283 , n29276 , n29094 );
or ( n29284 , n29281 , n29282 , n29283 );
and ( n29285 , n29268 , n29284 );
and ( n29286 , n26214 , n21779 );
and ( n29287 , n26107 , n21777 );
nor ( n29288 , n29286 , n29287 );
xnor ( n29289 , n29288 , n21789 );
and ( n29290 , n29284 , n29289 );
and ( n29291 , n29268 , n29289 );
or ( n29292 , n29285 , n29290 , n29291 );
and ( n29293 , n26107 , n21779 );
and ( n29294 , n25986 , n21777 );
nor ( n29295 , n29293 , n29294 );
xnor ( n29296 , n29295 , n21789 );
and ( n29297 , n29292 , n29296 );
xor ( n29298 , n29101 , n29105 );
xor ( n29299 , n29298 , n28861 );
and ( n29300 , n29296 , n29299 );
and ( n29301 , n29292 , n29299 );
or ( n29302 , n29297 , n29300 , n29301 );
and ( n29303 , n25427 , n22305 );
and ( n29304 , n25347 , n22303 );
nor ( n29305 , n29303 , n29304 );
xnor ( n29306 , n29305 , n22315 );
and ( n29307 , n29302 , n29306 );
xor ( n29308 , n29223 , n29227 );
xor ( n29309 , n29308 , n29230 );
and ( n29310 , n29306 , n29309 );
and ( n29311 , n29302 , n29309 );
or ( n29312 , n29307 , n29310 , n29311 );
and ( n29313 , n24753 , n21735 );
and ( n29314 , n24544 , n21732 );
nor ( n29315 , n29313 , n29314 );
xnor ( n29316 , n29315 , n21730 );
and ( n29317 , n29312 , n29316 );
and ( n29318 , n25004 , n22252 );
and ( n29319 , n24896 , n22250 );
nor ( n29320 , n29318 , n29319 );
xnor ( n29321 , n29320 , n22258 );
and ( n29322 , n29316 , n29321 );
and ( n29323 , n29312 , n29321 );
or ( n29324 , n29317 , n29322 , n29323 );
xor ( n29325 , n29243 , n29247 );
xor ( n29326 , n29325 , n29252 );
and ( n29327 , n29324 , n29326 );
xor ( n29328 , n29185 , n29189 );
xor ( n29329 , n29328 , n29192 );
and ( n29330 , n29326 , n29329 );
and ( n29331 , n29324 , n29329 );
or ( n29332 , n29327 , n29330 , n29331 );
and ( n29333 , n29267 , n29332 );
xor ( n29334 , n29267 , n29332 );
and ( n29335 , n25633 , n22305 );
and ( n29336 , n25427 , n22303 );
nor ( n29337 , n29335 , n29336 );
xnor ( n29338 , n29337 , n22315 );
and ( n29339 , n25833 , n21854 );
and ( n29340 , n25753 , n21852 );
nor ( n29341 , n29339 , n29340 );
xnor ( n29342 , n29341 , n21864 );
and ( n29343 , n29338 , n29342 );
xor ( n29344 , n29292 , n29296 );
xor ( n29345 , n29344 , n29299 );
and ( n29346 , n29342 , n29345 );
and ( n29347 , n29338 , n29345 );
or ( n29348 , n29343 , n29346 , n29347 );
and ( n29349 , n25337 , n22252 );
and ( n29350 , n25004 , n22250 );
nor ( n29351 , n29349 , n29350 );
xnor ( n29352 , n29351 , n22258 );
and ( n29353 , n29348 , n29352 );
xor ( n29354 , n29302 , n29306 );
xor ( n29355 , n29354 , n29309 );
and ( n29356 , n29352 , n29355 );
and ( n29357 , n29348 , n29355 );
or ( n29358 , n29353 , n29356 , n29357 );
xor ( n29359 , n29312 , n29316 );
xor ( n29360 , n29359 , n29321 );
and ( n29361 , n29358 , n29360 );
xor ( n29362 , n29233 , n29237 );
xor ( n29363 , n29362 , n29240 );
and ( n29364 , n29360 , n29363 );
and ( n29365 , n29358 , n29363 );
or ( n29366 , n29361 , n29364 , n29365 );
xor ( n29367 , n29324 , n29326 );
xor ( n29368 , n29367 , n29329 );
and ( n29369 , n29366 , n29368 );
xor ( n29370 , n29366 , n29368 );
xor ( n29371 , n29358 , n29360 );
xor ( n29372 , n29371 , n29363 );
and ( n29373 , n25753 , n22305 );
and ( n29374 , n25633 , n22303 );
nor ( n29375 , n29373 , n29374 );
xnor ( n29376 , n29375 , n22315 );
and ( n29377 , n25986 , n21854 );
and ( n29378 , n25833 , n21852 );
nor ( n29379 , n29377 , n29378 );
xnor ( n29380 , n29379 , n21864 );
and ( n29381 , n29376 , n29380 );
xor ( n29382 , n29268 , n29284 );
xor ( n29383 , n29382 , n29289 );
and ( n29384 , n29380 , n29383 );
and ( n29385 , n29376 , n29383 );
or ( n29386 , n29381 , n29384 , n29385 );
and ( n29387 , n25347 , n22252 );
and ( n29388 , n25337 , n22250 );
nor ( n29389 , n29387 , n29388 );
xnor ( n29390 , n29389 , n22258 );
and ( n29391 , n29386 , n29390 );
xor ( n29392 , n29338 , n29342 );
xor ( n29393 , n29392 , n29345 );
and ( n29394 , n29390 , n29393 );
and ( n29395 , n29386 , n29393 );
or ( n29396 , n29391 , n29394 , n29395 );
and ( n29397 , n24896 , n21735 );
and ( n29398 , n24753 , n21732 );
nor ( n29399 , n29397 , n29398 );
xnor ( n29400 , n29399 , n21730 );
and ( n29401 , n29396 , n29400 );
xor ( n29402 , n29348 , n29352 );
xor ( n29403 , n29402 , n29355 );
and ( n29404 , n29400 , n29403 );
and ( n29405 , n29396 , n29403 );
or ( n29406 , n29401 , n29404 , n29405 );
and ( n29407 , n29372 , n29406 );
xor ( n29408 , n29372 , n29406 );
xor ( n29409 , n29396 , n29400 );
xor ( n29410 , n29409 , n29403 );
xor ( n29411 , n29271 , n29275 );
and ( n29412 , n26360 , n21852 );
not ( n29413 , n29412 );
and ( n29414 , n29413 , n21864 );
and ( n29415 , n26360 , n21854 );
and ( n29416 , n26368 , n21852 );
nor ( n29417 , n29415 , n29416 );
xnor ( n29418 , n29417 , n21864 );
and ( n29419 , n29414 , n29418 );
and ( n29420 , n26368 , n21854 );
and ( n29421 , n26214 , n21852 );
nor ( n29422 , n29420 , n29421 );
xnor ( n29423 , n29422 , n21864 );
and ( n29424 , n29419 , n29423 );
and ( n29425 , n29423 , n29269 );
and ( n29426 , n29419 , n29269 );
or ( n29427 , n29424 , n29425 , n29426 );
and ( n29428 , n29411 , n29427 );
and ( n29429 , n26214 , n21854 );
and ( n29430 , n26107 , n21852 );
nor ( n29431 , n29429 , n29430 );
xnor ( n29432 , n29431 , n21864 );
and ( n29433 , n29427 , n29432 );
and ( n29434 , n29411 , n29432 );
or ( n29435 , n29428 , n29433 , n29434 );
and ( n29436 , n26107 , n21854 );
and ( n29437 , n25986 , n21852 );
nor ( n29438 , n29436 , n29437 );
xnor ( n29439 , n29438 , n21864 );
and ( n29440 , n29435 , n29439 );
xor ( n29441 , n29276 , n29280 );
xor ( n29442 , n29441 , n29094 );
and ( n29443 , n29439 , n29442 );
and ( n29444 , n29435 , n29442 );
or ( n29445 , n29440 , n29443 , n29444 );
and ( n29446 , n25427 , n22252 );
and ( n29447 , n25347 , n22250 );
nor ( n29448 , n29446 , n29447 );
xnor ( n29449 , n29448 , n22258 );
and ( n29450 , n29445 , n29449 );
xor ( n29451 , n29376 , n29380 );
xor ( n29452 , n29451 , n29383 );
and ( n29453 , n29449 , n29452 );
and ( n29454 , n29445 , n29452 );
or ( n29455 , n29450 , n29453 , n29454 );
and ( n29456 , n25004 , n21735 );
and ( n29457 , n24896 , n21732 );
nor ( n29458 , n29456 , n29457 );
xnor ( n29459 , n29458 , n21730 );
and ( n29460 , n29455 , n29459 );
xor ( n29461 , n29386 , n29390 );
xor ( n29462 , n29461 , n29393 );
and ( n29463 , n29459 , n29462 );
and ( n29464 , n29455 , n29462 );
or ( n29465 , n29460 , n29463 , n29464 );
and ( n29466 , n29410 , n29465 );
xor ( n29467 , n29410 , n29465 );
and ( n29468 , n25633 , n22252 );
and ( n29469 , n25427 , n22250 );
nor ( n29470 , n29468 , n29469 );
xnor ( n29471 , n29470 , n22258 );
and ( n29472 , n25833 , n22305 );
and ( n29473 , n25753 , n22303 );
nor ( n29474 , n29472 , n29473 );
xnor ( n29475 , n29474 , n22315 );
and ( n29476 , n29471 , n29475 );
xor ( n29477 , n29435 , n29439 );
xor ( n29478 , n29477 , n29442 );
and ( n29479 , n29475 , n29478 );
and ( n29480 , n29471 , n29478 );
or ( n29481 , n29476 , n29479 , n29480 );
and ( n29482 , n25337 , n21735 );
and ( n29483 , n25004 , n21732 );
nor ( n29484 , n29482 , n29483 );
xnor ( n29485 , n29484 , n21730 );
and ( n29486 , n29481 , n29485 );
xor ( n29487 , n29445 , n29449 );
xor ( n29488 , n29487 , n29452 );
and ( n29489 , n29485 , n29488 );
and ( n29490 , n29481 , n29488 );
or ( n29491 , n29486 , n29489 , n29490 );
xor ( n29492 , n29455 , n29459 );
xor ( n29493 , n29492 , n29462 );
and ( n29494 , n29491 , n29493 );
xor ( n29495 , n29491 , n29493 );
xor ( n29496 , n29481 , n29485 );
xor ( n29497 , n29496 , n29488 );
and ( n29498 , n25753 , n22252 );
and ( n29499 , n25633 , n22250 );
nor ( n29500 , n29498 , n29499 );
xnor ( n29501 , n29500 , n22258 );
and ( n29502 , n25986 , n22305 );
and ( n29503 , n25833 , n22303 );
nor ( n29504 , n29502 , n29503 );
xnor ( n29505 , n29504 , n22315 );
and ( n29506 , n29501 , n29505 );
xor ( n29507 , n29411 , n29427 );
xor ( n29508 , n29507 , n29432 );
and ( n29509 , n29505 , n29508 );
and ( n29510 , n29501 , n29508 );
or ( n29511 , n29506 , n29509 , n29510 );
and ( n29512 , n25347 , n21735 );
and ( n29513 , n25337 , n21732 );
nor ( n29514 , n29512 , n29513 );
xnor ( n29515 , n29514 , n21730 );
and ( n29516 , n29511 , n29515 );
xor ( n29517 , n29471 , n29475 );
xor ( n29518 , n29517 , n29478 );
and ( n29519 , n29515 , n29518 );
and ( n29520 , n29511 , n29518 );
or ( n29521 , n29516 , n29519 , n29520 );
and ( n29522 , n29497 , n29521 );
xor ( n29523 , n29497 , n29521 );
and ( n29524 , n25833 , n22252 );
and ( n29525 , n25753 , n22250 );
nor ( n29526 , n29524 , n29525 );
xnor ( n29527 , n29526 , n22258 );
and ( n29528 , n26107 , n22305 );
and ( n29529 , n25986 , n22303 );
nor ( n29530 , n29528 , n29529 );
xnor ( n29531 , n29530 , n22315 );
and ( n29532 , n29527 , n29531 );
xor ( n29533 , n29419 , n29423 );
xor ( n29534 , n29533 , n29269 );
and ( n29535 , n29531 , n29534 );
and ( n29536 , n29527 , n29534 );
or ( n29537 , n29532 , n29535 , n29536 );
and ( n29538 , n25427 , n21735 );
and ( n29539 , n25347 , n21732 );
nor ( n29540 , n29538 , n29539 );
xnor ( n29541 , n29540 , n21730 );
and ( n29542 , n29537 , n29541 );
xor ( n29543 , n29501 , n29505 );
xor ( n29544 , n29543 , n29508 );
and ( n29545 , n29541 , n29544 );
and ( n29546 , n29537 , n29544 );
or ( n29547 , n29542 , n29545 , n29546 );
xor ( n29548 , n29511 , n29515 );
xor ( n29549 , n29548 , n29518 );
and ( n29550 , n29547 , n29549 );
xor ( n29551 , n29547 , n29549 );
xor ( n29552 , n29414 , n29418 );
and ( n29553 , n26360 , n22303 );
not ( n29554 , n29553 );
and ( n29555 , n29554 , n22315 );
and ( n29556 , n26360 , n22305 );
and ( n29557 , n26368 , n22303 );
nor ( n29558 , n29556 , n29557 );
xnor ( n29559 , n29558 , n22315 );
and ( n29560 , n29555 , n29559 );
and ( n29561 , n26368 , n22305 );
and ( n29562 , n26214 , n22303 );
nor ( n29563 , n29561 , n29562 );
xnor ( n29564 , n29563 , n22315 );
and ( n29565 , n29560 , n29564 );
and ( n29566 , n29564 , n29412 );
and ( n29567 , n29560 , n29412 );
or ( n29568 , n29565 , n29566 , n29567 );
and ( n29569 , n29552 , n29568 );
and ( n29570 , n26214 , n22305 );
and ( n29571 , n26107 , n22303 );
nor ( n29572 , n29570 , n29571 );
xnor ( n29573 , n29572 , n22315 );
and ( n29574 , n29568 , n29573 );
and ( n29575 , n29552 , n29573 );
or ( n29576 , n29569 , n29574 , n29575 );
and ( n29577 , n25633 , n21735 );
and ( n29578 , n25427 , n21732 );
nor ( n29579 , n29577 , n29578 );
xnor ( n29580 , n29579 , n21730 );
and ( n29581 , n29576 , n29580 );
xor ( n29582 , n29527 , n29531 );
xor ( n29583 , n29582 , n29534 );
and ( n29584 , n29580 , n29583 );
and ( n29585 , n29576 , n29583 );
or ( n29586 , n29581 , n29584 , n29585 );
xor ( n29587 , n29537 , n29541 );
xor ( n29588 , n29587 , n29544 );
and ( n29589 , n29586 , n29588 );
xor ( n29590 , n29586 , n29588 );
xor ( n29591 , n29576 , n29580 );
xor ( n29592 , n29591 , n29583 );
and ( n29593 , n25753 , n21735 );
and ( n29594 , n25633 , n21732 );
nor ( n29595 , n29593 , n29594 );
xnor ( n29596 , n29595 , n21730 );
and ( n29597 , n25986 , n22252 );
and ( n29598 , n25833 , n22250 );
nor ( n29599 , n29597 , n29598 );
xnor ( n29600 , n29599 , n22258 );
and ( n29601 , n29596 , n29600 );
xor ( n29602 , n29552 , n29568 );
xor ( n29603 , n29602 , n29573 );
and ( n29604 , n29600 , n29603 );
and ( n29605 , n29596 , n29603 );
or ( n29606 , n29601 , n29604 , n29605 );
and ( n29607 , n29592 , n29606 );
xor ( n29608 , n29592 , n29606 );
and ( n29609 , n25833 , n21735 );
and ( n29610 , n25753 , n21732 );
nor ( n29611 , n29609 , n29610 );
xnor ( n29612 , n29611 , n21730 );
and ( n29613 , n26107 , n22252 );
and ( n29614 , n25986 , n22250 );
nor ( n29615 , n29613 , n29614 );
xnor ( n29616 , n29615 , n22258 );
and ( n29617 , n29612 , n29616 );
xor ( n29618 , n29560 , n29564 );
xor ( n29619 , n29618 , n29412 );
and ( n29620 , n29616 , n29619 );
and ( n29621 , n29612 , n29619 );
or ( n29622 , n29617 , n29620 , n29621 );
xor ( n29623 , n29596 , n29600 );
xor ( n29624 , n29623 , n29603 );
and ( n29625 , n29622 , n29624 );
xor ( n29626 , n29622 , n29624 );
xor ( n29627 , n29612 , n29616 );
xor ( n29628 , n29627 , n29619 );
xor ( n29629 , n29555 , n29559 );
and ( n29630 , n26360 , n22250 );
not ( n29631 , n29630 );
and ( n29632 , n29631 , n22258 );
and ( n29633 , n26360 , n22252 );
and ( n29634 , n26368 , n22250 );
nor ( n29635 , n29633 , n29634 );
xnor ( n29636 , n29635 , n22258 );
and ( n29637 , n29632 , n29636 );
and ( n29638 , n26368 , n22252 );
and ( n29639 , n26214 , n22250 );
nor ( n29640 , n29638 , n29639 );
xnor ( n29641 , n29640 , n22258 );
and ( n29642 , n29637 , n29641 );
and ( n29643 , n29641 , n29553 );
and ( n29644 , n29637 , n29553 );
or ( n29645 , n29642 , n29643 , n29644 );
and ( n29646 , n29629 , n29645 );
and ( n29647 , n26214 , n22252 );
and ( n29648 , n26107 , n22250 );
nor ( n29649 , n29647 , n29648 );
xnor ( n29650 , n29649 , n22258 );
and ( n29651 , n29645 , n29650 );
and ( n29652 , n29629 , n29650 );
or ( n29653 , n29646 , n29651 , n29652 );
and ( n29654 , n29628 , n29653 );
xor ( n29655 , n29628 , n29653 );
and ( n29656 , n25986 , n21735 );
and ( n29657 , n25833 , n21732 );
nor ( n29658 , n29656 , n29657 );
xnor ( n29659 , n29658 , n21730 );
xor ( n29660 , n29629 , n29645 );
xor ( n29661 , n29660 , n29650 );
and ( n29662 , n29659 , n29661 );
xor ( n29663 , n29659 , n29661 );
and ( n29664 , n26107 , n21735 );
and ( n29665 , n25986 , n21732 );
nor ( n29666 , n29664 , n29665 );
xnor ( n29667 , n29666 , n21730 );
xor ( n29668 , n29637 , n29641 );
xor ( n29669 , n29668 , n29553 );
and ( n29670 , n29667 , n29669 );
xor ( n29671 , n29667 , n29669 );
and ( n29672 , n26214 , n21735 );
and ( n29673 , n26107 , n21732 );
nor ( n29674 , n29672 , n29673 );
xnor ( n29675 , n29674 , n21730 );
xor ( n29676 , n29632 , n29636 );
and ( n29677 , n29675 , n29676 );
xor ( n29678 , n29675 , n29676 );
and ( n29679 , n26368 , n21735 );
and ( n29680 , n26214 , n21732 );
nor ( n29681 , n29679 , n29680 );
xnor ( n29682 , n29681 , n21730 );
and ( n29683 , n29682 , n29630 );
xor ( n29684 , n29682 , n29630 );
and ( n29685 , n26360 , n21735 );
and ( n29686 , n26368 , n21732 );
nor ( n29687 , n29685 , n29686 );
xnor ( n29688 , n29687 , n21730 );
and ( n29689 , n26360 , n21732 );
not ( n29690 , n29689 );
and ( n29691 , n29690 , n21730 );
and ( n29692 , n29688 , n29691 );
and ( n29693 , n29684 , n29692 );
or ( n29694 , n29683 , n29693 );
and ( n29695 , n29678 , n29694 );
or ( n29696 , n29677 , n29695 );
and ( n29697 , n29671 , n29696 );
or ( n29698 , n29670 , n29697 );
and ( n29699 , n29663 , n29698 );
or ( n29700 , n29662 , n29699 );
and ( n29701 , n29655 , n29700 );
or ( n29702 , n29654 , n29701 );
and ( n29703 , n29626 , n29702 );
or ( n29704 , n29625 , n29703 );
and ( n29705 , n29608 , n29704 );
or ( n29706 , n29607 , n29705 );
and ( n29707 , n29590 , n29706 );
or ( n29708 , n29589 , n29707 );
and ( n29709 , n29551 , n29708 );
or ( n29710 , n29550 , n29709 );
and ( n29711 , n29523 , n29710 );
or ( n29712 , n29522 , n29711 );
and ( n29713 , n29495 , n29712 );
or ( n29714 , n29494 , n29713 );
and ( n29715 , n29467 , n29714 );
or ( n29716 , n29466 , n29715 );
and ( n29717 , n29408 , n29716 );
or ( n29718 , n29407 , n29717 );
and ( n29719 , n29370 , n29718 );
or ( n29720 , n29369 , n29719 );
and ( n29721 , n29334 , n29720 );
or ( n29722 , n29333 , n29721 );
and ( n29723 , n29265 , n29722 );
or ( n29724 , n29264 , n29723 );
and ( n29725 , n29217 , n29724 );
or ( n29726 , n29216 , n29725 );
and ( n29727 , n29171 , n29726 );
or ( n29728 , n29170 , n29727 );
and ( n29729 , n29092 , n29728 );
or ( n29730 , n29091 , n29729 );
and ( n29731 , n29014 , n29730 );
or ( n29732 , n29013 , n29731 );
and ( n29733 , n28978 , n29732 );
or ( n29734 , n28977 , n29733 );
and ( n29735 , n28859 , n29734 );
or ( n29736 , n28858 , n29735 );
and ( n29737 , n28758 , n29736 );
or ( n29738 , n28757 , n29737 );
and ( n29739 , n28692 , n29738 );
or ( n29740 , n28691 , n29739 );
and ( n29741 , n28614 , n29740 );
or ( n29742 , n28613 , n29741 );
and ( n29743 , n28517 , n29742 );
or ( n29744 , n28516 , n29743 );
and ( n29745 , n28443 , n29744 );
or ( n29746 , n28442 , n29745 );
and ( n29747 , n28302 , n29746 );
or ( n29748 , n28301 , n29747 );
and ( n29749 , n28194 , n29748 );
or ( n29750 , n28193 , n29749 );
and ( n29751 , n28118 , n29750 );
or ( n29752 , n28117 , n29751 );
and ( n29753 , n27915 , n29752 );
or ( n29754 , n27914 , n29753 );
and ( n29755 , n27893 , n29754 );
or ( n29756 , n27892 , n29755 );
and ( n29757 , n27703 , n29756 );
or ( n29758 , n27702 , n29757 );
and ( n29759 , n27681 , n29758 );
or ( n29760 , n27680 , n29759 );
and ( n29761 , n27542 , n29760 );
or ( n29762 , n27541 , n29761 );
and ( n29763 , n27287 , n29762 );
or ( n29764 , n27286 , n29763 );
and ( n29765 , n27245 , n29764 );
or ( n29766 , n27244 , n29765 );
and ( n29767 , n27047 , n29766 );
or ( n29768 , n27046 , n29767 );
and ( n29769 , n26993 , n29768 );
and ( n29770 , n26991 , n29769 );
or ( n29771 , n26990 , n29770 );
and ( n29772 , n26557 , n29771 );
or ( n29773 , n26556 , n29772 );
and ( n29774 , n26297 , n29773 );
and ( n29775 , n26295 , n29774 );
and ( n29776 , n26293 , n29775 );
or ( n29777 , n26292 , n29776 );
and ( n29778 , n25941 , n29777 );
or ( n29779 , n25940 , n29778 );
and ( n29780 , n25818 , n29779 );
or ( n29781 , n25817 , n29780 );
and ( n29782 , n25492 , n29781 );
and ( n29783 , n25490 , n29782 );
or ( n29784 , n25489 , n29783 );
and ( n29785 , n25161 , n29784 );
and ( n29786 , n25159 , n29785 );
or ( n29787 , n25158 , n29786 );
and ( n29788 , n24987 , n29787 );
or ( n29789 , n24986 , n29788 );
and ( n29790 , n24872 , n29789 );
and ( n29791 , n24870 , n29790 );
and ( n29792 , n24868 , n29791 );
and ( n29793 , n24866 , n29792 );
and ( n29794 , n24864 , n29793 );
and ( n29795 , n24862 , n29794 );
and ( n29796 , n24860 , n29795 );
and ( n29797 , n24858 , n29796 );
and ( n29798 , n24856 , n29797 );
or ( n29799 , n24855 , n29798 );
and ( n29800 , n23386 , n29799 );
or ( n29801 , n23385 , n29800 );
xor ( n29802 , n23150 , n29801 );
buf ( n557067 , n29802 );
buf ( n557068 , n557067 );
xor ( n29805 , n23386 , n29799 );
buf ( n557070 , n29805 );
buf ( n557071 , n557070 );
xor ( n29808 , n24856 , n29797 );
buf ( n557073 , n29808 );
buf ( n557074 , n557073 );
xor ( n29811 , n24858 , n29796 );
buf ( n557076 , n29811 );
buf ( n557077 , n557076 );
xor ( n29814 , n24860 , n29795 );
buf ( n557079 , n29814 );
buf ( n557080 , n557079 );
xor ( n29817 , n24862 , n29794 );
buf ( n557082 , n29817 );
buf ( n557083 , n557082 );
xor ( n29820 , n24864 , n29793 );
buf ( n557085 , n29820 );
buf ( n557086 , n557085 );
xor ( n29823 , n24866 , n29792 );
buf ( n557088 , n29823 );
buf ( n557089 , n557088 );
xor ( n29826 , n24868 , n29791 );
buf ( n557091 , n29826 );
buf ( n557092 , n557091 );
xor ( n29829 , n24870 , n29790 );
buf ( n557094 , n29829 );
buf ( n557095 , n557094 );
xor ( n29832 , n24872 , n29789 );
buf ( n557097 , n29832 );
buf ( n557098 , n557097 );
xor ( n29835 , n24987 , n29787 );
buf ( n557100 , n29835 );
buf ( n557101 , n557100 );
xor ( n29838 , n25159 , n29785 );
buf ( n557103 , n29838 );
buf ( n557104 , n557103 );
xor ( n29841 , n25161 , n29784 );
buf ( n557106 , n29841 );
buf ( n557107 , n557106 );
xor ( n29844 , n25490 , n29782 );
buf ( n557109 , n29844 );
buf ( n557110 , n557109 );
xor ( n29847 , n25492 , n29781 );
buf ( n557112 , n29847 );
buf ( n557113 , n557112 );
xor ( n29850 , n25818 , n29779 );
buf ( n557115 , n29850 );
buf ( n557116 , n557115 );
xor ( n29853 , n25941 , n29777 );
buf ( n557118 , n29853 );
buf ( n557119 , n557118 );
xor ( n29856 , n26293 , n29775 );
buf ( n557121 , n29856 );
buf ( n557122 , n557121 );
xor ( n29859 , n26295 , n29774 );
buf ( n557124 , n29859 );
buf ( n557125 , n557124 );
xor ( n29862 , n26297 , n29773 );
buf ( n557127 , n29862 );
buf ( n557128 , n557127 );
xor ( n29865 , n26557 , n29771 );
buf ( n557130 , n29865 );
buf ( n557131 , n557130 );
xor ( n29868 , n26991 , n29769 );
buf ( n557133 , n29868 );
buf ( n557134 , n557133 );
xor ( n29871 , n26993 , n29768 );
buf ( n557136 , n29871 );
buf ( n557137 , n557136 );
xor ( n29874 , n27047 , n29766 );
buf ( n557139 , n29874 );
buf ( n557140 , n557139 );
xor ( n29877 , n27245 , n29764 );
buf ( n557142 , n29877 );
buf ( n557143 , n557142 );
xor ( n29880 , n27287 , n29762 );
buf ( n557145 , n29880 );
buf ( n557146 , n557145 );
xor ( n29883 , n27542 , n29760 );
buf ( n557148 , n29883 );
buf ( n557149 , n557148 );
xor ( n29886 , n27681 , n29758 );
buf ( n557151 , n29886 );
buf ( n557152 , n557151 );
xor ( n29889 , n27703 , n29756 );
buf ( n557154 , n29889 );
buf ( n557155 , n557154 );
xor ( n29892 , n27893 , n29754 );
buf ( n557157 , n29892 );
buf ( n557158 , n557157 );
xor ( n29895 , n27915 , n29752 );
buf ( n557160 , n29895 );
buf ( n557161 , n557160 );
xor ( n29898 , n28118 , n29750 );
buf ( n557163 , n29898 );
buf ( n557164 , n557163 );
xor ( n29901 , n28194 , n29748 );
buf ( n557166 , n29901 );
buf ( n557167 , n557166 );
xor ( n29904 , n28302 , n29746 );
buf ( n557169 , n29904 );
buf ( n557170 , n557169 );
xor ( n29907 , n28443 , n29744 );
buf ( n557172 , n29907 );
buf ( n557173 , n557172 );
xor ( n29910 , n28517 , n29742 );
buf ( n557175 , n29910 );
buf ( n557176 , n557175 );
xor ( n29913 , n28614 , n29740 );
buf ( n557178 , n29913 );
buf ( n557179 , n557178 );
xor ( n29916 , n28692 , n29738 );
buf ( n557181 , n29916 );
buf ( n557182 , n557181 );
xor ( n29919 , n28758 , n29736 );
buf ( n557184 , n29919 );
buf ( n557185 , n557184 );
xor ( n29922 , n28859 , n29734 );
buf ( n557187 , n29922 );
buf ( n557188 , n557187 );
xor ( n29925 , n28978 , n29732 );
buf ( n557190 , n29925 );
buf ( n557191 , n557190 );
xor ( n29928 , n29014 , n29730 );
buf ( n557193 , n29928 );
buf ( n557194 , n557193 );
xor ( n29931 , n29092 , n29728 );
buf ( n557196 , n29931 );
buf ( n557197 , n557196 );
xor ( n29934 , n29171 , n29726 );
buf ( n557199 , n29934 );
buf ( n557200 , n557199 );
xor ( n29937 , n29217 , n29724 );
buf ( n557202 , n29937 );
buf ( n557203 , n557202 );
xor ( n29940 , n29265 , n29722 );
buf ( n557205 , n29940 );
buf ( n557206 , n557205 );
xor ( n29943 , n29334 , n29720 );
buf ( n557208 , n29943 );
buf ( n557209 , n557208 );
xor ( n29946 , n29370 , n29718 );
buf ( n557211 , n29946 );
buf ( n557212 , n557211 );
xor ( n29949 , n29408 , n29716 );
buf ( n557214 , n29949 );
buf ( n557215 , n557214 );
xor ( n29952 , n29467 , n29714 );
buf ( n557217 , n29952 );
buf ( n557218 , n557217 );
xor ( n29955 , n29495 , n29712 );
buf ( n557220 , n29955 );
buf ( n557221 , n557220 );
xor ( n29958 , n29523 , n29710 );
buf ( n557223 , n29958 );
buf ( n557224 , n557223 );
xor ( n29961 , n29551 , n29708 );
buf ( n557226 , n29961 );
buf ( n557227 , n557226 );
xor ( n29964 , n29590 , n29706 );
buf ( n557229 , n29964 );
buf ( n557230 , n557229 );
xor ( n29967 , n29608 , n29704 );
buf ( n557232 , n29967 );
buf ( n557233 , n557232 );
xor ( n29970 , n29626 , n29702 );
buf ( n557235 , n29970 );
buf ( n557236 , n557235 );
xor ( n29973 , n29655 , n29700 );
buf ( n557238 , n29973 );
buf ( n557239 , n557238 );
xor ( n29976 , n29663 , n29698 );
buf ( n557241 , n29976 );
buf ( n557242 , n557241 );
xor ( n29979 , n29671 , n29696 );
buf ( n557244 , n29979 );
buf ( n557245 , n557244 );
xor ( n29982 , n29678 , n29694 );
buf ( n557247 , n29982 );
buf ( n557248 , n557247 );
xor ( n29985 , n29684 , n29692 );
buf ( n557250 , n29985 );
buf ( n557251 , n557250 );
xor ( n29988 , n29688 , n29691 );
buf ( n557253 , n29988 );
buf ( n557254 , n557253 );
buf ( n29991 , n29689 );
buf ( n557256 , n29991 );
buf ( n557257 , n557256 );
not ( n29994 , n557068 );
and ( n29995 , n543135 , n29994 );
not ( n29996 , n557071 );
and ( n29997 , n543138 , n29996 );
not ( n29998 , n557074 );
and ( n29999 , n543141 , n29998 );
not ( n30000 , n557077 );
and ( n30001 , n543144 , n30000 );
not ( n30002 , n557080 );
and ( n30003 , n543147 , n30002 );
not ( n30004 , n557083 );
and ( n30005 , n543150 , n30004 );
not ( n30006 , n557086 );
and ( n30007 , n543153 , n30006 );
not ( n30008 , n557089 );
and ( n30009 , n543156 , n30008 );
not ( n30010 , n557092 );
and ( n30011 , n543159 , n30010 );
not ( n30012 , n557095 );
and ( n30013 , n543162 , n30012 );
not ( n30014 , n557098 );
and ( n30015 , n543165 , n30014 );
not ( n30016 , n557101 );
and ( n30017 , n543168 , n30016 );
not ( n30018 , n557104 );
and ( n30019 , n543171 , n30018 );
not ( n30020 , n557107 );
and ( n30021 , n543174 , n30020 );
not ( n30022 , n557110 );
and ( n30023 , n543177 , n30022 );
not ( n30024 , n557113 );
and ( n30025 , n543180 , n30024 );
not ( n30026 , n557116 );
and ( n30027 , n543183 , n30026 );
not ( n30028 , n557119 );
and ( n30029 , n543186 , n30028 );
not ( n30030 , n557122 );
and ( n30031 , n543189 , n30030 );
not ( n30032 , n557125 );
and ( n30033 , n543192 , n30032 );
not ( n30034 , n557128 );
and ( n30035 , n543195 , n30034 );
not ( n30036 , n557131 );
and ( n30037 , n543198 , n30036 );
not ( n30038 , n557134 );
and ( n30039 , n543201 , n30038 );
not ( n30040 , n557137 );
and ( n30041 , n543204 , n30040 );
not ( n30042 , n557140 );
and ( n30043 , n543207 , n30042 );
not ( n30044 , n557143 );
and ( n30045 , n543210 , n30044 );
not ( n30046 , n557146 );
and ( n30047 , n543213 , n30046 );
not ( n30048 , n557149 );
and ( n30049 , n543216 , n30048 );
not ( n30050 , n557152 );
and ( n30051 , n543219 , n30050 );
not ( n30052 , n557155 );
and ( n30053 , n543222 , n30052 );
not ( n30054 , n557158 );
and ( n30055 , n543225 , n30054 );
not ( n30056 , n557161 );
and ( n30057 , n543228 , n30056 );
not ( n30058 , n557164 );
and ( n30059 , n543231 , n30058 );
not ( n30060 , n557167 );
and ( n30061 , n543234 , n30060 );
not ( n30062 , n557170 );
and ( n30063 , n543237 , n30062 );
not ( n30064 , n557173 );
and ( n30065 , n543240 , n30064 );
not ( n30066 , n557176 );
and ( n30067 , n543243 , n30066 );
not ( n30068 , n557179 );
and ( n30069 , n543246 , n30068 );
not ( n30070 , n557182 );
and ( n30071 , n543249 , n30070 );
not ( n30072 , n557185 );
and ( n30073 , n543252 , n30072 );
not ( n30074 , n557188 );
and ( n30075 , n543255 , n30074 );
not ( n30076 , n557191 );
and ( n30077 , n543258 , n30076 );
not ( n30078 , n557194 );
and ( n30079 , n543261 , n30078 );
not ( n30080 , n557197 );
and ( n30081 , n543264 , n30080 );
not ( n30082 , n557200 );
and ( n30083 , n543267 , n30082 );
not ( n30084 , n557203 );
and ( n30085 , n543270 , n30084 );
not ( n30086 , n557206 );
and ( n30087 , n543273 , n30086 );
not ( n30088 , n557209 );
and ( n30089 , n543276 , n30088 );
not ( n30090 , n557212 );
and ( n30091 , n543279 , n30090 );
not ( n30092 , n557215 );
and ( n30093 , n543282 , n30092 );
not ( n30094 , n557218 );
and ( n30095 , n543285 , n30094 );
not ( n30096 , n557221 );
and ( n30097 , n543288 , n30096 );
not ( n30098 , n557224 );
and ( n30099 , n543291 , n30098 );
not ( n30100 , n557227 );
and ( n30101 , n543294 , n30100 );
not ( n30102 , n557230 );
and ( n30103 , n543297 , n30102 );
not ( n30104 , n557233 );
and ( n30105 , n543300 , n30104 );
not ( n30106 , n557236 );
and ( n30107 , n543303 , n30106 );
not ( n30108 , n557239 );
and ( n30109 , n543306 , n30108 );
not ( n30110 , n557242 );
and ( n30111 , n543309 , n30110 );
not ( n30112 , n557245 );
and ( n30113 , n543312 , n30112 );
not ( n30114 , n557248 );
and ( n30115 , n543315 , n30114 );
not ( n30116 , n557251 );
and ( n30117 , n543318 , n30116 );
not ( n30118 , n557254 );
and ( n30119 , n543321 , n30118 );
not ( n30120 , n557257 );
or ( n30121 , n543324 , n30120 );
and ( n30122 , n30118 , n30121 );
and ( n30123 , n543321 , n30121 );
or ( n30124 , n30119 , n30122 , n30123 );
and ( n30125 , n30116 , n30124 );
and ( n30126 , n543318 , n30124 );
or ( n30127 , n30117 , n30125 , n30126 );
and ( n30128 , n30114 , n30127 );
and ( n30129 , n543315 , n30127 );
or ( n30130 , n30115 , n30128 , n30129 );
and ( n30131 , n30112 , n30130 );
and ( n30132 , n543312 , n30130 );
or ( n30133 , n30113 , n30131 , n30132 );
and ( n30134 , n30110 , n30133 );
and ( n30135 , n543309 , n30133 );
or ( n30136 , n30111 , n30134 , n30135 );
and ( n30137 , n30108 , n30136 );
and ( n30138 , n543306 , n30136 );
or ( n30139 , n30109 , n30137 , n30138 );
and ( n30140 , n30106 , n30139 );
and ( n30141 , n543303 , n30139 );
or ( n30142 , n30107 , n30140 , n30141 );
and ( n30143 , n30104 , n30142 );
and ( n30144 , n543300 , n30142 );
or ( n30145 , n30105 , n30143 , n30144 );
and ( n30146 , n30102 , n30145 );
and ( n30147 , n543297 , n30145 );
or ( n30148 , n30103 , n30146 , n30147 );
and ( n30149 , n30100 , n30148 );
and ( n30150 , n543294 , n30148 );
or ( n30151 , n30101 , n30149 , n30150 );
and ( n30152 , n30098 , n30151 );
and ( n30153 , n543291 , n30151 );
or ( n30154 , n30099 , n30152 , n30153 );
and ( n30155 , n30096 , n30154 );
and ( n30156 , n543288 , n30154 );
or ( n30157 , n30097 , n30155 , n30156 );
and ( n30158 , n30094 , n30157 );
and ( n30159 , n543285 , n30157 );
or ( n30160 , n30095 , n30158 , n30159 );
and ( n30161 , n30092 , n30160 );
and ( n30162 , n543282 , n30160 );
or ( n30163 , n30093 , n30161 , n30162 );
and ( n30164 , n30090 , n30163 );
and ( n30165 , n543279 , n30163 );
or ( n30166 , n30091 , n30164 , n30165 );
and ( n30167 , n30088 , n30166 );
and ( n30168 , n543276 , n30166 );
or ( n30169 , n30089 , n30167 , n30168 );
and ( n30170 , n30086 , n30169 );
and ( n30171 , n543273 , n30169 );
or ( n30172 , n30087 , n30170 , n30171 );
and ( n30173 , n30084 , n30172 );
and ( n30174 , n543270 , n30172 );
or ( n30175 , n30085 , n30173 , n30174 );
and ( n30176 , n30082 , n30175 );
and ( n30177 , n543267 , n30175 );
or ( n30178 , n30083 , n30176 , n30177 );
and ( n30179 , n30080 , n30178 );
and ( n30180 , n543264 , n30178 );
or ( n30181 , n30081 , n30179 , n30180 );
and ( n30182 , n30078 , n30181 );
and ( n30183 , n543261 , n30181 );
or ( n30184 , n30079 , n30182 , n30183 );
and ( n30185 , n30076 , n30184 );
and ( n30186 , n543258 , n30184 );
or ( n30187 , n30077 , n30185 , n30186 );
and ( n30188 , n30074 , n30187 );
and ( n30189 , n543255 , n30187 );
or ( n30190 , n30075 , n30188 , n30189 );
and ( n30191 , n30072 , n30190 );
and ( n30192 , n543252 , n30190 );
or ( n30193 , n30073 , n30191 , n30192 );
and ( n30194 , n30070 , n30193 );
and ( n30195 , n543249 , n30193 );
or ( n30196 , n30071 , n30194 , n30195 );
and ( n30197 , n30068 , n30196 );
and ( n30198 , n543246 , n30196 );
or ( n30199 , n30069 , n30197 , n30198 );
and ( n30200 , n30066 , n30199 );
and ( n30201 , n543243 , n30199 );
or ( n30202 , n30067 , n30200 , n30201 );
and ( n30203 , n30064 , n30202 );
and ( n30204 , n543240 , n30202 );
or ( n30205 , n30065 , n30203 , n30204 );
and ( n30206 , n30062 , n30205 );
and ( n30207 , n543237 , n30205 );
or ( n30208 , n30063 , n30206 , n30207 );
and ( n30209 , n30060 , n30208 );
and ( n30210 , n543234 , n30208 );
or ( n30211 , n30061 , n30209 , n30210 );
and ( n30212 , n30058 , n30211 );
and ( n30213 , n543231 , n30211 );
or ( n30214 , n30059 , n30212 , n30213 );
and ( n30215 , n30056 , n30214 );
and ( n30216 , n543228 , n30214 );
or ( n30217 , n30057 , n30215 , n30216 );
and ( n30218 , n30054 , n30217 );
and ( n30219 , n543225 , n30217 );
or ( n30220 , n30055 , n30218 , n30219 );
and ( n30221 , n30052 , n30220 );
and ( n30222 , n543222 , n30220 );
or ( n30223 , n30053 , n30221 , n30222 );
and ( n30224 , n30050 , n30223 );
and ( n30225 , n543219 , n30223 );
or ( n30226 , n30051 , n30224 , n30225 );
and ( n30227 , n30048 , n30226 );
and ( n30228 , n543216 , n30226 );
or ( n30229 , n30049 , n30227 , n30228 );
and ( n30230 , n30046 , n30229 );
and ( n30231 , n543213 , n30229 );
or ( n30232 , n30047 , n30230 , n30231 );
and ( n30233 , n30044 , n30232 );
and ( n30234 , n543210 , n30232 );
or ( n30235 , n30045 , n30233 , n30234 );
and ( n30236 , n30042 , n30235 );
and ( n30237 , n543207 , n30235 );
or ( n30238 , n30043 , n30236 , n30237 );
and ( n30239 , n30040 , n30238 );
and ( n30240 , n543204 , n30238 );
or ( n30241 , n30041 , n30239 , n30240 );
and ( n30242 , n30038 , n30241 );
and ( n30243 , n543201 , n30241 );
or ( n30244 , n30039 , n30242 , n30243 );
and ( n30245 , n30036 , n30244 );
and ( n30246 , n543198 , n30244 );
or ( n30247 , n30037 , n30245 , n30246 );
and ( n30248 , n30034 , n30247 );
and ( n30249 , n543195 , n30247 );
or ( n30250 , n30035 , n30248 , n30249 );
and ( n30251 , n30032 , n30250 );
and ( n30252 , n543192 , n30250 );
or ( n30253 , n30033 , n30251 , n30252 );
and ( n30254 , n30030 , n30253 );
and ( n30255 , n543189 , n30253 );
or ( n30256 , n30031 , n30254 , n30255 );
and ( n30257 , n30028 , n30256 );
and ( n30258 , n543186 , n30256 );
or ( n30259 , n30029 , n30257 , n30258 );
and ( n30260 , n30026 , n30259 );
and ( n30261 , n543183 , n30259 );
or ( n30262 , n30027 , n30260 , n30261 );
and ( n30263 , n30024 , n30262 );
and ( n30264 , n543180 , n30262 );
or ( n30265 , n30025 , n30263 , n30264 );
and ( n30266 , n30022 , n30265 );
and ( n30267 , n543177 , n30265 );
or ( n30268 , n30023 , n30266 , n30267 );
and ( n30269 , n30020 , n30268 );
and ( n30270 , n543174 , n30268 );
or ( n30271 , n30021 , n30269 , n30270 );
and ( n30272 , n30018 , n30271 );
and ( n30273 , n543171 , n30271 );
or ( n30274 , n30019 , n30272 , n30273 );
and ( n30275 , n30016 , n30274 );
and ( n30276 , n543168 , n30274 );
or ( n30277 , n30017 , n30275 , n30276 );
and ( n30278 , n30014 , n30277 );
and ( n30279 , n543165 , n30277 );
or ( n30280 , n30015 , n30278 , n30279 );
and ( n30281 , n30012 , n30280 );
and ( n30282 , n543162 , n30280 );
or ( n30283 , n30013 , n30281 , n30282 );
and ( n30284 , n30010 , n30283 );
and ( n30285 , n543159 , n30283 );
or ( n30286 , n30011 , n30284 , n30285 );
and ( n30287 , n30008 , n30286 );
and ( n30288 , n543156 , n30286 );
or ( n30289 , n30009 , n30287 , n30288 );
and ( n30290 , n30006 , n30289 );
and ( n30291 , n543153 , n30289 );
or ( n30292 , n30007 , n30290 , n30291 );
and ( n30293 , n30004 , n30292 );
and ( n30294 , n543150 , n30292 );
or ( n30295 , n30005 , n30293 , n30294 );
and ( n30296 , n30002 , n30295 );
and ( n30297 , n543147 , n30295 );
or ( n30298 , n30003 , n30296 , n30297 );
and ( n30299 , n30000 , n30298 );
and ( n30300 , n543144 , n30298 );
or ( n30301 , n30001 , n30299 , n30300 );
and ( n30302 , n29998 , n30301 );
and ( n30303 , n543141 , n30301 );
or ( n30304 , n29999 , n30302 , n30303 );
and ( n30305 , n29996 , n30304 );
and ( n30306 , n543138 , n30304 );
or ( n30307 , n29997 , n30305 , n30306 );
and ( n30308 , n29994 , n30307 );
and ( n30309 , n543135 , n30307 );
or ( n30310 , n29995 , n30308 , n30309 );
not ( n30311 , n30310 );
buf ( n557576 , n30311 );
xor ( n30313 , n543135 , n29994 );
xor ( n30314 , n30313 , n30307 );
buf ( n557579 , n30314 );
xor ( n30316 , n543138 , n29996 );
xor ( n30317 , n30316 , n30304 );
buf ( n557582 , n30317 );
xor ( n30319 , n543141 , n29998 );
xor ( n30320 , n30319 , n30301 );
buf ( n557585 , n30320 );
xor ( n30322 , n543144 , n30000 );
xor ( n30323 , n30322 , n30298 );
buf ( n557588 , n30323 );
xor ( n30325 , n543147 , n30002 );
xor ( n30326 , n30325 , n30295 );
buf ( n557591 , n30326 );
xor ( n30328 , n543150 , n30004 );
xor ( n30329 , n30328 , n30292 );
buf ( n557594 , n30329 );
xor ( n30331 , n543153 , n30006 );
xor ( n30332 , n30331 , n30289 );
buf ( n557597 , n30332 );
xor ( n30334 , n543156 , n30008 );
xor ( n30335 , n30334 , n30286 );
buf ( n557600 , n30335 );
xor ( n30337 , n543159 , n30010 );
xor ( n30338 , n30337 , n30283 );
buf ( n557603 , n30338 );
xor ( n30340 , n543162 , n30012 );
xor ( n30341 , n30340 , n30280 );
buf ( n557606 , n30341 );
xor ( n30343 , n543165 , n30014 );
xor ( n30344 , n30343 , n30277 );
buf ( n557609 , n30344 );
xor ( n30346 , n543168 , n30016 );
xor ( n30347 , n30346 , n30274 );
buf ( n557612 , n30347 );
xor ( n30349 , n543171 , n30018 );
xor ( n30350 , n30349 , n30271 );
buf ( n557615 , n30350 );
xor ( n30352 , n543174 , n30020 );
xor ( n30353 , n30352 , n30268 );
buf ( n557618 , n30353 );
xor ( n30355 , n543177 , n30022 );
xor ( n30356 , n30355 , n30265 );
buf ( n557621 , n30356 );
xor ( n30358 , n543180 , n30024 );
xor ( n30359 , n30358 , n30262 );
buf ( n557624 , n30359 );
xor ( n30361 , n543183 , n30026 );
xor ( n30362 , n30361 , n30259 );
buf ( n557627 , n30362 );
xor ( n30364 , n543186 , n30028 );
xor ( n30365 , n30364 , n30256 );
buf ( n557630 , n30365 );
xor ( n30367 , n543189 , n30030 );
xor ( n30368 , n30367 , n30253 );
buf ( n557633 , n30368 );
xor ( n30370 , n543192 , n30032 );
xor ( n30371 , n30370 , n30250 );
buf ( n557636 , n30371 );
xor ( n30373 , n543195 , n30034 );
xor ( n30374 , n30373 , n30247 );
buf ( n557639 , n30374 );
xor ( n30376 , n543198 , n30036 );
xor ( n30377 , n30376 , n30244 );
buf ( n557642 , n30377 );
xor ( n30379 , n543201 , n30038 );
xor ( n30380 , n30379 , n30241 );
buf ( n557645 , n30380 );
xor ( n30382 , n543204 , n30040 );
xor ( n30383 , n30382 , n30238 );
buf ( n557648 , n30383 );
xor ( n30385 , n543207 , n30042 );
xor ( n30386 , n30385 , n30235 );
buf ( n557651 , n30386 );
xor ( n30388 , n543210 , n30044 );
xor ( n30389 , n30388 , n30232 );
buf ( n557654 , n30389 );
xor ( n30391 , n543213 , n30046 );
xor ( n30392 , n30391 , n30229 );
buf ( n557657 , n30392 );
xor ( n30394 , n543216 , n30048 );
xor ( n30395 , n30394 , n30226 );
buf ( n557660 , n30395 );
xor ( n30397 , n543219 , n30050 );
xor ( n30398 , n30397 , n30223 );
buf ( n557663 , n30398 );
xor ( n30400 , n543222 , n30052 );
xor ( n30401 , n30400 , n30220 );
buf ( n557666 , n30401 );
xor ( n30403 , n543225 , n30054 );
xor ( n30404 , n30403 , n30217 );
buf ( n557669 , n30404 );
xor ( n30406 , n543228 , n30056 );
xor ( n30407 , n30406 , n30214 );
buf ( n557672 , n30407 );
xor ( n30409 , n543231 , n30058 );
xor ( n30410 , n30409 , n30211 );
buf ( n557675 , n30410 );
xor ( n30412 , n543234 , n30060 );
xor ( n30413 , n30412 , n30208 );
buf ( n557678 , n30413 );
xor ( n30415 , n543237 , n30062 );
xor ( n30416 , n30415 , n30205 );
buf ( n557681 , n30416 );
xor ( n30418 , n543240 , n30064 );
xor ( n30419 , n30418 , n30202 );
buf ( n557684 , n30419 );
xor ( n30421 , n543243 , n30066 );
xor ( n30422 , n30421 , n30199 );
buf ( n557687 , n30422 );
xor ( n30424 , n543246 , n30068 );
xor ( n30425 , n30424 , n30196 );
buf ( n557690 , n30425 );
xor ( n30427 , n543249 , n30070 );
xor ( n30428 , n30427 , n30193 );
buf ( n557693 , n30428 );
xor ( n30430 , n543252 , n30072 );
xor ( n30431 , n30430 , n30190 );
buf ( n557696 , n30431 );
xor ( n30433 , n543255 , n30074 );
xor ( n30434 , n30433 , n30187 );
buf ( n557699 , n30434 );
xor ( n30436 , n543258 , n30076 );
xor ( n30437 , n30436 , n30184 );
buf ( n557702 , n30437 );
xor ( n30439 , n543261 , n30078 );
xor ( n30440 , n30439 , n30181 );
buf ( n557705 , n30440 );
xor ( n30442 , n543264 , n30080 );
xor ( n30443 , n30442 , n30178 );
buf ( n557708 , n30443 );
xor ( n30445 , n543267 , n30082 );
xor ( n30446 , n30445 , n30175 );
buf ( n557711 , n30446 );
xor ( n30448 , n543270 , n30084 );
xor ( n30449 , n30448 , n30172 );
buf ( n557714 , n30449 );
xor ( n30451 , n543273 , n30086 );
xor ( n30452 , n30451 , n30169 );
buf ( n557717 , n30452 );
xor ( n30454 , n543276 , n30088 );
xor ( n30455 , n30454 , n30166 );
buf ( n557720 , n30455 );
xor ( n30457 , n543279 , n30090 );
xor ( n30458 , n30457 , n30163 );
buf ( n557723 , n30458 );
xor ( n30460 , n543282 , n30092 );
xor ( n30461 , n30460 , n30160 );
buf ( n557726 , n30461 );
xor ( n30463 , n543285 , n30094 );
xor ( n30464 , n30463 , n30157 );
buf ( n557729 , n30464 );
xor ( n30466 , n543288 , n30096 );
xor ( n30467 , n30466 , n30154 );
buf ( n557732 , n30467 );
xor ( n30469 , n543291 , n30098 );
xor ( n30470 , n30469 , n30151 );
buf ( n557735 , n30470 );
xor ( n30472 , n543294 , n30100 );
xor ( n30473 , n30472 , n30148 );
buf ( n557738 , n30473 );
xor ( n30475 , n543297 , n30102 );
xor ( n30476 , n30475 , n30145 );
buf ( n557741 , n30476 );
xor ( n30478 , n543300 , n30104 );
xor ( n30479 , n30478 , n30142 );
buf ( n557744 , n30479 );
xor ( n30481 , n543303 , n30106 );
xor ( n30482 , n30481 , n30139 );
buf ( n557747 , n30482 );
xor ( n30484 , n543306 , n30108 );
xor ( n30485 , n30484 , n30136 );
buf ( n557750 , n30485 );
xor ( n30487 , n543309 , n30110 );
xor ( n30488 , n30487 , n30133 );
buf ( n557753 , n30488 );
xor ( n30490 , n543312 , n30112 );
xor ( n30491 , n30490 , n30130 );
buf ( n557756 , n30491 );
xor ( n30493 , n543315 , n30114 );
xor ( n30494 , n30493 , n30127 );
buf ( n557759 , n30494 );
xor ( n30496 , n543318 , n30116 );
xor ( n30497 , n30496 , n30124 );
buf ( n557762 , n30497 );
xor ( n30499 , n543321 , n30118 );
xor ( n30500 , n30499 , n30121 );
buf ( n557765 , n30500 );
xor ( n30502 , n543324 , n557257 );
buf ( n557767 , n30502 );
buf ( n557768 , n557576 );
buf ( n557769 , n557579 );
buf ( n557770 , n557582 );
buf ( n557771 , n557585 );
buf ( n557772 , n557588 );
buf ( n557773 , n557591 );
buf ( n557774 , n557594 );
buf ( n557775 , n557597 );
buf ( n557776 , n557600 );
buf ( n557777 , n557603 );
buf ( n557778 , n557606 );
buf ( n557779 , n557609 );
buf ( n557780 , n557612 );
buf ( n557781 , n557615 );
buf ( n557782 , n557618 );
buf ( n557783 , n557621 );
buf ( n557784 , n557624 );
buf ( n557785 , n557627 );
buf ( n557786 , n557630 );
buf ( n557787 , n557633 );
buf ( n557788 , n557636 );
buf ( n557789 , n557639 );
buf ( n557790 , n557642 );
buf ( n557791 , n557645 );
buf ( n557792 , n557648 );
buf ( n557793 , n557651 );
buf ( n557794 , n557654 );
buf ( n557795 , n557657 );
buf ( n557796 , n557660 );
buf ( n557797 , n557663 );
buf ( n557798 , n557666 );
buf ( n557799 , n557669 );
buf ( n557800 , n557672 );
buf ( n557801 , n557675 );
buf ( n557802 , n557678 );
buf ( n557803 , n557681 );
buf ( n557804 , n557684 );
buf ( n557805 , n557687 );
buf ( n557806 , n557690 );
buf ( n557807 , n557693 );
buf ( n557808 , n557696 );
buf ( n557809 , n557699 );
buf ( n557810 , n557702 );
buf ( n557811 , n557705 );
buf ( n557812 , n557708 );
buf ( n557813 , n557711 );
buf ( n557814 , n557714 );
buf ( n557815 , n557717 );
buf ( n557816 , n557720 );
buf ( n557817 , n557723 );
buf ( n557818 , n557726 );
buf ( n557819 , n557729 );
buf ( n557820 , n557732 );
buf ( n557821 , n557735 );
buf ( n557822 , n557738 );
buf ( n557823 , n557741 );
buf ( n557824 , n557744 );
buf ( n557825 , n557747 );
buf ( n557826 , n557750 );
buf ( n557827 , n557753 );
buf ( n557828 , n557756 );
buf ( n557829 , n557759 );
buf ( n557830 , n557762 );
buf ( n557831 , n557765 );
buf ( n557832 , n557767 );
buf ( n557833 , n543134 );
buf ( n30570 , n557833 );
buf ( n557835 , n1218 );
buf ( n30572 , n557835 );
buf ( n30573 , n30572 );
buf ( n557838 , n543137 );
buf ( n30575 , n557838 );
and ( n30576 , n30573 , n30575 );
buf ( n557841 , n1219 );
buf ( n30578 , n557841 );
buf ( n557843 , n1218 );
buf ( n30580 , n557843 );
and ( n30581 , n30578 , n30580 );
buf ( n557846 , n1219 );
buf ( n30583 , n557846 );
and ( n30584 , n30572 , n30583 );
and ( n30585 , n30581 , n30584 );
buf ( n557850 , n543140 );
buf ( n30587 , n557850 );
and ( n30588 , n30584 , n30587 );
and ( n30589 , n30581 , n30587 );
or ( n30590 , n30585 , n30588 , n30589 );
and ( n30591 , n30575 , n30590 );
and ( n30592 , n30573 , n30590 );
or ( n30593 , n30576 , n30591 , n30592 );
and ( n30594 , n30570 , n30593 );
xor ( n30595 , n30573 , n30575 );
xor ( n30596 , n30595 , n30590 );
buf ( n557861 , n1220 );
buf ( n30598 , n557861 );
and ( n30599 , n30572 , n30598 );
buf ( n557864 , n1220 );
buf ( n30601 , n557864 );
and ( n30602 , n30601 , n30580 );
and ( n30603 , n30599 , n30602 );
xor ( n30604 , n30581 , n30584 );
xor ( n30605 , n30604 , n30587 );
and ( n30606 , n30603 , n30605 );
buf ( n30607 , n30578 );
buf ( n557872 , n543143 );
buf ( n30609 , n557872 );
and ( n30610 , n30607 , n30609 );
xor ( n30611 , n30599 , n30602 );
and ( n30612 , n30609 , n30611 );
and ( n30613 , n30607 , n30611 );
or ( n30614 , n30610 , n30612 , n30613 );
and ( n30615 , n30605 , n30614 );
and ( n30616 , n30603 , n30614 );
or ( n30617 , n30606 , n30615 , n30616 );
and ( n30618 , n30596 , n30617 );
buf ( n557883 , n1221 );
buf ( n30620 , n557883 );
and ( n30621 , n30572 , n30620 );
buf ( n557886 , n1221 );
buf ( n30623 , n557886 );
and ( n30624 , n30623 , n30580 );
and ( n30625 , n30621 , n30624 );
buf ( n557890 , n1222 );
buf ( n30627 , n557890 );
and ( n30628 , n30627 , n30580 );
and ( n30629 , n30623 , n30583 );
or ( n30630 , n30628 , n30629 );
buf ( n557895 , n1222 );
buf ( n30632 , n557895 );
and ( n30633 , n30572 , n30632 );
and ( n30634 , n30578 , n30620 );
or ( n30635 , n30633 , n30634 );
and ( n30636 , n30630 , n30635 );
and ( n30637 , n30625 , n30636 );
and ( n30638 , n30601 , n30583 );
and ( n30639 , n30578 , n30598 );
and ( n30640 , n30638 , n30639 );
xor ( n30641 , n30621 , n30624 );
and ( n30642 , n30639 , n30641 );
and ( n30643 , n30638 , n30641 );
or ( n30644 , n30640 , n30642 , n30643 );
and ( n30645 , n30636 , n30644 );
and ( n30646 , n30625 , n30644 );
or ( n30647 , n30637 , n30645 , n30646 );
xor ( n30648 , n30603 , n30605 );
xor ( n30649 , n30648 , n30614 );
and ( n30650 , n30647 , n30649 );
xor ( n30651 , n30607 , n30609 );
xor ( n30652 , n30651 , n30611 );
xnor ( n30653 , n30628 , n30629 );
xnor ( n30654 , n30633 , n30634 );
and ( n30655 , n30653 , n30654 );
not ( n30656 , n30655 );
buf ( n557921 , n543146 );
buf ( n30658 , n557921 );
and ( n30659 , n30656 , n30658 );
and ( n30660 , n30652 , n30659 );
buf ( n30661 , n30655 );
and ( n30662 , n30659 , n30661 );
and ( n30663 , n30652 , n30661 );
or ( n30664 , n30660 , n30662 , n30663 );
and ( n30665 , n30649 , n30664 );
and ( n30666 , n30647 , n30664 );
or ( n30667 , n30650 , n30665 , n30666 );
and ( n30668 , n30617 , n30667 );
and ( n30669 , n30596 , n30667 );
or ( n30670 , n30618 , n30668 , n30669 );
and ( n30671 , n30593 , n30670 );
and ( n30672 , n30570 , n30670 );
or ( n30673 , n30594 , n30671 , n30672 );
xor ( n30674 , n30570 , n30593 );
xor ( n30675 , n30674 , n30670 );
xor ( n30676 , n30596 , n30617 );
xor ( n30677 , n30676 , n30667 );
xor ( n30678 , n30630 , n30635 );
buf ( n557943 , n1223 );
buf ( n30680 , n557943 );
and ( n30681 , n30680 , n30580 );
and ( n30682 , n30627 , n30583 );
and ( n30683 , n30681 , n30682 );
buf ( n557948 , n1223 );
buf ( n30685 , n557948 );
and ( n30686 , n30572 , n30685 );
and ( n30687 , n30578 , n30632 );
and ( n30688 , n30686 , n30687 );
and ( n30689 , n30683 , n30688 );
and ( n30690 , n30678 , n30689 );
xor ( n30691 , n30638 , n30639 );
xor ( n30692 , n30691 , n30641 );
and ( n30693 , n30689 , n30692 );
and ( n30694 , n30678 , n30692 );
or ( n30695 , n30690 , n30693 , n30694 );
xor ( n30696 , n30625 , n30636 );
xor ( n30697 , n30696 , n30644 );
and ( n30698 , n30695 , n30697 );
xor ( n30699 , n30656 , n30658 );
buf ( n30700 , n30601 );
buf ( n557965 , n543149 );
buf ( n30702 , n557965 );
and ( n30703 , n30700 , n30702 );
xor ( n30704 , n30683 , n30688 );
and ( n30705 , n30702 , n30704 );
and ( n30706 , n30700 , n30704 );
or ( n30707 , n30703 , n30705 , n30706 );
and ( n30708 , n30699 , n30707 );
xor ( n30709 , n30653 , n30654 );
buf ( n557974 , n1224 );
buf ( n30711 , n557974 );
and ( n30712 , n30711 , n30580 );
and ( n30713 , n30627 , n30598 );
and ( n30714 , n30712 , n30713 );
buf ( n557979 , n1224 );
buf ( n30716 , n557979 );
and ( n30717 , n30572 , n30716 );
and ( n30718 , n30601 , n30632 );
and ( n30719 , n30717 , n30718 );
and ( n30720 , n30714 , n30719 );
and ( n30721 , n30709 , n30720 );
xor ( n30722 , n30681 , n30682 );
xor ( n30723 , n30686 , n30687 );
and ( n30724 , n30722 , n30723 );
and ( n30725 , n30720 , n30724 );
and ( n30726 , n30709 , n30724 );
or ( n30727 , n30721 , n30725 , n30726 );
and ( n30728 , n30707 , n30727 );
and ( n30729 , n30699 , n30727 );
or ( n30730 , n30708 , n30728 , n30729 );
and ( n30731 , n30697 , n30730 );
and ( n30732 , n30695 , n30730 );
or ( n30733 , n30698 , n30731 , n30732 );
xor ( n30734 , n30647 , n30649 );
xor ( n30735 , n30734 , n30664 );
and ( n30736 , n30733 , n30735 );
xor ( n30737 , n30652 , n30659 );
xor ( n30738 , n30737 , n30661 );
xor ( n30739 , n30678 , n30689 );
xor ( n30740 , n30739 , n30692 );
xor ( n30741 , n30712 , n30713 );
xor ( n30742 , n30717 , n30718 );
and ( n30743 , n30741 , n30742 );
buf ( n558008 , n543152 );
buf ( n30745 , n558008 );
and ( n30746 , n30743 , n30745 );
buf ( n558011 , n1225 );
buf ( n30748 , n558011 );
and ( n30749 , n30572 , n30748 );
and ( n30750 , n30578 , n30716 );
and ( n30751 , n30749 , n30750 );
and ( n30752 , n30601 , n30685 );
and ( n30753 , n30750 , n30752 );
and ( n30754 , n30749 , n30752 );
or ( n30755 , n30751 , n30753 , n30754 );
and ( n30756 , n30680 , n30583 );
and ( n30757 , n30755 , n30756 );
buf ( n558022 , n1225 );
buf ( n30759 , n558022 );
and ( n30760 , n30759 , n30580 );
and ( n30761 , n30711 , n30583 );
and ( n30762 , n30760 , n30761 );
and ( n30763 , n30680 , n30598 );
and ( n30764 , n30761 , n30763 );
and ( n30765 , n30760 , n30763 );
or ( n30766 , n30762 , n30764 , n30765 );
and ( n30767 , n30578 , n30685 );
and ( n30768 , n30766 , n30767 );
and ( n30769 , n30757 , n30768 );
and ( n30770 , n30746 , n30769 );
and ( n30771 , n30623 , n30598 );
and ( n30772 , n30601 , n30620 );
and ( n30773 , n30771 , n30772 );
xor ( n30774 , n30714 , n30719 );
and ( n30775 , n30772 , n30774 );
and ( n30776 , n30771 , n30774 );
or ( n30777 , n30773 , n30775 , n30776 );
and ( n30778 , n30769 , n30777 );
and ( n30779 , n30746 , n30777 );
or ( n30780 , n30770 , n30778 , n30779 );
and ( n30781 , n30740 , n30780 );
xor ( n30782 , n30699 , n30707 );
xor ( n30783 , n30782 , n30727 );
and ( n30784 , n30780 , n30783 );
and ( n30785 , n30740 , n30783 );
or ( n30786 , n30781 , n30784 , n30785 );
and ( n30787 , n30738 , n30786 );
xor ( n30788 , n30695 , n30697 );
xor ( n30789 , n30788 , n30730 );
and ( n30790 , n30786 , n30789 );
and ( n30791 , n30738 , n30789 );
or ( n30792 , n30787 , n30790 , n30791 );
and ( n30793 , n30735 , n30792 );
and ( n30794 , n30733 , n30792 );
or ( n30795 , n30736 , n30793 , n30794 );
and ( n30796 , n30677 , n30795 );
xor ( n30797 , n30733 , n30735 );
xor ( n30798 , n30797 , n30792 );
xor ( n30799 , n30738 , n30786 );
xor ( n30800 , n30799 , n30789 );
xor ( n30801 , n30700 , n30702 );
xor ( n30802 , n30801 , n30704 );
xor ( n30803 , n30709 , n30720 );
xor ( n30804 , n30803 , n30724 );
and ( n30805 , n30802 , n30804 );
xor ( n30806 , n30722 , n30723 );
xor ( n30807 , n30743 , n30745 );
and ( n30808 , n30806 , n30807 );
xor ( n30809 , n30757 , n30768 );
and ( n30810 , n30807 , n30809 );
and ( n30811 , n30806 , n30809 );
or ( n30812 , n30808 , n30810 , n30811 );
and ( n30813 , n30804 , n30812 );
and ( n30814 , n30802 , n30812 );
or ( n30815 , n30805 , n30813 , n30814 );
xor ( n30816 , n30740 , n30780 );
xor ( n30817 , n30816 , n30783 );
and ( n30818 , n30815 , n30817 );
xor ( n30819 , n30755 , n30756 );
xor ( n30820 , n30766 , n30767 );
and ( n30821 , n30819 , n30820 );
buf ( n30822 , n30623 );
buf ( n558087 , n543155 );
buf ( n30824 , n558087 );
and ( n30825 , n30822 , n30824 );
xor ( n30826 , n30741 , n30742 );
and ( n30827 , n30824 , n30826 );
and ( n30828 , n30822 , n30826 );
or ( n30829 , n30825 , n30827 , n30828 );
and ( n30830 , n30821 , n30829 );
xor ( n30831 , n30771 , n30772 );
xor ( n30832 , n30831 , n30774 );
and ( n30833 , n30829 , n30832 );
and ( n30834 , n30821 , n30832 );
or ( n30835 , n30830 , n30833 , n30834 );
xor ( n30836 , n30746 , n30769 );
xor ( n30837 , n30836 , n30777 );
and ( n30838 , n30835 , n30837 );
and ( n30839 , n30759 , n30583 );
and ( n30840 , n30680 , n30620 );
or ( n30841 , n30839 , n30840 );
and ( n30842 , n30578 , n30748 );
and ( n30843 , n30623 , n30685 );
or ( n30844 , n30842 , n30843 );
and ( n30845 , n30841 , n30844 );
xor ( n30846 , n30760 , n30761 );
xor ( n30847 , n30846 , n30763 );
xor ( n30848 , n30749 , n30750 );
xor ( n30849 , n30848 , n30752 );
and ( n30850 , n30847 , n30849 );
and ( n30851 , n30845 , n30850 );
xor ( n30852 , n30819 , n30820 );
and ( n30853 , n30850 , n30852 );
and ( n30854 , n30845 , n30852 );
or ( n30855 , n30851 , n30853 , n30854 );
xnor ( n30856 , n30839 , n30840 );
xnor ( n30857 , n30842 , n30843 );
and ( n30858 , n30856 , n30857 );
buf ( n558123 , n543158 );
buf ( n30860 , n558123 );
or ( n30861 , n30858 , n30860 );
buf ( n558126 , n1226 );
buf ( n30863 , n558126 );
and ( n30864 , n30578 , n30863 );
and ( n30865 , n30601 , n30748 );
and ( n30866 , n30864 , n30865 );
and ( n30867 , n30623 , n30716 );
and ( n30868 , n30865 , n30867 );
and ( n30869 , n30864 , n30867 );
or ( n30870 , n30866 , n30868 , n30869 );
buf ( n558135 , n1226 );
buf ( n30872 , n558135 );
and ( n30873 , n30872 , n30580 );
and ( n30874 , n30870 , n30873 );
and ( n30875 , n30711 , n30598 );
and ( n30876 , n30873 , n30875 );
and ( n30877 , n30870 , n30875 );
or ( n30878 , n30874 , n30876 , n30877 );
and ( n30879 , n30872 , n30583 );
and ( n30880 , n30759 , n30598 );
and ( n30881 , n30879 , n30880 );
and ( n30882 , n30711 , n30620 );
and ( n30883 , n30880 , n30882 );
and ( n30884 , n30879 , n30882 );
or ( n30885 , n30881 , n30883 , n30884 );
and ( n30886 , n30572 , n30863 );
and ( n30887 , n30885 , n30886 );
and ( n30888 , n30601 , n30716 );
and ( n30889 , n30886 , n30888 );
and ( n30890 , n30885 , n30888 );
or ( n30891 , n30887 , n30889 , n30890 );
and ( n30892 , n30878 , n30891 );
and ( n30893 , n30861 , n30892 );
and ( n30894 , n30627 , n30620 );
and ( n30895 , n30623 , n30632 );
and ( n30896 , n30894 , n30895 );
xor ( n30897 , n30841 , n30844 );
and ( n30898 , n30895 , n30897 );
and ( n30899 , n30894 , n30897 );
or ( n30900 , n30896 , n30898 , n30899 );
and ( n30901 , n30892 , n30900 );
and ( n30902 , n30861 , n30900 );
or ( n30903 , n30893 , n30901 , n30902 );
and ( n30904 , n30855 , n30903 );
xor ( n30905 , n30806 , n30807 );
xor ( n30906 , n30905 , n30809 );
and ( n30907 , n30903 , n30906 );
and ( n30908 , n30855 , n30906 );
or ( n30909 , n30904 , n30907 , n30908 );
and ( n30910 , n30837 , n30909 );
and ( n30911 , n30835 , n30909 );
or ( n30912 , n30838 , n30910 , n30911 );
and ( n30913 , n30817 , n30912 );
and ( n30914 , n30815 , n30912 );
or ( n30915 , n30818 , n30913 , n30914 );
and ( n30916 , n30800 , n30915 );
xor ( n30917 , n30802 , n30804 );
xor ( n30918 , n30917 , n30812 );
xor ( n30919 , n30821 , n30829 );
xor ( n30920 , n30919 , n30832 );
xor ( n30921 , n30822 , n30824 );
xor ( n30922 , n30921 , n30826 );
xor ( n30923 , n30847 , n30849 );
buf ( n30924 , n30627 );
buf ( n558189 , n543161 );
buf ( n30926 , n558189 );
and ( n30927 , n30924 , n30926 );
and ( n30928 , n30680 , n30632 );
and ( n30929 , n30627 , n30685 );
and ( n30930 , n30928 , n30929 );
buf ( n558195 , n543164 );
buf ( n30932 , n558195 );
and ( n30933 , n30929 , n30932 );
and ( n30934 , n30928 , n30932 );
or ( n30935 , n30930 , n30933 , n30934 );
and ( n30936 , n30926 , n30935 );
and ( n30937 , n30924 , n30935 );
or ( n30938 , n30927 , n30936 , n30937 );
and ( n30939 , n30923 , n30938 );
xnor ( n30940 , n30858 , n30860 );
and ( n30941 , n30938 , n30940 );
and ( n30942 , n30923 , n30940 );
or ( n30943 , n30939 , n30941 , n30942 );
and ( n30944 , n30922 , n30943 );
xor ( n30945 , n30878 , n30891 );
buf ( n558210 , n1228 );
buf ( n30947 , n558210 );
and ( n30948 , n30572 , n30947 );
buf ( n558213 , n1227 );
buf ( n30950 , n558213 );
and ( n30951 , n30578 , n30950 );
and ( n30952 , n30948 , n30951 );
and ( n30953 , n30623 , n30748 );
and ( n30954 , n30951 , n30953 );
and ( n30955 , n30948 , n30953 );
or ( n30956 , n30952 , n30954 , n30955 );
buf ( n558221 , n1227 );
buf ( n30958 , n558221 );
and ( n30959 , n30958 , n30580 );
or ( n30960 , n30956 , n30959 );
buf ( n558225 , n1228 );
buf ( n30962 , n558225 );
and ( n30963 , n30962 , n30580 );
and ( n30964 , n30958 , n30583 );
and ( n30965 , n30963 , n30964 );
and ( n30966 , n30759 , n30620 );
and ( n30967 , n30964 , n30966 );
and ( n30968 , n30963 , n30966 );
or ( n30969 , n30965 , n30967 , n30968 );
and ( n30970 , n30572 , n30950 );
or ( n30971 , n30969 , n30970 );
and ( n30972 , n30960 , n30971 );
and ( n30973 , n30945 , n30972 );
xor ( n30974 , n30870 , n30873 );
xor ( n30975 , n30974 , n30875 );
xor ( n30976 , n30885 , n30886 );
xor ( n30977 , n30976 , n30888 );
and ( n30978 , n30975 , n30977 );
and ( n30979 , n30972 , n30978 );
and ( n30980 , n30945 , n30978 );
or ( n30981 , n30973 , n30979 , n30980 );
and ( n30982 , n30943 , n30981 );
and ( n30983 , n30922 , n30981 );
or ( n30984 , n30944 , n30982 , n30983 );
and ( n30985 , n30920 , n30984 );
xor ( n30986 , n30855 , n30903 );
xor ( n30987 , n30986 , n30906 );
and ( n30988 , n30984 , n30987 );
and ( n30989 , n30920 , n30987 );
or ( n30990 , n30985 , n30988 , n30989 );
and ( n30991 , n30918 , n30990 );
xor ( n30992 , n30835 , n30837 );
xor ( n30993 , n30992 , n30909 );
and ( n30994 , n30990 , n30993 );
and ( n30995 , n30918 , n30993 );
or ( n30996 , n30991 , n30994 , n30995 );
xor ( n30997 , n30815 , n30817 );
xor ( n30998 , n30997 , n30912 );
and ( n30999 , n30996 , n30998 );
xor ( n31000 , n30918 , n30990 );
xor ( n31001 , n31000 , n30993 );
xor ( n31002 , n30845 , n30850 );
xor ( n31003 , n31002 , n30852 );
xor ( n31004 , n30861 , n30892 );
xor ( n31005 , n31004 , n30900 );
and ( n31006 , n31003 , n31005 );
xor ( n31007 , n30856 , n30857 );
and ( n31008 , n30872 , n30598 );
and ( n31009 , n30711 , n30632 );
or ( n31010 , n31008 , n31009 );
and ( n31011 , n30601 , n30863 );
and ( n31012 , n30627 , n30716 );
or ( n31013 , n31011 , n31012 );
and ( n31014 , n31010 , n31013 );
and ( n31015 , n31007 , n31014 );
xor ( n31016 , n30879 , n30880 );
xor ( n31017 , n31016 , n30882 );
xor ( n31018 , n30864 , n30865 );
xor ( n31019 , n31018 , n30867 );
and ( n31020 , n31017 , n31019 );
and ( n31021 , n31014 , n31020 );
and ( n31022 , n31007 , n31020 );
or ( n31023 , n31015 , n31021 , n31022 );
xor ( n31024 , n30894 , n30895 );
xor ( n31025 , n31024 , n30897 );
and ( n31026 , n31023 , n31025 );
xor ( n31027 , n30924 , n30926 );
xor ( n31028 , n31027 , n30935 );
xor ( n31029 , n30960 , n30971 );
and ( n31030 , n31028 , n31029 );
xor ( n31031 , n30975 , n30977 );
and ( n31032 , n31029 , n31031 );
and ( n31033 , n31028 , n31031 );
or ( n31034 , n31030 , n31032 , n31033 );
and ( n31035 , n31025 , n31034 );
and ( n31036 , n31023 , n31034 );
or ( n31037 , n31026 , n31035 , n31036 );
and ( n31038 , n31005 , n31037 );
and ( n31039 , n31003 , n31037 );
or ( n31040 , n31006 , n31038 , n31039 );
xor ( n31041 , n30920 , n30984 );
xor ( n31042 , n31041 , n30987 );
and ( n31043 , n31040 , n31042 );
xnor ( n31044 , n30956 , n30959 );
xnor ( n31045 , n30969 , n30970 );
and ( n31046 , n31044 , n31045 );
xor ( n31047 , n30928 , n30929 );
xor ( n31048 , n31047 , n30932 );
xor ( n31049 , n31010 , n31013 );
and ( n31050 , n31048 , n31049 );
xor ( n31051 , n31017 , n31019 );
and ( n31052 , n31049 , n31051 );
and ( n31053 , n31048 , n31051 );
or ( n31054 , n31050 , n31052 , n31053 );
and ( n31055 , n31046 , n31054 );
buf ( n558320 , n1229 );
buf ( n31057 , n558320 );
and ( n31058 , n31057 , n30580 );
and ( n31059 , n30872 , n30620 );
and ( n31060 , n31058 , n31059 );
and ( n31061 , n30759 , n30632 );
and ( n31062 , n31059 , n31061 );
and ( n31063 , n31058 , n31061 );
or ( n31064 , n31060 , n31062 , n31063 );
buf ( n558329 , n1229 );
buf ( n31066 , n558329 );
and ( n31067 , n30572 , n31066 );
and ( n31068 , n30623 , n30863 );
and ( n31069 , n31067 , n31068 );
and ( n31070 , n30627 , n30748 );
and ( n31071 , n31068 , n31070 );
and ( n31072 , n31067 , n31070 );
or ( n31073 , n31069 , n31071 , n31072 );
and ( n31074 , n31064 , n31073 );
and ( n31075 , n30962 , n30583 );
and ( n31076 , n30958 , n30598 );
or ( n31077 , n31075 , n31076 );
and ( n31078 , n30578 , n30947 );
and ( n31079 , n30601 , n30950 );
or ( n31080 , n31078 , n31079 );
and ( n31081 , n31077 , n31080 );
and ( n31082 , n31074 , n31081 );
xor ( n31083 , n30963 , n30964 );
xor ( n31084 , n31083 , n30966 );
xor ( n31085 , n30948 , n30951 );
xor ( n31086 , n31085 , n30953 );
and ( n31087 , n31084 , n31086 );
and ( n31088 , n31081 , n31087 );
and ( n31089 , n31074 , n31087 );
or ( n31090 , n31082 , n31088 , n31089 );
and ( n31091 , n31054 , n31090 );
and ( n31092 , n31046 , n31090 );
or ( n31093 , n31055 , n31091 , n31092 );
xor ( n31094 , n30923 , n30938 );
xor ( n31095 , n31094 , n30940 );
and ( n31096 , n31093 , n31095 );
xor ( n31097 , n30945 , n30972 );
xor ( n31098 , n31097 , n30978 );
and ( n31099 , n31095 , n31098 );
and ( n31100 , n31093 , n31098 );
or ( n31101 , n31096 , n31099 , n31100 );
xor ( n31102 , n30922 , n30943 );
xor ( n31103 , n31102 , n30981 );
and ( n31104 , n31101 , n31103 );
xor ( n31105 , n31007 , n31014 );
xor ( n31106 , n31105 , n31020 );
xnor ( n31107 , n31008 , n31009 );
xnor ( n31108 , n31011 , n31012 );
and ( n31109 , n31107 , n31108 );
xor ( n31110 , n31044 , n31045 );
and ( n31111 , n31109 , n31110 );
and ( n31112 , n30578 , n31066 );
and ( n31113 , n30601 , n30947 );
and ( n31114 , n31112 , n31113 );
and ( n31115 , n30627 , n30863 );
and ( n31116 , n31113 , n31115 );
and ( n31117 , n31112 , n31115 );
or ( n31118 , n31114 , n31116 , n31117 );
xor ( n31119 , n31067 , n31068 );
xor ( n31120 , n31119 , n31070 );
or ( n31121 , n31118 , n31120 );
and ( n31122 , n31057 , n30583 );
and ( n31123 , n30962 , n30598 );
and ( n31124 , n31122 , n31123 );
and ( n31125 , n30872 , n30632 );
and ( n31126 , n31123 , n31125 );
and ( n31127 , n31122 , n31125 );
or ( n31128 , n31124 , n31126 , n31127 );
xor ( n31129 , n31058 , n31059 );
xor ( n31130 , n31129 , n31061 );
or ( n31131 , n31128 , n31130 );
and ( n31132 , n31121 , n31131 );
and ( n31133 , n31110 , n31132 );
and ( n31134 , n31109 , n31132 );
or ( n31135 , n31111 , n31133 , n31134 );
and ( n31136 , n31106 , n31135 );
buf ( n31137 , n30680 );
buf ( n558402 , n543167 );
buf ( n31139 , n558402 );
and ( n31140 , n31137 , n31139 );
xor ( n31141 , n31064 , n31073 );
and ( n31142 , n31139 , n31141 );
and ( n31143 , n31137 , n31141 );
or ( n31144 , n31140 , n31142 , n31143 );
xor ( n31145 , n31077 , n31080 );
xor ( n31146 , n31084 , n31086 );
and ( n31147 , n31145 , n31146 );
xor ( n31148 , n31107 , n31108 );
and ( n31149 , n31146 , n31148 );
and ( n31150 , n31145 , n31148 );
or ( n31151 , n31147 , n31149 , n31150 );
and ( n31152 , n31144 , n31151 );
and ( n31153 , n30958 , n30620 );
and ( n31154 , n30759 , n30685 );
or ( n31155 , n31153 , n31154 );
and ( n31156 , n30623 , n30950 );
and ( n31157 , n30680 , n30748 );
or ( n31158 , n31156 , n31157 );
and ( n31159 , n31155 , n31158 );
xnor ( n31160 , n31075 , n31076 );
xnor ( n31161 , n31078 , n31079 );
and ( n31162 , n31160 , n31161 );
and ( n31163 , n31159 , n31162 );
and ( n31164 , n30711 , n30685 );
and ( n31165 , n30680 , n30716 );
and ( n31166 , n31164 , n31165 );
buf ( n558431 , n1230 );
buf ( n31168 , n558431 );
and ( n31169 , n30572 , n31168 );
buf ( n558434 , n1230 );
buf ( n31171 , n558434 );
and ( n31172 , n31171 , n30580 );
and ( n31173 , n31169 , n31172 );
and ( n31174 , n31165 , n31173 );
and ( n31175 , n31164 , n31173 );
or ( n31176 , n31166 , n31174 , n31175 );
and ( n31177 , n31162 , n31176 );
and ( n31178 , n31159 , n31176 );
or ( n31179 , n31163 , n31177 , n31178 );
and ( n31180 , n31151 , n31179 );
and ( n31181 , n31144 , n31179 );
or ( n31182 , n31152 , n31180 , n31181 );
and ( n31183 , n31135 , n31182 );
and ( n31184 , n31106 , n31182 );
or ( n31185 , n31136 , n31183 , n31184 );
xor ( n31186 , n31023 , n31025 );
xor ( n31187 , n31186 , n31034 );
and ( n31188 , n31185 , n31187 );
xor ( n31189 , n31093 , n31095 );
xor ( n31190 , n31189 , n31098 );
and ( n31191 , n31187 , n31190 );
and ( n31192 , n31185 , n31190 );
or ( n31193 , n31188 , n31191 , n31192 );
and ( n31194 , n31103 , n31193 );
and ( n31195 , n31101 , n31193 );
or ( n31196 , n31104 , n31194 , n31195 );
and ( n31197 , n31042 , n31196 );
and ( n31198 , n31040 , n31196 );
or ( n31199 , n31043 , n31197 , n31198 );
and ( n31200 , n31001 , n31199 );
xor ( n31201 , n31040 , n31042 );
xor ( n31202 , n31201 , n31196 );
xor ( n31203 , n31003 , n31005 );
xor ( n31204 , n31203 , n31037 );
xor ( n31205 , n31101 , n31103 );
xor ( n31206 , n31205 , n31193 );
and ( n31207 , n31204 , n31206 );
xor ( n31208 , n31028 , n31029 );
xor ( n31209 , n31208 , n31031 );
xor ( n31210 , n31046 , n31054 );
xor ( n31211 , n31210 , n31090 );
and ( n31212 , n31209 , n31211 );
xor ( n31213 , n31048 , n31049 );
xor ( n31214 , n31213 , n31051 );
xor ( n31215 , n31074 , n31081 );
xor ( n31216 , n31215 , n31087 );
and ( n31217 , n31214 , n31216 );
xor ( n31218 , n31121 , n31131 );
xnor ( n31219 , n31153 , n31154 );
xnor ( n31220 , n31156 , n31157 );
and ( n31221 , n31219 , n31220 );
not ( n31222 , n31221 );
buf ( n558487 , n543170 );
buf ( n31224 , n558487 );
and ( n31225 , n31222 , n31224 );
and ( n31226 , n31218 , n31225 );
buf ( n31227 , n31221 );
and ( n31228 , n31225 , n31227 );
and ( n31229 , n31218 , n31227 );
or ( n31230 , n31226 , n31228 , n31229 );
and ( n31231 , n31216 , n31230 );
and ( n31232 , n31214 , n31230 );
or ( n31233 , n31217 , n31231 , n31232 );
and ( n31234 , n31211 , n31233 );
and ( n31235 , n31209 , n31233 );
or ( n31236 , n31212 , n31234 , n31235 );
xor ( n31237 , n31185 , n31187 );
xor ( n31238 , n31237 , n31190 );
and ( n31239 , n31236 , n31238 );
and ( n31240 , n30601 , n31066 );
and ( n31241 , n30623 , n30947 );
and ( n31242 , n31240 , n31241 );
and ( n31243 , n30627 , n30950 );
and ( n31244 , n31241 , n31243 );
and ( n31245 , n31240 , n31243 );
or ( n31246 , n31242 , n31244 , n31245 );
xor ( n31247 , n31112 , n31113 );
xor ( n31248 , n31247 , n31115 );
or ( n31249 , n31246 , n31248 );
and ( n31250 , n31057 , n30598 );
and ( n31251 , n30962 , n30620 );
and ( n31252 , n31250 , n31251 );
and ( n31253 , n30958 , n30632 );
and ( n31254 , n31251 , n31253 );
and ( n31255 , n31250 , n31253 );
or ( n31256 , n31252 , n31254 , n31255 );
xor ( n31257 , n31122 , n31123 );
xor ( n31258 , n31257 , n31125 );
or ( n31259 , n31256 , n31258 );
and ( n31260 , n31249 , n31259 );
xnor ( n31261 , n31118 , n31120 );
xnor ( n31262 , n31128 , n31130 );
and ( n31263 , n31261 , n31262 );
and ( n31264 , n31260 , n31263 );
xor ( n31265 , n31155 , n31158 );
xor ( n31266 , n31160 , n31161 );
and ( n31267 , n31265 , n31266 );
buf ( n558532 , n1231 );
buf ( n31269 , n558532 );
and ( n31270 , n31269 , n30580 );
and ( n31271 , n31171 , n30583 );
and ( n31272 , n31270 , n31271 );
and ( n31273 , n30872 , n30685 );
and ( n31274 , n31271 , n31273 );
and ( n31275 , n31270 , n31273 );
or ( n31276 , n31272 , n31274 , n31275 );
buf ( n558541 , n1231 );
buf ( n31278 , n558541 );
and ( n31279 , n30572 , n31278 );
and ( n31280 , n30578 , n31168 );
and ( n31281 , n31279 , n31280 );
and ( n31282 , n30680 , n30863 );
and ( n31283 , n31280 , n31282 );
and ( n31284 , n31279 , n31282 );
or ( n31285 , n31281 , n31283 , n31284 );
and ( n31286 , n31276 , n31285 );
and ( n31287 , n31266 , n31286 );
and ( n31288 , n31265 , n31286 );
or ( n31289 , n31267 , n31287 , n31288 );
and ( n31290 , n31263 , n31289 );
and ( n31291 , n31260 , n31289 );
or ( n31292 , n31264 , n31290 , n31291 );
xor ( n31293 , n31137 , n31139 );
xor ( n31294 , n31293 , n31141 );
xor ( n31295 , n31145 , n31146 );
xor ( n31296 , n31295 , n31148 );
and ( n31297 , n31294 , n31296 );
xor ( n31298 , n31159 , n31162 );
xor ( n31299 , n31298 , n31176 );
and ( n31300 , n31296 , n31299 );
and ( n31301 , n31294 , n31299 );
or ( n31302 , n31297 , n31300 , n31301 );
and ( n31303 , n31292 , n31302 );
xor ( n31304 , n31109 , n31110 );
xor ( n31305 , n31304 , n31132 );
and ( n31306 , n31302 , n31305 );
and ( n31307 , n31292 , n31305 );
or ( n31308 , n31303 , n31306 , n31307 );
xor ( n31309 , n31106 , n31135 );
xor ( n31310 , n31309 , n31182 );
and ( n31311 , n31308 , n31310 );
xor ( n31312 , n31144 , n31151 );
xor ( n31313 , n31312 , n31179 );
buf ( n31314 , n30711 );
buf ( n558579 , n543173 );
buf ( n31316 , n558579 );
and ( n31317 , n31314 , n31316 );
xor ( n31318 , n31169 , n31172 );
and ( n31319 , n31316 , n31318 );
and ( n31320 , n31314 , n31318 );
or ( n31321 , n31317 , n31319 , n31320 );
xor ( n31322 , n31164 , n31165 );
xor ( n31323 , n31322 , n31173 );
and ( n31324 , n31321 , n31323 );
xor ( n31325 , n31222 , n31224 );
and ( n31326 , n31323 , n31325 );
and ( n31327 , n31321 , n31325 );
or ( n31328 , n31324 , n31326 , n31327 );
xor ( n31329 , n31249 , n31259 );
xor ( n31330 , n31261 , n31262 );
and ( n31331 , n31329 , n31330 );
xnor ( n31332 , n31246 , n31248 );
xnor ( n31333 , n31256 , n31258 );
and ( n31334 , n31332 , n31333 );
and ( n31335 , n31330 , n31334 );
and ( n31336 , n31329 , n31334 );
or ( n31337 , n31331 , n31335 , n31336 );
and ( n31338 , n31328 , n31337 );
xor ( n31339 , n31218 , n31225 );
xor ( n31340 , n31339 , n31227 );
and ( n31341 , n31337 , n31340 );
and ( n31342 , n31328 , n31340 );
or ( n31343 , n31338 , n31341 , n31342 );
and ( n31344 , n31313 , n31343 );
xor ( n31345 , n31214 , n31216 );
xor ( n31346 , n31345 , n31230 );
and ( n31347 , n31343 , n31346 );
and ( n31348 , n31313 , n31346 );
or ( n31349 , n31344 , n31347 , n31348 );
and ( n31350 , n31310 , n31349 );
and ( n31351 , n31308 , n31349 );
or ( n31352 , n31311 , n31350 , n31351 );
and ( n31353 , n31238 , n31352 );
and ( n31354 , n31236 , n31352 );
or ( n31355 , n31239 , n31353 , n31354 );
and ( n31356 , n31206 , n31355 );
and ( n31357 , n31204 , n31355 );
or ( n31358 , n31207 , n31356 , n31357 );
or ( n31359 , n31202 , n31358 );
and ( n31360 , n31199 , n31359 );
and ( n31361 , n31001 , n31359 );
or ( n31362 , n31200 , n31360 , n31361 );
and ( n31363 , n30998 , n31362 );
and ( n31364 , n30996 , n31362 );
or ( n31365 , n30999 , n31363 , n31364 );
and ( n31366 , n30915 , n31365 );
and ( n31367 , n30800 , n31365 );
or ( n31368 , n30916 , n31366 , n31367 );
or ( n31369 , n30798 , n31368 );
and ( n31370 , n30795 , n31369 );
and ( n31371 , n30677 , n31369 );
or ( n31372 , n30796 , n31370 , n31371 );
or ( n31373 , n30675 , n31372 );
xor ( n31374 , n30673 , n31373 );
not ( n31375 , n31374 );
xnor ( n31376 , n30675 , n31372 );
xor ( n31377 , n30677 , n30795 );
xor ( n31378 , n31377 , n31369 );
not ( n31379 , n31378 );
xnor ( n31380 , n30798 , n31368 );
xor ( n31381 , n30800 , n30915 );
xor ( n31382 , n31381 , n31365 );
xor ( n31383 , n30996 , n30998 );
xor ( n31384 , n31383 , n31362 );
not ( n31385 , n31384 );
xor ( n31386 , n31001 , n31199 );
xor ( n31387 , n31386 , n31359 );
not ( n31388 , n31387 );
xnor ( n31389 , n31202 , n31358 );
xor ( n31390 , n31204 , n31206 );
xor ( n31391 , n31390 , n31355 );
xor ( n31392 , n31209 , n31211 );
xor ( n31393 , n31392 , n31233 );
xor ( n31394 , n31292 , n31302 );
xor ( n31395 , n31394 , n31305 );
xor ( n31396 , n31260 , n31263 );
xor ( n31397 , n31396 , n31289 );
xor ( n31398 , n31294 , n31296 );
xor ( n31399 , n31398 , n31299 );
and ( n31400 , n31397 , n31399 );
xor ( n31401 , n31276 , n31285 );
xor ( n31402 , n31219 , n31220 );
and ( n31403 , n31401 , n31402 );
buf ( n558668 , n1232 );
buf ( n31405 , n558668 );
and ( n31406 , n31405 , n30580 );
and ( n31407 , n31057 , n30620 );
and ( n31408 , n31406 , n31407 );
and ( n31409 , n30958 , n30685 );
and ( n31410 , n31407 , n31409 );
and ( n31411 , n31406 , n31409 );
or ( n31412 , n31408 , n31410 , n31411 );
buf ( n558677 , n1232 );
buf ( n31414 , n558677 );
and ( n31415 , n30572 , n31414 );
and ( n31416 , n30623 , n31066 );
and ( n31417 , n31415 , n31416 );
and ( n31418 , n30680 , n30950 );
and ( n31419 , n31416 , n31418 );
and ( n31420 , n31415 , n31418 );
or ( n31421 , n31417 , n31419 , n31420 );
and ( n31422 , n31412 , n31421 );
and ( n31423 , n31402 , n31422 );
and ( n31424 , n31401 , n31422 );
or ( n31425 , n31403 , n31423 , n31424 );
xor ( n31426 , n31265 , n31266 );
xor ( n31427 , n31426 , n31286 );
and ( n31428 , n31425 , n31427 );
buf ( n558693 , n1233 );
buf ( n31430 , n558693 );
and ( n31431 , n31430 , n30580 );
and ( n31432 , n31057 , n30632 );
and ( n31433 , n31431 , n31432 );
and ( n31434 , n30962 , n30685 );
and ( n31435 , n31432 , n31434 );
and ( n31436 , n31431 , n31434 );
or ( n31437 , n31433 , n31435 , n31436 );
and ( n31438 , n30578 , n31278 );
and ( n31439 , n31437 , n31438 );
and ( n31440 , n30601 , n31168 );
and ( n31441 , n31438 , n31440 );
and ( n31442 , n31437 , n31440 );
or ( n31443 , n31439 , n31441 , n31442 );
xor ( n31444 , n31250 , n31251 );
xor ( n31445 , n31444 , n31253 );
and ( n31446 , n31443 , n31445 );
xor ( n31447 , n31270 , n31271 );
xor ( n31448 , n31447 , n31273 );
and ( n31449 , n31445 , n31448 );
and ( n31450 , n31443 , n31448 );
or ( n31451 , n31446 , n31449 , n31450 );
buf ( n558716 , n1233 );
buf ( n31453 , n558716 );
and ( n31454 , n30572 , n31453 );
and ( n31455 , n30627 , n31066 );
and ( n31456 , n31454 , n31455 );
and ( n31457 , n30680 , n30947 );
and ( n31458 , n31455 , n31457 );
and ( n31459 , n31454 , n31457 );
or ( n31460 , n31456 , n31458 , n31459 );
and ( n31461 , n31269 , n30583 );
and ( n31462 , n31460 , n31461 );
and ( n31463 , n31171 , n30598 );
and ( n31464 , n31461 , n31463 );
and ( n31465 , n31460 , n31463 );
or ( n31466 , n31462 , n31464 , n31465 );
xor ( n31467 , n31240 , n31241 );
xor ( n31468 , n31467 , n31243 );
and ( n31469 , n31466 , n31468 );
xor ( n31470 , n31279 , n31280 );
xor ( n31471 , n31470 , n31282 );
and ( n31472 , n31468 , n31471 );
and ( n31473 , n31466 , n31471 );
or ( n31474 , n31469 , n31472 , n31473 );
and ( n31475 , n31451 , n31474 );
and ( n31476 , n31427 , n31475 );
and ( n31477 , n31425 , n31475 );
or ( n31478 , n31428 , n31476 , n31477 );
and ( n31479 , n31399 , n31478 );
and ( n31480 , n31397 , n31478 );
or ( n31481 , n31400 , n31479 , n31480 );
and ( n31482 , n31395 , n31481 );
xor ( n31483 , n31313 , n31343 );
xor ( n31484 , n31483 , n31346 );
and ( n31485 , n31481 , n31484 );
and ( n31486 , n31395 , n31484 );
or ( n31487 , n31482 , n31485 , n31486 );
and ( n31488 , n31393 , n31487 );
xor ( n31489 , n31308 , n31310 );
xor ( n31490 , n31489 , n31349 );
and ( n31491 , n31487 , n31490 );
and ( n31492 , n31393 , n31490 );
or ( n31493 , n31488 , n31491 , n31492 );
xor ( n31494 , n31236 , n31238 );
xor ( n31495 , n31494 , n31352 );
and ( n31496 , n31493 , n31495 );
xor ( n31497 , n31393 , n31487 );
xor ( n31498 , n31497 , n31490 );
and ( n31499 , n30962 , n30632 );
and ( n31500 , n30872 , n30716 );
and ( n31501 , n31499 , n31500 );
and ( n31502 , n30627 , n30947 );
and ( n31503 , n30711 , n30863 );
and ( n31504 , n31502 , n31503 );
and ( n31505 , n31501 , n31504 );
xor ( n31506 , n31314 , n31316 );
xor ( n31507 , n31506 , n31318 );
and ( n31508 , n31505 , n31507 );
xor ( n31509 , n31332 , n31333 );
and ( n31510 , n31507 , n31509 );
and ( n31511 , n31505 , n31509 );
or ( n31512 , n31508 , n31510 , n31511 );
xor ( n31513 , n31499 , n31500 );
xor ( n31514 , n31502 , n31503 );
and ( n31515 , n31513 , n31514 );
buf ( n558780 , n543176 );
buf ( n31517 , n558780 );
and ( n31518 , n31515 , n31517 );
and ( n31519 , n30759 , n30716 );
and ( n31520 , n30711 , n30748 );
and ( n31521 , n31519 , n31520 );
xor ( n31522 , n31412 , n31421 );
and ( n31523 , n31520 , n31522 );
and ( n31524 , n31519 , n31522 );
or ( n31525 , n31521 , n31523 , n31524 );
and ( n31526 , n31518 , n31525 );
xor ( n31527 , n31501 , n31504 );
and ( n31528 , n31405 , n30583 );
and ( n31529 , n31269 , n30598 );
and ( n31530 , n31528 , n31529 );
and ( n31531 , n30958 , n30716 );
and ( n31532 , n31529 , n31531 );
and ( n31533 , n31528 , n31531 );
or ( n31534 , n31530 , n31532 , n31533 );
and ( n31535 , n30578 , n31414 );
and ( n31536 , n30601 , n31278 );
and ( n31537 , n31535 , n31536 );
and ( n31538 , n30711 , n30950 );
and ( n31539 , n31536 , n31538 );
and ( n31540 , n31535 , n31538 );
or ( n31541 , n31537 , n31539 , n31540 );
and ( n31542 , n31534 , n31541 );
and ( n31543 , n31527 , n31542 );
buf ( n31544 , n30759 );
buf ( n558809 , n543179 );
buf ( n31546 , n558809 );
and ( n31547 , n31544 , n31546 );
and ( n31548 , n30623 , n31168 );
and ( n31549 , n31171 , n30620 );
and ( n31550 , n31548 , n31549 );
and ( n31551 , n31546 , n31550 );
and ( n31552 , n31544 , n31550 );
or ( n31553 , n31547 , n31551 , n31552 );
and ( n31554 , n31542 , n31553 );
and ( n31555 , n31527 , n31553 );
or ( n31556 , n31543 , n31554 , n31555 );
and ( n31557 , n31525 , n31556 );
and ( n31558 , n31518 , n31556 );
or ( n31559 , n31526 , n31557 , n31558 );
and ( n31560 , n31512 , n31559 );
xor ( n31561 , n31321 , n31323 );
xor ( n31562 , n31561 , n31325 );
and ( n31563 , n31559 , n31562 );
and ( n31564 , n31512 , n31562 );
or ( n31565 , n31560 , n31563 , n31564 );
xor ( n31566 , n31328 , n31337 );
xor ( n31567 , n31566 , n31340 );
and ( n31568 , n31565 , n31567 );
xor ( n31569 , n31329 , n31330 );
xor ( n31570 , n31569 , n31334 );
xor ( n31571 , n31401 , n31402 );
xor ( n31572 , n31571 , n31422 );
xor ( n31573 , n31451 , n31474 );
and ( n31574 , n31572 , n31573 );
xor ( n31575 , n31415 , n31416 );
xor ( n31576 , n31575 , n31418 );
xor ( n31577 , n31437 , n31438 );
xor ( n31578 , n31577 , n31440 );
and ( n31579 , n31576 , n31578 );
xor ( n31580 , n31406 , n31407 );
xor ( n31581 , n31580 , n31409 );
xor ( n31582 , n31460 , n31461 );
xor ( n31583 , n31582 , n31463 );
and ( n31584 , n31581 , n31583 );
and ( n31585 , n31579 , n31584 );
and ( n31586 , n31573 , n31585 );
and ( n31587 , n31572 , n31585 );
or ( n31588 , n31574 , n31586 , n31587 );
and ( n31589 , n31570 , n31588 );
xor ( n31590 , n31443 , n31445 );
xor ( n31591 , n31590 , n31448 );
xor ( n31592 , n31466 , n31468 );
xor ( n31593 , n31592 , n31471 );
and ( n31594 , n31591 , n31593 );
xor ( n31595 , n31515 , n31517 );
buf ( n558860 , n1234 );
buf ( n31597 , n558860 );
and ( n31598 , n30572 , n31597 );
and ( n31599 , n30578 , n31453 );
and ( n31600 , n31598 , n31599 );
and ( n31601 , n30627 , n31168 );
and ( n31602 , n31599 , n31601 );
and ( n31603 , n31598 , n31601 );
or ( n31604 , n31600 , n31602 , n31603 );
and ( n31605 , n30601 , n31414 );
and ( n31606 , n30623 , n31278 );
and ( n31607 , n31605 , n31606 );
and ( n31608 , n30711 , n30947 );
and ( n31609 , n31606 , n31608 );
and ( n31610 , n31605 , n31608 );
or ( n31611 , n31607 , n31609 , n31610 );
and ( n31612 , n31604 , n31611 );
xor ( n31613 , n31528 , n31529 );
xor ( n31614 , n31613 , n31531 );
and ( n31615 , n31611 , n31614 );
and ( n31616 , n31604 , n31614 );
or ( n31617 , n31612 , n31615 , n31616 );
buf ( n558882 , n1234 );
buf ( n31619 , n558882 );
and ( n31620 , n31619 , n30580 );
and ( n31621 , n31430 , n30583 );
and ( n31622 , n31620 , n31621 );
and ( n31623 , n31171 , n30632 );
and ( n31624 , n31621 , n31623 );
and ( n31625 , n31620 , n31623 );
or ( n31626 , n31622 , n31624 , n31625 );
and ( n31627 , n31405 , n30598 );
and ( n31628 , n31269 , n30620 );
and ( n31629 , n31627 , n31628 );
and ( n31630 , n30962 , n30716 );
and ( n31631 , n31628 , n31630 );
and ( n31632 , n31627 , n31630 );
or ( n31633 , n31629 , n31631 , n31632 );
and ( n31634 , n31626 , n31633 );
xor ( n31635 , n31535 , n31536 );
xor ( n31636 , n31635 , n31538 );
and ( n31637 , n31633 , n31636 );
and ( n31638 , n31626 , n31636 );
or ( n31639 , n31634 , n31637 , n31638 );
and ( n31640 , n31617 , n31639 );
and ( n31641 , n31595 , n31640 );
xor ( n31642 , n31534 , n31541 );
xor ( n31643 , n31513 , n31514 );
and ( n31644 , n31642 , n31643 );
and ( n31645 , n31057 , n30685 );
and ( n31646 , n30958 , n30748 );
or ( n31647 , n31645 , n31646 );
and ( n31648 , n30680 , n31066 );
and ( n31649 , n30759 , n30950 );
or ( n31650 , n31648 , n31649 );
and ( n31651 , n31647 , n31650 );
and ( n31652 , n31643 , n31651 );
and ( n31653 , n31642 , n31651 );
or ( n31654 , n31644 , n31652 , n31653 );
and ( n31655 , n31640 , n31654 );
and ( n31656 , n31595 , n31654 );
or ( n31657 , n31641 , n31655 , n31656 );
and ( n31658 , n31594 , n31657 );
xor ( n31659 , n31431 , n31432 );
xor ( n31660 , n31659 , n31434 );
xor ( n31661 , n31454 , n31455 );
xor ( n31662 , n31661 , n31457 );
and ( n31663 , n31660 , n31662 );
and ( n31664 , n30872 , n30748 );
and ( n31665 , n30759 , n30863 );
and ( n31666 , n31664 , n31665 );
xor ( n31667 , n31548 , n31549 );
and ( n31668 , n31665 , n31667 );
and ( n31669 , n31664 , n31667 );
or ( n31670 , n31666 , n31668 , n31669 );
and ( n31671 , n31663 , n31670 );
xor ( n31672 , n31544 , n31546 );
xor ( n31673 , n31672 , n31550 );
and ( n31674 , n31670 , n31673 );
and ( n31675 , n31663 , n31673 );
or ( n31676 , n31671 , n31674 , n31675 );
xor ( n31677 , n31519 , n31520 );
xor ( n31678 , n31677 , n31522 );
and ( n31679 , n31676 , n31678 );
xor ( n31680 , n31527 , n31542 );
xor ( n31681 , n31680 , n31553 );
and ( n31682 , n31678 , n31681 );
and ( n31683 , n31676 , n31681 );
or ( n31684 , n31679 , n31682 , n31683 );
and ( n31685 , n31657 , n31684 );
and ( n31686 , n31594 , n31684 );
or ( n31687 , n31658 , n31685 , n31686 );
and ( n31688 , n31588 , n31687 );
and ( n31689 , n31570 , n31687 );
or ( n31690 , n31589 , n31688 , n31689 );
and ( n31691 , n31567 , n31690 );
and ( n31692 , n31565 , n31690 );
or ( n31693 , n31568 , n31691 , n31692 );
xor ( n31694 , n31395 , n31481 );
xor ( n31695 , n31694 , n31484 );
and ( n31696 , n31693 , n31695 );
xor ( n31697 , n31397 , n31399 );
xor ( n31698 , n31697 , n31478 );
xor ( n31699 , n31425 , n31427 );
xor ( n31700 , n31699 , n31475 );
xor ( n31701 , n31512 , n31559 );
xor ( n31702 , n31701 , n31562 );
and ( n31703 , n31700 , n31702 );
xor ( n31704 , n31505 , n31507 );
xor ( n31705 , n31704 , n31509 );
xor ( n31706 , n31518 , n31525 );
xor ( n31707 , n31706 , n31556 );
and ( n31708 , n31705 , n31707 );
xor ( n31709 , n31579 , n31584 );
xor ( n31710 , n31591 , n31593 );
and ( n31711 , n31709 , n31710 );
xor ( n31712 , n31576 , n31578 );
xor ( n31713 , n31581 , n31583 );
and ( n31714 , n31712 , n31713 );
and ( n31715 , n31710 , n31714 );
and ( n31716 , n31709 , n31714 );
or ( n31717 , n31711 , n31715 , n31716 );
and ( n31718 , n31707 , n31717 );
and ( n31719 , n31705 , n31717 );
or ( n31720 , n31708 , n31718 , n31719 );
and ( n31721 , n31702 , n31720 );
and ( n31722 , n31700 , n31720 );
or ( n31723 , n31703 , n31721 , n31722 );
and ( n31724 , n31698 , n31723 );
xor ( n31725 , n31565 , n31567 );
xor ( n31726 , n31725 , n31690 );
and ( n31727 , n31723 , n31726 );
and ( n31728 , n31698 , n31726 );
or ( n31729 , n31724 , n31727 , n31728 );
and ( n31730 , n31695 , n31729 );
and ( n31731 , n31693 , n31729 );
or ( n31732 , n31696 , n31730 , n31731 );
and ( n31733 , n31498 , n31732 );
xor ( n31734 , n31693 , n31695 );
xor ( n31735 , n31734 , n31729 );
xor ( n31736 , n31617 , n31639 );
xnor ( n31737 , n31645 , n31646 );
xnor ( n31738 , n31648 , n31649 );
and ( n31739 , n31737 , n31738 );
buf ( n559004 , n543182 );
buf ( n31741 , n559004 );
or ( n31742 , n31739 , n31741 );
and ( n31743 , n31736 , n31742 );
xor ( n31744 , n31598 , n31599 );
xor ( n31745 , n31744 , n31601 );
xor ( n31746 , n31605 , n31606 );
xor ( n31747 , n31746 , n31608 );
or ( n31748 , n31745 , n31747 );
xor ( n31749 , n31620 , n31621 );
xor ( n31750 , n31749 , n31623 );
xor ( n31751 , n31627 , n31628 );
xor ( n31752 , n31751 , n31630 );
or ( n31753 , n31750 , n31752 );
and ( n31754 , n31748 , n31753 );
and ( n31755 , n31742 , n31754 );
and ( n31756 , n31736 , n31754 );
or ( n31757 , n31743 , n31755 , n31756 );
and ( n31758 , n30601 , n31453 );
and ( n31759 , n30623 , n31414 );
and ( n31760 , n31758 , n31759 );
and ( n31761 , n30759 , n30947 );
and ( n31762 , n31759 , n31761 );
and ( n31763 , n31758 , n31761 );
or ( n31764 , n31760 , n31762 , n31763 );
buf ( n559029 , n1235 );
buf ( n31766 , n559029 );
and ( n31767 , n30572 , n31766 );
and ( n31768 , n30578 , n31597 );
and ( n31769 , n31767 , n31768 );
and ( n31770 , n30711 , n31066 );
and ( n31771 , n31768 , n31770 );
and ( n31772 , n31767 , n31770 );
or ( n31773 , n31769 , n31771 , n31772 );
or ( n31774 , n31764 , n31773 );
and ( n31775 , n31430 , n30598 );
and ( n31776 , n31405 , n30620 );
and ( n31777 , n31775 , n31776 );
and ( n31778 , n30962 , n30748 );
and ( n31779 , n31776 , n31778 );
and ( n31780 , n31775 , n31778 );
or ( n31781 , n31777 , n31779 , n31780 );
buf ( n559046 , n1235 );
buf ( n31783 , n559046 );
and ( n31784 , n31783 , n30580 );
and ( n31785 , n31619 , n30583 );
and ( n31786 , n31784 , n31785 );
and ( n31787 , n31057 , n30716 );
and ( n31788 , n31785 , n31787 );
and ( n31789 , n31784 , n31787 );
or ( n31790 , n31786 , n31788 , n31789 );
or ( n31791 , n31781 , n31790 );
and ( n31792 , n31774 , n31791 );
xor ( n31793 , n31604 , n31611 );
xor ( n31794 , n31793 , n31614 );
xor ( n31795 , n31626 , n31633 );
xor ( n31796 , n31795 , n31636 );
and ( n31797 , n31794 , n31796 );
and ( n31798 , n31792 , n31797 );
xor ( n31799 , n31647 , n31650 );
xor ( n31800 , n31660 , n31662 );
and ( n31801 , n31799 , n31800 );
and ( n31802 , n31269 , n30632 );
and ( n31803 , n31171 , n30685 );
or ( n31804 , n31802 , n31803 );
and ( n31805 , n30627 , n31278 );
and ( n31806 , n30680 , n31168 );
or ( n31807 , n31805 , n31806 );
and ( n31808 , n31804 , n31807 );
and ( n31809 , n31800 , n31808 );
and ( n31810 , n31799 , n31808 );
or ( n31811 , n31801 , n31809 , n31810 );
and ( n31812 , n31797 , n31811 );
and ( n31813 , n31792 , n31811 );
or ( n31814 , n31798 , n31812 , n31813 );
and ( n31815 , n31757 , n31814 );
xor ( n31816 , n31595 , n31640 );
xor ( n31817 , n31816 , n31654 );
and ( n31818 , n31814 , n31817 );
and ( n31819 , n31757 , n31817 );
or ( n31820 , n31815 , n31818 , n31819 );
xor ( n31821 , n31572 , n31573 );
xor ( n31822 , n31821 , n31585 );
and ( n31823 , n31820 , n31822 );
xor ( n31824 , n31594 , n31657 );
xor ( n31825 , n31824 , n31684 );
and ( n31826 , n31822 , n31825 );
and ( n31827 , n31820 , n31825 );
or ( n31828 , n31823 , n31826 , n31827 );
xor ( n31829 , n31570 , n31588 );
xor ( n31830 , n31829 , n31687 );
and ( n31831 , n31828 , n31830 );
xor ( n31832 , n31676 , n31678 );
xor ( n31833 , n31832 , n31681 );
xor ( n31834 , n31642 , n31643 );
xor ( n31835 , n31834 , n31651 );
xor ( n31836 , n31663 , n31670 );
xor ( n31837 , n31836 , n31673 );
and ( n31838 , n31835 , n31837 );
xor ( n31839 , n31712 , n31713 );
and ( n31840 , n31837 , n31839 );
and ( n31841 , n31835 , n31839 );
or ( n31842 , n31838 , n31840 , n31841 );
and ( n31843 , n31833 , n31842 );
xor ( n31844 , n31664 , n31665 );
xor ( n31845 , n31844 , n31667 );
xnor ( n31846 , n31739 , n31741 );
and ( n31847 , n31845 , n31846 );
xor ( n31848 , n31748 , n31753 );
and ( n31849 , n31846 , n31848 );
and ( n31850 , n31845 , n31848 );
or ( n31851 , n31847 , n31849 , n31850 );
xor ( n31852 , n31774 , n31791 );
xor ( n31853 , n31794 , n31796 );
and ( n31854 , n31852 , n31853 );
xor ( n31855 , n31758 , n31759 );
xor ( n31856 , n31855 , n31761 );
xor ( n31857 , n31767 , n31768 );
xor ( n31858 , n31857 , n31770 );
or ( n31859 , n31856 , n31858 );
xor ( n31860 , n31775 , n31776 );
xor ( n31861 , n31860 , n31778 );
xor ( n31862 , n31784 , n31785 );
xor ( n31863 , n31862 , n31787 );
or ( n31864 , n31861 , n31863 );
and ( n31865 , n31859 , n31864 );
and ( n31866 , n31853 , n31865 );
and ( n31867 , n31852 , n31865 );
or ( n31868 , n31854 , n31866 , n31867 );
and ( n31869 , n31851 , n31868 );
buf ( n559134 , n1236 );
buf ( n31871 , n559134 );
and ( n31872 , n30572 , n31871 );
and ( n31873 , n30627 , n31414 );
and ( n31874 , n31872 , n31873 );
and ( n31875 , n30759 , n31066 );
and ( n31876 , n31873 , n31875 );
and ( n31877 , n31872 , n31875 );
or ( n31878 , n31874 , n31876 , n31877 );
and ( n31879 , n30578 , n31766 );
and ( n31880 , n30601 , n31597 );
and ( n31881 , n31879 , n31880 );
and ( n31882 , n30680 , n31278 );
and ( n31883 , n31880 , n31882 );
and ( n31884 , n31879 , n31882 );
or ( n31885 , n31881 , n31883 , n31884 );
or ( n31886 , n31878 , n31885 );
buf ( n559151 , n1236 );
buf ( n31888 , n559151 );
and ( n31889 , n31888 , n30580 );
and ( n31890 , n31405 , n30632 );
and ( n31891 , n31889 , n31890 );
and ( n31892 , n31057 , n30748 );
and ( n31893 , n31890 , n31892 );
and ( n31894 , n31889 , n31892 );
or ( n31895 , n31891 , n31893 , n31894 );
and ( n31896 , n31783 , n30583 );
and ( n31897 , n31619 , n30598 );
and ( n31898 , n31896 , n31897 );
and ( n31899 , n31269 , n30685 );
and ( n31900 , n31897 , n31899 );
and ( n31901 , n31896 , n31899 );
or ( n31902 , n31898 , n31900 , n31901 );
or ( n31903 , n31895 , n31902 );
and ( n31904 , n31886 , n31903 );
xnor ( n31905 , n31745 , n31747 );
xnor ( n31906 , n31750 , n31752 );
and ( n31907 , n31905 , n31906 );
and ( n31908 , n31904 , n31907 );
xnor ( n31909 , n31764 , n31773 );
xnor ( n31910 , n31781 , n31790 );
and ( n31911 , n31909 , n31910 );
and ( n31912 , n31907 , n31911 );
and ( n31913 , n31904 , n31911 );
or ( n31914 , n31908 , n31912 , n31913 );
and ( n31915 , n31868 , n31914 );
and ( n31916 , n31851 , n31914 );
or ( n31917 , n31869 , n31915 , n31916 );
and ( n31918 , n31842 , n31917 );
and ( n31919 , n31833 , n31917 );
or ( n31920 , n31843 , n31918 , n31919 );
buf ( n31921 , n30872 );
buf ( n559186 , n543185 );
buf ( n31923 , n559186 );
and ( n31924 , n31921 , n31923 );
xor ( n31925 , n31804 , n31807 );
and ( n31926 , n31923 , n31925 );
and ( n31927 , n31921 , n31925 );
or ( n31928 , n31924 , n31926 , n31927 );
xor ( n31929 , n31737 , n31738 );
and ( n31930 , n31171 , n30716 );
and ( n31931 , n30962 , n30863 );
and ( n31932 , n31930 , n31931 );
and ( n31933 , n30711 , n31168 );
and ( n31934 , n30872 , n30947 );
and ( n31935 , n31933 , n31934 );
and ( n31936 , n31932 , n31935 );
and ( n31937 , n31929 , n31936 );
xnor ( n31938 , n31802 , n31803 );
xnor ( n31939 , n31805 , n31806 );
and ( n31940 , n31938 , n31939 );
and ( n31941 , n31936 , n31940 );
and ( n31942 , n31929 , n31940 );
or ( n31943 , n31937 , n31941 , n31942 );
and ( n31944 , n31928 , n31943 );
xor ( n31945 , n31799 , n31800 );
xor ( n31946 , n31945 , n31808 );
and ( n31947 , n31943 , n31946 );
and ( n31948 , n31928 , n31946 );
or ( n31949 , n31944 , n31947 , n31948 );
xor ( n31950 , n31736 , n31742 );
xor ( n31951 , n31950 , n31754 );
and ( n31952 , n31949 , n31951 );
xor ( n31953 , n31792 , n31797 );
xor ( n31954 , n31953 , n31811 );
and ( n31955 , n31951 , n31954 );
and ( n31956 , n31949 , n31954 );
or ( n31957 , n31952 , n31955 , n31956 );
xor ( n31958 , n31709 , n31710 );
xor ( n31959 , n31958 , n31714 );
and ( n31960 , n31957 , n31959 );
xor ( n31961 , n31757 , n31814 );
xor ( n31962 , n31961 , n31817 );
and ( n31963 , n31959 , n31962 );
and ( n31964 , n31957 , n31962 );
or ( n31965 , n31960 , n31963 , n31964 );
and ( n31966 , n31920 , n31965 );
xor ( n31967 , n31705 , n31707 );
xor ( n31968 , n31967 , n31717 );
and ( n31969 , n31965 , n31968 );
and ( n31970 , n31920 , n31968 );
or ( n31971 , n31966 , n31969 , n31970 );
and ( n31972 , n31830 , n31971 );
and ( n31973 , n31828 , n31971 );
or ( n31974 , n31831 , n31972 , n31973 );
xor ( n31975 , n31698 , n31723 );
xor ( n31976 , n31975 , n31726 );
and ( n31977 , n31974 , n31976 );
xor ( n31978 , n31700 , n31702 );
xor ( n31979 , n31978 , n31720 );
xor ( n31980 , n31820 , n31822 );
xor ( n31981 , n31980 , n31825 );
xor ( n31982 , n31859 , n31864 );
xor ( n31983 , n31886 , n31903 );
and ( n31984 , n31982 , n31983 );
xor ( n31985 , n31905 , n31906 );
and ( n31986 , n31983 , n31985 );
and ( n31987 , n31982 , n31985 );
or ( n31988 , n31984 , n31986 , n31987 );
xor ( n31989 , n31909 , n31910 );
xor ( n31990 , n31930 , n31931 );
xor ( n31991 , n31933 , n31934 );
and ( n31992 , n31990 , n31991 );
buf ( n559257 , n543188 );
buf ( n31993 , n559257 );
and ( n31994 , n31992 , n31993 );
and ( n31995 , n31989 , n31994 );
buf ( n559261 , n1237 );
buf ( n31997 , n559261 );
and ( n31998 , n30572 , n31997 );
and ( n31999 , n30680 , n31414 );
and ( n32000 , n31998 , n31999 );
and ( n32001 , n30711 , n31278 );
and ( n32002 , n31999 , n32001 );
and ( n32003 , n31998 , n32001 );
or ( n32004 , n32000 , n32002 , n32003 );
and ( n32005 , n30578 , n31871 );
and ( n32006 , n30601 , n31766 );
and ( n32007 , n32005 , n32006 );
and ( n32008 , n30759 , n31168 );
and ( n32009 , n32006 , n32008 );
and ( n32010 , n32005 , n32008 );
or ( n32011 , n32007 , n32009 , n32010 );
and ( n32012 , n32004 , n32011 );
xor ( n32013 , n31889 , n31890 );
xor ( n32014 , n32013 , n31892 );
and ( n32015 , n32011 , n32014 );
and ( n32016 , n32004 , n32014 );
or ( n32017 , n32012 , n32015 , n32016 );
buf ( n559283 , n1237 );
buf ( n32019 , n559283 );
and ( n32020 , n32019 , n30580 );
and ( n32021 , n31405 , n30685 );
and ( n32022 , n32020 , n32021 );
and ( n32023 , n31269 , n30716 );
and ( n32024 , n32021 , n32023 );
and ( n32025 , n32020 , n32023 );
or ( n32026 , n32022 , n32024 , n32025 );
and ( n32027 , n31888 , n30583 );
and ( n32028 , n31783 , n30598 );
and ( n32029 , n32027 , n32028 );
and ( n559295 , n31171 , n30748 );
and ( n559296 , n32028 , n559295 );
and ( n559297 , n32027 , n559295 );
or ( n559298 , n32029 , n559296 , n559297 );
and ( n559299 , n32026 , n559298 );
xor ( n559300 , n31872 , n31873 );
xor ( n32030 , n559300 , n31875 );
and ( n32031 , n559298 , n32030 );
and ( n32032 , n32026 , n32030 );
or ( n32033 , n559299 , n32031 , n32032 );
and ( n32034 , n32017 , n32033 );
and ( n32035 , n31994 , n32034 );
and ( n32036 , n31989 , n32034 );
or ( n32037 , n31995 , n32035 , n32036 );
and ( n32038 , n31988 , n32037 );
and ( n32039 , n30623 , n31597 );
and ( n559311 , n30627 , n31453 );
and ( n559312 , n32039 , n559311 );
and ( n32040 , n30872 , n31066 );
and ( n32041 , n559311 , n32040 );
and ( n32042 , n32039 , n32040 );
or ( n32043 , n559312 , n32041 , n32042 );
and ( n32044 , n31430 , n30620 );
or ( n32045 , n32043 , n32044 );
and ( n32046 , n31619 , n30620 );
and ( n32047 , n31430 , n30632 );
and ( n32048 , n32046 , n32047 );
and ( n32049 , n31057 , n30863 );
and ( n32050 , n32047 , n32049 );
and ( n32051 , n32046 , n32049 );
or ( n32052 , n32048 , n32050 , n32051 );
and ( n32053 , n30623 , n31453 );
or ( n32054 , n32052 , n32053 );
and ( n32055 , n32045 , n32054 );
xnor ( n32056 , n31856 , n31858 );
xnor ( n32057 , n31861 , n31863 );
and ( n32058 , n32056 , n32057 );
and ( n32059 , n32055 , n32058 );
xnor ( n32060 , n31878 , n31885 );
xnor ( n32061 , n31895 , n31902 );
and ( n32062 , n32060 , n32061 );
and ( n32063 , n32058 , n32062 );
and ( n32064 , n32055 , n32062 );
or ( n32065 , n32059 , n32063 , n32064 );
and ( n32066 , n32037 , n32065 );
and ( n32067 , n31988 , n32065 );
or ( n32068 , n32038 , n32066 , n32067 );
and ( n32069 , n30958 , n30863 );
and ( n32070 , n30872 , n30950 );
and ( n32071 , n32069 , n32070 );
xor ( n32072 , n31932 , n31935 );
and ( n32073 , n32070 , n32072 );
and ( n32074 , n32069 , n32072 );
or ( n32075 , n32071 , n32073 , n32074 );
xor ( n32076 , n31921 , n31923 );
xor ( n32077 , n32076 , n31925 );
and ( n32078 , n32075 , n32077 );
xor ( n32079 , n31929 , n31936 );
xor ( n32080 , n32079 , n31940 );
and ( n32081 , n32077 , n32080 );
and ( n32082 , n32075 , n32080 );
or ( n32083 , n32078 , n32081 , n32082 );
xor ( n32084 , n31845 , n31846 );
xor ( n32085 , n32084 , n31848 );
and ( n32086 , n32083 , n32085 );
xor ( n32087 , n31852 , n31853 );
xor ( n32088 , n32087 , n31865 );
and ( n32089 , n32085 , n32088 );
and ( n32090 , n32083 , n32088 );
or ( n32091 , n32086 , n32089 , n32090 );
and ( n32092 , n32068 , n32091 );
xor ( n32093 , n31835 , n31837 );
xor ( n32094 , n32093 , n31839 );
and ( n32095 , n32091 , n32094 );
and ( n32096 , n32068 , n32094 );
or ( n32097 , n32092 , n32095 , n32096 );
xor ( n32098 , n31833 , n31842 );
xor ( n32099 , n32098 , n31917 );
and ( n32100 , n32097 , n32099 );
xor ( n32101 , n31957 , n31959 );
xor ( n32102 , n32101 , n31962 );
and ( n32103 , n32099 , n32102 );
and ( n32104 , n32097 , n32102 );
or ( n32105 , n32100 , n32103 , n32104 );
and ( n32106 , n31981 , n32105 );
xor ( n32107 , n31920 , n31965 );
xor ( n32108 , n32107 , n31968 );
and ( n32109 , n32105 , n32108 );
and ( n32110 , n31981 , n32108 );
or ( n32111 , n32106 , n32109 , n32110 );
and ( n32112 , n31979 , n32111 );
xor ( n32113 , n31828 , n31830 );
xor ( n32114 , n32113 , n31971 );
and ( n32115 , n32111 , n32114 );
and ( n32116 , n31979 , n32114 );
or ( n32117 , n32112 , n32115 , n32116 );
and ( n32118 , n31976 , n32117 );
and ( n32119 , n31974 , n32117 );
or ( n32120 , n31977 , n32118 , n32119 );
or ( n32121 , n31735 , n32120 );
and ( n32122 , n31732 , n32121 );
and ( n32123 , n31498 , n32121 );
or ( n32124 , n31733 , n32122 , n32123 );
and ( n32125 , n31495 , n32124 );
and ( n32126 , n31493 , n32124 );
or ( n32127 , n31496 , n32125 , n32126 );
and ( n32128 , n31391 , n32127 );
xor ( n32129 , n31391 , n32127 );
xor ( n32130 , n31493 , n31495 );
xor ( n32131 , n32130 , n32124 );
xor ( n32132 , n31498 , n31732 );
xor ( n32133 , n32132 , n32121 );
not ( n32134 , n32133 );
xnor ( n32135 , n31735 , n32120 );
xor ( n32136 , n31974 , n31976 );
xor ( n32137 , n32136 , n32117 );
xor ( n32138 , n31979 , n32111 );
xor ( n32139 , n32138 , n32114 );
xor ( n32140 , n31981 , n32105 );
xor ( n32141 , n32140 , n32108 );
xor ( n32142 , n31851 , n31868 );
xor ( n32143 , n32142 , n31914 );
xor ( n32144 , n31949 , n31951 );
xor ( n32145 , n32144 , n31954 );
and ( n32146 , n32143 , n32145 );
xor ( n32147 , n31904 , n31907 );
xor ( n32148 , n32147 , n31911 );
xor ( n32149 , n31928 , n31943 );
xor ( n32150 , n32149 , n31946 );
and ( n32151 , n32148 , n32150 );
xor ( n32152 , n31896 , n31897 );
xor ( n32153 , n32152 , n31899 );
xor ( n32154 , n31879 , n31880 );
xor ( n32155 , n32154 , n31882 );
and ( n32156 , n32153 , n32155 );
xor ( n32157 , n31992 , n31993 );
and ( n32158 , n32156 , n32157 );
and ( n32159 , n31888 , n30598 );
and ( n32160 , n31783 , n30620 );
and ( n32161 , n32159 , n32160 );
and ( n32162 , n31405 , n30716 );
and ( n32163 , n32160 , n32162 );
and ( n32164 , n32159 , n32162 );
or ( n32165 , n32161 , n32163 , n32164 );
xor ( n32166 , n32005 , n32006 );
xor ( n32167 , n32166 , n32008 );
and ( n32168 , n32165 , n32167 );
xor ( n32169 , n32039 , n559311 );
xor ( n32170 , n32169 , n32040 );
and ( n32171 , n32167 , n32170 );
and ( n32172 , n32165 , n32170 );
or ( n32173 , n32168 , n32171 , n32172 );
xor ( n32174 , n32026 , n559298 );
xor ( n32175 , n32174 , n32030 );
and ( n32176 , n32173 , n32175 );
and ( n32177 , n30601 , n31871 );
and ( n32178 , n30623 , n31766 );
and ( n32179 , n32177 , n32178 );
and ( n32180 , n30711 , n31414 );
and ( n32181 , n32178 , n32180 );
and ( n32182 , n32177 , n32180 );
or ( n32183 , n32179 , n32181 , n32182 );
xor ( n32184 , n32027 , n32028 );
xor ( n32185 , n32184 , n559295 );
and ( n32186 , n32183 , n32185 );
xor ( n32187 , n32046 , n32047 );
xor ( n32188 , n32187 , n32049 );
and ( n32189 , n32185 , n32188 );
and ( n32190 , n32183 , n32188 );
or ( n32191 , n32186 , n32189 , n32190 );
xor ( n32192 , n32004 , n32011 );
xor ( n32193 , n32192 , n32014 );
and ( n32194 , n32191 , n32193 );
and ( n32195 , n32176 , n32194 );
and ( n32196 , n32158 , n32195 );
xor ( n32197 , n31938 , n31939 );
xor ( n32198 , n32017 , n32033 );
and ( n32199 , n32197 , n32198 );
xor ( n32200 , n32045 , n32054 );
and ( n32201 , n32198 , n32200 );
and ( n32202 , n32197 , n32200 );
or ( n32203 , n32199 , n32201 , n32202 );
and ( n32204 , n32195 , n32203 );
and ( n32205 , n32158 , n32203 );
or ( n32206 , n32196 , n32204 , n32205 );
and ( n32207 , n32150 , n32206 );
and ( n32208 , n32148 , n32206 );
or ( n32209 , n32151 , n32207 , n32208 );
and ( n32210 , n32145 , n32209 );
and ( n32211 , n32143 , n32209 );
or ( n32212 , n32146 , n32210 , n32211 );
xor ( n32213 , n32097 , n32099 );
xor ( n32214 , n32213 , n32102 );
and ( n32215 , n32212 , n32214 );
xor ( n32216 , n32056 , n32057 );
xor ( n32217 , n32060 , n32061 );
and ( n32218 , n32216 , n32217 );
xnor ( n32219 , n32043 , n32044 );
xnor ( n32220 , n32052 , n32053 );
and ( n32221 , n32219 , n32220 );
and ( n32222 , n32217 , n32221 );
and ( n32223 , n32216 , n32221 );
or ( n32224 , n32218 , n32222 , n32223 );
buf ( n32225 , n30958 );
buf ( n559499 , n543191 );
buf ( n32227 , n559499 );
and ( n32228 , n32225 , n32227 );
xor ( n32229 , n32153 , n32155 );
and ( n32230 , n32227 , n32229 );
and ( n32231 , n32225 , n32229 );
or ( n32232 , n32228 , n32230 , n32231 );
xor ( n32233 , n31990 , n31991 );
buf ( n559507 , n1238 );
buf ( n32235 , n559507 );
and ( n32236 , n32235 , n30580 );
and ( n32237 , n32019 , n30583 );
and ( n32238 , n32236 , n32237 );
and ( n32239 , n31171 , n30863 );
and ( n32240 , n32237 , n32239 );
and ( n32241 , n32236 , n32239 );
or ( n32242 , n32238 , n32240 , n32241 );
buf ( n559516 , n1238 );
buf ( n32244 , n559516 );
and ( n32245 , n30572 , n32244 );
and ( n32246 , n30578 , n31997 );
and ( n32247 , n32245 , n32246 );
and ( n32248 , n30872 , n31168 );
and ( n32249 , n32246 , n32248 );
and ( n32250 , n32245 , n32248 );
or ( n32251 , n32247 , n32249 , n32250 );
and ( n32252 , n32242 , n32251 );
and ( n32253 , n32233 , n32252 );
and ( n32254 , n31269 , n30748 );
not ( n32255 , n32254 );
and ( n32256 , n31057 , n30950 );
and ( n32257 , n32255 , n32256 );
and ( n32258 , n30759 , n31278 );
not ( n32259 , n32258 );
and ( n32260 , n30958 , n31066 );
and ( n32261 , n32259 , n32260 );
and ( n32262 , n32257 , n32261 );
and ( n32263 , n32252 , n32262 );
and ( n32264 , n32233 , n32262 );
or ( n32265 , n32253 , n32263 , n32264 );
and ( n32266 , n32232 , n32265 );
xor ( n32267 , n32069 , n32070 );
xor ( n32268 , n32267 , n32072 );
and ( n32269 , n32265 , n32268 );
and ( n32270 , n32232 , n32268 );
or ( n32271 , n32266 , n32269 , n32270 );
and ( n32272 , n32224 , n32271 );
xor ( n32273 , n31982 , n31983 );
xor ( n32274 , n32273 , n31985 );
and ( n32275 , n32271 , n32274 );
and ( n32276 , n32224 , n32274 );
or ( n32277 , n32272 , n32275 , n32276 );
xor ( n32278 , n31989 , n31994 );
xor ( n32279 , n32278 , n32034 );
xor ( n32280 , n32055 , n32058 );
xor ( n32281 , n32280 , n32062 );
and ( n32282 , n32279 , n32281 );
xor ( n32283 , n32075 , n32077 );
xor ( n32284 , n32283 , n32080 );
and ( n32285 , n32281 , n32284 );
and ( n32286 , n32279 , n32284 );
or ( n32287 , n32282 , n32285 , n32286 );
and ( n32288 , n32277 , n32287 );
xor ( n32289 , n31988 , n32037 );
xor ( n32290 , n32289 , n32065 );
and ( n32291 , n32287 , n32290 );
and ( n32292 , n32277 , n32290 );
or ( n32293 , n32288 , n32291 , n32292 );
xor ( n32294 , n32068 , n32091 );
xor ( n32295 , n32294 , n32094 );
and ( n559569 , n32293 , n32295 );
xor ( n32296 , n32083 , n32085 );
xor ( n32297 , n32296 , n32088 );
xor ( n32298 , n32156 , n32157 );
xor ( n32299 , n32176 , n32194 );
and ( n32300 , n32298 , n32299 );
buf ( n559575 , n1239 );
buf ( n32302 , n559575 );
and ( n32303 , n32302 , n30580 );
and ( n32304 , n32235 , n30583 );
and ( n32305 , n32303 , n32304 );
and ( n32306 , n31405 , n30748 );
and ( n32307 , n32304 , n32306 );
and ( n32308 , n32303 , n32306 );
or ( n32309 , n32305 , n32307 , n32308 );
and ( n32310 , n30627 , n31597 );
and ( n32311 , n32309 , n32310 );
and ( n32312 , n30680 , n31453 );
and ( n32313 , n32310 , n32312 );
and ( n32314 , n32309 , n32312 );
or ( n32315 , n32311 , n32313 , n32314 );
xor ( n32316 , n31998 , n31999 );
xor ( n32317 , n32316 , n32001 );
or ( n32318 , n32315 , n32317 );
buf ( n559593 , n1239 );
buf ( n32320 , n559593 );
and ( n32321 , n30572 , n32320 );
and ( n32322 , n30578 , n32244 );
and ( n32323 , n32321 , n32322 );
and ( n32324 , n30759 , n31414 );
and ( n32325 , n32322 , n32324 );
and ( n32326 , n32321 , n32324 );
or ( n32327 , n32323 , n32325 , n32326 );
and ( n32328 , n31619 , n30632 );
and ( n32329 , n32327 , n32328 );
and ( n32330 , n31430 , n30685 );
and ( n32331 , n32328 , n32330 );
and ( n32332 , n32327 , n32330 );
or ( n32333 , n32329 , n32331 , n32332 );
xor ( n32334 , n32020 , n32021 );
xor ( n32335 , n32334 , n32023 );
or ( n32336 , n32333 , n32335 );
and ( n32337 , n32318 , n32336 );
and ( n32338 , n32299 , n32337 );
and ( n32339 , n32298 , n32337 );
or ( n32340 , n32300 , n32338 , n32339 );
xor ( n32341 , n32173 , n32175 );
xor ( n32342 , n32191 , n32193 );
and ( n32343 , n32341 , n32342 );
buf ( n32344 , n32254 );
buf ( n32345 , n32258 );
and ( n32346 , n32344 , n32345 );
xor ( n32347 , n32219 , n32220 );
and ( n32348 , n32346 , n32347 );
xor ( n32349 , n32245 , n32246 );
xor ( n32350 , n32349 , n32248 );
xor ( n32351 , n32177 , n32178 );
xor ( n32352 , n32351 , n32180 );
or ( n32353 , n32350 , n32352 );
xor ( n32354 , n32236 , n32237 );
xor ( n32355 , n32354 , n32239 );
xor ( n32356 , n32159 , n32160 );
xor ( n32357 , n32356 , n32162 );
or ( n32358 , n32355 , n32357 );
and ( n32359 , n32353 , n32358 );
and ( n32360 , n32347 , n32359 );
and ( n32361 , n32346 , n32359 );
or ( n32362 , n32348 , n32360 , n32361 );
and ( n32363 , n32343 , n32362 );
xor ( n32364 , n32183 , n32185 );
xor ( n32365 , n32364 , n32188 );
xor ( n32366 , n32165 , n32167 );
xor ( n32367 , n32366 , n32170 );
and ( n32368 , n32365 , n32367 );
and ( n32369 , n30962 , n30950 );
and ( n32370 , n30958 , n30947 );
and ( n32371 , n32369 , n32370 );
xor ( n32372 , n32242 , n32251 );
and ( n32373 , n32370 , n32372 );
and ( n32374 , n32369 , n32372 );
or ( n32375 , n32371 , n32373 , n32374 );
and ( n32376 , n32368 , n32375 );
xor ( n32377 , n32257 , n32261 );
xor ( n32378 , n32344 , n32345 );
and ( n32379 , n32377 , n32378 );
and ( n32380 , n31783 , n30632 );
and ( n32381 , n31619 , n30685 );
and ( n32382 , n32380 , n32381 );
and ( n32383 , n31171 , n30950 );
and ( n32384 , n32381 , n32383 );
and ( n32385 , n32380 , n32383 );
or ( n32386 , n32382 , n32384 , n32385 );
and ( n32387 , n30627 , n31766 );
and ( n32388 , n30680 , n31597 );
and ( n32389 , n32387 , n32388 );
and ( n32390 , n30958 , n31168 );
and ( n32391 , n32388 , n32390 );
and ( n32392 , n32387 , n32390 );
or ( n32393 , n32389 , n32391 , n32392 );
and ( n32394 , n32386 , n32393 );
and ( n32395 , n32378 , n32394 );
and ( n32396 , n32377 , n32394 );
or ( n32397 , n32379 , n32395 , n32396 );
and ( n32398 , n32375 , n32397 );
and ( n32399 , n32368 , n32397 );
or ( n32400 , n32376 , n32398 , n32399 );
and ( n32401 , n32362 , n32400 );
and ( n32402 , n32343 , n32400 );
or ( n32403 , n32363 , n32401 , n32402 );
and ( n32404 , n32340 , n32403 );
xor ( n32405 , n32197 , n32198 );
xor ( n32406 , n32405 , n32200 );
xor ( n32407 , n32216 , n32217 );
xor ( n32408 , n32407 , n32221 );
and ( n32409 , n32406 , n32408 );
xor ( n32410 , n32232 , n32265 );
xor ( n32411 , n32410 , n32268 );
and ( n32412 , n32408 , n32411 );
and ( n32413 , n32406 , n32411 );
or ( n32414 , n32409 , n32412 , n32413 );
and ( n32415 , n32403 , n32414 );
and ( n32416 , n32340 , n32414 );
or ( n32417 , n32404 , n32415 , n32416 );
and ( n32418 , n32297 , n32417 );
xor ( n32419 , n32158 , n32195 );
xor ( n32420 , n32419 , n32203 );
xor ( n32421 , n32224 , n32271 );
xor ( n32422 , n32421 , n32274 );
and ( n32423 , n32420 , n32422 );
xor ( n32424 , n32279 , n32281 );
xor ( n32425 , n32424 , n32284 );
and ( n32426 , n32422 , n32425 );
and ( n32427 , n32420 , n32425 );
or ( n32428 , n32423 , n32426 , n32427 );
and ( n32429 , n32417 , n32428 );
and ( n32430 , n32297 , n32428 );
or ( n32431 , n32418 , n32429 , n32430 );
and ( n32432 , n32295 , n32431 );
and ( n32433 , n32293 , n32431 );
or ( n32434 , n559569 , n32432 , n32433 );
and ( n32435 , n32214 , n32434 );
and ( n32436 , n32212 , n32434 );
or ( n32437 , n32215 , n32435 , n32436 );
and ( n32438 , n32141 , n32437 );
xor ( n32439 , n32143 , n32145 );
xor ( n32440 , n32439 , n32209 );
xor ( n32441 , n32148 , n32150 );
xor ( n32442 , n32441 , n32206 );
xor ( n32443 , n32277 , n32287 );
xor ( n32444 , n32443 , n32290 );
and ( n32445 , n32442 , n32444 );
xor ( n32446 , n32225 , n32227 );
xor ( n32447 , n32446 , n32229 );
xor ( n32448 , n32233 , n32252 );
xor ( n32449 , n32448 , n32262 );
and ( n32450 , n32447 , n32449 );
xor ( n32451 , n32318 , n32336 );
and ( n32452 , n32449 , n32451 );
and ( n32453 , n32447 , n32451 );
or ( n32454 , n32450 , n32452 , n32453 );
xor ( n32455 , n32341 , n32342 );
xnor ( n32456 , n32355 , n32357 );
xor ( n32457 , n32255 , n32256 );
or ( n32458 , n32456 , n32457 );
xnor ( n32459 , n32350 , n32352 );
xor ( n32460 , n32259 , n32260 );
or ( n32461 , n32459 , n32460 );
and ( n32462 , n32458 , n32461 );
and ( n32463 , n32455 , n32462 );
xnor ( n32464 , n32315 , n32317 );
xnor ( n32465 , n32333 , n32335 );
and ( n32466 , n32464 , n32465 );
and ( n32467 , n32462 , n32466 );
and ( n32468 , n32455 , n32466 );
or ( n32469 , n32463 , n32467 , n32468 );
and ( n32470 , n32454 , n32469 );
and ( n32471 , n32019 , n30598 );
and ( n32472 , n31888 , n30620 );
and ( n32473 , n32471 , n32472 );
and ( n32474 , n31269 , n30863 );
and ( n32475 , n32472 , n32474 );
and ( n32476 , n32471 , n32474 );
or ( n32477 , n32473 , n32475 , n32476 );
and ( n32478 , n30601 , n31997 );
and ( n32479 , n30623 , n31871 );
and ( n32480 , n32478 , n32479 );
and ( n32481 , n30872 , n31278 );
and ( n32482 , n32479 , n32481 );
and ( n32483 , n32478 , n32481 );
or ( n32484 , n32480 , n32482 , n32483 );
and ( n32485 , n32477 , n32484 );
buf ( n32486 , n30962 );
buf ( n559761 , n543197 );
buf ( n32488 , n559761 );
and ( n32489 , n32486 , n32488 );
and ( n32490 , n31057 , n30947 );
and ( n32491 , n30962 , n31066 );
and ( n32492 , n32490 , n32491 );
buf ( n559767 , n543200 );
buf ( n32494 , n559767 );
and ( n32495 , n32491 , n32494 );
and ( n32496 , n32490 , n32494 );
or ( n32497 , n32492 , n32495 , n32496 );
and ( n32498 , n32488 , n32497 );
and ( n32499 , n32486 , n32497 );
or ( n32500 , n32489 , n32498 , n32499 );
and ( n32501 , n32485 , n32500 );
xor ( n32502 , n32353 , n32358 );
and ( n32503 , n32500 , n32502 );
and ( n32504 , n32485 , n32502 );
or ( n32505 , n32501 , n32503 , n32504 );
xor ( n32506 , n32365 , n32367 );
buf ( n559781 , n1240 );
buf ( n32508 , n559781 );
and ( n32509 , n30572 , n32508 );
and ( n32510 , n30680 , n31766 );
and ( n32511 , n32509 , n32510 );
and ( n32512 , n30711 , n31597 );
and ( n32513 , n32510 , n32512 );
and ( n32514 , n32509 , n32512 );
or ( n32515 , n32511 , n32513 , n32514 );
and ( n32516 , n30623 , n31997 );
and ( n32517 , n30627 , n31871 );
and ( n32518 , n32516 , n32517 );
and ( n32519 , n30759 , n31453 );
and ( n32520 , n32517 , n32519 );
and ( n32521 , n32516 , n32519 );
or ( n32522 , n32518 , n32520 , n32521 );
or ( n32523 , n32515 , n32522 );
buf ( n559798 , n1240 );
buf ( n32525 , n559798 );
and ( n32526 , n32525 , n30580 );
and ( n32527 , n31783 , n30685 );
and ( n32528 , n32526 , n32527 );
and ( n32529 , n31619 , n30716 );
and ( n32530 , n32527 , n32529 );
and ( n32531 , n32526 , n32529 );
or ( n32532 , n32528 , n32530 , n32531 );
and ( n32533 , n32019 , n30620 );
and ( n32534 , n31888 , n30632 );
and ( n32535 , n32533 , n32534 );
and ( n32536 , n31430 , n30748 );
and ( n32537 , n32534 , n32536 );
and ( n32538 , n32533 , n32536 );
or ( n32539 , n32535 , n32537 , n32538 );
or ( n32540 , n32532 , n32539 );
and ( n32541 , n32523 , n32540 );
and ( n32542 , n32506 , n32541 );
and ( n32543 , n30578 , n32320 );
and ( n32544 , n30601 , n32244 );
and ( n32545 , n32543 , n32544 );
and ( n32546 , n30958 , n31278 );
and ( n32547 , n32544 , n32546 );
and ( n32548 , n32543 , n32546 );
or ( n32549 , n32545 , n32547 , n32548 );
and ( n32550 , n31430 , n30716 );
or ( n32551 , n32549 , n32550 );
and ( n32552 , n32302 , n30583 );
and ( n32553 , n32235 , n30598 );
and ( n32554 , n32552 , n32553 );
and ( n32555 , n31269 , n30950 );
and ( n32556 , n32553 , n32555 );
and ( n32557 , n32552 , n32555 );
or ( n32558 , n32554 , n32556 , n32557 );
and ( n32559 , n30711 , n31453 );
or ( n32560 , n32558 , n32559 );
and ( n32561 , n32551 , n32560 );
and ( n32562 , n32541 , n32561 );
and ( n32563 , n32506 , n32561 );
or ( n32564 , n32542 , n32562 , n32563 );
and ( n32565 , n32505 , n32564 );
xor ( n32566 , n32327 , n32328 );
xor ( n32567 , n32566 , n32330 );
xor ( n32568 , n32309 , n32310 );
xor ( n32569 , n32568 , n32312 );
and ( n32570 , n32567 , n32569 );
xor ( n32571 , n32386 , n32393 );
xor ( n32572 , n32477 , n32484 );
and ( n32573 , n32571 , n32572 );
and ( n32574 , n31405 , n30863 );
and ( n32575 , n31171 , n30947 );
or ( n32576 , n32574 , n32575 );
and ( n32577 , n30872 , n31414 );
and ( n32578 , n30962 , n31168 );
or ( n32579 , n32577 , n32578 );
and ( n32580 , n32576 , n32579 );
and ( n32581 , n32572 , n32580 );
and ( n32582 , n32571 , n32580 );
or ( n32583 , n32573 , n32581 , n32582 );
and ( n32584 , n32570 , n32583 );
xor ( n32585 , n32380 , n32381 );
xor ( n32586 , n32585 , n32383 );
xor ( n32587 , n32387 , n32388 );
xor ( n32588 , n32587 , n32390 );
and ( n32589 , n32586 , n32588 );
xor ( n32590 , n32471 , n32472 );
xor ( n32591 , n32590 , n32474 );
xor ( n32592 , n32478 , n32479 );
xor ( n32593 , n32592 , n32481 );
and ( n32594 , n32591 , n32593 );
and ( n32595 , n32589 , n32594 );
xor ( n32596 , n32303 , n32304 );
xor ( n32597 , n32596 , n32306 );
xor ( n32598 , n32321 , n32322 );
xor ( n32599 , n32598 , n32324 );
and ( n32600 , n32597 , n32599 );
and ( n32601 , n32594 , n32600 );
and ( n32602 , n32589 , n32600 );
or ( n32603 , n32595 , n32601 , n32602 );
and ( n32604 , n32583 , n32603 );
and ( n32605 , n32570 , n32603 );
or ( n32606 , n32584 , n32604 , n32605 );
and ( n32607 , n32564 , n32606 );
and ( n32608 , n32505 , n32606 );
or ( n32609 , n32565 , n32607 , n32608 );
and ( n32610 , n32469 , n32609 );
and ( n32611 , n32454 , n32609 );
or ( n32612 , n32470 , n32610 , n32611 );
xor ( n32613 , n32298 , n32299 );
xor ( n32614 , n32613 , n32337 );
xor ( n32615 , n32343 , n32362 );
xor ( n32616 , n32615 , n32400 );
and ( n32617 , n32614 , n32616 );
xor ( n32618 , n32406 , n32408 );
xor ( n32619 , n32618 , n32411 );
and ( n32620 , n32616 , n32619 );
and ( n32621 , n32614 , n32619 );
or ( n32622 , n32617 , n32620 , n32621 );
and ( n32623 , n32612 , n32622 );
xor ( n32624 , n32340 , n32403 );
xor ( n32625 , n32624 , n32414 );
and ( n32626 , n32622 , n32625 );
and ( n32627 , n32612 , n32625 );
or ( n32628 , n32623 , n32626 , n32627 );
and ( n32629 , n32444 , n32628 );
and ( n32630 , n32442 , n32628 );
or ( n32631 , n32445 , n32629 , n32630 );
and ( n32632 , n32440 , n32631 );
xor ( n32633 , n32293 , n32295 );
xor ( n32634 , n32633 , n32431 );
and ( n32635 , n32631 , n32634 );
and ( n32636 , n32440 , n32634 );
or ( n32637 , n32632 , n32635 , n32636 );
xor ( n32638 , n32212 , n32214 );
xor ( n32639 , n32638 , n32434 );
and ( n32640 , n32637 , n32639 );
xor ( n32641 , n32297 , n32417 );
xor ( n32642 , n32641 , n32428 );
xor ( n32643 , n32420 , n32422 );
xor ( n32644 , n32643 , n32425 );
xor ( n32645 , n32346 , n32347 );
xor ( n32646 , n32645 , n32359 );
xor ( n32647 , n32368 , n32375 );
xor ( n32648 , n32647 , n32397 );
and ( n32649 , n32646 , n32648 );
xnor ( n32650 , n32456 , n32457 );
xnor ( n32651 , n32459 , n32460 );
and ( n32652 , n32650 , n32651 );
not ( n32653 , n32652 );
buf ( n559928 , n543194 );
buf ( n32655 , n559928 );
and ( n32656 , n32653 , n32655 );
and ( n32657 , n32648 , n32656 );
and ( n32658 , n32646 , n32656 );
or ( n32659 , n32649 , n32657 , n32658 );
buf ( n32660 , n32652 );
xor ( n32661 , n32369 , n32370 );
xor ( n32662 , n32661 , n32372 );
xor ( n32663 , n32377 , n32378 );
xor ( n32664 , n32663 , n32394 );
and ( n32665 , n32662 , n32664 );
xor ( n32666 , n32458 , n32461 );
and ( n32667 , n32664 , n32666 );
and ( n32668 , n32662 , n32666 );
or ( n32669 , n32665 , n32667 , n32668 );
and ( n32670 , n32660 , n32669 );
xor ( n32671 , n32464 , n32465 );
xor ( n32672 , n32486 , n32488 );
xor ( n32673 , n32672 , n32497 );
xor ( n32674 , n32523 , n32540 );
and ( n32675 , n32673 , n32674 );
xor ( n32676 , n32551 , n32560 );
and ( n32677 , n32674 , n32676 );
and ( n32678 , n32673 , n32676 );
or ( n32679 , n32675 , n32677 , n32678 );
and ( n32680 , n32671 , n32679 );
xor ( n32681 , n32567 , n32569 );
and ( n32682 , n30623 , n32244 );
and ( n32683 , n30627 , n31997 );
and ( n32684 , n32682 , n32683 );
and ( n32685 , n30958 , n31414 );
and ( n32686 , n32683 , n32685 );
and ( n32687 , n32682 , n32685 );
or ( n32688 , n32684 , n32686 , n32687 );
xor ( n32689 , n32526 , n32527 );
xor ( n32690 , n32689 , n32529 );
and ( n32691 , n32688 , n32690 );
xor ( n32692 , n32552 , n32553 );
xor ( n32693 , n32692 , n32555 );
and ( n32694 , n32690 , n32693 );
and ( n32695 , n32688 , n32693 );
or ( n32696 , n32691 , n32694 , n32695 );
and ( n32697 , n32235 , n30620 );
and ( n32698 , n32019 , n30632 );
and ( n32699 , n32697 , n32698 );
and ( n32700 , n31405 , n30950 );
and ( n32701 , n32698 , n32700 );
and ( n32702 , n32697 , n32700 );
or ( n32703 , n32699 , n32701 , n32702 );
xor ( n32704 , n32509 , n32510 );
xor ( n32705 , n32704 , n32512 );
and ( n32706 , n32703 , n32705 );
xor ( n32707 , n32543 , n32544 );
xor ( n32708 , n32707 , n32546 );
and ( n32709 , n32705 , n32708 );
and ( n32710 , n32703 , n32708 );
or ( n32711 , n32706 , n32709 , n32710 );
and ( n32712 , n32696 , n32711 );
and ( n32713 , n32681 , n32712 );
and ( n32714 , n30578 , n32508 );
and ( n32715 , n30601 , n32320 );
and ( n32716 , n32714 , n32715 );
and ( n32717 , n30872 , n31453 );
and ( n32718 , n32715 , n32717 );
and ( n32719 , n32714 , n32717 );
or ( n32720 , n32716 , n32718 , n32719 );
and ( n32721 , n30680 , n31871 );
and ( n32722 , n30711 , n31766 );
and ( n32723 , n32721 , n32722 );
and ( n32724 , n30962 , n31278 );
and ( n32725 , n32722 , n32724 );
and ( n32726 , n32721 , n32724 );
or ( n32727 , n32723 , n32725 , n32726 );
or ( n32728 , n32720 , n32727 );
and ( n32729 , n32525 , n30583 );
and ( n32730 , n32302 , n30598 );
and ( n32731 , n32729 , n32730 );
and ( n32732 , n31430 , n30863 );
and ( n32733 , n32730 , n32732 );
and ( n32734 , n32729 , n32732 );
or ( n32735 , n32731 , n32733 , n32734 );
and ( n32736 , n31888 , n30685 );
and ( n32737 , n31783 , n30716 );
and ( n32738 , n32736 , n32737 );
and ( n32739 , n31269 , n30947 );
and ( n32740 , n32737 , n32739 );
and ( n32741 , n32736 , n32739 );
or ( n32742 , n32738 , n32740 , n32741 );
or ( n32743 , n32735 , n32742 );
and ( n32744 , n32728 , n32743 );
and ( n32745 , n32712 , n32744 );
and ( n32746 , n32681 , n32744 );
or ( n32747 , n32713 , n32745 , n32746 );
and ( n32748 , n32679 , n32747 );
and ( n32749 , n32671 , n32747 );
or ( n32750 , n32680 , n32748 , n32749 );
and ( n32751 , n32669 , n32750 );
and ( n32752 , n32660 , n32750 );
or ( n32753 , n32670 , n32751 , n32752 );
and ( n32754 , n32659 , n32753 );
xnor ( n32755 , n32515 , n32522 );
xnor ( n32756 , n32532 , n32539 );
and ( n32757 , n32755 , n32756 );
xnor ( n32758 , n32549 , n32550 );
xnor ( n32759 , n32558 , n32559 );
and ( n32760 , n32758 , n32759 );
and ( n32761 , n32757 , n32760 );
xor ( n32762 , n32490 , n32491 );
xor ( n32763 , n32762 , n32494 );
xor ( n32764 , n32576 , n32579 );
and ( n32765 , n32763 , n32764 );
xor ( n32766 , n32586 , n32588 );
and ( n32767 , n32764 , n32766 );
and ( n32768 , n32763 , n32766 );
or ( n32769 , n32765 , n32767 , n32768 );
and ( n32770 , n32760 , n32769 );
and ( n32771 , n32757 , n32769 );
or ( n32772 , n32761 , n32770 , n32771 );
xor ( n32773 , n32591 , n32593 );
xor ( n32774 , n32597 , n32599 );
and ( n32775 , n32773 , n32774 );
xnor ( n32776 , n32574 , n32575 );
xnor ( n32777 , n32577 , n32578 );
and ( n32778 , n32776 , n32777 );
and ( n32779 , n32774 , n32778 );
and ( n32780 , n32773 , n32778 );
or ( n32781 , n32775 , n32779 , n32780 );
xor ( n32782 , n32571 , n32572 );
xor ( n32783 , n32782 , n32580 );
and ( n32784 , n32781 , n32783 );
xor ( n32785 , n32589 , n32594 );
xor ( n32786 , n32785 , n32600 );
and ( n32787 , n32783 , n32786 );
and ( n32788 , n32781 , n32786 );
or ( n32789 , n32784 , n32787 , n32788 );
and ( n32790 , n32772 , n32789 );
xor ( n32791 , n32485 , n32500 );
xor ( n32792 , n32791 , n32502 );
and ( n32793 , n32789 , n32792 );
and ( n32794 , n32772 , n32792 );
or ( n32795 , n32790 , n32793 , n32794 );
xor ( n32796 , n32447 , n32449 );
xor ( n32797 , n32796 , n32451 );
and ( n32798 , n32795 , n32797 );
xor ( n32799 , n32455 , n32462 );
xor ( n32800 , n32799 , n32466 );
and ( n32801 , n32797 , n32800 );
and ( n32802 , n32795 , n32800 );
or ( n32803 , n32798 , n32801 , n32802 );
and ( n32804 , n32753 , n32803 );
and ( n32805 , n32659 , n32803 );
or ( n32806 , n32754 , n32804 , n32805 );
and ( n32807 , n32644 , n32806 );
xor ( n32808 , n32612 , n32622 );
xor ( n32809 , n32808 , n32625 );
and ( n32810 , n32806 , n32809 );
and ( n32811 , n32644 , n32809 );
or ( n32812 , n32807 , n32810 , n32811 );
and ( n32813 , n32642 , n32812 );
xor ( n32814 , n32442 , n32444 );
xor ( n32815 , n32814 , n32628 );
and ( n32816 , n32812 , n32815 );
and ( n32817 , n32642 , n32815 );
or ( n32818 , n32813 , n32816 , n32817 );
xor ( n32819 , n32440 , n32631 );
xor ( n32820 , n32819 , n32634 );
and ( n32821 , n32818 , n32820 );
xor ( n32822 , n32642 , n32812 );
xor ( n32823 , n32822 , n32815 );
xor ( n32824 , n32454 , n32469 );
xor ( n32825 , n32824 , n32609 );
xor ( n32826 , n32614 , n32616 );
xor ( n32827 , n32826 , n32619 );
and ( n32828 , n32825 , n32827 );
xor ( n32829 , n32505 , n32564 );
xor ( n32830 , n32829 , n32606 );
xor ( n32831 , n32506 , n32541 );
xor ( n32832 , n32831 , n32561 );
xor ( n32833 , n32570 , n32583 );
xor ( n32834 , n32833 , n32603 );
and ( n32835 , n32832 , n32834 );
xor ( n32836 , n32653 , n32655 );
and ( n32837 , n32834 , n32836 );
and ( n32838 , n32832 , n32836 );
or ( n32839 , n32835 , n32837 , n32838 );
and ( n32840 , n32830 , n32839 );
xor ( n32841 , n32650 , n32651 );
and ( n32842 , n32235 , n30632 );
and ( n32843 , n32019 , n30685 );
and ( n32844 , n32842 , n32843 );
and ( n32845 , n31619 , n30863 );
and ( n32846 , n32843 , n32845 );
and ( n32847 , n32842 , n32845 );
or ( n32848 , n32844 , n32846 , n32847 );
buf ( n560123 , n1241 );
buf ( n32850 , n560123 );
and ( n32851 , n30572 , n32850 );
and ( n32852 , n32848 , n32851 );
and ( n32853 , n30759 , n31597 );
and ( n32854 , n32851 , n32853 );
and ( n32855 , n32848 , n32853 );
or ( n32856 , n32852 , n32854 , n32855 );
xor ( n32857 , n32516 , n32517 );
xor ( n32858 , n32857 , n32519 );
or ( n32859 , n32856 , n32858 );
and ( n32860 , n30627 , n32244 );
and ( n32861 , n30680 , n31997 );
and ( n32862 , n32860 , n32861 );
and ( n32863 , n30872 , n31597 );
and ( n32864 , n32861 , n32863 );
and ( n32865 , n32860 , n32863 );
or ( n32866 , n32862 , n32864 , n32865 );
buf ( n560141 , n1241 );
buf ( n32868 , n560141 );
and ( n32869 , n32868 , n30580 );
and ( n32870 , n32866 , n32869 );
and ( n32871 , n31619 , n30748 );
and ( n32872 , n32869 , n32871 );
and ( n32873 , n32866 , n32871 );
or ( n32874 , n32870 , n32872 , n32873 );
xor ( n32875 , n32533 , n32534 );
xor ( n32876 , n32875 , n32536 );
or ( n32877 , n32874 , n32876 );
and ( n32878 , n32859 , n32877 );
and ( n32879 , n32841 , n32878 );
buf ( n32880 , n31057 );
buf ( n560155 , n543203 );
buf ( n32882 , n560155 );
and ( n32883 , n32880 , n32882 );
and ( n32884 , n31171 , n31066 );
and ( n32885 , n31057 , n31168 );
and ( n32886 , n32884 , n32885 );
buf ( n560161 , n543206 );
buf ( n32888 , n560161 );
and ( n32889 , n32885 , n32888 );
and ( n32890 , n32884 , n32888 );
or ( n32891 , n32886 , n32889 , n32890 );
and ( n32892 , n32882 , n32891 );
and ( n32893 , n32880 , n32891 );
or ( n32894 , n32883 , n32892 , n32893 );
xor ( n32895 , n32696 , n32711 );
and ( n32896 , n32894 , n32895 );
xor ( n32897 , n32728 , n32743 );
and ( n32898 , n32895 , n32897 );
and ( n32899 , n32894 , n32897 );
or ( n32900 , n32896 , n32898 , n32899 );
and ( n32901 , n32878 , n32900 );
and ( n32902 , n32841 , n32900 );
or ( n32903 , n32879 , n32901 , n32902 );
xor ( n32904 , n32755 , n32756 );
xor ( n32905 , n32758 , n32759 );
and ( n32906 , n32904 , n32905 );
xor ( n32907 , n32721 , n32722 );
xor ( n32908 , n32907 , n32724 );
xor ( n32909 , n32682 , n32683 );
xor ( n32910 , n32909 , n32685 );
or ( n32911 , n32908 , n32910 );
xor ( n32912 , n32736 , n32737 );
xor ( n32913 , n32912 , n32739 );
xor ( n32914 , n32697 , n32698 );
xor ( n32915 , n32914 , n32700 );
or ( n32916 , n32913 , n32915 );
and ( n32917 , n32911 , n32916 );
and ( n32918 , n32905 , n32917 );
and ( n32919 , n32904 , n32917 );
or ( n32920 , n32906 , n32918 , n32919 );
buf ( n560195 , n1242 );
buf ( n32922 , n560195 );
and ( n32923 , n30572 , n32922 );
and ( n32924 , n30578 , n32850 );
and ( n32925 , n32923 , n32924 );
and ( n32926 , n30759 , n31766 );
and ( n32927 , n32924 , n32926 );
and ( n32928 , n32923 , n32926 );
or ( n32929 , n32925 , n32927 , n32928 );
not ( n32930 , n32929 );
and ( n32931 , n30601 , n32508 );
and ( n32932 , n30623 , n32320 );
and ( n32933 , n32931 , n32932 );
and ( n32934 , n30962 , n31414 );
and ( n32935 , n32932 , n32934 );
and ( n32936 , n32931 , n32934 );
or ( n32937 , n32933 , n32935 , n32936 );
and ( n32938 , n32930 , n32937 );
buf ( n560213 , n1242 );
buf ( n32940 , n560213 );
and ( n32941 , n32940 , n30580 );
and ( n32942 , n32868 , n30583 );
and ( n32943 , n32941 , n32942 );
and ( n32944 , n31783 , n30748 );
and ( n32945 , n32942 , n32944 );
and ( n32946 , n32941 , n32944 );
or ( n32947 , n32943 , n32945 , n32946 );
not ( n32948 , n32947 );
and ( n32949 , n32525 , n30598 );
and ( n32950 , n32302 , n30620 );
and ( n32951 , n32949 , n32950 );
and ( n32952 , n31405 , n30947 );
and ( n32953 , n32950 , n32952 );
and ( n32954 , n32949 , n32952 );
or ( n32955 , n32951 , n32953 , n32954 );
and ( n32956 , n32948 , n32955 );
and ( n32957 , n32938 , n32956 );
buf ( n32958 , n32929 );
buf ( n32959 , n32947 );
and ( n32960 , n32958 , n32959 );
and ( n32961 , n32957 , n32960 );
xor ( n32962 , n32688 , n32690 );
xor ( n32963 , n32962 , n32693 );
xor ( n32964 , n32703 , n32705 );
xor ( n32965 , n32964 , n32708 );
and ( n32966 , n32963 , n32965 );
and ( n32967 , n32960 , n32966 );
and ( n32968 , n32957 , n32966 );
or ( n32969 , n32961 , n32967 , n32968 );
and ( n32970 , n32920 , n32969 );
xnor ( n32971 , n32720 , n32727 );
xnor ( n32972 , n32735 , n32742 );
and ( n32973 , n32971 , n32972 );
xor ( n32974 , n32776 , n32777 );
and ( n32975 , n30958 , n31453 );
and ( n32976 , n31430 , n30950 );
and ( n32977 , n32975 , n32976 );
and ( n32978 , n31057 , n31278 );
and ( n32979 , n31269 , n31066 );
and ( n32980 , n32978 , n32979 );
and ( n32981 , n32977 , n32980 );
xor ( n32982 , n32884 , n32885 );
xor ( n32983 , n32982 , n32888 );
and ( n32984 , n32980 , n32983 );
and ( n32985 , n32977 , n32983 );
or ( n32986 , n32981 , n32984 , n32985 );
and ( n32987 , n32974 , n32986 );
xor ( n32988 , n32880 , n32882 );
xor ( n32989 , n32988 , n32891 );
and ( n32990 , n32986 , n32989 );
and ( n32991 , n32974 , n32989 );
or ( n32992 , n32987 , n32990 , n32991 );
and ( n32993 , n32973 , n32992 );
xor ( n32994 , n32763 , n32764 );
xor ( n32995 , n32994 , n32766 );
and ( n32996 , n32992 , n32995 );
and ( n32997 , n32973 , n32995 );
or ( n32998 , n32993 , n32996 , n32997 );
and ( n32999 , n32969 , n32998 );
and ( n33000 , n32920 , n32998 );
or ( n33001 , n32970 , n32999 , n33000 );
and ( n33002 , n32903 , n33001 );
xor ( n33003 , n32673 , n32674 );
xor ( n33004 , n33003 , n32676 );
xor ( n33005 , n32681 , n32712 );
xor ( n33006 , n33005 , n32744 );
and ( n33007 , n33004 , n33006 );
xor ( n33008 , n32757 , n32760 );
xor ( n33009 , n33008 , n32769 );
and ( n33010 , n33006 , n33009 );
and ( n33011 , n33004 , n33009 );
or ( n33012 , n33007 , n33010 , n33011 );
and ( n33013 , n33001 , n33012 );
and ( n33014 , n32903 , n33012 );
or ( n33015 , n33002 , n33013 , n33014 );
and ( n33016 , n32839 , n33015 );
and ( n33017 , n32830 , n33015 );
or ( n33018 , n32840 , n33016 , n33017 );
and ( n33019 , n32827 , n33018 );
and ( n33020 , n32825 , n33018 );
or ( n33021 , n32828 , n33019 , n33020 );
xor ( n33022 , n32644 , n32806 );
xor ( n33023 , n33022 , n32809 );
and ( n33024 , n33021 , n33023 );
xor ( n33025 , n32662 , n32664 );
xor ( n33026 , n33025 , n32666 );
xor ( n33027 , n32671 , n32679 );
xor ( n33028 , n33027 , n32747 );
and ( n33029 , n33026 , n33028 );
xor ( n33030 , n32772 , n32789 );
xor ( n33031 , n33030 , n32792 );
and ( n33032 , n33028 , n33031 );
and ( n33033 , n33026 , n33031 );
or ( n33034 , n33029 , n33032 , n33033 );
xor ( n33035 , n32646 , n32648 );
xor ( n33036 , n33035 , n32656 );
and ( n33037 , n33034 , n33036 );
xor ( n33038 , n32660 , n32669 );
xor ( n33039 , n33038 , n32750 );
and ( n33040 , n33036 , n33039 );
and ( n33041 , n33034 , n33039 );
or ( n33042 , n33037 , n33040 , n33041 );
xor ( n33043 , n32659 , n32753 );
xor ( n33044 , n33043 , n32803 );
and ( n33045 , n33042 , n33044 );
xor ( n33046 , n32795 , n32797 );
xor ( n33047 , n33046 , n32800 );
xor ( n33048 , n32781 , n32783 );
xor ( n33049 , n33048 , n32786 );
xor ( n33050 , n32773 , n32774 );
xor ( n33051 , n33050 , n32778 );
xor ( n33052 , n32859 , n32877 );
and ( n33053 , n33051 , n33052 );
xor ( n33054 , n32714 , n32715 );
xor ( n33055 , n33054 , n32717 );
xor ( n33056 , n32848 , n32851 );
xor ( n33057 , n33056 , n32853 );
or ( n33058 , n33055 , n33057 );
xor ( n33059 , n32729 , n32730 );
xor ( n33060 , n33059 , n32732 );
xor ( n33061 , n32866 , n32869 );
xor ( n33062 , n33061 , n32871 );
or ( n33063 , n33060 , n33062 );
and ( n33064 , n33058 , n33063 );
and ( n33065 , n33052 , n33064 );
and ( n33066 , n33051 , n33064 );
or ( n33067 , n33053 , n33065 , n33066 );
and ( n33068 , n33049 , n33067 );
xnor ( n33069 , n32856 , n32858 );
xnor ( n33070 , n32874 , n32876 );
and ( n33071 , n33069 , n33070 );
xor ( n33072 , n32911 , n32916 );
xor ( n33073 , n32938 , n32956 );
and ( n33074 , n33072 , n33073 );
xor ( n33075 , n32958 , n32959 );
and ( n33076 , n33073 , n33075 );
and ( n33077 , n33072 , n33075 );
or ( n33078 , n33074 , n33076 , n33077 );
and ( n33079 , n33071 , n33078 );
xor ( n33080 , n32963 , n32965 );
xor ( n33081 , n32971 , n32972 );
and ( n33082 , n33080 , n33081 );
and ( n33083 , n30601 , n32850 );
and ( n33084 , n30623 , n32508 );
and ( n33085 , n33083 , n33084 );
and ( n33086 , n30958 , n31597 );
and ( n33087 , n33084 , n33086 );
and ( n33088 , n33083 , n33086 );
or ( n33089 , n33085 , n33087 , n33088 );
and ( n33090 , n30627 , n32320 );
and ( n33091 , n30680 , n32244 );
and ( n33092 , n33090 , n33091 );
and ( n33093 , n30962 , n31453 );
and ( n33094 , n33091 , n33093 );
and ( n33095 , n33090 , n33093 );
or ( n33096 , n33092 , n33094 , n33095 );
and ( n33097 , n33089 , n33096 );
and ( n33098 , n31888 , n30716 );
and ( n33099 , n33096 , n33098 );
and ( n33100 , n33089 , n33098 );
or ( n33101 , n33097 , n33099 , n33100 );
and ( n33102 , n32868 , n30598 );
and ( n33103 , n32525 , n30620 );
and ( n33104 , n33102 , n33103 );
and ( n33105 , n31619 , n30950 );
and ( n33106 , n33103 , n33105 );
and ( n33107 , n33102 , n33105 );
or ( n33108 , n33104 , n33106 , n33107 );
and ( n33109 , n32302 , n30632 );
and ( n33110 , n32235 , n30685 );
and ( n33111 , n33109 , n33110 );
and ( n33112 , n31430 , n30947 );
and ( n33113 , n33110 , n33112 );
and ( n33114 , n33109 , n33112 );
or ( n33115 , n33111 , n33113 , n33114 );
and ( n33116 , n33108 , n33115 );
and ( n33117 , n30711 , n31871 );
and ( n33118 , n33115 , n33117 );
and ( n33119 , n33108 , n33117 );
or ( n33120 , n33116 , n33118 , n33119 );
and ( n33121 , n33101 , n33120 );
and ( n33122 , n33081 , n33121 );
and ( n33123 , n33080 , n33121 );
or ( n33124 , n33082 , n33122 , n33123 );
and ( n33125 , n33078 , n33124 );
and ( n33126 , n33071 , n33124 );
or ( n33127 , n33079 , n33125 , n33126 );
and ( n33128 , n33067 , n33127 );
and ( n33129 , n33049 , n33127 );
or ( n33130 , n33068 , n33128 , n33129 );
xor ( n33131 , n32923 , n32924 );
xor ( n33132 , n33131 , n32926 );
xor ( n33133 , n32931 , n32932 );
xor ( n33134 , n33133 , n32934 );
or ( n33135 , n33132 , n33134 );
xor ( n33136 , n32941 , n32942 );
xor ( n33137 , n33136 , n32944 );
xor ( n33138 , n32949 , n32950 );
xor ( n33139 , n33138 , n32952 );
or ( n33140 , n33137 , n33139 );
and ( n33141 , n33135 , n33140 );
xnor ( n33142 , n32908 , n32910 );
xnor ( n33143 , n32913 , n32915 );
and ( n33144 , n33142 , n33143 );
and ( n33145 , n33141 , n33144 );
xor ( n33146 , n32930 , n32937 );
xor ( n33147 , n32948 , n32955 );
and ( n33148 , n33146 , n33147 );
and ( n33149 , n33144 , n33148 );
and ( n33150 , n33141 , n33148 );
or ( n33151 , n33145 , n33149 , n33150 );
xor ( n33152 , n32894 , n32895 );
xor ( n33153 , n33152 , n32897 );
and ( n33154 , n33151 , n33153 );
xor ( n33155 , n32904 , n32905 );
xor ( n33156 , n33155 , n32917 );
and ( n33157 , n33153 , n33156 );
and ( n33158 , n33151 , n33156 );
or ( n33159 , n33154 , n33157 , n33158 );
xor ( n33160 , n32841 , n32878 );
xor ( n33161 , n33160 , n32900 );
and ( n33162 , n33159 , n33161 );
xor ( n33163 , n32920 , n32969 );
xor ( n33164 , n33163 , n32998 );
and ( n33165 , n33161 , n33164 );
and ( n33166 , n33159 , n33164 );
or ( n33167 , n33162 , n33165 , n33166 );
and ( n33168 , n33130 , n33167 );
xor ( n33169 , n32832 , n32834 );
xor ( n33170 , n33169 , n32836 );
and ( n33171 , n33167 , n33170 );
and ( n33172 , n33130 , n33170 );
or ( n33173 , n33168 , n33171 , n33172 );
and ( n33174 , n33047 , n33173 );
xor ( n33175 , n32830 , n32839 );
xor ( n33176 , n33175 , n33015 );
and ( n33177 , n33173 , n33176 );
and ( n33178 , n33047 , n33176 );
or ( n33179 , n33174 , n33177 , n33178 );
and ( n33180 , n33044 , n33179 );
and ( n33181 , n33042 , n33179 );
or ( n33182 , n33045 , n33180 , n33181 );
and ( n33183 , n33023 , n33182 );
and ( n33184 , n33021 , n33182 );
or ( n33185 , n33024 , n33183 , n33184 );
and ( n33186 , n32823 , n33185 );
xor ( n33187 , n32825 , n32827 );
xor ( n33188 , n33187 , n33018 );
xor ( n33189 , n33034 , n33036 );
xor ( n33190 , n33189 , n33039 );
xor ( n33191 , n32903 , n33001 );
xor ( n33192 , n33191 , n33012 );
xor ( n33193 , n33026 , n33028 );
xor ( n33194 , n33193 , n33031 );
and ( n33195 , n33192 , n33194 );
xor ( n33196 , n33004 , n33006 );
xor ( n33197 , n33196 , n33009 );
xor ( n33198 , n32957 , n32960 );
xor ( n33199 , n33198 , n32966 );
xor ( n33200 , n32973 , n32992 );
xor ( n33201 , n33200 , n32995 );
and ( n33202 , n33199 , n33201 );
buf ( n560477 , n1243 );
buf ( n33204 , n560477 );
and ( n33205 , n33204 , n30580 );
and ( n33206 , n32940 , n30583 );
and ( n33207 , n33205 , n33206 );
and ( n33208 , n31783 , n30863 );
and ( n33209 , n33206 , n33208 );
and ( n33210 , n33205 , n33208 );
or ( n33211 , n33207 , n33209 , n33210 );
buf ( n560486 , n1243 );
buf ( n33213 , n560486 );
and ( n33214 , n30572 , n33213 );
and ( n33215 , n30578 , n32922 );
and ( n33216 , n33214 , n33215 );
and ( n33217 , n30872 , n31766 );
and ( n33218 , n33215 , n33217 );
and ( n33219 , n33214 , n33217 );
or ( n33220 , n33216 , n33218 , n33219 );
and ( n33221 , n33211 , n33220 );
and ( n33222 , n32019 , n30716 );
and ( n33223 , n31888 , n30748 );
and ( n33224 , n33222 , n33223 );
and ( n33225 , n31405 , n31066 );
and ( n33226 , n33223 , n33225 );
and ( n33227 , n33222 , n33225 );
or ( n33228 , n33224 , n33226 , n33227 );
and ( n33229 , n30711 , n31997 );
and ( n33230 , n30759 , n31871 );
and ( n33231 , n33229 , n33230 );
and ( n33232 , n31057 , n31414 );
and ( n33233 , n33230 , n33232 );
and ( n33234 , n33229 , n33232 );
or ( n33235 , n33231 , n33233 , n33234 );
and ( n33236 , n33228 , n33235 );
and ( n33237 , n33221 , n33236 );
buf ( n33238 , n31171 );
buf ( n560513 , n543209 );
buf ( n33240 , n560513 );
and ( n33241 , n33238 , n33240 );
xor ( n33242 , n32975 , n32976 );
and ( n33243 , n33240 , n33242 );
and ( n33244 , n33238 , n33242 );
or ( n33245 , n33241 , n33243 , n33244 );
and ( n33246 , n33236 , n33245 );
and ( n33247 , n33221 , n33245 );
or ( n33248 , n33237 , n33246 , n33247 );
xor ( n33249 , n32974 , n32986 );
xor ( n33250 , n33249 , n32989 );
and ( n33251 , n33248 , n33250 );
xor ( n33252 , n33058 , n33063 );
and ( n33253 , n33250 , n33252 );
and ( n33254 , n33248 , n33252 );
or ( n33255 , n33251 , n33253 , n33254 );
and ( n33256 , n33201 , n33255 );
and ( n33257 , n33199 , n33255 );
or ( n33258 , n33202 , n33256 , n33257 );
and ( n33259 , n33197 , n33258 );
xor ( n33260 , n33069 , n33070 );
xor ( n33261 , n33083 , n33084 );
xor ( n33262 , n33261 , n33086 );
xor ( n33263 , n33229 , n33230 );
xor ( n33264 , n33263 , n33232 );
and ( n33265 , n33262 , n33264 );
xor ( n33266 , n33090 , n33091 );
xor ( n33267 , n33266 , n33093 );
and ( n33268 , n33264 , n33267 );
and ( n33269 , n33262 , n33267 );
or ( n33270 , n33265 , n33268 , n33269 );
xor ( n33271 , n32860 , n32861 );
xor ( n33272 , n33271 , n32863 );
or ( n33273 , n33270 , n33272 );
xor ( n33274 , n33102 , n33103 );
xor ( n33275 , n33274 , n33105 );
xor ( n33276 , n33222 , n33223 );
xor ( n33277 , n33276 , n33225 );
and ( n33278 , n33275 , n33277 );
xor ( n33279 , n33109 , n33110 );
xor ( n33280 , n33279 , n33112 );
and ( n33281 , n33277 , n33280 );
and ( n33282 , n33275 , n33280 );
or ( n33283 , n33278 , n33281 , n33282 );
xor ( n33284 , n32842 , n32843 );
xor ( n33285 , n33284 , n32845 );
or ( n33286 , n33283 , n33285 );
and ( n33287 , n33273 , n33286 );
and ( n33288 , n33260 , n33287 );
and ( n33289 , n33204 , n30583 );
and ( n33290 , n32940 , n30598 );
and ( n33291 , n33289 , n33290 );
and ( n33292 , n31888 , n30863 );
and ( n33293 , n33290 , n33292 );
and ( n33294 , n33289 , n33292 );
or ( n33295 , n33291 , n33293 , n33294 );
and ( n33296 , n32868 , n30620 );
and ( n33297 , n32525 , n30632 );
and ( n33298 , n33296 , n33297 );
and ( n33299 , n31430 , n31066 );
and ( n33300 , n33297 , n33299 );
and ( n33301 , n33296 , n33299 );
or ( n33302 , n33298 , n33300 , n33301 );
and ( n33303 , n33295 , n33302 );
xor ( n33304 , n33214 , n33215 );
xor ( n33305 , n33304 , n33217 );
and ( n33306 , n33302 , n33305 );
and ( n33307 , n33295 , n33305 );
or ( n33308 , n33303 , n33306 , n33307 );
not ( n33309 , n33308 );
xor ( n33310 , n33108 , n33115 );
xor ( n33311 , n33310 , n33117 );
and ( n33312 , n33309 , n33311 );
and ( n33313 , n30578 , n33213 );
and ( n33314 , n30601 , n32922 );
and ( n33315 , n33313 , n33314 );
and ( n33316 , n30872 , n31871 );
and ( n33317 , n33314 , n33316 );
and ( n33318 , n33313 , n33316 );
or ( n33319 , n33315 , n33317 , n33318 );
and ( n33320 , n30623 , n32850 );
and ( n33321 , n30627 , n32508 );
and ( n33322 , n33320 , n33321 );
and ( n33323 , n31057 , n31453 );
and ( n33324 , n33321 , n33323 );
and ( n33325 , n33320 , n33323 );
or ( n33326 , n33322 , n33324 , n33325 );
and ( n33327 , n33319 , n33326 );
xor ( n33328 , n33205 , n33206 );
xor ( n33329 , n33328 , n33208 );
and ( n33330 , n33326 , n33329 );
and ( n33331 , n33319 , n33329 );
or ( n33332 , n33327 , n33330 , n33331 );
not ( n33333 , n33332 );
xor ( n33334 , n33089 , n33096 );
xor ( n33335 , n33334 , n33098 );
and ( n33336 , n33333 , n33335 );
and ( n33337 , n33312 , n33336 );
and ( n33338 , n33287 , n33337 );
and ( n33339 , n33260 , n33337 );
or ( n33340 , n33288 , n33338 , n33339 );
buf ( n33341 , n33308 );
buf ( n33342 , n33332 );
and ( n33343 , n33341 , n33342 );
xnor ( n33344 , n33055 , n33057 );
xnor ( n33345 , n33060 , n33062 );
and ( n33346 , n33344 , n33345 );
and ( n33347 , n33343 , n33346 );
xor ( n33348 , n32977 , n32980 );
xor ( n33349 , n33348 , n32983 );
xor ( n33350 , n33101 , n33120 );
and ( n33351 , n33349 , n33350 );
xor ( n33352 , n33135 , n33140 );
and ( n33353 , n33350 , n33352 );
and ( n33354 , n33349 , n33352 );
or ( n33355 , n33351 , n33353 , n33354 );
and ( n33356 , n33346 , n33355 );
and ( n33357 , n33343 , n33355 );
or ( n33358 , n33347 , n33356 , n33357 );
and ( n33359 , n33340 , n33358 );
xor ( n33360 , n33142 , n33143 );
xor ( n33361 , n33146 , n33147 );
and ( n33362 , n33360 , n33361 );
xnor ( n33363 , n33132 , n33134 );
xnor ( n33364 , n33137 , n33139 );
and ( n33365 , n33363 , n33364 );
and ( n33366 , n33361 , n33365 );
and ( n33367 , n33360 , n33365 );
or ( n33368 , n33362 , n33366 , n33367 );
xor ( n33369 , n32978 , n32979 );
and ( n33370 , n31269 , n31168 );
and ( n33371 , n31171 , n31278 );
and ( n33372 , n33370 , n33371 );
buf ( n560647 , n543212 );
buf ( n33374 , n560647 );
and ( n33375 , n33371 , n33374 );
and ( n33376 , n33370 , n33374 );
or ( n33377 , n33372 , n33375 , n33376 );
and ( n33378 , n33369 , n33377 );
xor ( n33379 , n33211 , n33220 );
and ( n33380 , n33377 , n33379 );
and ( n33381 , n33369 , n33379 );
or ( n33382 , n33378 , n33380 , n33381 );
xor ( n33383 , n33228 , n33235 );
and ( n33384 , n32302 , n30685 );
and ( n33385 , n32235 , n30716 );
and ( n33386 , n33384 , n33385 );
and ( n33387 , n31783 , n30950 );
and ( n33388 , n33385 , n33387 );
and ( n33389 , n33384 , n33387 );
or ( n33390 , n33386 , n33388 , n33389 );
and ( n33391 , n30680 , n32320 );
and ( n33392 , n30711 , n32244 );
and ( n33393 , n33391 , n33392 );
and ( n33394 , n30958 , n31766 );
and ( n33395 , n33392 , n33394 );
and ( n33396 , n33391 , n33394 );
or ( n33397 , n33393 , n33395 , n33396 );
and ( n33398 , n33390 , n33397 );
and ( n33399 , n33383 , n33398 );
and ( n33400 , n31619 , n30947 );
and ( n33401 , n31405 , n31168 );
or ( n33402 , n33400 , n33401 );
and ( n33403 , n30962 , n31597 );
and ( n33404 , n31171 , n31414 );
or ( n33405 , n33403 , n33404 );
and ( n33406 , n33402 , n33405 );
and ( n33407 , n33398 , n33406 );
and ( n33408 , n33383 , n33406 );
or ( n33409 , n33399 , n33407 , n33408 );
and ( n33410 , n33382 , n33409 );
xor ( n33411 , n33221 , n33236 );
xor ( n33412 , n33411 , n33245 );
and ( n33413 , n33409 , n33412 );
and ( n33414 , n33382 , n33412 );
or ( n33415 , n33410 , n33413 , n33414 );
and ( n33416 , n33368 , n33415 );
xor ( n33417 , n33072 , n33073 );
xor ( n33418 , n33417 , n33075 );
and ( n33419 , n33415 , n33418 );
and ( n33420 , n33368 , n33418 );
or ( n33421 , n33416 , n33419 , n33420 );
and ( n33422 , n33358 , n33421 );
and ( n33423 , n33340 , n33421 );
or ( n33424 , n33359 , n33422 , n33423 );
and ( n33425 , n33258 , n33424 );
and ( n33426 , n33197 , n33424 );
or ( n33427 , n33259 , n33425 , n33426 );
and ( n33428 , n33194 , n33427 );
and ( n33429 , n33192 , n33427 );
or ( n33430 , n33195 , n33428 , n33429 );
and ( n33431 , n33190 , n33430 );
xor ( n33432 , n33047 , n33173 );
xor ( n33433 , n33432 , n33176 );
and ( n33434 , n33430 , n33433 );
and ( n33435 , n33190 , n33433 );
or ( n33436 , n33431 , n33434 , n33435 );
and ( n33437 , n33188 , n33436 );
xor ( n33438 , n33042 , n33044 );
xor ( n33439 , n33438 , n33179 );
and ( n33440 , n33436 , n33439 );
and ( n33441 , n33188 , n33439 );
or ( n33442 , n33437 , n33440 , n33441 );
xor ( n33443 , n33021 , n33023 );
xor ( n33444 , n33443 , n33182 );
and ( n33445 , n33442 , n33444 );
xor ( n33446 , n33188 , n33436 );
xor ( n33447 , n33446 , n33439 );
xor ( n33448 , n33051 , n33052 );
xor ( n33449 , n33448 , n33064 );
xor ( n33450 , n33071 , n33078 );
xor ( n33451 , n33450 , n33124 );
and ( n33452 , n33449 , n33451 );
xor ( n33453 , n33151 , n33153 );
xor ( n33454 , n33453 , n33156 );
and ( n33455 , n33451 , n33454 );
and ( n33456 , n33449 , n33454 );
or ( n33457 , n33452 , n33455 , n33456 );
xor ( n33458 , n33049 , n33067 );
xor ( n33459 , n33458 , n33127 );
and ( n33460 , n33457 , n33459 );
xor ( n33461 , n33159 , n33161 );
xor ( n33462 , n33461 , n33164 );
and ( n33463 , n33459 , n33462 );
and ( n33464 , n33457 , n33462 );
or ( n33465 , n33460 , n33463 , n33464 );
xor ( n33466 , n33130 , n33167 );
xor ( n33467 , n33466 , n33170 );
and ( n33468 , n33465 , n33467 );
xor ( n33469 , n33080 , n33081 );
xor ( n33470 , n33469 , n33121 );
xor ( n33471 , n33141 , n33144 );
xor ( n33472 , n33471 , n33148 );
and ( n33473 , n33470 , n33472 );
xor ( n33474 , n33273 , n33286 );
xor ( n33475 , n33312 , n33336 );
and ( n33476 , n33474 , n33475 );
xor ( n33477 , n33341 , n33342 );
and ( n33478 , n33475 , n33477 );
and ( n33479 , n33474 , n33477 );
or ( n33480 , n33476 , n33478 , n33479 );
and ( n33481 , n33472 , n33480 );
and ( n33482 , n33470 , n33480 );
or ( n33483 , n33473 , n33481 , n33482 );
xor ( n33484 , n33344 , n33345 );
xor ( n33485 , n33295 , n33302 );
xor ( n33486 , n33485 , n33305 );
xor ( n33487 , n33262 , n33264 );
xor ( n33488 , n33487 , n33267 );
or ( n33489 , n33486 , n33488 );
xor ( n33490 , n33319 , n33326 );
xor ( n33491 , n33490 , n33329 );
xor ( n33492 , n33275 , n33277 );
xor ( n33493 , n33492 , n33280 );
or ( n33494 , n33491 , n33493 );
and ( n33495 , n33489 , n33494 );
and ( n33496 , n33484 , n33495 );
and ( n33497 , n32868 , n30632 );
and ( n33498 , n32525 , n30685 );
and ( n33499 , n33497 , n33498 );
and ( n33500 , n31783 , n30947 );
and ( n33501 , n33498 , n33500 );
and ( n33502 , n33497 , n33500 );
or ( n33503 , n33499 , n33501 , n33502 );
and ( n33504 , n32302 , n30716 );
and ( n33505 , n32235 , n30748 );
and ( n33506 , n33504 , n33505 );
and ( n33507 , n31619 , n31066 );
and ( n33508 , n33505 , n33507 );
and ( n33509 , n33504 , n33507 );
or ( n33510 , n33506 , n33508 , n33509 );
and ( n33511 , n33503 , n33510 );
buf ( n560786 , n1245 );
buf ( n33513 , n560786 );
and ( n33514 , n33513 , n30580 );
and ( n33515 , n32019 , n30863 );
and ( n33516 , n33514 , n33515 );
and ( n33517 , n31430 , n31168 );
and ( n33518 , n33515 , n33517 );
and ( n33519 , n33514 , n33517 );
or ( n33520 , n33516 , n33518 , n33519 );
and ( n33521 , n33510 , n33520 );
and ( n33522 , n33503 , n33520 );
or ( n33523 , n33511 , n33521 , n33522 );
and ( n33524 , n33204 , n30598 );
and ( n33525 , n32940 , n30620 );
and ( n33526 , n33524 , n33525 );
and ( n33527 , n31888 , n30950 );
and ( n33528 , n33525 , n33527 );
and ( n33529 , n33524 , n33527 );
or ( n33530 , n33526 , n33528 , n33529 );
buf ( n560805 , n1244 );
buf ( n33532 , n560805 );
and ( n33533 , n30572 , n33532 );
and ( n33534 , n33530 , n33533 );
and ( n33535 , n30759 , n31997 );
and ( n33536 , n33533 , n33535 );
and ( n33537 , n33530 , n33535 );
or ( n33538 , n33534 , n33536 , n33537 );
or ( n33539 , n33523 , n33538 );
and ( n33540 , n30627 , n32850 );
and ( n33541 , n30680 , n32508 );
and ( n33542 , n33540 , n33541 );
and ( n33543 , n30962 , n31766 );
and ( n33544 , n33541 , n33543 );
and ( n33545 , n33540 , n33543 );
or ( n33546 , n33542 , n33544 , n33545 );
and ( n33547 , n30711 , n32320 );
and ( n33548 , n30759 , n32244 );
and ( n33549 , n33547 , n33548 );
and ( n33550 , n31057 , n31597 );
and ( n33551 , n33548 , n33550 );
and ( n33552 , n33547 , n33550 );
or ( n33553 , n33549 , n33551 , n33552 );
and ( n33554 , n33546 , n33553 );
buf ( n560829 , n1245 );
buf ( n33556 , n560829 );
and ( n33557 , n30572 , n33556 );
and ( n33558 , n30872 , n31997 );
and ( n33559 , n33557 , n33558 );
and ( n33560 , n31171 , n31453 );
and ( n33561 , n33558 , n33560 );
and ( n33562 , n33557 , n33560 );
or ( n33563 , n33559 , n33561 , n33562 );
and ( n33564 , n33553 , n33563 );
and ( n33565 , n33546 , n33563 );
or ( n33566 , n33554 , n33564 , n33565 );
and ( n33567 , n30601 , n33213 );
and ( n33568 , n30623 , n32922 );
and ( n33569 , n33567 , n33568 );
and ( n33570 , n30958 , n31871 );
and ( n33571 , n33568 , n33570 );
and ( n33572 , n33567 , n33570 );
or ( n33573 , n33569 , n33571 , n33572 );
buf ( n560848 , n1244 );
buf ( n33575 , n560848 );
and ( n33576 , n33575 , n30580 );
and ( n33577 , n33573 , n33576 );
and ( n33578 , n32019 , n30748 );
and ( n33579 , n33576 , n33578 );
and ( n33580 , n33573 , n33578 );
or ( n33581 , n33577 , n33579 , n33580 );
or ( n33582 , n33566 , n33581 );
and ( n33583 , n33539 , n33582 );
and ( n33584 , n33495 , n33583 );
and ( n33585 , n33484 , n33583 );
or ( n33586 , n33496 , n33584 , n33585 );
xnor ( n33587 , n33270 , n33272 );
xnor ( n33588 , n33283 , n33285 );
and ( n33589 , n33587 , n33588 );
xor ( n33590 , n33309 , n33311 );
xor ( n33591 , n33333 , n33335 );
and ( n33592 , n33590 , n33591 );
and ( n33593 , n33589 , n33592 );
xor ( n33594 , n33238 , n33240 );
xor ( n33595 , n33594 , n33242 );
xor ( n33596 , n33363 , n33364 );
and ( n33597 , n33595 , n33596 );
xor ( n33598 , n33370 , n33371 );
xor ( n33599 , n33598 , n33374 );
xor ( n33600 , n33390 , n33397 );
and ( n33601 , n33599 , n33600 );
xor ( n33602 , n33402 , n33405 );
and ( n33603 , n33600 , n33602 );
and ( n33604 , n33599 , n33602 );
or ( n33605 , n33601 , n33603 , n33604 );
and ( n33606 , n33596 , n33605 );
and ( n33607 , n33595 , n33605 );
or ( n33608 , n33597 , n33606 , n33607 );
and ( n33609 , n33592 , n33608 );
and ( n33610 , n33589 , n33608 );
or ( n33611 , n33593 , n33609 , n33610 );
and ( n33612 , n33586 , n33611 );
xor ( n33613 , n33384 , n33385 );
xor ( n33614 , n33613 , n33387 );
xor ( n33615 , n33391 , n33392 );
xor ( n33616 , n33615 , n33394 );
and ( n33617 , n33614 , n33616 );
xnor ( n33618 , n33400 , n33401 );
xnor ( n33619 , n33403 , n33404 );
and ( n33620 , n33618 , n33619 );
and ( n33621 , n33617 , n33620 );
buf ( n33622 , n31269 );
buf ( n560897 , n543215 );
buf ( n33624 , n560897 );
and ( n33625 , n33622 , n33624 );
and ( n33626 , n30578 , n33532 );
and ( n33627 , n33575 , n30583 );
and ( n33628 , n33626 , n33627 );
and ( n33629 , n33624 , n33628 );
and ( n33630 , n33622 , n33628 );
or ( n33631 , n33625 , n33629 , n33630 );
and ( n33632 , n33620 , n33631 );
and ( n33633 , n33617 , n33631 );
or ( n33634 , n33621 , n33632 , n33633 );
xor ( n33635 , n33369 , n33377 );
xor ( n33636 , n33635 , n33379 );
and ( n33637 , n33634 , n33636 );
xor ( n33638 , n33383 , n33398 );
xor ( n33639 , n33638 , n33406 );
and ( n33640 , n33636 , n33639 );
and ( n33641 , n33634 , n33639 );
or ( n33642 , n33637 , n33640 , n33641 );
xor ( n33643 , n33349 , n33350 );
xor ( n33644 , n33643 , n33352 );
and ( n33645 , n33642 , n33644 );
xor ( n33646 , n33360 , n33361 );
xor ( n33647 , n33646 , n33365 );
and ( n33648 , n33644 , n33647 );
and ( n33649 , n33642 , n33647 );
or ( n33650 , n33645 , n33648 , n33649 );
and ( n33651 , n33611 , n33650 );
and ( n33652 , n33586 , n33650 );
or ( n33653 , n33612 , n33651 , n33652 );
and ( n33654 , n33483 , n33653 );
xor ( n33655 , n33248 , n33250 );
xor ( n33656 , n33655 , n33252 );
xor ( n33657 , n33260 , n33287 );
xor ( n33658 , n33657 , n33337 );
and ( n33659 , n33656 , n33658 );
xor ( n33660 , n33343 , n33346 );
xor ( n33661 , n33660 , n33355 );
and ( n33662 , n33658 , n33661 );
and ( n33663 , n33656 , n33661 );
or ( n33664 , n33659 , n33662 , n33663 );
and ( n33665 , n33653 , n33664 );
and ( n33666 , n33483 , n33664 );
or ( n33667 , n33654 , n33665 , n33666 );
xor ( n33668 , n33199 , n33201 );
xor ( n33669 , n33668 , n33255 );
xor ( n33670 , n33340 , n33358 );
xor ( n33671 , n33670 , n33421 );
and ( n33672 , n33669 , n33671 );
xor ( n33673 , n33449 , n33451 );
xor ( n33674 , n33673 , n33454 );
and ( n33675 , n33671 , n33674 );
and ( n33676 , n33669 , n33674 );
or ( n33677 , n33672 , n33675 , n33676 );
and ( n33678 , n33667 , n33677 );
xor ( n33679 , n33197 , n33258 );
xor ( n33680 , n33679 , n33424 );
and ( n33681 , n33677 , n33680 );
and ( n33682 , n33667 , n33680 );
or ( n33683 , n33678 , n33681 , n33682 );
and ( n33684 , n33467 , n33683 );
and ( n33685 , n33465 , n33683 );
or ( n33686 , n33468 , n33684 , n33685 );
xor ( n33687 , n33190 , n33430 );
xor ( n33688 , n33687 , n33433 );
and ( n33689 , n33686 , n33688 );
xor ( n33690 , n33192 , n33194 );
xor ( n33691 , n33690 , n33427 );
xor ( n33692 , n33457 , n33459 );
xor ( n33693 , n33692 , n33462 );
xor ( n33694 , n33368 , n33415 );
xor ( n33695 , n33694 , n33418 );
xor ( n33696 , n33382 , n33409 );
xor ( n33697 , n33696 , n33412 );
xor ( n33698 , n33489 , n33494 );
xor ( n33699 , n33539 , n33582 );
and ( n33700 , n33698 , n33699 );
xor ( n33701 , n33587 , n33588 );
and ( n33702 , n33699 , n33701 );
and ( n33703 , n33698 , n33701 );
or ( n33704 , n33700 , n33702 , n33703 );
and ( n33705 , n33697 , n33704 );
xor ( n33706 , n33590 , n33591 );
xor ( n33707 , n33289 , n33290 );
xor ( n33708 , n33707 , n33292 );
xor ( n33709 , n33296 , n33297 );
xor ( n33710 , n33709 , n33299 );
and ( n33711 , n33708 , n33710 );
xor ( n33712 , n33573 , n33576 );
xor ( n33713 , n33712 , n33578 );
and ( n33714 , n33710 , n33713 );
and ( n33715 , n33708 , n33713 );
or ( n33716 , n33711 , n33714 , n33715 );
xor ( n33717 , n33313 , n33314 );
xor ( n33718 , n33717 , n33316 );
xor ( n33719 , n33320 , n33321 );
xor ( n33720 , n33719 , n33323 );
and ( n33721 , n33718 , n33720 );
xor ( n33722 , n33530 , n33533 );
xor ( n33723 , n33722 , n33535 );
and ( n33724 , n33720 , n33723 );
and ( n33725 , n33718 , n33723 );
or ( n33726 , n33721 , n33724 , n33725 );
and ( n33727 , n33716 , n33726 );
and ( n33728 , n33706 , n33727 );
and ( n33729 , n32525 , n30716 );
and ( n33730 , n32302 , n30748 );
and ( n33731 , n33729 , n33730 );
and ( n33732 , n31888 , n30947 );
and ( n33733 , n33730 , n33732 );
and ( n33734 , n33729 , n33732 );
or ( n33735 , n33731 , n33733 , n33734 );
and ( n33736 , n33575 , n30598 );
and ( n33737 , n33204 , n30620 );
and ( n33738 , n33736 , n33737 );
and ( n33739 , n32019 , n30950 );
and ( n33740 , n33737 , n33739 );
and ( n33741 , n33736 , n33739 );
or ( n33742 , n33738 , n33740 , n33741 );
and ( n33743 , n33735 , n33742 );
and ( n33744 , n32940 , n30632 );
and ( n33745 , n32868 , n30685 );
and ( n33746 , n33744 , n33745 );
and ( n33747 , n31619 , n31168 );
and ( n33748 , n33745 , n33747 );
and ( n33749 , n33744 , n33747 );
or ( n33750 , n33746 , n33748 , n33749 );
and ( n33751 , n33742 , n33750 );
and ( n33752 , n33735 , n33750 );
or ( n33753 , n33743 , n33751 , n33752 );
xor ( n33754 , n33503 , n33510 );
xor ( n33755 , n33754 , n33520 );
or ( n33756 , n33753 , n33755 );
and ( n33757 , n30711 , n32508 );
and ( n33758 , n30759 , n32320 );
and ( n33759 , n33757 , n33758 );
and ( n33760 , n30962 , n31871 );
and ( n33761 , n33758 , n33760 );
and ( n33762 , n33757 , n33760 );
or ( n33763 , n33759 , n33761 , n33762 );
and ( n33764 , n30601 , n33532 );
and ( n33765 , n30623 , n33213 );
and ( n33766 , n33764 , n33765 );
and ( n33767 , n30958 , n31997 );
and ( n33768 , n33765 , n33767 );
and ( n33769 , n33764 , n33767 );
or ( n33770 , n33766 , n33768 , n33769 );
and ( n33771 , n33763 , n33770 );
and ( n33772 , n30627 , n32922 );
and ( n33773 , n30680 , n32850 );
and ( n33774 , n33772 , n33773 );
and ( n33775 , n31171 , n31597 );
and ( n33776 , n33773 , n33775 );
and ( n33777 , n33772 , n33775 );
or ( n33778 , n33774 , n33776 , n33777 );
and ( n33779 , n33770 , n33778 );
and ( n33780 , n33763 , n33778 );
or ( n33781 , n33771 , n33779 , n33780 );
xor ( n33782 , n33546 , n33553 );
xor ( n33783 , n33782 , n33563 );
or ( n33784 , n33781 , n33783 );
and ( n33785 , n33756 , n33784 );
and ( n33786 , n33727 , n33785 );
and ( n33787 , n33706 , n33785 );
or ( n33788 , n33728 , n33786 , n33787 );
and ( n33789 , n33704 , n33788 );
and ( n33790 , n33697 , n33788 );
or ( n33791 , n33705 , n33789 , n33790 );
and ( n33792 , n33695 , n33791 );
xnor ( n33793 , n33486 , n33488 );
xnor ( n33794 , n33491 , n33493 );
and ( n33795 , n33793 , n33794 );
xnor ( n33796 , n33523 , n33538 );
xnor ( n33797 , n33566 , n33581 );
and ( n33798 , n33796 , n33797 );
and ( n33799 , n33795 , n33798 );
xor ( n33800 , n33540 , n33541 );
xor ( n33801 , n33800 , n33543 );
xor ( n33802 , n33547 , n33548 );
xor ( n33803 , n33802 , n33550 );
or ( n33804 , n33801 , n33803 );
xor ( n33805 , n33497 , n33498 );
xor ( n33806 , n33805 , n33500 );
xor ( n33807 , n33504 , n33505 );
xor ( n33808 , n33807 , n33507 );
or ( n33809 , n33806 , n33808 );
and ( n33810 , n33804 , n33809 );
and ( n33811 , n31405 , n31278 );
and ( n33812 , n31269 , n31414 );
and ( n33813 , n33811 , n33812 );
buf ( n561088 , n543218 );
buf ( n33815 , n561088 );
and ( n33816 , n33812 , n33815 );
and ( n33817 , n33811 , n33815 );
or ( n33818 , n33813 , n33816 , n33817 );
xor ( n33819 , n33614 , n33616 );
and ( n33820 , n33818 , n33819 );
xor ( n33821 , n33618 , n33619 );
and ( n33822 , n33819 , n33821 );
and ( n33823 , n33818 , n33821 );
or ( n33824 , n33820 , n33822 , n33823 );
and ( n33825 , n33810 , n33824 );
xor ( n33826 , n33599 , n33600 );
xor ( n33827 , n33826 , n33602 );
and ( n33828 , n33824 , n33827 );
and ( n33829 , n33810 , n33827 );
or ( n33830 , n33825 , n33828 , n33829 );
and ( n33831 , n33798 , n33830 );
and ( n33832 , n33795 , n33830 );
or ( n33833 , n33799 , n33831 , n33832 );
xor ( n33834 , n33474 , n33475 );
xor ( n33835 , n33834 , n33477 );
and ( n33836 , n33833 , n33835 );
xor ( n33837 , n33484 , n33495 );
xor ( n33838 , n33837 , n33583 );
and ( n33839 , n33835 , n33838 );
and ( n33840 , n33833 , n33838 );
or ( n33841 , n33836 , n33839 , n33840 );
and ( n33842 , n33791 , n33841 );
and ( n33843 , n33695 , n33841 );
or ( n33844 , n33792 , n33842 , n33843 );
xor ( n33845 , n33470 , n33472 );
xor ( n33846 , n33845 , n33480 );
xor ( n33847 , n33586 , n33611 );
xor ( n33848 , n33847 , n33650 );
and ( n33849 , n33846 , n33848 );
xor ( n33850 , n33656 , n33658 );
xor ( n33851 , n33850 , n33661 );
and ( n33852 , n33848 , n33851 );
and ( n33853 , n33846 , n33851 );
or ( n33854 , n33849 , n33852 , n33853 );
and ( n33855 , n33844 , n33854 );
xor ( n33856 , n33483 , n33653 );
xor ( n33857 , n33856 , n33664 );
and ( n33858 , n33854 , n33857 );
and ( n33859 , n33844 , n33857 );
or ( n33860 , n33855 , n33858 , n33859 );
and ( n33861 , n33693 , n33860 );
xor ( n33862 , n33667 , n33677 );
xor ( n33863 , n33862 , n33680 );
and ( n33864 , n33860 , n33863 );
and ( n33865 , n33693 , n33863 );
or ( n33866 , n33861 , n33864 , n33865 );
and ( n33867 , n33691 , n33866 );
xor ( n33868 , n33465 , n33467 );
xor ( n33869 , n33868 , n33683 );
and ( n33870 , n33866 , n33869 );
and ( n33871 , n33691 , n33869 );
or ( n33872 , n33867 , n33870 , n33871 );
and ( n33873 , n33688 , n33872 );
and ( n33874 , n33686 , n33872 );
or ( n33875 , n33689 , n33873 , n33874 );
and ( n33876 , n33447 , n33875 );
xor ( n33877 , n33686 , n33688 );
xor ( n33878 , n33877 , n33872 );
xor ( n33879 , n33691 , n33866 );
xor ( n33880 , n33879 , n33869 );
xor ( n33881 , n33669 , n33671 );
xor ( n33882 , n33881 , n33674 );
xor ( n33883 , n33589 , n33592 );
xor ( n33884 , n33883 , n33608 );
xor ( n33885 , n33642 , n33644 );
xor ( n33886 , n33885 , n33647 );
and ( n33887 , n33884 , n33886 );
xor ( n33888 , n33595 , n33596 );
xor ( n33889 , n33888 , n33605 );
xor ( n33890 , n33634 , n33636 );
xor ( n33891 , n33890 , n33639 );
and ( n33892 , n33889 , n33891 );
buf ( n561167 , n1246 );
buf ( n33894 , n561167 );
and ( n33895 , n33894 , n30580 );
and ( n33896 , n33513 , n30583 );
and ( n33897 , n33895 , n33896 );
and ( n33898 , n32235 , n30863 );
and ( n33899 , n33896 , n33898 );
and ( n33900 , n33895 , n33898 );
or ( n33901 , n33897 , n33899 , n33900 );
xor ( n33902 , n33567 , n33568 );
xor ( n33903 , n33902 , n33570 );
and ( n33904 , n33901 , n33903 );
xor ( n33905 , n33557 , n33558 );
xor ( n33906 , n33905 , n33560 );
and ( n33907 , n33903 , n33906 );
and ( n33908 , n33901 , n33906 );
or ( n33909 , n33904 , n33907 , n33908 );
xor ( n33910 , n33718 , n33720 );
xor ( n33911 , n33910 , n33723 );
or ( n33912 , n33909 , n33911 );
buf ( n561187 , n1246 );
buf ( n33914 , n561187 );
and ( n33915 , n30572 , n33914 );
and ( n33916 , n30578 , n33556 );
and ( n33917 , n33915 , n33916 );
and ( n33918 , n30872 , n32244 );
and ( n33919 , n33916 , n33918 );
and ( n33920 , n33915 , n33918 );
or ( n33921 , n33917 , n33919 , n33920 );
xor ( n33922 , n33524 , n33525 );
xor ( n33923 , n33922 , n33527 );
and ( n33924 , n33921 , n33923 );
xor ( n33925 , n33514 , n33515 );
xor ( n33926 , n33925 , n33517 );
and ( n33927 , n33923 , n33926 );
and ( n33928 , n33921 , n33926 );
or ( n33929 , n33924 , n33927 , n33928 );
xor ( n33930 , n33708 , n33710 );
xor ( n33931 , n33930 , n33713 );
or ( n33932 , n33929 , n33931 );
and ( n33933 , n33912 , n33932 );
and ( n33934 , n33891 , n33933 );
and ( n33935 , n33889 , n33933 );
or ( n33936 , n33892 , n33934 , n33935 );
and ( n33937 , n33886 , n33936 );
and ( n33938 , n33884 , n33936 );
or ( n33939 , n33887 , n33937 , n33938 );
xor ( n33940 , n33617 , n33620 );
xor ( n33941 , n33940 , n33631 );
xor ( n33942 , n33716 , n33726 );
and ( n33943 , n33941 , n33942 );
xor ( n33944 , n33756 , n33784 );
and ( n33945 , n33942 , n33944 );
and ( n33946 , n33941 , n33944 );
or ( n33947 , n33943 , n33945 , n33946 );
xor ( n33948 , n33793 , n33794 );
xor ( n33949 , n33796 , n33797 );
and ( n33950 , n33948 , n33949 );
and ( n33951 , n32868 , n30716 );
and ( n33952 , n32525 , n30748 );
and ( n33953 , n33951 , n33952 );
and ( n33954 , n31888 , n31066 );
and ( n33955 , n33952 , n33954 );
and ( n33956 , n33951 , n33954 );
or ( n33957 , n33953 , n33955 , n33956 );
and ( n33958 , n33204 , n30632 );
and ( n33959 , n32940 , n30685 );
and ( n33960 , n33958 , n33959 );
and ( n33961 , n32019 , n30947 );
and ( n33962 , n33959 , n33961 );
and ( n33963 , n33958 , n33961 );
or ( n33964 , n33960 , n33962 , n33963 );
and ( n33965 , n33957 , n33964 );
xor ( n33966 , n33757 , n33758 );
xor ( n33967 , n33966 , n33760 );
and ( n33968 , n33964 , n33967 );
and ( n33969 , n33957 , n33967 );
or ( n33970 , n33965 , n33968 , n33969 );
xor ( n33971 , n33901 , n33903 );
xor ( n33972 , n33971 , n33906 );
or ( n33973 , n33970 , n33972 );
and ( n33974 , n30711 , n32850 );
and ( n33975 , n30759 , n32508 );
and ( n33976 , n33974 , n33975 );
and ( n33977 , n31057 , n31871 );
and ( n33978 , n33975 , n33977 );
and ( n33979 , n33974 , n33977 );
or ( n33980 , n33976 , n33978 , n33979 );
and ( n33981 , n30627 , n33213 );
and ( n33982 , n30680 , n32922 );
and ( n33983 , n33981 , n33982 );
and ( n33984 , n30962 , n31997 );
and ( n33985 , n33982 , n33984 );
and ( n33986 , n33981 , n33984 );
or ( n33987 , n33983 , n33985 , n33986 );
and ( n33988 , n33980 , n33987 );
xor ( n33989 , n33729 , n33730 );
xor ( n33990 , n33989 , n33732 );
and ( n33991 , n33987 , n33990 );
and ( n33992 , n33980 , n33990 );
or ( n33993 , n33988 , n33991 , n33992 );
xor ( n33994 , n33921 , n33923 );
xor ( n33995 , n33994 , n33926 );
or ( n33996 , n33993 , n33995 );
and ( n33997 , n33973 , n33996 );
and ( n33998 , n33949 , n33997 );
and ( n33999 , n33948 , n33997 );
or ( n34000 , n33950 , n33998 , n33999 );
and ( n34001 , n33947 , n34000 );
xnor ( n34002 , n33753 , n33755 );
xnor ( n34003 , n33781 , n33783 );
and ( n34004 , n34002 , n34003 );
and ( n34005 , n31783 , n31066 );
and ( n34006 , n31430 , n31278 );
or ( n34007 , n34005 , n34006 );
and ( n34008 , n31057 , n31766 );
and ( n34009 , n31269 , n31453 );
or ( n34010 , n34008 , n34009 );
and ( n34011 , n34007 , n34010 );
xor ( n34012 , n33622 , n33624 );
xor ( n34013 , n34012 , n33628 );
and ( n34014 , n34011 , n34013 );
xor ( n34015 , n33804 , n33809 );
and ( n34016 , n34013 , n34015 );
and ( n34017 , n34011 , n34015 );
or ( n34018 , n34014 , n34016 , n34017 );
and ( n34019 , n34004 , n34018 );
xor ( n34020 , n33915 , n33916 );
xor ( n34021 , n34020 , n33918 );
xor ( n34022 , n33764 , n33765 );
xor ( n34023 , n34022 , n33767 );
or ( n34024 , n34021 , n34023 );
xor ( n34025 , n33895 , n33896 );
xor ( n34026 , n34025 , n33898 );
xor ( n34027 , n33736 , n33737 );
xor ( n34028 , n34027 , n33739 );
or ( n34029 , n34026 , n34028 );
and ( n34030 , n34024 , n34029 );
buf ( n561305 , n1247 );
buf ( n34032 , n561305 );
and ( n34033 , n30572 , n34032 );
and ( n34034 , n30872 , n32320 );
and ( n34035 , n34033 , n34034 );
and ( n34036 , n31171 , n31766 );
and ( n34037 , n34034 , n34036 );
and ( n34038 , n34033 , n34036 );
or ( n34039 , n34035 , n34037 , n34038 );
and ( n34040 , n30578 , n33914 );
and ( n34041 , n30958 , n32244 );
and ( n34042 , n34040 , n34041 );
and ( n34043 , n31269 , n31597 );
and ( n34044 , n34041 , n34043 );
and ( n34045 , n34040 , n34043 );
or ( n34046 , n34042 , n34044 , n34045 );
or ( n34047 , n34039 , n34046 );
buf ( n561322 , n1247 );
buf ( n34049 , n561322 );
and ( n34050 , n34049 , n30580 );
and ( n34051 , n32302 , n30863 );
and ( n34052 , n34050 , n34051 );
and ( n34053 , n31783 , n31168 );
and ( n34054 , n34051 , n34053 );
and ( n34055 , n34050 , n34053 );
or ( n34056 , n34052 , n34054 , n34055 );
and ( n34057 , n33894 , n30583 );
and ( n34058 , n32235 , n30950 );
and ( n34059 , n34057 , n34058 );
and ( n34060 , n31619 , n31278 );
and ( n34061 , n34058 , n34060 );
and ( n34062 , n34057 , n34060 );
or ( n34063 , n34059 , n34061 , n34062 );
or ( n34064 , n34056 , n34063 );
and ( n34065 , n34047 , n34064 );
and ( n34066 , n34030 , n34065 );
xor ( n34067 , n33763 , n33770 );
xor ( n34068 , n34067 , n33778 );
xor ( n34069 , n33735 , n33742 );
xor ( n34070 , n34069 , n33750 );
and ( n34071 , n34068 , n34070 );
and ( n34072 , n34065 , n34071 );
and ( n34073 , n34030 , n34071 );
or ( n34074 , n34066 , n34072 , n34073 );
and ( n34075 , n34018 , n34074 );
and ( n34076 , n34004 , n34074 );
or ( n34077 , n34019 , n34075 , n34076 );
and ( n34078 , n34000 , n34077 );
and ( n34079 , n33947 , n34077 );
or ( n34080 , n34001 , n34078 , n34079 );
xor ( n34081 , n33698 , n33699 );
xor ( n34082 , n34081 , n33701 );
xor ( n34083 , n33706 , n33727 );
xor ( n34084 , n34083 , n33785 );
and ( n34085 , n34082 , n34084 );
xor ( n34086 , n33795 , n33798 );
xor ( n34087 , n34086 , n33830 );
and ( n34088 , n34084 , n34087 );
and ( n34089 , n34082 , n34087 );
or ( n34090 , n34085 , n34088 , n34089 );
and ( n34091 , n34080 , n34090 );
xor ( n34092 , n33697 , n33704 );
xor ( n34093 , n34092 , n33788 );
and ( n34094 , n34090 , n34093 );
and ( n34095 , n34080 , n34093 );
or ( n34096 , n34091 , n34094 , n34095 );
and ( n34097 , n33939 , n34096 );
xor ( n34098 , n33695 , n33791 );
xor ( n34099 , n34098 , n33841 );
and ( n34100 , n34096 , n34099 );
and ( n34101 , n33939 , n34099 );
or ( n34102 , n34097 , n34100 , n34101 );
and ( n34103 , n33882 , n34102 );
xor ( n34104 , n33844 , n33854 );
xor ( n34105 , n34104 , n33857 );
and ( n34106 , n34102 , n34105 );
and ( n34107 , n33882 , n34105 );
or ( n34108 , n34103 , n34106 , n34107 );
xor ( n34109 , n33693 , n33860 );
xor ( n34110 , n34109 , n33863 );
and ( n34111 , n34108 , n34110 );
xor ( n34112 , n33846 , n33848 );
xor ( n34113 , n34112 , n33851 );
xor ( n34114 , n33833 , n33835 );
xor ( n34115 , n34114 , n33838 );
xnor ( n34116 , n33801 , n33803 );
xnor ( n34117 , n33806 , n33808 );
and ( n34118 , n34116 , n34117 );
xor ( n34119 , n33626 , n33627 );
xor ( n34120 , n33811 , n33812 );
xor ( n34121 , n34120 , n33815 );
and ( n34122 , n34119 , n34121 );
xor ( n34123 , n34007 , n34010 );
and ( n34124 , n34121 , n34123 );
and ( n34125 , n34119 , n34123 );
or ( n34126 , n34122 , n34124 , n34125 );
and ( n34127 , n34118 , n34126 );
and ( n34128 , n33513 , n30598 );
and ( n34129 , n33575 , n30620 );
and ( n34130 , n34128 , n34129 );
and ( n34131 , n30601 , n33556 );
and ( n34132 , n30623 , n33532 );
and ( n34133 , n34131 , n34132 );
and ( n34134 , n34130 , n34133 );
xor ( n34135 , n33744 , n33745 );
xor ( n34136 , n34135 , n33747 );
xor ( n34137 , n33772 , n33773 );
xor ( n34138 , n34137 , n33775 );
and ( n34139 , n34136 , n34138 );
and ( n34140 , n34134 , n34139 );
buf ( n34141 , n31405 );
buf ( n561416 , n543221 );
buf ( n34143 , n561416 );
and ( n34144 , n34141 , n34143 );
and ( n34145 , n31430 , n31414 );
and ( n34146 , n31405 , n31453 );
and ( n34147 , n34145 , n34146 );
buf ( n561422 , n543224 );
buf ( n34149 , n561422 );
and ( n34150 , n34146 , n34149 );
and ( n34151 , n34145 , n34149 );
or ( n34152 , n34147 , n34150 , n34151 );
and ( n34153 , n34143 , n34152 );
and ( n34154 , n34141 , n34152 );
or ( n34155 , n34144 , n34153 , n34154 );
and ( n34156 , n34139 , n34155 );
and ( n34157 , n34134 , n34155 );
or ( n34158 , n34140 , n34156 , n34157 );
and ( n34159 , n34126 , n34158 );
and ( n34160 , n34118 , n34158 );
or ( n34161 , n34127 , n34159 , n34160 );
xor ( n34162 , n33810 , n33824 );
xor ( n34163 , n34162 , n33827 );
and ( n34164 , n34161 , n34163 );
xor ( n34165 , n33912 , n33932 );
and ( n34166 , n34163 , n34165 );
and ( n34167 , n34161 , n34165 );
or ( n34168 , n34164 , n34166 , n34167 );
xnor ( n34169 , n33909 , n33911 );
xnor ( n34170 , n33929 , n33931 );
and ( n34171 , n34169 , n34170 );
xor ( n34172 , n33818 , n33819 );
xor ( n34173 , n34172 , n33821 );
xor ( n34174 , n33973 , n33996 );
and ( n34175 , n34173 , n34174 );
xor ( n34176 , n34002 , n34003 );
and ( n34177 , n34174 , n34176 );
and ( n34178 , n34173 , n34176 );
or ( n34179 , n34175 , n34177 , n34178 );
and ( n34180 , n34171 , n34179 );
xnor ( n34181 , n34008 , n34009 );
not ( n34182 , n34181 );
xnor ( n34183 , n34026 , n34028 );
and ( n34184 , n34182 , n34183 );
xnor ( n34185 , n34005 , n34006 );
not ( n34186 , n34185 );
xnor ( n34187 , n34021 , n34023 );
and ( n34188 , n34186 , n34187 );
and ( n34189 , n34184 , n34188 );
buf ( n34190 , n34181 );
buf ( n34191 , n34185 );
and ( n34192 , n34190 , n34191 );
and ( n34193 , n34189 , n34192 );
and ( n34194 , n33575 , n30632 );
and ( n34195 , n32235 , n30947 );
and ( n34196 , n34194 , n34195 );
and ( n34197 , n31783 , n31278 );
and ( n34198 , n34195 , n34197 );
and ( n34199 , n34194 , n34197 );
or ( n34200 , n34196 , n34198 , n34199 );
and ( n34201 , n33894 , n30598 );
and ( n34202 , n33513 , n30620 );
and ( n34203 , n34201 , n34202 );
and ( n34204 , n32302 , n30950 );
and ( n34205 , n34202 , n34204 );
and ( n34206 , n34201 , n34204 );
or ( n34207 , n34203 , n34205 , n34206 );
and ( n34208 , n34200 , n34207 );
xor ( n34209 , n34040 , n34041 );
xor ( n34210 , n34209 , n34043 );
and ( n34211 , n34207 , n34210 );
and ( n34212 , n34200 , n34210 );
or ( n34213 , n34208 , n34211 , n34212 );
not ( n34214 , n34213 );
xor ( n34215 , n33957 , n33964 );
xor ( n34216 , n34215 , n33967 );
and ( n34217 , n34214 , n34216 );
and ( n34218 , n30627 , n33532 );
and ( n34219 , n30962 , n32244 );
and ( n34220 , n34218 , n34219 );
and ( n34221 , n31269 , n31766 );
and ( n34222 , n34219 , n34221 );
and ( n34223 , n34218 , n34221 );
or ( n34224 , n34220 , n34222 , n34223 );
and ( n34225 , n30601 , n33914 );
and ( n34226 , n30623 , n33556 );
and ( n34227 , n34225 , n34226 );
and ( n34228 , n30958 , n32320 );
and ( n34229 , n34226 , n34228 );
and ( n34230 , n34225 , n34228 );
or ( n34231 , n34227 , n34229 , n34230 );
and ( n34232 , n34224 , n34231 );
xor ( n34233 , n34057 , n34058 );
xor ( n34234 , n34233 , n34060 );
and ( n34235 , n34231 , n34234 );
and ( n34236 , n34224 , n34234 );
or ( n34237 , n34232 , n34235 , n34236 );
not ( n34238 , n34237 );
xor ( n34239 , n33980 , n33987 );
xor ( n34240 , n34239 , n33990 );
and ( n34241 , n34238 , n34240 );
and ( n34242 , n34217 , n34241 );
and ( n34243 , n34192 , n34242 );
and ( n34244 , n34189 , n34242 );
or ( n34245 , n34193 , n34243 , n34244 );
and ( n34246 , n34179 , n34245 );
and ( n34247 , n34171 , n34245 );
or ( n34248 , n34180 , n34246 , n34247 );
and ( n34249 , n34168 , n34248 );
buf ( n34250 , n34213 );
buf ( n34251 , n34237 );
and ( n34252 , n34250 , n34251 );
xnor ( n34253 , n33970 , n33972 );
xnor ( n34254 , n33993 , n33995 );
and ( n34255 , n34253 , n34254 );
and ( n34256 , n34252 , n34255 );
xor ( n34257 , n34024 , n34029 );
xor ( n34258 , n34047 , n34064 );
and ( n34259 , n34257 , n34258 );
xor ( n34260 , n34068 , n34070 );
and ( n34261 , n34258 , n34260 );
and ( n34262 , n34257 , n34260 );
or ( n34263 , n34259 , n34261 , n34262 );
and ( n34264 , n34255 , n34263 );
and ( n34265 , n34252 , n34263 );
or ( n34266 , n34256 , n34264 , n34265 );
xor ( n34267 , n34116 , n34117 );
xor ( n34268 , n34050 , n34051 );
xor ( n34269 , n34268 , n34053 );
xor ( n34270 , n33951 , n33952 );
xor ( n34271 , n34270 , n33954 );
and ( n34272 , n34269 , n34271 );
xor ( n34273 , n33958 , n33959 );
xor ( n34274 , n34273 , n33961 );
and ( n34275 , n34271 , n34274 );
and ( n34276 , n34269 , n34274 );
or ( n34277 , n34272 , n34275 , n34276 );
xor ( n34278 , n34033 , n34034 );
xor ( n34279 , n34278 , n34036 );
xor ( n34280 , n33974 , n33975 );
xor ( n34281 , n34280 , n33977 );
and ( n34282 , n34279 , n34281 );
xor ( n34283 , n33981 , n33982 );
xor ( n34284 , n34283 , n33984 );
and ( n34285 , n34281 , n34284 );
and ( n34286 , n34279 , n34284 );
or ( n34287 , n34282 , n34285 , n34286 );
and ( n34288 , n34277 , n34287 );
and ( n34289 , n34267 , n34288 );
and ( n34290 , n30680 , n33213 );
and ( n34291 , n30711 , n32922 );
and ( n34292 , n34290 , n34291 );
and ( n34293 , n31057 , n31997 );
and ( n34294 , n34291 , n34293 );
and ( n34295 , n34290 , n34293 );
or ( n34296 , n34292 , n34294 , n34295 );
buf ( n561571 , n1248 );
buf ( n34298 , n561571 );
and ( n34299 , n30572 , n34298 );
and ( n34300 , n30759 , n32850 );
and ( n34301 , n34299 , n34300 );
and ( n34302 , n30872 , n32508 );
and ( n34303 , n34300 , n34302 );
and ( n34304 , n34299 , n34302 );
or ( n34305 , n34301 , n34303 , n34304 );
or ( n34306 , n34296 , n34305 );
and ( n34307 , n33204 , n30685 );
and ( n34308 , n32940 , n30716 );
and ( n34309 , n34307 , n34308 );
and ( n34310 , n32019 , n31066 );
and ( n34311 , n34308 , n34310 );
and ( n34312 , n34307 , n34310 );
or ( n34313 , n34309 , n34311 , n34312 );
buf ( n561588 , n1248 );
buf ( n34315 , n561588 );
and ( n34316 , n34315 , n30580 );
and ( n34317 , n32868 , n30748 );
and ( n34318 , n34316 , n34317 );
and ( n34319 , n32525 , n30863 );
and ( n34320 , n34317 , n34319 );
and ( n34321 , n34316 , n34319 );
or ( n34322 , n34318 , n34320 , n34321 );
or ( n34323 , n34313 , n34322 );
and ( n34324 , n34306 , n34323 );
and ( n34325 , n34288 , n34324 );
and ( n34326 , n34267 , n34324 );
or ( n34327 , n34289 , n34325 , n34326 );
xnor ( n34328 , n34039 , n34046 );
xnor ( n34329 , n34056 , n34063 );
and ( n34330 , n34328 , n34329 );
xor ( n34331 , n34130 , n34133 );
xor ( n34332 , n34136 , n34138 );
and ( n34333 , n34331 , n34332 );
and ( n34334 , n31888 , n31168 );
and ( n34335 , n31619 , n31414 );
or ( n34336 , n34334 , n34335 );
and ( n34337 , n31171 , n31871 );
and ( n34338 , n31405 , n31597 );
or ( n34339 , n34337 , n34338 );
and ( n34340 , n34336 , n34339 );
and ( n34341 , n34332 , n34340 );
and ( n34342 , n34331 , n34340 );
or ( n34343 , n34333 , n34341 , n34342 );
and ( n34344 , n34330 , n34343 );
xor ( n34345 , n34119 , n34121 );
xor ( n34346 , n34345 , n34123 );
and ( n34347 , n34343 , n34346 );
and ( n34348 , n34330 , n34346 );
or ( n34349 , n34344 , n34347 , n34348 );
and ( n34350 , n34327 , n34349 );
xor ( n34351 , n34011 , n34013 );
xor ( n34352 , n34351 , n34015 );
and ( n34353 , n34349 , n34352 );
and ( n34354 , n34327 , n34352 );
or ( n34355 , n34350 , n34353 , n34354 );
and ( n34356 , n34266 , n34355 );
xor ( n34357 , n33941 , n33942 );
xor ( n34358 , n34357 , n33944 );
and ( n34359 , n34355 , n34358 );
and ( n34360 , n34266 , n34358 );
or ( n34361 , n34356 , n34359 , n34360 );
and ( n34362 , n34248 , n34361 );
and ( n34363 , n34168 , n34361 );
or ( n34364 , n34249 , n34362 , n34363 );
and ( n34365 , n34115 , n34364 );
xor ( n34366 , n33889 , n33891 );
xor ( n34367 , n34366 , n33933 );
xor ( n34368 , n33947 , n34000 );
xor ( n34369 , n34368 , n34077 );
and ( n34370 , n34367 , n34369 );
xor ( n34371 , n34082 , n34084 );
xor ( n34372 , n34371 , n34087 );
and ( n34373 , n34369 , n34372 );
and ( n34374 , n34367 , n34372 );
or ( n34375 , n34370 , n34373 , n34374 );
and ( n34376 , n34364 , n34375 );
and ( n34377 , n34115 , n34375 );
or ( n34378 , n34365 , n34376 , n34377 );
and ( n34379 , n34113 , n34378 );
xor ( n34380 , n33939 , n34096 );
xor ( n34381 , n34380 , n34099 );
and ( n34382 , n34378 , n34381 );
and ( n34383 , n34113 , n34381 );
or ( n34384 , n34379 , n34382 , n34383 );
xor ( n34385 , n33882 , n34102 );
xor ( n34386 , n34385 , n34105 );
and ( n34387 , n34384 , n34386 );
xor ( n34388 , n33884 , n33886 );
xor ( n34389 , n34388 , n33936 );
xor ( n34390 , n34080 , n34090 );
xor ( n34391 , n34390 , n34093 );
and ( n34392 , n34389 , n34391 );
xor ( n34393 , n33948 , n33949 );
xor ( n34394 , n34393 , n33997 );
xor ( n34395 , n34004 , n34018 );
xor ( n34396 , n34395 , n34074 );
and ( n34397 , n34394 , n34396 );
xor ( n34398 , n34030 , n34065 );
xor ( n34399 , n34398 , n34071 );
xor ( n34400 , n34118 , n34126 );
xor ( n34401 , n34400 , n34158 );
and ( n34402 , n34399 , n34401 );
xor ( n34403 , n34169 , n34170 );
and ( n34404 , n34401 , n34403 );
and ( n34405 , n34399 , n34403 );
or ( n34406 , n34402 , n34404 , n34405 );
and ( n34407 , n34396 , n34406 );
and ( n34408 , n34394 , n34406 );
or ( n34409 , n34397 , n34407 , n34408 );
xor ( n34410 , n34134 , n34139 );
xor ( n34411 , n34410 , n34155 );
xor ( n34412 , n34184 , n34188 );
and ( n34413 , n34411 , n34412 );
xor ( n34414 , n34190 , n34191 );
and ( n34415 , n34412 , n34414 );
and ( n34416 , n34411 , n34414 );
or ( n34417 , n34413 , n34415 , n34416 );
xor ( n34418 , n34217 , n34241 );
xor ( n34419 , n34250 , n34251 );
and ( n34420 , n34418 , n34419 );
xor ( n34421 , n34253 , n34254 );
and ( n34422 , n34419 , n34421 );
and ( n34423 , n34418 , n34421 );
or ( n34424 , n34420 , n34422 , n34423 );
and ( n34425 , n34417 , n34424 );
xor ( n34426 , n34182 , n34183 );
xor ( n34427 , n34186 , n34187 );
and ( n34428 , n34426 , n34427 );
xor ( n34429 , n34214 , n34216 );
xor ( n34430 , n34238 , n34240 );
and ( n34431 , n34429 , n34430 );
and ( n34432 , n34428 , n34431 );
xor ( n34433 , n34128 , n34129 );
xor ( n34434 , n34131 , n34132 );
and ( n34435 , n34433 , n34434 );
xor ( n34436 , n34141 , n34143 );
xor ( n34437 , n34436 , n34152 );
and ( n34438 , n34435 , n34437 );
xor ( n34439 , n34277 , n34287 );
and ( n34440 , n34437 , n34439 );
and ( n34441 , n34435 , n34439 );
or ( n34442 , n34438 , n34440 , n34441 );
and ( n34443 , n34431 , n34442 );
and ( n34444 , n34428 , n34442 );
or ( n34445 , n34432 , n34443 , n34444 );
and ( n34446 , n34424 , n34445 );
and ( n34447 , n34417 , n34445 );
or ( n34448 , n34425 , n34446 , n34447 );
xor ( n34449 , n34306 , n34323 );
xor ( n34450 , n34328 , n34329 );
and ( n34451 , n34449 , n34450 );
buf ( n561726 , n1249 );
buf ( n34453 , n561726 );
and ( n34454 , n30572 , n34453 );
and ( n34455 , n30872 , n32850 );
and ( n34456 , n34454 , n34455 );
and ( n34457 , n31269 , n31871 );
and ( n34458 , n34455 , n34457 );
and ( n34459 , n34454 , n34457 );
or ( n34460 , n34456 , n34458 , n34459 );
and ( n34461 , n30711 , n33213 );
and ( n34462 , n30759 , n32922 );
and ( n34463 , n34461 , n34462 );
and ( n34464 , n31171 , n31997 );
and ( n34465 , n34462 , n34464 );
and ( n34466 , n34461 , n34464 );
or ( n34467 , n34463 , n34465 , n34466 );
and ( n34468 , n34460 , n34467 );
and ( n34469 , n30578 , n34298 );
and ( n34470 , n30601 , n34032 );
and ( n34471 , n34469 , n34470 );
and ( n34472 , n30958 , n32508 );
and ( n34473 , n34470 , n34472 );
and ( n34474 , n34469 , n34472 );
or ( n34475 , n34471 , n34473 , n34474 );
and ( n34476 , n34467 , n34475 );
and ( n34477 , n34460 , n34475 );
or ( n34478 , n34468 , n34476 , n34477 );
buf ( n561753 , n1249 );
buf ( n34480 , n561753 );
and ( n34481 , n34480 , n30580 );
and ( n34482 , n32868 , n30863 );
and ( n34483 , n34481 , n34482 );
and ( n34484 , n31888 , n31278 );
and ( n34485 , n34482 , n34484 );
and ( n34486 , n34481 , n34484 );
or ( n34487 , n34483 , n34485 , n34486 );
and ( n34488 , n33204 , n30716 );
and ( n34489 , n32940 , n30748 );
and ( n34490 , n34488 , n34489 );
and ( n34491 , n32019 , n31168 );
and ( n34492 , n34489 , n34491 );
and ( n34493 , n34488 , n34491 );
or ( n34494 , n34490 , n34492 , n34493 );
and ( n34495 , n34487 , n34494 );
and ( n34496 , n34315 , n30583 );
and ( n34497 , n34049 , n30598 );
and ( n34498 , n34496 , n34497 );
and ( n34499 , n32525 , n30950 );
and ( n34500 , n34497 , n34499 );
and ( n34501 , n34496 , n34499 );
or ( n34502 , n34498 , n34500 , n34501 );
and ( n34503 , n34494 , n34502 );
and ( n34504 , n34487 , n34502 );
or ( n34505 , n34495 , n34503 , n34504 );
and ( n34506 , n34478 , n34505 );
and ( n34507 , n34450 , n34506 );
and ( n34508 , n34449 , n34506 );
or ( n34509 , n34451 , n34507 , n34508 );
xor ( n34510 , n34194 , n34195 );
xor ( n34511 , n34510 , n34197 );
xor ( n34512 , n34307 , n34308 );
xor ( n34513 , n34512 , n34310 );
and ( n34514 , n34511 , n34513 );
xor ( n34515 , n34201 , n34202 );
xor ( n34516 , n34515 , n34204 );
and ( n34517 , n34513 , n34516 );
and ( n34518 , n34511 , n34516 );
or ( n34519 , n34514 , n34517 , n34518 );
xor ( n34520 , n34218 , n34219 );
xor ( n34521 , n34520 , n34221 );
xor ( n34522 , n34290 , n34291 );
xor ( n34523 , n34522 , n34293 );
and ( n34524 , n34521 , n34523 );
xor ( n34525 , n34225 , n34226 );
xor ( n34526 , n34525 , n34228 );
and ( n34527 , n34523 , n34526 );
and ( n34528 , n34521 , n34526 );
or ( n34529 , n34524 , n34527 , n34528 );
and ( n34530 , n34519 , n34529 );
and ( n34531 , n30962 , n32320 );
and ( n34532 , n31405 , n31766 );
and ( n34533 , n34531 , n34532 );
and ( n34534 , n31430 , n31597 );
and ( n34535 , n34532 , n34534 );
and ( n34536 , n34531 , n34534 );
or ( n34537 , n34533 , n34535 , n34536 );
and ( n34538 , n34049 , n30583 );
or ( n34539 , n34537 , n34538 );
and ( n34540 , n32302 , n30947 );
and ( n34541 , n31783 , n31414 );
and ( n34542 , n34540 , n34541 );
and ( n34543 , n31619 , n31453 );
and ( n34544 , n34541 , n34543 );
and ( n34545 , n34540 , n34543 );
or ( n34546 , n34542 , n34544 , n34545 );
and ( n34547 , n30578 , n34032 );
or ( n34548 , n34546 , n34547 );
and ( n34549 , n34539 , n34548 );
and ( n34550 , n34530 , n34549 );
and ( n34551 , n30627 , n33556 );
and ( n34552 , n30680 , n33532 );
and ( n34553 , n34551 , n34552 );
and ( n34554 , n31057 , n32244 );
and ( n34555 , n34552 , n34554 );
and ( n34556 , n34551 , n34554 );
or ( n34557 , n34553 , n34555 , n34556 );
xor ( n34558 , n34299 , n34300 );
xor ( n34559 , n34558 , n34302 );
or ( n34560 , n34557 , n34559 );
and ( n34561 , n33513 , n30632 );
and ( n34562 , n33575 , n30685 );
and ( n34563 , n34561 , n34562 );
and ( n34564 , n32235 , n31066 );
and ( n34565 , n34562 , n34564 );
and ( n34566 , n34561 , n34564 );
or ( n34567 , n34563 , n34565 , n34566 );
xor ( n34568 , n34316 , n34317 );
xor ( n34569 , n34568 , n34319 );
or ( n34570 , n34567 , n34569 );
and ( n34571 , n34560 , n34570 );
and ( n34572 , n34549 , n34571 );
and ( n34573 , n34530 , n34571 );
or ( n34574 , n34550 , n34572 , n34573 );
and ( n34575 , n34509 , n34574 );
xor ( n34576 , n34224 , n34231 );
xor ( n34577 , n34576 , n34234 );
xor ( n34578 , n34200 , n34207 );
xor ( n34579 , n34578 , n34210 );
and ( n34580 , n34577 , n34579 );
xor ( n34581 , n34269 , n34271 );
xor ( n34582 , n34581 , n34274 );
xor ( n34583 , n34279 , n34281 );
xor ( n34584 , n34583 , n34284 );
and ( n34585 , n34582 , n34584 );
and ( n34586 , n34580 , n34585 );
xnor ( n34587 , n34296 , n34305 );
xnor ( n34588 , n34313 , n34322 );
and ( n34589 , n34587 , n34588 );
and ( n34590 , n34585 , n34589 );
and ( n34591 , n34580 , n34589 );
or ( n34592 , n34586 , n34590 , n34591 );
and ( n34593 , n34574 , n34592 );
and ( n34594 , n34509 , n34592 );
or ( n34595 , n34575 , n34593 , n34594 );
xor ( n34596 , n34257 , n34258 );
xor ( n34597 , n34596 , n34260 );
xor ( n34598 , n34267 , n34288 );
xor ( n34599 , n34598 , n34324 );
and ( n34600 , n34597 , n34599 );
xor ( n34601 , n34330 , n34343 );
xor ( n34602 , n34601 , n34346 );
and ( n34603 , n34599 , n34602 );
and ( n34604 , n34597 , n34602 );
or ( n34605 , n34600 , n34603 , n34604 );
and ( n34606 , n34595 , n34605 );
xor ( n34607 , n34173 , n34174 );
xor ( n34608 , n34607 , n34176 );
and ( n34609 , n34605 , n34608 );
and ( n34610 , n34595 , n34608 );
or ( n34611 , n34606 , n34609 , n34610 );
and ( n34612 , n34448 , n34611 );
xor ( n34613 , n34189 , n34192 );
xor ( n34614 , n34613 , n34242 );
xor ( n34615 , n34252 , n34255 );
xor ( n34616 , n34615 , n34263 );
and ( n34617 , n34614 , n34616 );
xor ( n34618 , n34327 , n34349 );
xor ( n34619 , n34618 , n34352 );
and ( n34620 , n34616 , n34619 );
and ( n34621 , n34614 , n34619 );
or ( n34622 , n34617 , n34620 , n34621 );
and ( n34623 , n34611 , n34622 );
and ( n34624 , n34448 , n34622 );
or ( n34625 , n34612 , n34623 , n34624 );
and ( n34626 , n34409 , n34625 );
xor ( n34627 , n34161 , n34163 );
xor ( n34628 , n34627 , n34165 );
xor ( n34629 , n34171 , n34179 );
xor ( n34630 , n34629 , n34245 );
and ( n34631 , n34628 , n34630 );
xor ( n34632 , n34266 , n34355 );
xor ( n34633 , n34632 , n34358 );
and ( n34634 , n34630 , n34633 );
and ( n34635 , n34628 , n34633 );
or ( n34636 , n34631 , n34634 , n34635 );
and ( n34637 , n34625 , n34636 );
and ( n34638 , n34409 , n34636 );
or ( n34639 , n34626 , n34637 , n34638 );
and ( n34640 , n34391 , n34639 );
and ( n34641 , n34389 , n34639 );
or ( n34642 , n34392 , n34640 , n34641 );
xor ( n34643 , n34113 , n34378 );
xor ( n34644 , n34643 , n34381 );
and ( n34645 , n34642 , n34644 );
xor ( n34646 , n34115 , n34364 );
xor ( n34647 , n34646 , n34375 );
xor ( n34648 , n34168 , n34248 );
xor ( n34649 , n34648 , n34361 );
xor ( n34650 , n34367 , n34369 );
xor ( n34651 , n34650 , n34372 );
and ( n34652 , n34649 , n34651 );
xor ( n34653 , n34145 , n34146 );
xor ( n34654 , n34653 , n34149 );
xor ( n34655 , n34336 , n34339 );
and ( n34656 , n34654 , n34655 );
xor ( n34657 , n34433 , n34434 );
and ( n34658 , n34655 , n34657 );
and ( n34659 , n34654 , n34657 );
or ( n34660 , n34656 , n34658 , n34659 );
xor ( n34661 , n34331 , n34332 );
xor ( n34662 , n34661 , n34340 );
and ( n34663 , n34660 , n34662 );
xor ( n34664 , n34426 , n34427 );
and ( n34665 , n34662 , n34664 );
and ( n34666 , n34660 , n34664 );
or ( n34667 , n34663 , n34665 , n34666 );
xor ( n34668 , n34429 , n34430 );
and ( n34669 , n33894 , n30632 );
and ( n34670 , n33513 , n30685 );
and ( n34671 , n34669 , n34670 );
and ( n34672 , n32525 , n30947 );
and ( n34673 , n34670 , n34672 );
and ( n34674 , n34669 , n34672 );
or ( n34675 , n34671 , n34673 , n34674 );
xor ( n34676 , n34551 , n34552 );
xor ( n34677 , n34676 , n34554 );
and ( n34678 , n34675 , n34677 );
xor ( n34679 , n34531 , n34532 );
xor ( n34680 , n34679 , n34534 );
and ( n34681 , n34677 , n34680 );
and ( n34682 , n34675 , n34680 );
or ( n34683 , n34678 , n34681 , n34682 );
xor ( n34684 , n34487 , n34494 );
xor ( n34685 , n34684 , n34502 );
or ( n34686 , n34683 , n34685 );
and ( n34687 , n30627 , n33914 );
and ( n34688 , n30680 , n33556 );
and ( n34689 , n34687 , n34688 );
and ( n34690 , n30962 , n32508 );
and ( n34691 , n34688 , n34690 );
and ( n34692 , n34687 , n34690 );
or ( n34693 , n34689 , n34691 , n34692 );
xor ( n34694 , n34561 , n34562 );
xor ( n34695 , n34694 , n34564 );
and ( n34696 , n34693 , n34695 );
xor ( n34697 , n34540 , n34541 );
xor ( n34698 , n34697 , n34543 );
and ( n34699 , n34695 , n34698 );
and ( n34700 , n34693 , n34698 );
or ( n34701 , n34696 , n34699 , n34700 );
xor ( n34702 , n34460 , n34467 );
xor ( n34703 , n34702 , n34475 );
or ( n34704 , n34701 , n34703 );
and ( n34705 , n34686 , n34704 );
and ( n34706 , n34668 , n34705 );
xnor ( n34707 , n34334 , n34335 );
xnor ( n34708 , n34337 , n34338 );
and ( n34709 , n34707 , n34708 );
buf ( n34710 , n31430 );
buf ( n561985 , n543227 );
buf ( n34712 , n561985 );
and ( n34713 , n34710 , n34712 );
and ( n34714 , n30623 , n33914 );
and ( n34715 , n33894 , n30620 );
and ( n34716 , n34714 , n34715 );
and ( n34717 , n34712 , n34716 );
and ( n34718 , n34710 , n34716 );
or ( n34719 , n34713 , n34717 , n34718 );
and ( n34720 , n34709 , n34719 );
xor ( n34721 , n34478 , n34505 );
and ( n34722 , n34719 , n34721 );
and ( n34723 , n34709 , n34721 );
or ( n34724 , n34720 , n34722 , n34723 );
and ( n34725 , n34705 , n34724 );
and ( n34726 , n34668 , n34724 );
or ( n34727 , n34706 , n34725 , n34726 );
and ( n34728 , n34667 , n34727 );
xor ( n34729 , n34519 , n34529 );
xor ( n34730 , n34539 , n34548 );
and ( n34731 , n34729 , n34730 );
xor ( n34732 , n34560 , n34570 );
and ( n34733 , n34730 , n34732 );
and ( n34734 , n34729 , n34732 );
or ( n34735 , n34731 , n34733 , n34734 );
xor ( n34736 , n34577 , n34579 );
xor ( n34737 , n34582 , n34584 );
and ( n34738 , n34736 , n34737 );
xor ( n34739 , n34587 , n34588 );
and ( n34740 , n34737 , n34739 );
and ( n34741 , n34736 , n34739 );
or ( n34742 , n34738 , n34740 , n34741 );
and ( n34743 , n34735 , n34742 );
and ( n34744 , n30711 , n33532 );
and ( n34745 , n31057 , n32320 );
and ( n34746 , n34744 , n34745 );
and ( n34747 , n31405 , n31871 );
and ( n34748 , n34745 , n34747 );
and ( n34749 , n34744 , n34747 );
or ( n34750 , n34746 , n34748 , n34749 );
and ( n34751 , n30578 , n34453 );
and ( n34752 , n30958 , n32850 );
and ( n34753 , n34751 , n34752 );
and ( n34754 , n31269 , n31997 );
and ( n34755 , n34752 , n34754 );
and ( n34756 , n34751 , n34754 );
or ( n34757 , n34753 , n34755 , n34756 );
and ( n34758 , n34750 , n34757 );
and ( n34759 , n30759 , n33213 );
and ( n34760 , n30872 , n32922 );
and ( n34761 , n34759 , n34760 );
and ( n34762 , n31171 , n32244 );
and ( n34763 , n34760 , n34762 );
and ( n34764 , n34759 , n34762 );
or ( n34765 , n34761 , n34763 , n34764 );
and ( n34766 , n34757 , n34765 );
and ( n34767 , n34750 , n34765 );
or ( n34768 , n34758 , n34766 , n34767 );
and ( n34769 , n33575 , n30716 );
and ( n34770 , n32302 , n31066 );
and ( n34771 , n34769 , n34770 );
and ( n34772 , n31888 , n31414 );
and ( n34773 , n34770 , n34772 );
and ( n34774 , n34769 , n34772 );
or ( n34775 , n34771 , n34773 , n34774 );
and ( n34776 , n34480 , n30583 );
and ( n34777 , n32868 , n30950 );
and ( n34778 , n34776 , n34777 );
and ( n34779 , n32019 , n31278 );
and ( n34780 , n34777 , n34779 );
and ( n34781 , n34776 , n34779 );
or ( n34782 , n34778 , n34780 , n34781 );
and ( n34783 , n34775 , n34782 );
and ( n34784 , n33204 , n30748 );
and ( n34785 , n32940 , n30863 );
and ( n34786 , n34784 , n34785 );
and ( n34787 , n32235 , n31168 );
and ( n34788 , n34785 , n34787 );
and ( n34789 , n34784 , n34787 );
or ( n34790 , n34786 , n34788 , n34789 );
and ( n34791 , n34782 , n34790 );
and ( n34792 , n34775 , n34790 );
or ( n34793 , n34783 , n34791 , n34792 );
and ( n34794 , n34768 , n34793 );
xor ( n34795 , n34454 , n34455 );
xor ( n34796 , n34795 , n34457 );
xor ( n34797 , n34461 , n34462 );
xor ( n34798 , n34797 , n34464 );
or ( n34799 , n34796 , n34798 );
xor ( n34800 , n34481 , n34482 );
xor ( n34801 , n34800 , n34484 );
xor ( n34802 , n34488 , n34489 );
xor ( n34803 , n34802 , n34491 );
or ( n34804 , n34801 , n34803 );
and ( n34805 , n34799 , n34804 );
and ( n34806 , n34794 , n34805 );
xor ( n34807 , n34511 , n34513 );
xor ( n34808 , n34807 , n34516 );
xor ( n34809 , n34521 , n34523 );
xor ( n34810 , n34809 , n34526 );
and ( n34811 , n34808 , n34810 );
and ( n34812 , n34805 , n34811 );
and ( n34813 , n34794 , n34811 );
or ( n34814 , n34806 , n34812 , n34813 );
and ( n34815 , n34742 , n34814 );
and ( n34816 , n34735 , n34814 );
or ( n34817 , n34743 , n34815 , n34816 );
and ( n34818 , n34727 , n34817 );
and ( n34819 , n34667 , n34817 );
or ( n34820 , n34728 , n34818 , n34819 );
xnor ( n34821 , n34537 , n34538 );
xnor ( n34822 , n34546 , n34547 );
and ( n34823 , n34821 , n34822 );
xnor ( n34824 , n34557 , n34559 );
xnor ( n34825 , n34567 , n34569 );
and ( n34826 , n34824 , n34825 );
and ( n34827 , n34823 , n34826 );
xor ( n34828 , n34707 , n34708 );
and ( n34829 , n31430 , n31766 );
and ( n34830 , n31783 , n31453 );
and ( n34831 , n34829 , n34830 );
buf ( n562106 , n543230 );
buf ( n34833 , n562106 );
and ( n34834 , n34831 , n34833 );
and ( n34835 , n34828 , n34834 );
and ( n34836 , n34315 , n30598 );
and ( n34837 , n34049 , n30620 );
or ( n34838 , n34836 , n34837 );
and ( n34839 , n30601 , n34298 );
and ( n34840 , n30623 , n34032 );
or ( n34841 , n34839 , n34840 );
and ( n34842 , n34838 , n34841 );
and ( n34843 , n34834 , n34842 );
and ( n34844 , n34828 , n34842 );
or ( n34845 , n34835 , n34843 , n34844 );
and ( n34846 , n34826 , n34845 );
and ( n34847 , n34823 , n34845 );
or ( n34848 , n34827 , n34846 , n34847 );
xor ( n34849 , n34435 , n34437 );
xor ( n34850 , n34849 , n34439 );
and ( n34851 , n34848 , n34850 );
xor ( n34852 , n34449 , n34450 );
xor ( n34853 , n34852 , n34506 );
and ( n34854 , n34850 , n34853 );
and ( n34855 , n34848 , n34853 );
or ( n34856 , n34851 , n34854 , n34855 );
xor ( n34857 , n34411 , n34412 );
xor ( n34858 , n34857 , n34414 );
and ( n34859 , n34856 , n34858 );
xor ( n34860 , n34418 , n34419 );
xor ( n34861 , n34860 , n34421 );
and ( n34862 , n34858 , n34861 );
and ( n34863 , n34856 , n34861 );
or ( n34864 , n34859 , n34862 , n34863 );
and ( n34865 , n34820 , n34864 );
xor ( n34866 , n34428 , n34431 );
xor ( n34867 , n34866 , n34442 );
xor ( n34868 , n34509 , n34574 );
xor ( n34869 , n34868 , n34592 );
and ( n34870 , n34867 , n34869 );
xor ( n34871 , n34597 , n34599 );
xor ( n34872 , n34871 , n34602 );
and ( n34873 , n34869 , n34872 );
and ( n34874 , n34867 , n34872 );
or ( n34875 , n34870 , n34873 , n34874 );
and ( n34876 , n34864 , n34875 );
and ( n34877 , n34820 , n34875 );
or ( n34878 , n34865 , n34876 , n34877 );
xor ( n34879 , n34399 , n34401 );
xor ( n34880 , n34879 , n34403 );
xor ( n34881 , n34417 , n34424 );
xor ( n34882 , n34881 , n34445 );
and ( n34883 , n34880 , n34882 );
xor ( n34884 , n34595 , n34605 );
xor ( n34885 , n34884 , n34608 );
and ( n34886 , n34882 , n34885 );
and ( n34887 , n34880 , n34885 );
or ( n34888 , n34883 , n34886 , n34887 );
and ( n34889 , n34878 , n34888 );
xor ( n34890 , n34394 , n34396 );
xor ( n34891 , n34890 , n34406 );
and ( n34892 , n34888 , n34891 );
and ( n34893 , n34878 , n34891 );
or ( n34894 , n34889 , n34892 , n34893 );
and ( n34895 , n34651 , n34894 );
and ( n34896 , n34649 , n34894 );
or ( n34897 , n34652 , n34895 , n34896 );
and ( n34898 , n34647 , n34897 );
xor ( n34899 , n34389 , n34391 );
xor ( n34900 , n34899 , n34639 );
and ( n34901 , n34897 , n34900 );
and ( n34902 , n34647 , n34900 );
or ( n34903 , n34898 , n34901 , n34902 );
and ( n34904 , n34644 , n34903 );
and ( n34905 , n34642 , n34903 );
or ( n34906 , n34645 , n34904 , n34905 );
and ( n34907 , n34386 , n34906 );
and ( n34908 , n34384 , n34906 );
or ( n34909 , n34387 , n34907 , n34908 );
and ( n34910 , n34110 , n34909 );
and ( n34911 , n34108 , n34909 );
or ( n34912 , n34111 , n34910 , n34911 );
or ( n34913 , n33880 , n34912 );
or ( n34914 , n33878 , n34913 );
and ( n34915 , n33875 , n34914 );
and ( n34916 , n33447 , n34914 );
or ( n34917 , n33876 , n34915 , n34916 );
and ( n34918 , n33444 , n34917 );
and ( n34919 , n33442 , n34917 );
or ( n34920 , n33445 , n34918 , n34919 );
and ( n34921 , n33185 , n34920 );
and ( n34922 , n32823 , n34920 );
or ( n34923 , n33186 , n34921 , n34922 );
and ( n34924 , n32820 , n34923 );
and ( n34925 , n32818 , n34923 );
or ( n34926 , n32821 , n34924 , n34925 );
and ( n34927 , n32639 , n34926 );
and ( n34928 , n32637 , n34926 );
or ( n34929 , n32640 , n34927 , n34928 );
and ( n34930 , n32437 , n34929 );
and ( n34931 , n32141 , n34929 );
or ( n34932 , n32438 , n34930 , n34931 );
and ( n34933 , n32139 , n34932 );
xor ( n34934 , n32139 , n34932 );
xor ( n34935 , n32141 , n32437 );
xor ( n34936 , n34935 , n34929 );
not ( n34937 , n34936 );
xor ( n34938 , n32637 , n32639 );
xor ( n34939 , n34938 , n34926 );
xor ( n34940 , n32818 , n32820 );
xor ( n34941 , n34940 , n34923 );
xor ( n34942 , n32823 , n33185 );
xor ( n34943 , n34942 , n34920 );
not ( n34944 , n34943 );
xor ( n34945 , n33442 , n33444 );
xor ( n34946 , n34945 , n34917 );
not ( n34947 , n34946 );
xor ( n34948 , n33447 , n33875 );
xor ( n34949 , n34948 , n34914 );
xnor ( n34950 , n33878 , n34913 );
xnor ( n34951 , n33880 , n34912 );
xor ( n34952 , n34108 , n34110 );
xor ( n34953 , n34952 , n34909 );
not ( n34954 , n34953 );
xor ( n34955 , n34384 , n34386 );
xor ( n34956 , n34955 , n34906 );
xor ( n34957 , n34642 , n34644 );
xor ( n34958 , n34957 , n34903 );
xor ( n34959 , n34409 , n34625 );
xor ( n34960 , n34959 , n34636 );
xor ( n34961 , n34448 , n34611 );
xor ( n34962 , n34961 , n34622 );
xor ( n34963 , n34628 , n34630 );
xor ( n34964 , n34963 , n34633 );
and ( n34965 , n34962 , n34964 );
xor ( n34966 , n34614 , n34616 );
xor ( n34967 , n34966 , n34619 );
xor ( n34968 , n34530 , n34549 );
xor ( n34969 , n34968 , n34571 );
xor ( n34970 , n34580 , n34585 );
xor ( n34971 , n34970 , n34589 );
and ( n34972 , n34969 , n34971 );
xor ( n34973 , n34654 , n34655 );
xor ( n34974 , n34973 , n34657 );
xor ( n34975 , n34686 , n34704 );
and ( n34976 , n34974 , n34975 );
and ( n34977 , n34049 , n30632 );
and ( n34978 , n33894 , n30685 );
and ( n34979 , n34977 , n34978 );
and ( n34980 , n32302 , n31168 );
and ( n34981 , n34978 , n34980 );
and ( n34982 , n34977 , n34980 );
or ( n34983 , n34979 , n34981 , n34982 );
and ( n34984 , n33204 , n30863 );
and ( n34985 , n32940 , n30950 );
and ( n34986 , n34984 , n34985 );
and ( n34987 , n32019 , n31414 );
and ( n34988 , n34985 , n34987 );
and ( n34989 , n34984 , n34987 );
or ( n34990 , n34986 , n34988 , n34989 );
and ( n34991 , n34983 , n34990 );
and ( n34992 , n33513 , n30716 );
and ( n34993 , n33575 , n30748 );
and ( n34994 , n34992 , n34993 );
and ( n34995 , n32235 , n31278 );
and ( n34996 , n34993 , n34995 );
and ( n34997 , n34992 , n34995 );
or ( n34998 , n34994 , n34996 , n34997 );
and ( n34999 , n34990 , n34998 );
and ( n35000 , n34983 , n34998 );
or ( n35001 , n34991 , n34999 , n35000 );
xor ( n35002 , n34469 , n34470 );
xor ( n35003 , n35002 , n34472 );
or ( n35004 , n35001 , n35003 );
and ( n35005 , n30627 , n34032 );
and ( n35006 , n30680 , n33914 );
and ( n35007 , n35005 , n35006 );
and ( n35008 , n31171 , n32320 );
and ( n35009 , n35006 , n35008 );
and ( n35010 , n35005 , n35008 );
or ( n35011 , n35007 , n35009 , n35010 );
and ( n35012 , n30872 , n33213 );
and ( n35013 , n30958 , n32922 );
and ( n35014 , n35012 , n35013 );
and ( n35015 , n31405 , n31997 );
and ( n35016 , n35013 , n35015 );
and ( n35017 , n35012 , n35015 );
or ( n35018 , n35014 , n35016 , n35017 );
and ( n35019 , n35011 , n35018 );
and ( n35020 , n30711 , n33556 );
and ( n35021 , n30759 , n33532 );
and ( n35022 , n35020 , n35021 );
and ( n35023 , n31269 , n32244 );
and ( n35024 , n35021 , n35023 );
and ( n35025 , n35020 , n35023 );
or ( n35026 , n35022 , n35024 , n35025 );
and ( n35027 , n35018 , n35026 );
and ( n35028 , n35011 , n35026 );
or ( n35029 , n35019 , n35027 , n35028 );
xor ( n35030 , n34496 , n34497 );
xor ( n35031 , n35030 , n34499 );
or ( n35032 , n35029 , n35031 );
and ( n35033 , n35004 , n35032 );
and ( n35034 , n34975 , n35033 );
and ( n35035 , n34974 , n35033 );
or ( n35036 , n34976 , n35034 , n35035 );
and ( n35037 , n34971 , n35036 );
and ( n35038 , n34969 , n35036 );
or ( n35039 , n34972 , n35037 , n35038 );
xor ( n35040 , n34675 , n34677 );
xor ( n35041 , n35040 , n34680 );
not ( n35042 , n35041 );
xnor ( n35043 , n34801 , n34803 );
and ( n35044 , n35042 , n35043 );
xor ( n35045 , n34693 , n34695 );
xor ( n35046 , n35045 , n34698 );
not ( n35047 , n35046 );
xnor ( n35048 , n34796 , n34798 );
and ( n35049 , n35047 , n35048 );
and ( n35050 , n35044 , n35049 );
buf ( n35051 , n35041 );
buf ( n35052 , n35046 );
and ( n35053 , n35051 , n35052 );
and ( n35054 , n35050 , n35053 );
xnor ( n35055 , n34683 , n34685 );
xnor ( n35056 , n34701 , n34703 );
and ( n35057 , n35055 , n35056 );
and ( n35058 , n35053 , n35057 );
and ( n35059 , n35050 , n35057 );
or ( n35060 , n35054 , n35058 , n35059 );
xor ( n35061 , n34710 , n34712 );
xor ( n35062 , n35061 , n34716 );
xor ( n35063 , n34768 , n34793 );
and ( n35064 , n35062 , n35063 );
xor ( n35065 , n34799 , n34804 );
and ( n35066 , n35063 , n35065 );
and ( n35067 , n35062 , n35065 );
or ( n35068 , n35064 , n35066 , n35067 );
xor ( n35069 , n34808 , n34810 );
xor ( n35070 , n34821 , n34822 );
and ( n35071 , n35069 , n35070 );
xor ( n35072 , n34824 , n34825 );
and ( n35073 , n35070 , n35072 );
and ( n35074 , n35069 , n35072 );
or ( n35075 , n35071 , n35073 , n35074 );
and ( n35076 , n35068 , n35075 );
xor ( n35077 , n34744 , n34745 );
xor ( n35078 , n35077 , n34747 );
xor ( n35079 , n34751 , n34752 );
xor ( n35080 , n35079 , n34754 );
or ( n35081 , n35078 , n35080 );
xor ( n35082 , n34769 , n34770 );
xor ( n35083 , n35082 , n34772 );
xor ( n35084 , n34776 , n34777 );
xor ( n35085 , n35084 , n34779 );
or ( n35086 , n35083 , n35085 );
and ( n35087 , n35081 , n35086 );
xor ( n35088 , n34759 , n34760 );
xor ( n35089 , n35088 , n34762 );
xor ( n35090 , n34687 , n34688 );
xor ( n35091 , n35090 , n34690 );
or ( n35092 , n35089 , n35091 );
xor ( n35093 , n34784 , n34785 );
xor ( n35094 , n35093 , n34787 );
xor ( n35095 , n34669 , n34670 );
xor ( n35096 , n35095 , n34672 );
or ( n35097 , n35094 , n35096 );
and ( n35098 , n35092 , n35097 );
and ( n35099 , n35087 , n35098 );
and ( n35100 , n31057 , n32508 );
and ( n35101 , n31430 , n31871 );
and ( n35102 , n35100 , n35101 );
and ( n35103 , n31619 , n31766 );
and ( n35104 , n35101 , n35103 );
and ( n35105 , n35100 , n35103 );
or ( n35106 , n35102 , n35104 , n35105 );
not ( n35107 , n35106 );
and ( n35108 , n30601 , n34453 );
and ( n35109 , n30623 , n34298 );
and ( n35110 , n35108 , n35109 );
and ( n35111 , n30962 , n32850 );
and ( n35112 , n35109 , n35111 );
and ( n35113 , n35108 , n35111 );
or ( n35114 , n35110 , n35112 , n35113 );
and ( n35115 , n35107 , n35114 );
and ( n35116 , n32525 , n31066 );
and ( n35117 , n31888 , n31453 );
and ( n35118 , n35116 , n35117 );
and ( n35119 , n31783 , n31597 );
and ( n35120 , n35117 , n35119 );
and ( n35121 , n35116 , n35119 );
or ( n35122 , n35118 , n35120 , n35121 );
not ( n35123 , n35122 );
and ( n35124 , n34480 , n30598 );
and ( n35125 , n34315 , n30620 );
and ( n35126 , n35124 , n35125 );
and ( n35127 , n32868 , n30947 );
and ( n35128 , n35125 , n35127 );
and ( n35129 , n35124 , n35127 );
or ( n35130 , n35126 , n35128 , n35129 );
and ( n35131 , n35123 , n35130 );
and ( n35132 , n35115 , n35131 );
and ( n35133 , n35098 , n35132 );
and ( n35134 , n35087 , n35132 );
or ( n35135 , n35099 , n35133 , n35134 );
and ( n35136 , n35075 , n35135 );
and ( n35137 , n35068 , n35135 );
or ( n35138 , n35076 , n35136 , n35137 );
and ( n35139 , n35060 , n35138 );
buf ( n35140 , n35106 );
buf ( n35141 , n35122 );
and ( n35142 , n35140 , n35141 );
xor ( n35143 , n34750 , n34757 );
xor ( n35144 , n35143 , n34765 );
xor ( n35145 , n34775 , n34782 );
xor ( n35146 , n35145 , n34790 );
and ( n35147 , n35144 , n35146 );
and ( n35148 , n35142 , n35147 );
xor ( n35149 , n34714 , n34715 );
buf ( n35150 , n31619 );
buf ( n562425 , n543233 );
buf ( n35152 , n562425 );
or ( n35153 , n35150 , n35152 );
and ( n35154 , n35149 , n35153 );
xor ( n35155 , n34831 , n34833 );
and ( n35156 , n35153 , n35155 );
and ( n35157 , n35149 , n35155 );
or ( n35158 , n35154 , n35156 , n35157 );
and ( n35159 , n35147 , n35158 );
and ( n35160 , n35142 , n35158 );
or ( n35161 , n35148 , n35159 , n35160 );
xor ( n35162 , n34709 , n34719 );
xor ( n35163 , n35162 , n34721 );
and ( n35164 , n35161 , n35163 );
xor ( n35165 , n34729 , n34730 );
xor ( n35166 , n35165 , n34732 );
and ( n35167 , n35163 , n35166 );
and ( n35168 , n35161 , n35166 );
or ( n35169 , n35164 , n35167 , n35168 );
and ( n35170 , n35138 , n35169 );
and ( n35171 , n35060 , n35169 );
or ( n35172 , n35139 , n35170 , n35171 );
and ( n35173 , n35039 , n35172 );
xor ( n35174 , n34736 , n34737 );
xor ( n35175 , n35174 , n34739 );
xor ( n35176 , n34794 , n34805 );
xor ( n35177 , n35176 , n34811 );
and ( n35178 , n35175 , n35177 );
xor ( n35179 , n34823 , n34826 );
xor ( n35180 , n35179 , n34845 );
and ( n35181 , n35177 , n35180 );
and ( n35182 , n35175 , n35180 );
or ( n35183 , n35178 , n35181 , n35182 );
xor ( n35184 , n34660 , n34662 );
xor ( n35185 , n35184 , n34664 );
and ( n35186 , n35183 , n35185 );
xor ( n35187 , n34668 , n34705 );
xor ( n35188 , n35187 , n34724 );
and ( n35189 , n35185 , n35188 );
and ( n35190 , n35183 , n35188 );
or ( n35191 , n35186 , n35189 , n35190 );
and ( n35192 , n35172 , n35191 );
and ( n35193 , n35039 , n35191 );
or ( n35194 , n35173 , n35192 , n35193 );
and ( n35195 , n34967 , n35194 );
xor ( n35196 , n34667 , n34727 );
xor ( n35197 , n35196 , n34817 );
xor ( n35198 , n34856 , n34858 );
xor ( n35199 , n35198 , n34861 );
and ( n35200 , n35197 , n35199 );
xor ( n35201 , n34867 , n34869 );
xor ( n35202 , n35201 , n34872 );
and ( n35203 , n35199 , n35202 );
and ( n35204 , n35197 , n35202 );
or ( n35205 , n35200 , n35203 , n35204 );
and ( n35206 , n35194 , n35205 );
and ( n35207 , n34967 , n35205 );
or ( n35208 , n35195 , n35206 , n35207 );
and ( n35209 , n34964 , n35208 );
and ( n35210 , n34962 , n35208 );
or ( n35211 , n34965 , n35209 , n35210 );
and ( n35212 , n34960 , n35211 );
xor ( n35213 , n34649 , n34651 );
xor ( n35214 , n35213 , n34894 );
and ( n35215 , n35211 , n35214 );
and ( n35216 , n34960 , n35214 );
or ( n35217 , n35212 , n35215 , n35216 );
xor ( n35218 , n34647 , n34897 );
xor ( n35219 , n35218 , n34900 );
and ( n35220 , n35217 , n35219 );
xor ( n35221 , n34878 , n34888 );
xor ( n35222 , n35221 , n34891 );
xor ( n35223 , n34820 , n34864 );
xor ( n35224 , n35223 , n34875 );
xor ( n35225 , n34880 , n34882 );
xor ( n35226 , n35225 , n34885 );
and ( n35227 , n35224 , n35226 );
xor ( n35228 , n34735 , n34742 );
xor ( n35229 , n35228 , n34814 );
xor ( n35230 , n34848 , n34850 );
xor ( n35231 , n35230 , n34853 );
and ( n35232 , n35229 , n35231 );
xor ( n35233 , n34828 , n34834 );
xor ( n35234 , n35233 , n34842 );
xor ( n35235 , n35004 , n35032 );
and ( n35236 , n35234 , n35235 );
xor ( n35237 , n35044 , n35049 );
and ( n35238 , n35235 , n35237 );
and ( n35239 , n35234 , n35237 );
or ( n35240 , n35236 , n35238 , n35239 );
xor ( n35241 , n35051 , n35052 );
xor ( n35242 , n35055 , n35056 );
and ( n35243 , n35241 , n35242 );
xnor ( n35244 , n34839 , n34840 );
xnor ( n35245 , n35094 , n35096 );
or ( n35246 , n35244 , n35245 );
xnor ( n35247 , n34836 , n34837 );
xnor ( n35248 , n35089 , n35091 );
or ( n35249 , n35247 , n35248 );
and ( n35250 , n35246 , n35249 );
and ( n35251 , n35242 , n35250 );
and ( n35252 , n35241 , n35250 );
or ( n35253 , n35243 , n35251 , n35252 );
and ( n35254 , n35240 , n35253 );
and ( n35255 , n34315 , n30632 );
and ( n35256 , n34049 , n30685 );
and ( n35257 , n35255 , n35256 );
and ( n35258 , n32868 , n31066 );
and ( n35259 , n35256 , n35258 );
and ( n35260 , n35255 , n35258 );
or ( n35261 , n35257 , n35259 , n35260 );
and ( n35262 , n33513 , n30748 );
and ( n35263 , n33575 , n30863 );
and ( n35264 , n35262 , n35263 );
and ( n35265 , n32302 , n31278 );
and ( n35266 , n35263 , n35265 );
and ( n35267 , n35262 , n35265 );
or ( n35268 , n35264 , n35266 , n35267 );
and ( n35269 , n35261 , n35268 );
and ( n35270 , n33894 , n30716 );
and ( n35271 , n32525 , n31168 );
and ( n35272 , n35270 , n35271 );
and ( n35273 , n32019 , n31453 );
and ( n35274 , n35271 , n35273 );
and ( n35275 , n35270 , n35273 );
or ( n35276 , n35272 , n35274 , n35275 );
and ( n35277 , n35268 , n35276 );
and ( n35278 , n35261 , n35276 );
or ( n35279 , n35269 , n35277 , n35278 );
xor ( n35280 , n34983 , n34990 );
xor ( n35281 , n35280 , n34998 );
and ( n35282 , n35279 , n35281 );
and ( n35283 , n30627 , n34298 );
and ( n35284 , n30680 , n34032 );
and ( n35285 , n35283 , n35284 );
and ( n35286 , n31057 , n32850 );
and ( n35287 , n35284 , n35286 );
and ( n35288 , n35283 , n35286 );
or ( n35289 , n35285 , n35287 , n35288 );
and ( n35290 , n30759 , n33556 );
and ( n35291 , n30872 , n33532 );
and ( n35292 , n35290 , n35291 );
and ( n35293 , n31269 , n32320 );
and ( n35294 , n35291 , n35293 );
and ( n35295 , n35290 , n35293 );
or ( n35296 , n35292 , n35294 , n35295 );
and ( n35297 , n35289 , n35296 );
and ( n35298 , n30711 , n33914 );
and ( n35299 , n31171 , n32508 );
and ( n35300 , n35298 , n35299 );
and ( n35301 , n31430 , n31997 );
and ( n35302 , n35299 , n35301 );
and ( n35303 , n35298 , n35301 );
or ( n35304 , n35300 , n35302 , n35303 );
and ( n35305 , n35296 , n35304 );
and ( n35306 , n35289 , n35304 );
or ( n35307 , n35297 , n35305 , n35306 );
xor ( n35308 , n35011 , n35018 );
xor ( n35309 , n35308 , n35026 );
and ( n35310 , n35307 , n35309 );
and ( n35311 , n35282 , n35310 );
xnor ( n35312 , n35001 , n35003 );
xnor ( n35313 , n35029 , n35031 );
and ( n35314 , n35312 , n35313 );
and ( n35315 , n35311 , n35314 );
xor ( n35316 , n35042 , n35043 );
xor ( n35317 , n35047 , n35048 );
and ( n35318 , n35316 , n35317 );
and ( n35319 , n35314 , n35318 );
and ( n35320 , n35311 , n35318 );
or ( n35321 , n35315 , n35319 , n35320 );
and ( n35322 , n35253 , n35321 );
and ( n35323 , n35240 , n35321 );
or ( n35324 , n35254 , n35322 , n35323 );
and ( n35325 , n35231 , n35324 );
and ( n35326 , n35229 , n35324 );
or ( n35327 , n35232 , n35325 , n35326 );
xor ( n35328 , n34838 , n34841 );
xor ( n35329 , n35081 , n35086 );
and ( n35330 , n35328 , n35329 );
xor ( n35331 , n35092 , n35097 );
and ( n35332 , n35329 , n35331 );
and ( n35333 , n35328 , n35331 );
or ( n35334 , n35330 , n35332 , n35333 );
xor ( n35335 , n35115 , n35131 );
xor ( n35336 , n35140 , n35141 );
and ( n35337 , n35335 , n35336 );
xor ( n35338 , n35144 , n35146 );
and ( n35339 , n35336 , n35338 );
and ( n35340 , n35335 , n35338 );
or ( n35341 , n35337 , n35339 , n35340 );
and ( n35342 , n35334 , n35341 );
xor ( n35343 , n34977 , n34978 );
xor ( n35344 , n35343 , n34980 );
xor ( n35345 , n35116 , n35117 );
xor ( n35346 , n35345 , n35119 );
and ( n35347 , n35344 , n35346 );
xor ( n35348 , n35124 , n35125 );
xor ( n35349 , n35348 , n35127 );
and ( n35350 , n35346 , n35349 );
and ( n35351 , n35344 , n35349 );
or ( n35352 , n35347 , n35350 , n35351 );
xor ( n35353 , n35005 , n35006 );
xor ( n35354 , n35353 , n35008 );
xor ( n35355 , n35100 , n35101 );
xor ( n35356 , n35355 , n35103 );
and ( n35357 , n35354 , n35356 );
xor ( n35358 , n35108 , n35109 );
xor ( n35359 , n35358 , n35111 );
and ( n35360 , n35356 , n35359 );
and ( n35361 , n35354 , n35359 );
or ( n35362 , n35357 , n35360 , n35361 );
and ( n35363 , n35352 , n35362 );
xor ( n35364 , n35012 , n35013 );
xor ( n35365 , n35364 , n35015 );
xor ( n35366 , n35020 , n35021 );
xor ( n35367 , n35366 , n35023 );
or ( n35368 , n35365 , n35367 );
xor ( n35369 , n34984 , n34985 );
xor ( n35370 , n35369 , n34987 );
xor ( n35371 , n34992 , n34993 );
xor ( n35372 , n35371 , n34995 );
or ( n35373 , n35370 , n35372 );
and ( n35374 , n35368 , n35373 );
and ( n35375 , n35363 , n35374 );
xnor ( n35376 , n35078 , n35080 );
xnor ( n35377 , n35083 , n35085 );
and ( n35378 , n35376 , n35377 );
and ( n35379 , n35374 , n35378 );
and ( n35380 , n35363 , n35378 );
or ( n35381 , n35375 , n35379 , n35380 );
and ( n35382 , n35341 , n35381 );
and ( n35383 , n35334 , n35381 );
or ( n35384 , n35342 , n35382 , n35383 );
xor ( n35385 , n35107 , n35114 );
xor ( n35386 , n35123 , n35130 );
and ( n35387 , n35385 , n35386 );
xnor ( n35388 , n35150 , n35152 );
xor ( n35389 , n34829 , n34830 );
and ( n35390 , n35388 , n35389 );
and ( n35391 , n33204 , n30950 );
and ( n35392 , n32940 , n30947 );
and ( n35393 , n35391 , n35392 );
and ( n35394 , n32235 , n31414 );
and ( n35395 , n35392 , n35394 );
and ( n35396 , n35391 , n35394 );
or ( n35397 , n35393 , n35395 , n35396 );
and ( n35398 , n30958 , n33213 );
and ( n35399 , n30962 , n32922 );
and ( n35400 , n35398 , n35399 );
and ( n35401 , n31405 , n32244 );
and ( n35402 , n35399 , n35401 );
and ( n35403 , n35398 , n35401 );
or ( n35404 , n35400 , n35402 , n35403 );
and ( n35405 , n35397 , n35404 );
and ( n35406 , n35389 , n35405 );
and ( n35407 , n35388 , n35405 );
or ( n35408 , n35390 , n35406 , n35407 );
and ( n35409 , n35387 , n35408 );
xor ( n35410 , n35149 , n35153 );
xor ( n35411 , n35410 , n35155 );
and ( n35412 , n35408 , n35411 );
and ( n35413 , n35387 , n35411 );
or ( n35414 , n35409 , n35412 , n35413 );
xor ( n35415 , n35062 , n35063 );
xor ( n35416 , n35415 , n35065 );
and ( n35417 , n35414 , n35416 );
xor ( n35418 , n35069 , n35070 );
xor ( n35419 , n35418 , n35072 );
and ( n35420 , n35416 , n35419 );
and ( n35421 , n35414 , n35419 );
or ( n35422 , n35417 , n35420 , n35421 );
and ( n35423 , n35384 , n35422 );
xor ( n35424 , n34974 , n34975 );
xor ( n35425 , n35424 , n35033 );
and ( n35426 , n35422 , n35425 );
and ( n35427 , n35384 , n35425 );
or ( n35428 , n35423 , n35426 , n35427 );
xor ( n35429 , n35050 , n35053 );
xor ( n35430 , n35429 , n35057 );
xor ( n35431 , n35068 , n35075 );
xor ( n35432 , n35431 , n35135 );
and ( n35433 , n35430 , n35432 );
xor ( n35434 , n35161 , n35163 );
xor ( n35435 , n35434 , n35166 );
and ( n35436 , n35432 , n35435 );
and ( n35437 , n35430 , n35435 );
or ( n35438 , n35433 , n35436 , n35437 );
and ( n35439 , n35428 , n35438 );
xor ( n35440 , n34969 , n34971 );
xor ( n35441 , n35440 , n35036 );
and ( n35442 , n35438 , n35441 );
and ( n35443 , n35428 , n35441 );
or ( n35444 , n35439 , n35442 , n35443 );
and ( n35445 , n35327 , n35444 );
xor ( n35446 , n35039 , n35172 );
xor ( n35447 , n35446 , n35191 );
and ( n35448 , n35444 , n35447 );
and ( n35449 , n35327 , n35447 );
or ( n35450 , n35445 , n35448 , n35449 );
and ( n35451 , n35226 , n35450 );
and ( n35452 , n35224 , n35450 );
or ( n35453 , n35227 , n35451 , n35452 );
and ( n35454 , n35222 , n35453 );
xor ( n35455 , n34962 , n34964 );
xor ( n35456 , n35455 , n35208 );
and ( n35457 , n35453 , n35456 );
and ( n35458 , n35222 , n35456 );
or ( n35459 , n35454 , n35457 , n35458 );
xor ( n35460 , n34960 , n35211 );
xor ( n35461 , n35460 , n35214 );
and ( n35462 , n35459 , n35461 );
xor ( n35463 , n34967 , n35194 );
xor ( n35464 , n35463 , n35205 );
xor ( n35465 , n35197 , n35199 );
xor ( n35466 , n35465 , n35202 );
xor ( n35467 , n35060 , n35138 );
xor ( n35468 , n35467 , n35169 );
xor ( n35469 , n35183 , n35185 );
xor ( n35470 , n35469 , n35188 );
and ( n35471 , n35468 , n35470 );
xor ( n35472 , n35175 , n35177 );
xor ( n35473 , n35472 , n35180 );
xor ( n35474 , n35087 , n35098 );
xor ( n35475 , n35474 , n35132 );
xor ( n35476 , n35142 , n35147 );
xor ( n35477 , n35476 , n35158 );
and ( n35478 , n35475 , n35477 );
xor ( n35479 , n35246 , n35249 );
xor ( n35480 , n35282 , n35310 );
and ( n35481 , n35479 , n35480 );
xor ( n35482 , n35312 , n35313 );
and ( n35483 , n35480 , n35482 );
and ( n35484 , n35479 , n35482 );
or ( n35485 , n35481 , n35483 , n35484 );
and ( n35486 , n35477 , n35485 );
and ( n35487 , n35475 , n35485 );
or ( n35488 , n35478 , n35486 , n35487 );
and ( n35489 , n35473 , n35488 );
xor ( n35490 , n35316 , n35317 );
and ( n35491 , n33575 , n30950 );
and ( n35492 , n33204 , n30947 );
and ( n35493 , n35491 , n35492 );
and ( n35494 , n32302 , n31414 );
and ( n35495 , n35492 , n35494 );
and ( n35496 , n35491 , n35494 );
or ( n35497 , n35493 , n35495 , n35496 );
and ( n35498 , n34480 , n30632 );
and ( n35499 , n32940 , n31066 );
and ( n35500 , n35498 , n35499 );
and ( n35501 , n32235 , n31453 );
and ( n35502 , n35499 , n35501 );
and ( n35503 , n35498 , n35501 );
or ( n35504 , n35500 , n35502 , n35503 );
and ( n35505 , n35497 , n35504 );
and ( n35506 , n32868 , n31168 );
and ( n35507 , n32019 , n31597 );
and ( n35508 , n35506 , n35507 );
and ( n35509 , n31888 , n31766 );
and ( n35510 , n35507 , n35509 );
and ( n35511 , n35506 , n35509 );
or ( n35512 , n35508 , n35510 , n35511 );
and ( n35513 , n35504 , n35512 );
and ( n35514 , n35497 , n35512 );
or ( n35515 , n35505 , n35513 , n35514 );
xor ( n35516 , n35261 , n35268 );
xor ( n35517 , n35516 , n35276 );
or ( n35518 , n35515 , n35517 );
and ( n35519 , n30958 , n33532 );
and ( n35520 , n30962 , n33213 );
and ( n35521 , n35519 , n35520 );
and ( n35522 , n31405 , n32320 );
and ( n35523 , n35520 , n35522 );
and ( n35524 , n35519 , n35522 );
or ( n35525 , n35521 , n35523 , n35524 );
and ( n35526 , n30627 , n34453 );
and ( n35527 , n31057 , n32922 );
and ( n35528 , n35526 , n35527 );
and ( n35529 , n31430 , n32244 );
and ( n35530 , n35527 , n35529 );
and ( n35531 , n35526 , n35529 );
or ( n35532 , n35528 , n35530 , n35531 );
and ( n35533 , n35525 , n35532 );
and ( n35534 , n31171 , n32850 );
and ( n35535 , n31619 , n31997 );
and ( n35536 , n35534 , n35535 );
and ( n35537 , n31783 , n31871 );
and ( n35538 , n35535 , n35537 );
and ( n35539 , n35534 , n35537 );
or ( n35540 , n35536 , n35538 , n35539 );
and ( n35541 , n35532 , n35540 );
and ( n35542 , n35525 , n35540 );
or ( n35543 , n35533 , n35541 , n35542 );
xor ( n35544 , n35289 , n35296 );
xor ( n35545 , n35544 , n35304 );
or ( n35546 , n35543 , n35545 );
and ( n35547 , n35518 , n35546 );
and ( n35548 , n35490 , n35547 );
xnor ( n35549 , n35244 , n35245 );
xnor ( n35550 , n35247 , n35248 );
and ( n35551 , n35549 , n35550 );
and ( n35552 , n35547 , n35551 );
and ( n35553 , n35490 , n35551 );
or ( n35554 , n35548 , n35552 , n35553 );
xor ( n35555 , n35279 , n35281 );
xor ( n35556 , n35307 , n35309 );
and ( n35557 , n35555 , n35556 );
buf ( n562832 , n543236 );
buf ( n35559 , n562832 );
buf ( n35560 , n31783 );
buf ( n562835 , n543239 );
buf ( n35562 , n562835 );
or ( n35563 , n35560 , n35562 );
and ( n35564 , n35559 , n35563 );
and ( n35565 , n30623 , n34453 );
and ( n35566 , n34480 , n30620 );
and ( n35567 , n35565 , n35566 );
and ( n35568 , n35563 , n35567 );
and ( n35569 , n35559 , n35567 );
or ( n35570 , n35564 , n35568 , n35569 );
xor ( n35571 , n35352 , n35362 );
and ( n35572 , n35570 , n35571 );
xor ( n35573 , n35368 , n35373 );
and ( n35574 , n35571 , n35573 );
and ( n35575 , n35570 , n35573 );
or ( n35576 , n35572 , n35574 , n35575 );
and ( n35577 , n35557 , n35576 );
xor ( n35578 , n35376 , n35377 );
xor ( n35579 , n35385 , n35386 );
and ( n35580 , n35578 , n35579 );
and ( n35581 , n30759 , n33914 );
and ( n35582 , n30872 , n33556 );
and ( n35583 , n35581 , n35582 );
and ( n35584 , n31269 , n32508 );
and ( n35585 , n35582 , n35584 );
and ( n35586 , n35581 , n35584 );
or ( n35587 , n35583 , n35585 , n35586 );
xor ( n35588 , n35391 , n35392 );
xor ( n35589 , n35588 , n35394 );
and ( n35590 , n35587 , n35589 );
xor ( n35591 , n35255 , n35256 );
xor ( n35592 , n35591 , n35258 );
and ( n35593 , n35589 , n35592 );
and ( n35594 , n35587 , n35592 );
or ( n35595 , n35590 , n35593 , n35594 );
and ( n35596 , n33894 , n30748 );
and ( n35597 , n33513 , n30863 );
and ( n35598 , n35596 , n35597 );
and ( n35599 , n32525 , n31278 );
and ( n35600 , n35597 , n35599 );
and ( n35601 , n35596 , n35599 );
or ( n35602 , n35598 , n35600 , n35601 );
xor ( n35603 , n35398 , n35399 );
xor ( n35604 , n35603 , n35401 );
and ( n35605 , n35602 , n35604 );
xor ( n35606 , n35283 , n35284 );
xor ( n35607 , n35606 , n35286 );
and ( n35608 , n35604 , n35607 );
and ( n35609 , n35602 , n35607 );
or ( n35610 , n35605 , n35608 , n35609 );
and ( n35611 , n35595 , n35610 );
and ( n35612 , n35579 , n35611 );
and ( n35613 , n35578 , n35611 );
or ( n35614 , n35580 , n35612 , n35613 );
and ( n35615 , n35576 , n35614 );
and ( n35616 , n35557 , n35614 );
or ( n35617 , n35577 , n35615 , n35616 );
and ( n35618 , n35554 , n35617 );
xor ( n35619 , n35290 , n35291 );
xor ( n35620 , n35619 , n35293 );
xor ( n35621 , n35298 , n35299 );
xor ( n35622 , n35621 , n35301 );
or ( n35623 , n35620 , n35622 );
xor ( n35624 , n35262 , n35263 );
xor ( n35625 , n35624 , n35265 );
xor ( n35626 , n35270 , n35271 );
xor ( n35627 , n35626 , n35273 );
or ( n35628 , n35625 , n35627 );
and ( n35629 , n35623 , n35628 );
xor ( n35630 , n35344 , n35346 );
xor ( n35631 , n35630 , n35349 );
xor ( n35632 , n35354 , n35356 );
xor ( n35633 , n35632 , n35359 );
and ( n35634 , n35631 , n35633 );
and ( n35635 , n35629 , n35634 );
xnor ( n35636 , n35365 , n35367 );
xnor ( n35637 , n35370 , n35372 );
and ( n35638 , n35636 , n35637 );
and ( n35639 , n35634 , n35638 );
and ( n35640 , n35629 , n35638 );
or ( n35641 , n35635 , n35639 , n35640 );
xor ( n35642 , n35328 , n35329 );
xor ( n35643 , n35642 , n35331 );
and ( n35644 , n35641 , n35643 );
xor ( n35645 , n35335 , n35336 );
xor ( n35646 , n35645 , n35338 );
and ( n35647 , n35643 , n35646 );
and ( n35648 , n35641 , n35646 );
or ( n35649 , n35644 , n35647 , n35648 );
and ( n35650 , n35617 , n35649 );
and ( n35651 , n35554 , n35649 );
or ( n35652 , n35618 , n35650 , n35651 );
and ( n35653 , n35488 , n35652 );
and ( n35654 , n35473 , n35652 );
or ( n35655 , n35489 , n35653 , n35654 );
and ( n35656 , n35470 , n35655 );
and ( n35657 , n35468 , n35655 );
or ( n35658 , n35471 , n35656 , n35657 );
and ( n35659 , n35466 , n35658 );
xor ( n35660 , n35234 , n35235 );
xor ( n35661 , n35660 , n35237 );
xor ( n35662 , n35241 , n35242 );
xor ( n35663 , n35662 , n35250 );
and ( n35664 , n35661 , n35663 );
xor ( n35665 , n35311 , n35314 );
xor ( n35666 , n35665 , n35318 );
and ( n35667 , n35663 , n35666 );
and ( n35668 , n35661 , n35666 );
or ( n35669 , n35664 , n35667 , n35668 );
xor ( n35670 , n35240 , n35253 );
xor ( n35671 , n35670 , n35321 );
and ( n35672 , n35669 , n35671 );
xor ( n35673 , n35384 , n35422 );
xor ( n35674 , n35673 , n35425 );
and ( n35675 , n35671 , n35674 );
and ( n35676 , n35669 , n35674 );
or ( n35677 , n35672 , n35675 , n35676 );
xor ( n35678 , n35229 , n35231 );
xor ( n35679 , n35678 , n35324 );
and ( n35680 , n35677 , n35679 );
xor ( n35681 , n35428 , n35438 );
xor ( n35682 , n35681 , n35441 );
and ( n35683 , n35679 , n35682 );
and ( n35684 , n35677 , n35682 );
or ( n35685 , n35680 , n35683 , n35684 );
and ( n35686 , n35658 , n35685 );
and ( n35687 , n35466 , n35685 );
or ( n35688 , n35659 , n35686 , n35687 );
and ( n35689 , n35464 , n35688 );
xor ( n35690 , n35224 , n35226 );
xor ( n35691 , n35690 , n35450 );
and ( n35692 , n35688 , n35691 );
and ( n35693 , n35464 , n35691 );
or ( n35694 , n35689 , n35692 , n35693 );
xor ( n35695 , n35222 , n35453 );
xor ( n35696 , n35695 , n35456 );
and ( n35697 , n35694 , n35696 );
xor ( n35698 , n35327 , n35444 );
xor ( n35699 , n35698 , n35447 );
xor ( n35700 , n35430 , n35432 );
xor ( n35701 , n35700 , n35435 );
xor ( n35702 , n35334 , n35341 );
xor ( n35703 , n35702 , n35381 );
xor ( n35704 , n35414 , n35416 );
xor ( n35705 , n35704 , n35419 );
and ( n35706 , n35703 , n35705 );
xor ( n35707 , n35363 , n35374 );
xor ( n35708 , n35707 , n35378 );
xor ( n35709 , n35387 , n35408 );
xor ( n35710 , n35709 , n35411 );
and ( n35711 , n35708 , n35710 );
and ( n35712 , n31619 , n31871 );
and ( n35713 , n31888 , n31597 );
and ( n35714 , n35712 , n35713 );
xor ( n35715 , n35397 , n35404 );
and ( n35716 , n35714 , n35715 );
and ( n35717 , n34315 , n30685 );
and ( n35718 , n34049 , n30716 );
or ( n35719 , n35717 , n35718 );
and ( n35720 , n30680 , n34298 );
and ( n35721 , n30711 , n34032 );
or ( n35722 , n35720 , n35721 );
and ( n35723 , n35719 , n35722 );
and ( n35724 , n35715 , n35723 );
and ( n35725 , n35714 , n35723 );
or ( n35726 , n35716 , n35724 , n35725 );
xor ( n35727 , n35388 , n35389 );
xor ( n35728 , n35727 , n35405 );
and ( n35729 , n35726 , n35728 );
xor ( n35730 , n35518 , n35546 );
and ( n35731 , n35728 , n35730 );
and ( n35732 , n35726 , n35730 );
or ( n35733 , n35729 , n35731 , n35732 );
and ( n35734 , n35710 , n35733 );
and ( n35735 , n35708 , n35733 );
or ( n35736 , n35711 , n35734 , n35735 );
and ( n35737 , n35705 , n35736 );
and ( n35738 , n35703 , n35736 );
or ( n35739 , n35706 , n35737 , n35738 );
and ( n35740 , n35701 , n35739 );
xor ( n35741 , n35549 , n35550 );
xor ( n35742 , n35555 , n35556 );
and ( n35743 , n35741 , n35742 );
xnor ( n35744 , n35515 , n35517 );
xnor ( n35745 , n35543 , n35545 );
and ( n35746 , n35744 , n35745 );
and ( n35747 , n35742 , n35746 );
and ( n35748 , n35741 , n35746 );
or ( n35749 , n35743 , n35747 , n35748 );
xnor ( n35750 , n35560 , n35562 );
xor ( n35751 , n35565 , n35566 );
and ( n35752 , n35750 , n35751 );
xor ( n35753 , n35712 , n35713 );
and ( n35754 , n35751 , n35753 );
and ( n35755 , n35750 , n35753 );
or ( n35756 , n35752 , n35754 , n35755 );
xor ( n35757 , n35559 , n35563 );
xor ( n35758 , n35757 , n35567 );
and ( n35759 , n35756 , n35758 );
xor ( n35760 , n35595 , n35610 );
and ( n35761 , n35758 , n35760 );
and ( n35762 , n35756 , n35760 );
or ( n35763 , n35759 , n35761 , n35762 );
xor ( n35764 , n35623 , n35628 );
xor ( n35765 , n35631 , n35633 );
and ( n35766 , n35764 , n35765 );
xor ( n35767 , n35636 , n35637 );
and ( n35768 , n35765 , n35767 );
and ( n35769 , n35764 , n35767 );
or ( n35770 , n35766 , n35768 , n35769 );
and ( n35771 , n35763 , n35770 );
xor ( n35772 , n35596 , n35597 );
xor ( n35773 , n35772 , n35599 );
xor ( n35774 , n35491 , n35492 );
xor ( n35775 , n35774 , n35494 );
and ( n35776 , n35773 , n35775 );
xor ( n35777 , n35498 , n35499 );
xor ( n35778 , n35777 , n35501 );
and ( n35779 , n35775 , n35778 );
and ( n35780 , n35773 , n35778 );
or ( n35781 , n35776 , n35779 , n35780 );
xor ( n35782 , n35581 , n35582 );
xor ( n35783 , n35782 , n35584 );
xor ( n35784 , n35519 , n35520 );
xor ( n35785 , n35784 , n35522 );
and ( n35786 , n35783 , n35785 );
xor ( n35787 , n35526 , n35527 );
xor ( n35788 , n35787 , n35529 );
and ( n35789 , n35785 , n35788 );
and ( n35790 , n35783 , n35788 );
or ( n35791 , n35786 , n35789 , n35790 );
and ( n35792 , n35781 , n35791 );
and ( n35793 , n30680 , n34453 );
and ( n35794 , n30711 , n34298 );
and ( n35795 , n35793 , n35794 );
and ( n35796 , n31171 , n32922 );
and ( n35797 , n35794 , n35796 );
and ( n35798 , n35793 , n35796 );
or ( n35799 , n35795 , n35797 , n35798 );
and ( n35800 , n30759 , n34032 );
and ( n35801 , n31269 , n32850 );
and ( n35802 , n35800 , n35801 );
and ( n35803 , n31619 , n32244 );
and ( n35804 , n35801 , n35803 );
and ( n35805 , n35800 , n35803 );
or ( n35806 , n35802 , n35804 , n35805 );
or ( n35807 , n35799 , n35806 );
and ( n35808 , n34480 , n30685 );
and ( n35809 , n34315 , n30716 );
and ( n35810 , n35808 , n35809 );
and ( n35811 , n32940 , n31168 );
and ( n35812 , n35809 , n35811 );
and ( n35813 , n35808 , n35811 );
or ( n35814 , n35810 , n35812 , n35813 );
and ( n35815 , n34049 , n30748 );
and ( n35816 , n32868 , n31278 );
and ( n35817 , n35815 , n35816 );
and ( n35818 , n32235 , n31597 );
and ( n35819 , n35816 , n35818 );
and ( n35820 , n35815 , n35818 );
or ( n35821 , n35817 , n35819 , n35820 );
or ( n35822 , n35814 , n35821 );
and ( n35823 , n35807 , n35822 );
and ( n35824 , n35792 , n35823 );
and ( n563099 , n30962 , n33532 );
and ( n35825 , n31057 , n33213 );
and ( n35826 , n563099 , n35825 );
and ( n35827 , n31430 , n32320 );
and ( n35828 , n35825 , n35827 );
and ( n35829 , n563099 , n35827 );
or ( n35830 , n35826 , n35828 , n35829 );
not ( n35831 , n35830 );
and ( n35832 , n30872 , n33914 );
and ( n35833 , n30958 , n33556 );
and ( n35834 , n35832 , n35833 );
and ( n35835 , n31405 , n32508 );
and ( n35836 , n35833 , n35835 );
and ( n35837 , n35832 , n35835 );
or ( n35838 , n35834 , n35836 , n35837 );
and ( n35839 , n35831 , n35838 );
and ( n35840 , n33575 , n30947 );
and ( n35841 , n33204 , n31066 );
and ( n35842 , n35840 , n35841 );
and ( n35843 , n32302 , n31453 );
and ( n35844 , n35841 , n35843 );
and ( n35845 , n35840 , n35843 );
or ( n35846 , n35842 , n35844 , n35845 );
not ( n35847 , n35846 );
and ( n35848 , n33894 , n30863 );
and ( n35849 , n33513 , n30950 );
and ( n35850 , n35848 , n35849 );
and ( n35851 , n32525 , n31414 );
and ( n35852 , n35849 , n35851 );
and ( n35853 , n35848 , n35851 );
or ( n35854 , n35850 , n35852 , n35853 );
and ( n35855 , n35847 , n35854 );
and ( n35856 , n35839 , n35855 );
and ( n35857 , n35823 , n35856 );
and ( n35858 , n35792 , n35856 );
or ( n35859 , n35824 , n35857 , n35858 );
and ( n35860 , n35770 , n35859 );
and ( n35861 , n35763 , n35859 );
or ( n35862 , n35771 , n35860 , n35861 );
and ( n35863 , n35749 , n35862 );
buf ( n35864 , n35830 );
buf ( n35865 , n35846 );
and ( n35866 , n35864 , n35865 );
xor ( n35867 , n35525 , n35532 );
xor ( n35868 , n35867 , n35540 );
xor ( n35869 , n35497 , n35504 );
xor ( n35870 , n35869 , n35512 );
and ( n35871 , n35868 , n35870 );
and ( n35872 , n35866 , n35871 );
xor ( n35873 , n35587 , n35589 );
xor ( n35874 , n35873 , n35592 );
xor ( n35875 , n35602 , n35604 );
xor ( n35876 , n35875 , n35607 );
and ( n35877 , n35874 , n35876 );
and ( n35878 , n35871 , n35877 );
and ( n35879 , n35866 , n35877 );
or ( n35880 , n35872 , n35878 , n35879 );
xnor ( n35881 , n35620 , n35622 );
xnor ( n35882 , n35625 , n35627 );
and ( n35883 , n35881 , n35882 );
xor ( n35884 , n35719 , n35722 );
and ( n35885 , n31783 , n31997 );
and ( n35886 , n32019 , n31766 );
and ( n35887 , n35885 , n35886 );
buf ( n563163 , n543242 );
buf ( n35889 , n563163 );
and ( n35890 , n35887 , n35889 );
and ( n35891 , n35884 , n35890 );
xnor ( n35892 , n35717 , n35718 );
xnor ( n35893 , n35720 , n35721 );
and ( n35894 , n35892 , n35893 );
and ( n35895 , n35890 , n35894 );
and ( n35896 , n35884 , n35894 );
or ( n35897 , n35891 , n35895 , n35896 );
and ( n35898 , n35883 , n35897 );
xor ( n35899 , n35714 , n35715 );
xor ( n35900 , n35899 , n35723 );
and ( n35901 , n35897 , n35900 );
and ( n35902 , n35883 , n35900 );
or ( n35903 , n35898 , n35901 , n35902 );
and ( n35904 , n35880 , n35903 );
xor ( n35905 , n35570 , n35571 );
xor ( n35906 , n35905 , n35573 );
and ( n35907 , n35903 , n35906 );
and ( n35908 , n35880 , n35906 );
or ( n35909 , n35904 , n35907 , n35908 );
and ( n35910 , n35862 , n35909 );
and ( n35911 , n35749 , n35909 );
or ( n35912 , n35863 , n35910 , n35911 );
xor ( n35913 , n35479 , n35480 );
xor ( n35914 , n35913 , n35482 );
xor ( n35915 , n35490 , n35547 );
xor ( n35916 , n35915 , n35551 );
and ( n35917 , n35914 , n35916 );
xor ( n35918 , n35557 , n35576 );
xor ( n35919 , n35918 , n35614 );
and ( n35920 , n35916 , n35919 );
and ( n35921 , n35914 , n35919 );
or ( n35922 , n35917 , n35920 , n35921 );
and ( n35923 , n35912 , n35922 );
xor ( n35924 , n35475 , n35477 );
xor ( n35925 , n35924 , n35485 );
and ( n35926 , n35922 , n35925 );
and ( n35927 , n35912 , n35925 );
or ( n35928 , n35923 , n35926 , n35927 );
and ( n35929 , n35739 , n35928 );
and ( n35930 , n35701 , n35928 );
or ( n35931 , n35740 , n35929 , n35930 );
xor ( n35932 , n35468 , n35470 );
xor ( n35933 , n35932 , n35655 );
and ( n35934 , n35931 , n35933 );
xor ( n35935 , n35677 , n35679 );
xor ( n35936 , n35935 , n35682 );
and ( n35937 , n35933 , n35936 );
and ( n35938 , n35931 , n35936 );
or ( n35939 , n35934 , n35937 , n35938 );
and ( n35940 , n35699 , n35939 );
xor ( n35941 , n35466 , n35658 );
xor ( n35942 , n35941 , n35685 );
and ( n35943 , n35939 , n35942 );
and ( n35944 , n35699 , n35942 );
or ( n35945 , n35940 , n35943 , n35944 );
xor ( n35946 , n35464 , n35688 );
xor ( n35947 , n35946 , n35691 );
and ( n35948 , n35945 , n35947 );
xor ( n35949 , n35699 , n35939 );
xor ( n35950 , n35949 , n35942 );
xor ( n35951 , n35473 , n35488 );
xor ( n35952 , n35951 , n35652 );
xor ( n35953 , n35669 , n35671 );
xor ( n35954 , n35953 , n35674 );
and ( n35955 , n35952 , n35954 );
xor ( n35956 , n35554 , n35617 );
xor ( n35957 , n35956 , n35649 );
xor ( n35958 , n35661 , n35663 );
xor ( n35959 , n35958 , n35666 );
and ( n35960 , n35957 , n35959 );
xor ( n35961 , n35641 , n35643 );
xor ( n35962 , n35961 , n35646 );
xor ( n35963 , n35578 , n35579 );
xor ( n35964 , n35963 , n35611 );
xor ( n35965 , n35629 , n35634 );
xor ( n35966 , n35965 , n35638 );
and ( n35967 , n35964 , n35966 );
xor ( n35968 , n35744 , n35745 );
and ( n35969 , n33894 , n30950 );
and ( n35970 , n33513 , n30947 );
and ( n563246 , n35969 , n35970 );
and ( n35971 , n32525 , n31453 );
and ( n35972 , n35970 , n35971 );
and ( n35973 , n35969 , n35971 );
or ( n35974 , n563246 , n35972 , n35973 );
and ( n35975 , n34315 , n30748 );
and ( n35976 , n34049 , n30863 );
and ( n35977 , n35975 , n35976 );
and ( n35978 , n32868 , n31414 );
and ( n35979 , n35976 , n35978 );
and ( n35980 , n35975 , n35978 );
or ( n35981 , n35977 , n35979 , n35980 );
and ( n35982 , n35974 , n35981 );
and ( n35983 , n33575 , n31066 );
and ( n35984 , n33204 , n31168 );
and ( n35985 , n35983 , n35984 );
and ( n35986 , n32302 , n31597 );
and ( n35987 , n35984 , n35986 );
and ( n35988 , n35983 , n35986 );
or ( n35989 , n35985 , n35987 , n35988 );
and ( n35990 , n35981 , n35989 );
and ( n35991 , n35974 , n35989 );
or ( n35992 , n35982 , n35990 , n35991 );
xor ( n35993 , n35534 , n35535 );
xor ( n35994 , n35993 , n35537 );
or ( n35995 , n35992 , n35994 );
and ( n35996 , n30958 , n33914 );
and ( n35997 , n30962 , n33556 );
and ( n35998 , n35996 , n35997 );
and ( n35999 , n31430 , n32508 );
and ( n36000 , n35997 , n35999 );
and ( n36001 , n35996 , n35999 );
or ( n36002 , n35998 , n36000 , n36001 );
and ( n36003 , n30759 , n34298 );
and ( n36004 , n30872 , n34032 );
and ( n36005 , n36003 , n36004 );
and ( n36006 , n31405 , n32850 );
and ( n36007 , n36004 , n36006 );
and ( n36008 , n36003 , n36006 );
or ( n36009 , n36005 , n36007 , n36008 );
and ( n36010 , n36002 , n36009 );
and ( n36011 , n31057 , n33532 );
and ( n36012 , n31171 , n33213 );
and ( n36013 , n36011 , n36012 );
and ( n36014 , n31619 , n32320 );
and ( n36015 , n36012 , n36014 );
and ( n36016 , n36011 , n36014 );
or ( n36017 , n36013 , n36015 , n36016 );
and ( n36018 , n36009 , n36017 );
and ( n36019 , n36002 , n36017 );
or ( n36020 , n36010 , n36018 , n36019 );
xor ( n36021 , n35506 , n35507 );
xor ( n36022 , n36021 , n35509 );
or ( n36023 , n36020 , n36022 );
and ( n36024 , n35995 , n36023 );
and ( n36025 , n35968 , n36024 );
xor ( n36026 , n35750 , n35751 );
xor ( n36027 , n36026 , n35753 );
xor ( n36028 , n35781 , n35791 );
and ( n36029 , n36027 , n36028 );
xor ( n36030 , n35807 , n35822 );
and ( n36031 , n36028 , n36030 );
and ( n36032 , n36027 , n36030 );
or ( n36033 , n36029 , n36031 , n36032 );
and ( n36034 , n36024 , n36033 );
and ( n36035 , n35968 , n36033 );
or ( n36036 , n36025 , n36034 , n36035 );
and ( n36037 , n35966 , n36036 );
and ( n36038 , n35964 , n36036 );
or ( n563315 , n35967 , n36037 , n36038 );
and ( n36039 , n35962 , n563315 );
xor ( n36040 , n35839 , n35855 );
xor ( n36041 , n35864 , n35865 );
and ( n36042 , n36040 , n36041 );
xor ( n36043 , n35868 , n35870 );
and ( n36044 , n36041 , n36043 );
and ( n36045 , n36040 , n36043 );
or ( n36046 , n36042 , n36044 , n36045 );
xor ( n36047 , n35874 , n35876 );
xor ( n36048 , n35881 , n35882 );
and ( n36049 , n36047 , n36048 );
xor ( n36050 , n35887 , n35889 );
buf ( n36051 , n31888 );
buf ( n563329 , n543245 );
buf ( n36053 , n563329 );
and ( n36054 , n36051 , n36053 );
and ( n36055 , n36050 , n36054 );
and ( n36056 , n32940 , n31278 );
and ( n36057 , n32235 , n31766 );
and ( n36058 , n36056 , n36057 );
and ( n36059 , n32019 , n31871 );
and ( n36060 , n36057 , n36059 );
and ( n36061 , n36056 , n36059 );
or ( n36062 , n36058 , n36060 , n36061 );
and ( n36063 , n31269 , n32922 );
and ( n36064 , n31783 , n32244 );
and ( n36065 , n36063 , n36064 );
and ( n36066 , n31888 , n31997 );
and ( n36067 , n36064 , n36066 );
and ( n36068 , n36063 , n36066 );
or ( n36069 , n36065 , n36067 , n36068 );
and ( n36070 , n36062 , n36069 );
and ( n36071 , n36054 , n36070 );
and ( n36072 , n36050 , n36070 );
or ( n36073 , n36055 , n36071 , n36072 );
and ( n36074 , n36048 , n36073 );
and ( n36075 , n36047 , n36073 );
or ( n36076 , n36049 , n36074 , n36075 );
and ( n36077 , n36046 , n36076 );
xor ( n36078 , n35808 , n35809 );
xor ( n36079 , n36078 , n35811 );
xor ( n36080 , n35815 , n35816 );
xor ( n36081 , n36080 , n35818 );
and ( n36082 , n36079 , n36081 );
xor ( n36083 , n35840 , n35841 );
xor ( n36084 , n36083 , n35843 );
and ( n36085 , n36081 , n36084 );
and ( n36086 , n36079 , n36084 );
or ( n36087 , n36082 , n36085 , n36086 );
xor ( n36088 , n35793 , n35794 );
xor ( n36089 , n36088 , n35796 );
xor ( n36090 , n35800 , n35801 );
xor ( n36091 , n36090 , n35803 );
and ( n36092 , n36089 , n36091 );
xor ( n36093 , n563099 , n35825 );
xor ( n36094 , n36093 , n35827 );
and ( n36095 , n36091 , n36094 );
and ( n36096 , n36089 , n36094 );
or ( n36097 , n36092 , n36095 , n36096 );
and ( n36098 , n36087 , n36097 );
xor ( n36099 , n35773 , n35775 );
xor ( n36100 , n36099 , n35778 );
xor ( n36101 , n35783 , n35785 );
xor ( n36102 , n36101 , n35788 );
and ( n36103 , n36100 , n36102 );
and ( n36104 , n36098 , n36103 );
xnor ( n36105 , n35799 , n35806 );
xnor ( n36106 , n35814 , n35821 );
and ( n36107 , n36105 , n36106 );
and ( n36108 , n36103 , n36107 );
and ( n36109 , n36098 , n36107 );
or ( n36110 , n36104 , n36108 , n36109 );
and ( n36111 , n36076 , n36110 );
and ( n36112 , n36046 , n36110 );
or ( n36113 , n36077 , n36111 , n36112 );
xor ( n36114 , n35756 , n35758 );
xor ( n36115 , n36114 , n35760 );
xor ( n36116 , n35764 , n35765 );
xor ( n36117 , n36116 , n35767 );
and ( n36118 , n36115 , n36117 );
xor ( n36119 , n35792 , n35823 );
xor ( n36120 , n36119 , n35856 );
and ( n36121 , n36117 , n36120 );
and ( n36122 , n36115 , n36120 );
or ( n36123 , n36118 , n36121 , n36122 );
and ( n36124 , n36113 , n36123 );
xor ( n36125 , n35726 , n35728 );
xor ( n36126 , n36125 , n35730 );
and ( n36127 , n36123 , n36126 );
and ( n36128 , n36113 , n36126 );
or ( n36129 , n36124 , n36127 , n36128 );
and ( n36130 , n563315 , n36129 );
and ( n36131 , n35962 , n36129 );
or ( n36132 , n36039 , n36130 , n36131 );
and ( n36133 , n35959 , n36132 );
and ( n36134 , n35957 , n36132 );
or ( n36135 , n35960 , n36133 , n36134 );
and ( n36136 , n35954 , n36135 );
and ( n36137 , n35952 , n36135 );
or ( n36138 , n35955 , n36136 , n36137 );
xor ( n36139 , n35931 , n35933 );
xor ( n36140 , n36139 , n35936 );
and ( n36141 , n36138 , n36140 );
xor ( n36142 , n35741 , n35742 );
xor ( n36143 , n36142 , n35746 );
xor ( n36144 , n35763 , n35770 );
xor ( n36145 , n36144 , n35859 );
and ( n36146 , n36143 , n36145 );
xor ( n36147 , n35880 , n35903 );
xor ( n36148 , n36147 , n35906 );
and ( n36149 , n36145 , n36148 );
and ( n36150 , n36143 , n36148 );
or ( n36151 , n36146 , n36149 , n36150 );
xor ( n36152 , n35708 , n35710 );
xor ( n36153 , n36152 , n35733 );
and ( n36154 , n36151 , n36153 );
xor ( n36155 , n35749 , n35862 );
xor ( n36156 , n36155 , n35909 );
and ( n36157 , n36153 , n36156 );
and ( n36158 , n36151 , n36156 );
or ( n36159 , n36154 , n36157 , n36158 );
xor ( n36160 , n35703 , n35705 );
xor ( n36161 , n36160 , n35736 );
and ( n36162 , n36159 , n36161 );
xor ( n36163 , n35912 , n35922 );
xor ( n36164 , n36163 , n35925 );
and ( n36165 , n36161 , n36164 );
and ( n36166 , n36159 , n36164 );
or ( n36167 , n36162 , n36165 , n36166 );
xor ( n36168 , n35701 , n35739 );
xor ( n36169 , n36168 , n35928 );
and ( n36170 , n36167 , n36169 );
xor ( n36171 , n35914 , n35916 );
xor ( n36172 , n36171 , n35919 );
xor ( n36173 , n35866 , n35871 );
xor ( n36174 , n36173 , n35877 );
xor ( n36175 , n35883 , n35897 );
xor ( n36176 , n36175 , n35900 );
and ( n36177 , n36174 , n36176 );
xor ( n36178 , n35831 , n35838 );
xor ( n36179 , n35847 , n35854 );
and ( n36180 , n36178 , n36179 );
xor ( n36181 , n35884 , n35890 );
xor ( n36182 , n36181 , n35894 );
and ( n36183 , n36180 , n36182 );
xor ( n36184 , n35995 , n36023 );
and ( n36185 , n36182 , n36184 );
and ( n36186 , n36180 , n36184 );
or ( n36187 , n36183 , n36185 , n36186 );
and ( n36188 , n36176 , n36187 );
and ( n36189 , n36174 , n36187 );
or ( n36190 , n36177 , n36188 , n36189 );
xor ( n36191 , n36051 , n36053 );
and ( n36192 , n31888 , n32244 );
and ( n36193 , n32235 , n31871 );
and ( n36194 , n36192 , n36193 );
buf ( n563472 , n543248 );
buf ( n36196 , n563472 );
and ( n36197 , n36194 , n36196 );
and ( n36198 , n36191 , n36197 );
and ( n36199 , n30711 , n34453 );
and ( n36200 , n34480 , n30716 );
and ( n36201 , n36199 , n36200 );
and ( n36202 , n36197 , n36201 );
and ( n36203 , n36191 , n36201 );
or ( n36204 , n36198 , n36202 , n36203 );
xor ( n36205 , n35848 , n35849 );
xor ( n563483 , n36205 , n35851 );
xor ( n36206 , n35832 , n35833 );
xor ( n36207 , n36206 , n35835 );
and ( n36208 , n563483 , n36207 );
and ( n36209 , n36204 , n36208 );
xor ( n36210 , n36050 , n36054 );
xor ( n36211 , n36210 , n36070 );
and ( n36212 , n36208 , n36211 );
and ( n36213 , n36204 , n36211 );
or ( n36214 , n36209 , n36212 , n36213 );
and ( n36215 , n33513 , n31066 );
and ( n36216 , n33575 , n31168 );
and ( n36217 , n36215 , n36216 );
and ( n36218 , n32525 , n31597 );
and ( n36219 , n36216 , n36218 );
and ( n36220 , n36215 , n36218 );
or ( n36221 , n36217 , n36219 , n36220 );
and ( n36222 , n34049 , n30950 );
and ( n36223 , n33894 , n30947 );
and ( n36224 , n36222 , n36223 );
and ( n36225 , n32868 , n31453 );
and ( n36226 , n36223 , n36225 );
and ( n36227 , n36222 , n36225 );
or ( n36228 , n36224 , n36226 , n36227 );
and ( n36229 , n36221 , n36228 );
and ( n36230 , n34315 , n30863 );
and ( n36231 , n32940 , n31414 );
and ( n36232 , n36230 , n36231 );
and ( n36233 , n32302 , n31766 );
and ( n36234 , n36231 , n36233 );
and ( n36235 , n36230 , n36233 );
or ( n36236 , n36232 , n36234 , n36235 );
and ( n36237 , n36228 , n36236 );
and ( n36238 , n36221 , n36236 );
or ( n36239 , n36229 , n36237 , n36238 );
xor ( n36240 , n35974 , n35981 );
xor ( n36241 , n36240 , n35989 );
or ( n36242 , n36239 , n36241 );
and ( n36243 , n31057 , n33556 );
and ( n36244 , n31171 , n33532 );
and ( n36245 , n36243 , n36244 );
and ( n36246 , n31619 , n32508 );
and ( n36247 , n36244 , n36246 );
and ( n36248 , n36243 , n36246 );
or ( n36249 , n36245 , n36247 , n36248 );
and ( n36250 , n30958 , n34032 );
and ( n36251 , n30962 , n33914 );
and ( n36252 , n36250 , n36251 );
and ( n36253 , n31430 , n32850 );
and ( n36254 , n36251 , n36253 );
and ( n36255 , n36250 , n36253 );
or ( n36256 , n36252 , n36254 , n36255 );
and ( n36257 , n36249 , n36256 );
and ( n36258 , n30872 , n34298 );
and ( n36259 , n31405 , n32922 );
and ( n36260 , n36258 , n36259 );
and ( n36261 , n31783 , n32320 );
and ( n36262 , n36259 , n36261 );
and ( n36263 , n36258 , n36261 );
or ( n36264 , n36260 , n36262 , n36263 );
and ( n36265 , n36256 , n36264 );
and ( n36266 , n36249 , n36264 );
or ( n36267 , n36257 , n36265 , n36266 );
xor ( n36268 , n36002 , n36009 );
xor ( n36269 , n36268 , n36017 );
or ( n36270 , n36267 , n36269 );
and ( n36271 , n36242 , n36270 );
and ( n36272 , n36214 , n36271 );
xnor ( n36273 , n35992 , n35994 );
xnor ( n36274 , n36020 , n36022 );
and ( n36275 , n36273 , n36274 );
and ( n36276 , n36271 , n36275 );
and ( n36277 , n36214 , n36275 );
or ( n36278 , n36272 , n36276 , n36277 );
xor ( n36279 , n35892 , n35893 );
xor ( n36280 , n36087 , n36097 );
and ( n36281 , n36279 , n36280 );
xor ( n36282 , n36100 , n36102 );
and ( n36283 , n36280 , n36282 );
and ( n36284 , n36279 , n36282 );
or ( n36285 , n36281 , n36283 , n36284 );
xor ( n36286 , n36105 , n36106 );
xor ( n36287 , n36178 , n36179 );
and ( n36288 , n36286 , n36287 );
xor ( n36289 , n35996 , n35997 );
xor ( n36290 , n36289 , n35999 );
xor ( n36291 , n36003 , n36004 );
xor ( n36292 , n36291 , n36006 );
and ( n36293 , n36290 , n36292 );
xor ( n36294 , n35969 , n35970 );
xor ( n36295 , n36294 , n35971 );
xor ( n36296 , n35975 , n35976 );
xor ( n36297 , n36296 , n35978 );
and ( n36298 , n36295 , n36297 );
and ( n36299 , n36293 , n36298 );
and ( n36300 , n36287 , n36299 );
and ( n36301 , n36286 , n36299 );
or ( n36302 , n36288 , n36300 , n36301 );
and ( n36303 , n36285 , n36302 );
xor ( n36304 , n36063 , n36064 );
xor ( n36305 , n36304 , n36066 );
xor ( n36306 , n36011 , n36012 );
xor ( n36307 , n36306 , n36014 );
and ( n36308 , n36305 , n36307 );
xor ( n36309 , n36056 , n36057 );
xor ( n36310 , n36309 , n36059 );
xor ( n36311 , n35983 , n35984 );
xor ( n36312 , n36311 , n35986 );
and ( n36313 , n36310 , n36312 );
and ( n36314 , n36308 , n36313 );
xor ( n36315 , n36079 , n36081 );
xor ( n36316 , n36315 , n36084 );
xor ( n36317 , n36089 , n36091 );
xor ( n36318 , n36317 , n36094 );
and ( n36319 , n36316 , n36318 );
and ( n36320 , n36314 , n36319 );
xor ( n36321 , n35885 , n35886 );
xor ( n36322 , n36062 , n36069 );
and ( n36323 , n36321 , n36322 );
xor ( n36324 , n563483 , n36207 );
and ( n36325 , n36322 , n36324 );
and ( n36326 , n36321 , n36324 );
or ( n36327 , n36323 , n36325 , n36326 );
and ( n36328 , n36319 , n36327 );
and ( n36329 , n36314 , n36327 );
or ( n36330 , n36320 , n36328 , n36329 );
and ( n36331 , n36302 , n36330 );
and ( n36332 , n36285 , n36330 );
or ( n36333 , n36303 , n36331 , n36332 );
and ( n36334 , n36278 , n36333 );
xor ( n36335 , n36027 , n36028 );
xor ( n36336 , n36335 , n36030 );
xor ( n36337 , n36040 , n36041 );
xor ( n36338 , n36337 , n36043 );
and ( n36339 , n36336 , n36338 );
xor ( n36340 , n36047 , n36048 );
xor ( n36341 , n36340 , n36073 );
and ( n36342 , n36338 , n36341 );
and ( n36343 , n36336 , n36341 );
or ( n36344 , n36339 , n36342 , n36343 );
and ( n36345 , n36333 , n36344 );
and ( n36346 , n36278 , n36344 );
or ( n36347 , n36334 , n36345 , n36346 );
and ( n36348 , n36190 , n36347 );
xor ( n36349 , n35968 , n36024 );
xor ( n36350 , n36349 , n36033 );
xor ( n36351 , n36046 , n36076 );
xor ( n36352 , n36351 , n36110 );
and ( n36353 , n36350 , n36352 );
xor ( n36354 , n36115 , n36117 );
xor ( n36355 , n36354 , n36120 );
and ( n36356 , n36352 , n36355 );
and ( n36357 , n36350 , n36355 );
or ( n36358 , n36353 , n36356 , n36357 );
and ( n36359 , n36347 , n36358 );
and ( n36360 , n36190 , n36358 );
or ( n36361 , n36348 , n36359 , n36360 );
and ( n36362 , n36172 , n36361 );
xor ( n36363 , n35964 , n35966 );
xor ( n36364 , n36363 , n36036 );
xor ( n36365 , n36113 , n36123 );
xor ( n36366 , n36365 , n36126 );
and ( n36367 , n36364 , n36366 );
xor ( n36368 , n36143 , n36145 );
xor ( n36369 , n36368 , n36148 );
and ( n36370 , n36366 , n36369 );
and ( n36371 , n36364 , n36369 );
or ( n36372 , n36367 , n36370 , n36371 );
and ( n36373 , n36361 , n36372 );
and ( n36374 , n36172 , n36372 );
or ( n36375 , n36362 , n36373 , n36374 );
xor ( n36376 , n35957 , n35959 );
xor ( n36377 , n36376 , n36132 );
and ( n36378 , n36375 , n36377 );
xor ( n36379 , n36159 , n36161 );
xor ( n36380 , n36379 , n36164 );
and ( n36381 , n36377 , n36380 );
and ( n36382 , n36375 , n36380 );
or ( n36383 , n36378 , n36381 , n36382 );
and ( n36384 , n36169 , n36383 );
and ( n36385 , n36167 , n36383 );
or ( n36386 , n36170 , n36384 , n36385 );
and ( n36387 , n36140 , n36386 );
and ( n36388 , n36138 , n36386 );
or ( n36389 , n36141 , n36387 , n36388 );
and ( n36390 , n35950 , n36389 );
xor ( n36391 , n36138 , n36140 );
xor ( n36392 , n36391 , n36386 );
xor ( n36393 , n35952 , n35954 );
xor ( n36394 , n36393 , n36135 );
xor ( n36395 , n36167 , n36169 );
xor ( n36396 , n36395 , n36383 );
and ( n36397 , n36394 , n36396 );
xor ( n36398 , n35962 , n563315 );
xor ( n36399 , n36398 , n36129 );
xor ( n36400 , n36151 , n36153 );
xor ( n36401 , n36400 , n36156 );
and ( n36402 , n36399 , n36401 );
xor ( n36403 , n36098 , n36103 );
xor ( n36404 , n36403 , n36107 );
xor ( n36405 , n36204 , n36208 );
xor ( n36406 , n36405 , n36211 );
xor ( n36407 , n36242 , n36270 );
and ( n36408 , n36406 , n36407 );
xor ( n36409 , n36273 , n36274 );
and ( n36410 , n36407 , n36409 );
and ( n36411 , n36406 , n36409 );
or ( n36412 , n36408 , n36410 , n36411 );
and ( n36413 , n36404 , n36412 );
xor ( n36414 , n36305 , n36307 );
xor ( n36415 , n36310 , n36312 );
and ( n36416 , n36414 , n36415 );
xor ( n36417 , n36191 , n36197 );
xor ( n36418 , n36417 , n36201 );
and ( n36419 , n36416 , n36418 );
xnor ( n36420 , n36239 , n36241 );
xnor ( n36421 , n36267 , n36269 );
and ( n36422 , n36420 , n36421 );
and ( n36423 , n36419 , n36422 );
and ( n36424 , n34480 , n30748 );
and ( n36425 , n33204 , n31278 );
or ( n36426 , n36424 , n36425 );
and ( n36427 , n30759 , n34453 );
and ( n36428 , n31269 , n33213 );
or ( n36429 , n36427 , n36428 );
and ( n36430 , n36426 , n36429 );
xor ( n36431 , n36293 , n36298 );
and ( n36432 , n36430 , n36431 );
xor ( n36433 , n36308 , n36313 );
and ( n36434 , n36431 , n36433 );
and ( n36435 , n36430 , n36433 );
or ( n36436 , n36432 , n36434 , n36435 );
and ( n36437 , n36422 , n36436 );
and ( n36438 , n36419 , n36436 );
or ( n36439 , n36423 , n36437 , n36438 );
and ( n36440 , n36412 , n36439 );
and ( n36441 , n36404 , n36439 );
or ( n36442 , n36413 , n36440 , n36441 );
xor ( n36443 , n36316 , n36318 );
xor ( n36444 , n36215 , n36216 );
xor ( n36445 , n36444 , n36218 );
xor ( n36446 , n36222 , n36223 );
xor ( n36447 , n36446 , n36225 );
and ( n36448 , n36445 , n36447 );
xor ( n36449 , n36230 , n36231 );
xor ( n36450 , n36449 , n36233 );
and ( n36451 , n36447 , n36450 );
and ( n36452 , n36445 , n36450 );
or ( n36453 , n36448 , n36451 , n36452 );
xor ( n36454 , n36243 , n36244 );
xor ( n36455 , n36454 , n36246 );
xor ( n36456 , n36250 , n36251 );
xor ( n36457 , n36456 , n36253 );
and ( n36458 , n36455 , n36457 );
xor ( n36459 , n36258 , n36259 );
xor ( n36460 , n36459 , n36261 );
and ( n36461 , n36457 , n36460 );
and ( n36462 , n36455 , n36460 );
or ( n36463 , n36458 , n36461 , n36462 );
and ( n36464 , n36453 , n36463 );
and ( n36465 , n36443 , n36464 );
and ( n36466 , n31171 , n33556 );
and ( n36467 , n31269 , n33532 );
and ( n36468 , n36466 , n36467 );
and ( n563747 , n31783 , n32508 );
and ( n36469 , n36467 , n563747 );
and ( n563749 , n36466 , n563747 );
or ( n563750 , n36468 , n36469 , n563749 );
and ( n36470 , n30962 , n34032 );
and ( n36471 , n31057 , n33914 );
and ( n36472 , n36470 , n36471 );
and ( n36473 , n31619 , n32850 );
and ( n36474 , n36471 , n36473 );
and ( n36475 , n36470 , n36473 );
or ( n36476 , n36472 , n36474 , n36475 );
or ( n36477 , n563750 , n36476 );
and ( n36478 , n33513 , n31168 );
and ( n36479 , n33575 , n31278 );
and ( n36480 , n36478 , n36479 );
and ( n36481 , n32525 , n31766 );
and ( n36482 , n36479 , n36481 );
and ( n36483 , n36478 , n36481 );
or ( n36484 , n36480 , n36482 , n36483 );
and ( n36485 , n34049 , n30947 );
and ( n36486 , n33894 , n31066 );
and ( n36487 , n36485 , n36486 );
and ( n36488 , n32868 , n31597 );
and ( n36489 , n36486 , n36488 );
and ( n36490 , n36485 , n36488 );
or ( n36491 , n36487 , n36489 , n36490 );
or ( n36492 , n36484 , n36491 );
and ( n36493 , n36477 , n36492 );
and ( n36494 , n36464 , n36493 );
and ( n36495 , n36443 , n36493 );
or ( n36496 , n36465 , n36494 , n36495 );
and ( n36497 , n30872 , n34453 );
and ( n36498 , n30958 , n34298 );
and ( n36499 , n36497 , n36498 );
and ( n36500 , n31430 , n32922 );
and ( n36501 , n36498 , n36500 );
and ( n36502 , n36497 , n36500 );
or ( n36503 , n36499 , n36501 , n36502 );
and ( n36504 , n31405 , n33213 );
and ( n36505 , n31888 , n32320 );
and ( n36506 , n36504 , n36505 );
and ( n36507 , n32019 , n32244 );
and ( n36508 , n36505 , n36507 );
and ( n36509 , n36504 , n36507 );
or ( n36510 , n36506 , n36508 , n36509 );
or ( n36511 , n36503 , n36510 );
and ( n36512 , n34480 , n30863 );
and ( n36513 , n34315 , n30950 );
and ( n36514 , n36512 , n36513 );
and ( n36515 , n32940 , n31453 );
and ( n36516 , n36513 , n36515 );
and ( n36517 , n36512 , n36515 );
or ( n36518 , n36514 , n36516 , n36517 );
and ( n36519 , n33204 , n31414 );
and ( n36520 , n32302 , n31871 );
and ( n36521 , n36519 , n36520 );
and ( n36522 , n32235 , n31997 );
and ( n36523 , n36520 , n36522 );
and ( n36524 , n36519 , n36522 );
or ( n36525 , n36521 , n36523 , n36524 );
or ( n36526 , n36518 , n36525 );
and ( n36527 , n36511 , n36526 );
xor ( n36528 , n36249 , n36256 );
xor ( n36529 , n36528 , n36264 );
xor ( n36530 , n36221 , n36228 );
xor ( n36531 , n36530 , n36236 );
and ( n36532 , n36529 , n36531 );
and ( n36533 , n36527 , n36532 );
xor ( n36534 , n36290 , n36292 );
xor ( n36535 , n36295 , n36297 );
and ( n36536 , n36534 , n36535 );
and ( n36537 , n36532 , n36536 );
and ( n36538 , n36527 , n36536 );
or ( n36539 , n36533 , n36537 , n36538 );
and ( n36540 , n36496 , n36539 );
xor ( n36541 , n36279 , n36280 );
xor ( n36542 , n36541 , n36282 );
and ( n36543 , n36539 , n36542 );
and ( n36544 , n36496 , n36542 );
or ( n36545 , n36540 , n36543 , n36544 );
xor ( n36546 , n36180 , n36182 );
xor ( n36547 , n36546 , n36184 );
and ( n36548 , n36545 , n36547 );
xor ( n36549 , n36214 , n36271 );
xor ( n36550 , n36549 , n36275 );
and ( n36551 , n36547 , n36550 );
and ( n36552 , n36545 , n36550 );
or ( n36553 , n36548 , n36551 , n36552 );
and ( n36554 , n36442 , n36553 );
xor ( n36555 , n36174 , n36176 );
xor ( n36556 , n36555 , n36187 );
and ( n36557 , n36553 , n36556 );
and ( n36558 , n36442 , n36556 );
or ( n36559 , n36554 , n36557 , n36558 );
xor ( n36560 , n36190 , n36347 );
xor ( n36561 , n36560 , n36358 );
and ( n36562 , n36559 , n36561 );
xor ( n36563 , n36364 , n36366 );
xor ( n36564 , n36563 , n36369 );
and ( n36565 , n36561 , n36564 );
and ( n36566 , n36559 , n36564 );
or ( n36567 , n36562 , n36565 , n36566 );
and ( n36568 , n36401 , n36567 );
and ( n36569 , n36399 , n36567 );
or ( n36570 , n36402 , n36568 , n36569 );
xor ( n36571 , n36375 , n36377 );
xor ( n36572 , n36571 , n36380 );
and ( n36573 , n36570 , n36572 );
xor ( n36574 , n36172 , n36361 );
xor ( n36575 , n36574 , n36372 );
xor ( n36576 , n36399 , n36401 );
xor ( n36577 , n36576 , n36567 );
and ( n36578 , n36575 , n36577 );
xor ( n36579 , n36278 , n36333 );
xor ( n36580 , n36579 , n36344 );
xor ( n36581 , n36350 , n36352 );
xor ( n36582 , n36581 , n36355 );
and ( n36583 , n36580 , n36582 );
xor ( n36584 , n36285 , n36302 );
xor ( n36585 , n36584 , n36330 );
xor ( n36586 , n36336 , n36338 );
xor ( n36587 , n36586 , n36341 );
and ( n36588 , n36585 , n36587 );
xor ( n563870 , n36286 , n36287 );
xor ( n36589 , n563870 , n36299 );
xor ( n36590 , n36314 , n36319 );
xor ( n36591 , n36590 , n36327 );
and ( n36592 , n36589 , n36591 );
xor ( n36593 , n36199 , n36200 );
xor ( n36594 , n36194 , n36196 );
and ( n36595 , n36593 , n36594 );
xor ( n36596 , n36426 , n36429 );
and ( n36597 , n36594 , n36596 );
and ( n36598 , n36593 , n36596 );
or ( n36599 , n36595 , n36597 , n36598 );
xor ( n36600 , n36321 , n36322 );
xor ( n36601 , n36600 , n36324 );
and ( n36602 , n36599 , n36601 );
xor ( n36603 , n36416 , n36418 );
and ( n36604 , n36601 , n36603 );
and ( n36605 , n36599 , n36603 );
or ( n36606 , n36602 , n36604 , n36605 );
and ( n36607 , n36591 , n36606 );
and ( n36608 , n36589 , n36606 );
or ( n36609 , n36592 , n36607 , n36608 );
and ( n36610 , n36587 , n36609 );
and ( n36611 , n36585 , n36609 );
or ( n36612 , n36588 , n36610 , n36611 );
and ( n36613 , n36582 , n36612 );
and ( n36614 , n36580 , n36612 );
or ( n36615 , n36583 , n36613 , n36614 );
xor ( n36616 , n36559 , n36561 );
xor ( n36617 , n36616 , n36564 );
and ( n36618 , n36615 , n36617 );
xor ( n36619 , n36420 , n36421 );
xnor ( n36620 , n36427 , n36428 );
xnor ( n36621 , n36518 , n36525 );
or ( n36622 , n36620 , n36621 );
xnor ( n36623 , n36424 , n36425 );
xnor ( n36624 , n36503 , n36510 );
or ( n36625 , n36623 , n36624 );
and ( n36626 , n36622 , n36625 );
and ( n36627 , n36619 , n36626 );
and ( n36628 , n34480 , n30950 );
and ( n36629 , n33204 , n31453 );
and ( n36630 , n36628 , n36629 );
and ( n36631 , n32525 , n31871 );
and ( n36632 , n36629 , n36631 );
and ( n36633 , n36628 , n36631 );
or ( n36634 , n36630 , n36632 , n36633 );
and ( n36635 , n34315 , n30947 );
and ( n36636 , n34049 , n31066 );
and ( n36637 , n36635 , n36636 );
and ( n36638 , n32940 , n31597 );
and ( n36639 , n36636 , n36638 );
and ( n36640 , n36635 , n36638 );
or ( n36641 , n36637 , n36639 , n36640 );
and ( n36642 , n36634 , n36641 );
xor ( n36643 , n36497 , n36498 );
xor ( n36644 , n36643 , n36500 );
and ( n36645 , n36641 , n36644 );
and ( n36646 , n36634 , n36644 );
or ( n36647 , n36642 , n36645 , n36646 );
xor ( n36648 , n36455 , n36457 );
xor ( n36649 , n36648 , n36460 );
and ( n36650 , n36647 , n36649 );
and ( n36651 , n30958 , n34453 );
and ( n36652 , n31430 , n33213 );
and ( n36653 , n36651 , n36652 );
and ( n36654 , n31888 , n32508 );
and ( n36655 , n36652 , n36654 );
and ( n36656 , n36651 , n36654 );
or ( n36657 , n36653 , n36655 , n36656 );
and ( n36658 , n30962 , n34298 );
and ( n36659 , n31057 , n34032 );
and ( n36660 , n36658 , n36659 );
and ( n36661 , n31619 , n32922 );
and ( n36662 , n36659 , n36661 );
and ( n36663 , n36658 , n36661 );
or ( n36664 , n36660 , n36662 , n36663 );
and ( n36665 , n36657 , n36664 );
xor ( n36666 , n36512 , n36513 );
xor ( n36667 , n36666 , n36515 );
and ( n36668 , n36664 , n36667 );
and ( n36669 , n36657 , n36667 );
or ( n36670 , n36665 , n36668 , n36669 );
xor ( n36671 , n36445 , n36447 );
xor ( n36672 , n36671 , n36450 );
and ( n36673 , n36670 , n36672 );
and ( n36674 , n36650 , n36673 );
and ( n36675 , n36626 , n36674 );
and ( n36676 , n36619 , n36674 );
or ( n36677 , n36627 , n36675 , n36676 );
xor ( n36678 , n36453 , n36463 );
xor ( n36679 , n36477 , n36492 );
and ( n36680 , n36678 , n36679 );
xor ( n36681 , n36511 , n36526 );
and ( n36682 , n36679 , n36681 );
and ( n36683 , n36678 , n36681 );
or ( n36684 , n36680 , n36682 , n36683 );
xor ( n36685 , n36529 , n36531 );
xor ( n36686 , n36534 , n36535 );
and ( n36687 , n36685 , n36686 );
xor ( n36688 , n36414 , n36415 );
and ( n36689 , n36686 , n36688 );
and ( n36690 , n36685 , n36688 );
or ( n36691 , n36687 , n36689 , n36690 );
and ( n36692 , n36684 , n36691 );
xor ( n36693 , n36430 , n36431 );
xor ( n36694 , n36693 , n36433 );
and ( n36695 , n36691 , n36694 );
and ( n36696 , n36684 , n36694 );
or ( n36697 , n36692 , n36695 , n36696 );
and ( n36698 , n36677 , n36697 );
xor ( n36699 , n36406 , n36407 );
xor ( n36700 , n36699 , n36409 );
and ( n36701 , n36697 , n36700 );
and ( n36702 , n36677 , n36700 );
or ( n36703 , n36698 , n36701 , n36702 );
xor ( n36704 , n36404 , n36412 );
xor ( n36705 , n36704 , n36439 );
and ( n36706 , n36703 , n36705 );
xor ( n36707 , n36545 , n36547 );
xor ( n36708 , n36707 , n36550 );
and ( n36709 , n36705 , n36708 );
and ( n36710 , n36703 , n36708 );
or ( n36711 , n36706 , n36709 , n36710 );
xor ( n36712 , n36442 , n36553 );
xor ( n36713 , n36712 , n36556 );
and ( n36714 , n36711 , n36713 );
xor ( n36715 , n36419 , n36422 );
xor ( n36716 , n36715 , n36436 );
xor ( n36717 , n36496 , n36539 );
xor ( n36718 , n36717 , n36542 );
and ( n36719 , n36716 , n36718 );
xor ( n36720 , n36443 , n36464 );
xor ( n36721 , n36720 , n36493 );
xor ( n36722 , n36527 , n36532 );
xor ( n36723 , n36722 , n36536 );
and ( n36724 , n36721 , n36723 );
buf ( n36725 , n32019 );
buf ( n564008 , n543251 );
buf ( n36727 , n564008 );
and ( n36728 , n36725 , n36727 );
xnor ( n36729 , n36620 , n36621 );
xnor ( n36730 , n36623 , n36624 );
and ( n36731 , n36729 , n36730 );
or ( n36732 , n36728 , n36731 );
and ( n36733 , n36723 , n36732 );
and ( n36734 , n36721 , n36732 );
or ( n36735 , n36724 , n36733 , n36734 );
and ( n36736 , n36718 , n36735 );
and ( n36737 , n36716 , n36735 );
or ( n36738 , n36719 , n36736 , n36737 );
xnor ( n36739 , n563750 , n36476 );
xnor ( n36740 , n36484 , n36491 );
and ( n36741 , n36739 , n36740 );
xor ( n36742 , n36593 , n36594 );
xor ( n36743 , n36742 , n36596 );
and ( n36744 , n36741 , n36743 );
xor ( n36745 , n36622 , n36625 );
and ( n36746 , n36743 , n36745 );
and ( n36747 , n36741 , n36745 );
or ( n36748 , n36744 , n36746 , n36747 );
xor ( n36749 , n36650 , n36673 );
and ( n36750 , n32019 , n32320 );
and ( n36751 , n32302 , n31997 );
and ( n36752 , n36750 , n36751 );
buf ( n564035 , n543254 );
buf ( n36754 , n564035 );
xor ( n36755 , n36752 , n36754 );
buf ( n36756 , n32235 );
buf ( n564039 , n543257 );
buf ( n36758 , n564039 );
and ( n36759 , n36756 , n36758 );
and ( n36760 , n36755 , n36759 );
and ( n36761 , n31405 , n33532 );
and ( n36762 , n33575 , n31414 );
and ( n36763 , n36761 , n36762 );
and ( n36764 , n36759 , n36763 );
and ( n36765 , n36755 , n36763 );
or ( n36766 , n36760 , n36764 , n36765 );
and ( n36767 , n31269 , n33914 );
and ( n36768 , n31405 , n33556 );
and ( n36769 , n36767 , n36768 );
and ( n36770 , n31888 , n32850 );
and ( n36771 , n36768 , n36770 );
and ( n36772 , n36767 , n36770 );
or ( n36773 , n36769 , n36771 , n36772 );
and ( n36774 , n31057 , n34298 );
and ( n36775 , n31171 , n34032 );
and ( n36776 , n36774 , n36775 );
and ( n36777 , n31783 , n32922 );
and ( n36778 , n36775 , n36777 );
and ( n36779 , n36774 , n36777 );
or ( n36780 , n36776 , n36778 , n36779 );
and ( n36781 , n36773 , n36780 );
and ( n36782 , n31430 , n33532 );
and ( n36783 , n32019 , n32508 );
and ( n36784 , n36782 , n36783 );
and ( n36785 , n32235 , n32320 );
and ( n36786 , n36783 , n36785 );
and ( n36787 , n36782 , n36785 );
or ( n36788 , n36784 , n36786 , n36787 );
and ( n36789 , n36780 , n36788 );
and ( n36790 , n36773 , n36788 );
or ( n36791 , n36781 , n36789 , n36790 );
and ( n36792 , n33894 , n31278 );
and ( n36793 , n33513 , n31414 );
and ( n36794 , n36792 , n36793 );
and ( n36795 , n32868 , n31871 );
and ( n36796 , n36793 , n36795 );
and ( n36797 , n36792 , n36795 );
or ( n36798 , n36794 , n36796 , n36797 );
and ( n36799 , n34315 , n31066 );
and ( n36800 , n34049 , n31168 );
and ( n36801 , n36799 , n36800 );
and ( n36802 , n32940 , n31766 );
and ( n36803 , n36800 , n36802 );
and ( n36804 , n36799 , n36802 );
or ( n36805 , n36801 , n36803 , n36804 );
and ( n36806 , n36798 , n36805 );
and ( n36807 , n33575 , n31453 );
and ( n36808 , n32525 , n31997 );
and ( n36809 , n36807 , n36808 );
and ( n36810 , n32302 , n32244 );
and ( n36811 , n36808 , n36810 );
and ( n36812 , n36807 , n36810 );
or ( n36813 , n36809 , n36811 , n36812 );
and ( n36814 , n36805 , n36813 );
and ( n36815 , n36798 , n36813 );
or ( n36816 , n36806 , n36814 , n36815 );
and ( n36817 , n36791 , n36816 );
and ( n36818 , n36766 , n36817 );
xor ( n36819 , n36725 , n36727 );
and ( n36820 , n36752 , n36754 );
xor ( n36821 , n36819 , n36820 );
and ( n36822 , n33894 , n31168 );
and ( n36823 , n33513 , n31278 );
and ( n36824 , n36822 , n36823 );
and ( n36825 , n32868 , n31766 );
and ( n36826 , n36823 , n36825 );
and ( n36827 , n36822 , n36825 );
or ( n36828 , n36824 , n36826 , n36827 );
and ( n36829 , n31171 , n33914 );
and ( n36830 , n31269 , n33556 );
and ( n36831 , n36829 , n36830 );
and ( n36832 , n31783 , n32850 );
and ( n36833 , n36830 , n36832 );
and ( n36834 , n36829 , n36832 );
or ( n36835 , n36831 , n36833 , n36834 );
and ( n36836 , n36828 , n36835 );
xor ( n36837 , n36821 , n36836 );
and ( n36838 , n36817 , n36837 );
and ( n36839 , n36766 , n36837 );
or ( n36840 , n36818 , n36838 , n36839 );
and ( n36841 , n36749 , n36840 );
xor ( n36842 , n36634 , n36641 );
xor ( n36843 , n36842 , n36644 );
xor ( n36844 , n36466 , n36467 );
xor ( n36845 , n36844 , n563747 );
xor ( n36846 , n36470 , n36471 );
xor ( n36847 , n36846 , n36473 );
xor ( n36848 , n36845 , n36847 );
xor ( n36849 , n36504 , n36505 );
xor ( n36850 , n36849 , n36507 );
xor ( n36851 , n36848 , n36850 );
and ( n36852 , n36843 , n36851 );
xor ( n36853 , n36657 , n36664 );
xor ( n36854 , n36853 , n36667 );
xor ( n36855 , n36478 , n36479 );
xor ( n36856 , n36855 , n36481 );
xor ( n36857 , n36485 , n36486 );
xor ( n36858 , n36857 , n36488 );
xor ( n36859 , n36856 , n36858 );
xor ( n36860 , n36519 , n36520 );
xor ( n36861 , n36860 , n36522 );
xor ( n36862 , n36859 , n36861 );
and ( n36863 , n36854 , n36862 );
and ( n36864 , n36852 , n36863 );
and ( n36865 , n36840 , n36864 );
and ( n36866 , n36749 , n36864 );
or ( n36867 , n36841 , n36865 , n36866 );
and ( n36868 , n36748 , n36867 );
xor ( n36869 , n36647 , n36649 );
xor ( n36870 , n36670 , n36672 );
and ( n36871 , n36869 , n36870 );
xor ( n36872 , n36192 , n36193 );
and ( n36873 , n36856 , n36858 );
and ( n36874 , n36858 , n36861 );
and ( n36875 , n36856 , n36861 );
or ( n36876 , n36873 , n36874 , n36875 );
and ( n36877 , n36845 , n36847 );
and ( n36878 , n36847 , n36850 );
and ( n36879 , n36845 , n36850 );
or ( n36880 , n36877 , n36878 , n36879 );
xor ( n36881 , n36876 , n36880 );
and ( n36882 , n36872 , n36881 );
xor ( n36883 , n36739 , n36740 );
and ( n36884 , n36881 , n36883 );
and ( n36885 , n36872 , n36883 );
or ( n36886 , n36882 , n36884 , n36885 );
and ( n36887 , n36871 , n36886 );
xor ( n36888 , n36678 , n36679 );
xor ( n36889 , n36888 , n36681 );
and ( n36890 , n36886 , n36889 );
and ( n36891 , n36871 , n36889 );
or ( n36892 , n36887 , n36890 , n36891 );
and ( n36893 , n36867 , n36892 );
and ( n36894 , n36748 , n36892 );
or ( n36895 , n36868 , n36893 , n36894 );
xor ( n564178 , n36599 , n36601 );
xor ( n36896 , n564178 , n36603 );
xor ( n564180 , n36619 , n36626 );
xor ( n36897 , n564180 , n36674 );
and ( n36898 , n36896 , n36897 );
xor ( n36899 , n36684 , n36691 );
xor ( n36900 , n36899 , n36694 );
and ( n36901 , n36897 , n36900 );
and ( n564186 , n36896 , n36900 );
or ( n36902 , n36898 , n36901 , n564186 );
and ( n36903 , n36895 , n36902 );
xor ( n36904 , n36589 , n36591 );
xor ( n36905 , n36904 , n36606 );
and ( n36906 , n36902 , n36905 );
and ( n36907 , n36895 , n36905 );
or ( n36908 , n36903 , n36906 , n36907 );
and ( n36909 , n36738 , n36908 );
xor ( n36910 , n36585 , n36587 );
xor ( n36911 , n36910 , n36609 );
and ( n36912 , n36908 , n36911 );
and ( n36913 , n36738 , n36911 );
or ( n36914 , n36909 , n36912 , n36913 );
and ( n36915 , n36713 , n36914 );
and ( n36916 , n36711 , n36914 );
or ( n36917 , n36714 , n36915 , n36916 );
and ( n36918 , n36617 , n36917 );
and ( n36919 , n36615 , n36917 );
or ( n36920 , n36618 , n36918 , n36919 );
and ( n36921 , n36577 , n36920 );
and ( n36922 , n36575 , n36920 );
or ( n36923 , n36578 , n36921 , n36922 );
and ( n36924 , n36572 , n36923 );
and ( n36925 , n36570 , n36923 );
or ( n36926 , n36573 , n36924 , n36925 );
and ( n36927 , n36396 , n36926 );
and ( n36928 , n36394 , n36926 );
or ( n36929 , n36397 , n36927 , n36928 );
or ( n36930 , n36392 , n36929 );
and ( n36931 , n36389 , n36930 );
and ( n36932 , n35950 , n36930 );
or ( n36933 , n36390 , n36931 , n36932 );
and ( n36934 , n35947 , n36933 );
and ( n36935 , n35945 , n36933 );
or ( n36936 , n35948 , n36934 , n36935 );
and ( n36937 , n35696 , n36936 );
and ( n36938 , n35694 , n36936 );
or ( n36939 , n35697 , n36937 , n36938 );
and ( n36940 , n35461 , n36939 );
and ( n36941 , n35459 , n36939 );
or ( n36942 , n35462 , n36940 , n36941 );
and ( n36943 , n35219 , n36942 );
and ( n36944 , n35217 , n36942 );
or ( n36945 , n35220 , n36943 , n36944 );
and ( n36946 , n34958 , n36945 );
xor ( n36947 , n34958 , n36945 );
xor ( n36948 , n35217 , n35219 );
xor ( n36949 , n36948 , n36942 );
xor ( n36950 , n35459 , n35461 );
xor ( n36951 , n36950 , n36939 );
not ( n36952 , n36951 );
xor ( n36953 , n35694 , n35696 );
xor ( n36954 , n36953 , n36936 );
xor ( n36955 , n35945 , n35947 );
xor ( n36956 , n36955 , n36933 );
xor ( n36957 , n35950 , n36389 );
xor ( n36958 , n36957 , n36930 );
xnor ( n36959 , n36392 , n36929 );
xor ( n36960 , n36394 , n36396 );
xor ( n36961 , n36960 , n36926 );
xor ( n36962 , n36570 , n36572 );
xor ( n36963 , n36962 , n36923 );
not ( n36964 , n36963 );
xor ( n36965 , n36575 , n36577 );
xor ( n36966 , n36965 , n36920 );
xor ( n36967 , n36580 , n36582 );
xor ( n36968 , n36967 , n36612 );
xor ( n36969 , n36703 , n36705 );
xor ( n36970 , n36969 , n36708 );
xor ( n36971 , n36677 , n36697 );
xor ( n36972 , n36971 , n36700 );
xnor ( n36973 , n36728 , n36731 );
and ( n36974 , n36819 , n36820 );
and ( n36975 , n36820 , n36836 );
and ( n36976 , n36819 , n36836 );
or ( n36977 , n36974 , n36975 , n36976 );
and ( n36978 , n36973 , n36977 );
and ( n36979 , n36876 , n36880 );
and ( n36980 , n36977 , n36979 );
and ( n36981 , n36973 , n36979 );
or ( n36982 , n36978 , n36980 , n36981 );
xor ( n36983 , n36685 , n36686 );
xor ( n36984 , n36983 , n36688 );
xor ( n36985 , n36651 , n36652 );
xor ( n36986 , n36985 , n36654 );
xor ( n36987 , n36658 , n36659 );
xor ( n36988 , n36987 , n36661 );
and ( n36989 , n36986 , n36988 );
xor ( n36990 , n36628 , n36629 );
xor ( n36991 , n36990 , n36631 );
xor ( n36992 , n36635 , n36636 );
xor ( n36993 , n36992 , n36638 );
and ( n36994 , n36991 , n36993 );
and ( n36995 , n36989 , n36994 );
xor ( n36996 , n36828 , n36835 );
and ( n36997 , n34480 , n30947 );
and ( n36998 , n33204 , n31597 );
and ( n36999 , n36997 , n36998 );
and ( n37000 , n30962 , n34453 );
and ( n37001 , n31619 , n33213 );
and ( n37002 , n37000 , n37001 );
and ( n37003 , n36999 , n37002 );
and ( n37004 , n36996 , n37003 );
xor ( n37005 , n36822 , n36823 );
xor ( n37006 , n37005 , n36825 );
xor ( n37007 , n36829 , n36830 );
xor ( n37008 , n37007 , n36832 );
and ( n37009 , n37006 , n37008 );
and ( n37010 , n37003 , n37009 );
and ( n37011 , n36996 , n37009 );
or ( n37012 , n37004 , n37010 , n37011 );
and ( n37013 , n36995 , n37012 );
xor ( n37014 , n36766 , n36817 );
xor ( n37015 , n37014 , n36837 );
and ( n37016 , n37012 , n37015 );
and ( n37017 , n36995 , n37015 );
or ( n37018 , n37013 , n37016 , n37017 );
and ( n37019 , n36984 , n37018 );
xor ( n37020 , n36852 , n36863 );
xor ( n37021 , n36729 , n36730 );
and ( n37022 , n37020 , n37021 );
xor ( n37023 , n36869 , n36870 );
and ( n37024 , n37021 , n37023 );
and ( n37025 , n37020 , n37023 );
or ( n37026 , n37022 , n37024 , n37025 );
and ( n37027 , n37018 , n37026 );
and ( n37028 , n36984 , n37026 );
or ( n37029 , n37019 , n37027 , n37028 );
and ( n37030 , n36982 , n37029 );
and ( n37031 , n34049 , n31278 );
and ( n37032 , n33894 , n31414 );
and ( n37033 , n37031 , n37032 );
and ( n37034 , n32940 , n31871 );
and ( n37035 , n37032 , n37034 );
and ( n37036 , n37031 , n37034 );
or ( n37037 , n37033 , n37035 , n37036 );
xor ( n37038 , n36767 , n36768 );
xor ( n37039 , n37038 , n36770 );
and ( n37040 , n37037 , n37039 );
xor ( n37041 , n36774 , n36775 );
xor ( n37042 , n37041 , n36777 );
and ( n37043 , n37039 , n37042 );
and ( n37044 , n37037 , n37042 );
or ( n37045 , n37040 , n37043 , n37044 );
xor ( n37046 , n36798 , n36805 );
xor ( n37047 , n37046 , n36813 );
or ( n37048 , n37045 , n37047 );
and ( n37049 , n31269 , n34032 );
and ( n37050 , n31405 , n33914 );
and ( n37051 , n37049 , n37050 );
and ( n37052 , n31888 , n32922 );
and ( n37053 , n37050 , n37052 );
and ( n37054 , n37049 , n37052 );
or ( n37055 , n37051 , n37053 , n37054 );
xor ( n37056 , n36792 , n36793 );
xor ( n37057 , n37056 , n36795 );
and ( n37058 , n37055 , n37057 );
xor ( n37059 , n36799 , n36800 );
xor ( n37060 , n37059 , n36802 );
and ( n37061 , n37057 , n37060 );
and ( n37062 , n37055 , n37060 );
or ( n37063 , n37058 , n37061 , n37062 );
xor ( n37064 , n36773 , n36780 );
xor ( n37065 , n37064 , n36788 );
or ( n37066 , n37063 , n37065 );
and ( n37067 , n37048 , n37066 );
xor ( n37068 , n36843 , n36851 );
xor ( n37069 , n36854 , n36862 );
and ( n37070 , n37068 , n37069 );
and ( n37071 , n37067 , n37070 );
xor ( n37072 , n36755 , n36759 );
xor ( n37073 , n37072 , n36763 );
xor ( n37074 , n36791 , n36816 );
and ( n37075 , n37073 , n37074 );
xor ( n37076 , n36989 , n36994 );
and ( n37077 , n37074 , n37076 );
and ( n37078 , n37073 , n37076 );
or ( n37079 , n37075 , n37077 , n37078 );
and ( n37080 , n37070 , n37079 );
and ( n37081 , n37067 , n37079 );
or ( n37082 , n37071 , n37080 , n37081 );
xor ( n37083 , n36997 , n36998 );
xor ( n37084 , n37000 , n37001 );
and ( n37085 , n37083 , n37084 );
xor ( n37086 , n36756 , n36758 );
and ( n37087 , n37085 , n37086 );
and ( n37088 , n31430 , n33556 );
and ( n37089 , n31619 , n33532 );
and ( n37090 , n37088 , n37089 );
and ( n37091 , n32019 , n32850 );
and ( n37092 , n37089 , n37091 );
and ( n37093 , n37088 , n37091 );
or ( n37094 , n37090 , n37092 , n37093 );
not ( n37095 , n37094 );
and ( n37096 , n31057 , n34453 );
and ( n37097 , n31171 , n34298 );
and ( n37098 , n37096 , n37097 );
and ( n37099 , n31783 , n33213 );
and ( n37100 , n37097 , n37099 );
and ( n37101 , n37096 , n37099 );
or ( n37102 , n37098 , n37100 , n37101 );
and ( n37103 , n37095 , n37102 );
and ( n37104 , n33513 , n31453 );
and ( n37105 , n33575 , n31597 );
and ( n37106 , n37104 , n37105 );
and ( n37107 , n32868 , n31997 );
and ( n37108 , n37105 , n37107 );
and ( n37109 , n37104 , n37107 );
or ( n37110 , n37106 , n37108 , n37109 );
not ( n37111 , n37110 );
and ( n37112 , n34480 , n31066 );
and ( n37113 , n34315 , n31168 );
and ( n37114 , n37112 , n37113 );
and ( n37115 , n33204 , n31766 );
and ( n37116 , n37113 , n37115 );
and ( n37117 , n37112 , n37115 );
or ( n37118 , n37114 , n37116 , n37117 );
and ( n37119 , n37111 , n37118 );
and ( n37120 , n37103 , n37119 );
and ( n37121 , n37087 , n37120 );
buf ( n37122 , n37094 );
buf ( n37123 , n37110 );
and ( n37124 , n37122 , n37123 );
and ( n37125 , n37120 , n37124 );
and ( n37126 , n37087 , n37124 );
or ( n37127 , n37121 , n37125 , n37126 );
xor ( n37128 , n36986 , n36988 );
xor ( n37129 , n36991 , n36993 );
and ( n37130 , n37128 , n37129 );
xor ( n37131 , n36761 , n36762 );
xor ( n37132 , n36750 , n36751 );
and ( n37133 , n37131 , n37132 );
xor ( n37134 , n36999 , n37002 );
and ( n37135 , n37132 , n37134 );
and ( n37136 , n37131 , n37134 );
or ( n37137 , n37133 , n37135 , n37136 );
and ( n37138 , n37130 , n37137 );
xor ( n37139 , n36996 , n37003 );
xor ( n37140 , n37139 , n37009 );
and ( n37141 , n37137 , n37140 );
and ( n37142 , n37130 , n37140 );
or ( n37143 , n37138 , n37141 , n37142 );
and ( n37144 , n37127 , n37143 );
xor ( n37145 , n36872 , n36881 );
xor ( n37146 , n37145 , n36883 );
and ( n37147 , n37143 , n37146 );
and ( n37148 , n37127 , n37146 );
or ( n37149 , n37144 , n37147 , n37148 );
and ( n37150 , n37082 , n37149 );
xor ( n37151 , n36741 , n36743 );
xor ( n37152 , n37151 , n36745 );
and ( n37153 , n37149 , n37152 );
and ( n37154 , n37082 , n37152 );
or ( n37155 , n37150 , n37153 , n37154 );
and ( n37156 , n37029 , n37155 );
and ( n37157 , n36982 , n37155 );
or ( n37158 , n37030 , n37156 , n37157 );
and ( n37159 , n36972 , n37158 );
xor ( n37160 , n36721 , n36723 );
xor ( n37161 , n37160 , n36732 );
xor ( n37162 , n36748 , n36867 );
xor ( n37163 , n37162 , n36892 );
and ( n37164 , n37161 , n37163 );
xor ( n37165 , n36896 , n36897 );
xor ( n37166 , n37165 , n36900 );
and ( n37167 , n37163 , n37166 );
and ( n37168 , n37161 , n37166 );
or ( n37169 , n37164 , n37167 , n37168 );
and ( n37170 , n37158 , n37169 );
and ( n37171 , n36972 , n37169 );
or ( n37172 , n37159 , n37170 , n37171 );
and ( n37173 , n36970 , n37172 );
xor ( n37174 , n36738 , n36908 );
xor ( n37175 , n37174 , n36911 );
and ( n37176 , n37172 , n37175 );
and ( n37177 , n36970 , n37175 );
or ( n37178 , n37173 , n37176 , n37177 );
and ( n37179 , n36968 , n37178 );
xor ( n37180 , n36711 , n36713 );
xor ( n37181 , n37180 , n36914 );
and ( n37182 , n37178 , n37181 );
and ( n37183 , n36968 , n37181 );
or ( n37184 , n37179 , n37182 , n37183 );
xor ( n37185 , n36615 , n36617 );
xor ( n37186 , n37185 , n36917 );
and ( n37187 , n37184 , n37186 );
xor ( n37188 , n36968 , n37178 );
xor ( n37189 , n37188 , n37181 );
xor ( n37190 , n36716 , n36718 );
xor ( n37191 , n37190 , n36735 );
xor ( n37192 , n36895 , n36902 );
xor ( n37193 , n37192 , n36905 );
and ( n37194 , n37191 , n37193 );
xor ( n37195 , n36749 , n36840 );
xor ( n37196 , n37195 , n36864 );
xor ( n37197 , n36871 , n36886 );
xor ( n37198 , n37197 , n36889 );
and ( n37199 , n37196 , n37198 );
xor ( n37200 , n36973 , n36977 );
xor ( n37201 , n37200 , n36979 );
and ( n37202 , n37198 , n37201 );
and ( n37203 , n37196 , n37201 );
or ( n37204 , n37199 , n37202 , n37203 );
xor ( n37205 , n37048 , n37066 );
xor ( n37206 , n37068 , n37069 );
and ( n37207 , n37205 , n37206 );
xor ( n37208 , n36807 , n36808 );
xor ( n37209 , n37208 , n36810 );
xor ( n37210 , n36782 , n36783 );
xor ( n37211 , n37210 , n36785 );
and ( n37212 , n37209 , n37211 );
xor ( n37213 , n37085 , n37086 );
and ( n37214 , n37212 , n37213 );
and ( n37215 , n37206 , n37214 );
and ( n37216 , n37205 , n37214 );
or ( n37217 , n37207 , n37215 , n37216 );
xnor ( n37218 , n37045 , n37047 );
xnor ( n37219 , n37063 , n37065 );
and ( n37220 , n37218 , n37219 );
xor ( n37221 , n37006 , n37008 );
xor ( n37222 , n37103 , n37119 );
and ( n37223 , n37221 , n37222 );
xor ( n37224 , n37122 , n37123 );
and ( n37225 , n37222 , n37224 );
and ( n37226 , n37221 , n37224 );
or ( n37227 , n37223 , n37225 , n37226 );
and ( n37228 , n37220 , n37227 );
xor ( n37229 , n37128 , n37129 );
buf ( n37230 , n32302 );
buf ( n564516 , n543263 );
buf ( n37232 , n564516 );
and ( n37233 , n37230 , n37232 );
and ( n37234 , n34480 , n31168 );
and ( n37235 , n34315 , n31278 );
and ( n37236 , n37234 , n37235 );
and ( n37237 , n33204 , n31871 );
and ( n37238 , n37235 , n37237 );
and ( n37239 , n37234 , n37237 );
or ( n37240 , n37236 , n37238 , n37239 );
and ( n37241 , n31171 , n34453 );
and ( n37242 , n31269 , n34298 );
and ( n37243 , n37241 , n37242 );
and ( n37244 , n31888 , n33213 );
and ( n37245 , n37242 , n37244 );
and ( n37246 , n37241 , n37244 );
or ( n37247 , n37243 , n37245 , n37246 );
and ( n37248 , n37240 , n37247 );
or ( n37249 , n37233 , n37248 );
and ( n37250 , n37229 , n37249 );
and ( n37251 , n31619 , n33556 );
and ( n37252 , n32235 , n32850 );
and ( n37253 , n37251 , n37252 );
and ( n37254 , n32302 , n32508 );
and ( n37255 , n37252 , n37254 );
and ( n37256 , n37251 , n37254 );
or ( n37257 , n37253 , n37255 , n37256 );
and ( n37258 , n31405 , n34032 );
and ( n37259 , n31430 , n33914 );
and ( n37260 , n37258 , n37259 );
and ( n37261 , n32019 , n32922 );
and ( n37262 , n37259 , n37261 );
and ( n37263 , n37258 , n37261 );
or ( n37264 , n37260 , n37262 , n37263 );
and ( n37265 , n37257 , n37264 );
xor ( n37266 , n37104 , n37105 );
xor ( n37267 , n37266 , n37107 );
and ( n37268 , n37264 , n37267 );
and ( n37269 , n37257 , n37267 );
or ( n37270 , n37265 , n37268 , n37269 );
and ( n37271 , n33513 , n31597 );
and ( n37272 , n32868 , n32244 );
and ( n37273 , n37271 , n37272 );
and ( n37274 , n32525 , n32320 );
and ( n37275 , n37272 , n37274 );
and ( n37276 , n37271 , n37274 );
or ( n37277 , n37273 , n37275 , n37276 );
and ( n37278 , n34049 , n31414 );
and ( n37279 , n33894 , n31453 );
and ( n37280 , n37278 , n37279 );
and ( n37281 , n32940 , n31997 );
and ( n37282 , n37279 , n37281 );
and ( n37283 , n37278 , n37281 );
or ( n37284 , n37280 , n37282 , n37283 );
and ( n37285 , n37277 , n37284 );
xor ( n37286 , n37088 , n37089 );
xor ( n37287 , n37286 , n37091 );
and ( n37288 , n37284 , n37287 );
and ( n37289 , n37277 , n37287 );
or ( n37290 , n37285 , n37288 , n37289 );
and ( n37291 , n37270 , n37290 );
and ( n37292 , n37249 , n37291 );
and ( n37293 , n37229 , n37291 );
or ( n37294 , n37250 , n37292 , n37293 );
and ( n37295 , n37227 , n37294 );
and ( n37296 , n37220 , n37294 );
or ( n37297 , n37228 , n37295 , n37296 );
and ( n37298 , n37217 , n37297 );
xor ( n37299 , n37049 , n37050 );
xor ( n37300 , n37299 , n37052 );
xor ( n37301 , n37096 , n37097 );
xor ( n37302 , n37301 , n37099 );
and ( n37303 , n37300 , n37302 );
xor ( n37304 , n37031 , n37032 );
xor ( n37305 , n37304 , n37034 );
xor ( n37306 , n37112 , n37113 );
xor ( n37307 , n37306 , n37115 );
and ( n37308 , n37305 , n37307 );
and ( n37309 , n37303 , n37308 );
xor ( n37310 , n37055 , n37057 );
xor ( n37311 , n37310 , n37060 );
xor ( n37312 , n37037 , n37039 );
xor ( n37313 , n37312 , n37042 );
and ( n37314 , n37311 , n37313 );
and ( n37315 , n37309 , n37314 );
xor ( n37316 , n37095 , n37102 );
xor ( n37317 , n37111 , n37118 );
and ( n37318 , n37316 , n37317 );
and ( n37319 , n37314 , n37318 );
and ( n37320 , n37309 , n37318 );
or ( n37321 , n37315 , n37319 , n37320 );
xor ( n37322 , n37073 , n37074 );
xor ( n37323 , n37322 , n37076 );
and ( n37324 , n37321 , n37323 );
xor ( n37325 , n37087 , n37120 );
xor ( n37326 , n37325 , n37124 );
and ( n37327 , n37323 , n37326 );
and ( n37328 , n37321 , n37326 );
or ( n37329 , n37324 , n37327 , n37328 );
and ( n37330 , n37297 , n37329 );
and ( n37331 , n37217 , n37329 );
or ( n37332 , n37298 , n37330 , n37331 );
xor ( n37333 , n36995 , n37012 );
xor ( n37334 , n37333 , n37015 );
xor ( n37335 , n37020 , n37021 );
xor ( n37336 , n37335 , n37023 );
and ( n37337 , n37334 , n37336 );
xor ( n37338 , n37067 , n37070 );
xor ( n37339 , n37338 , n37079 );
and ( n37340 , n37336 , n37339 );
and ( n37341 , n37334 , n37339 );
or ( n37342 , n37337 , n37340 , n37341 );
and ( n37343 , n37332 , n37342 );
xor ( n37344 , n36984 , n37018 );
xor ( n37345 , n37344 , n37026 );
and ( n37346 , n37342 , n37345 );
and ( n37347 , n37332 , n37345 );
or ( n37348 , n37343 , n37346 , n37347 );
and ( n37349 , n37204 , n37348 );
xor ( n37350 , n36982 , n37029 );
xor ( n37351 , n37350 , n37155 );
and ( n37352 , n37348 , n37351 );
and ( n37353 , n37204 , n37351 );
or ( n37354 , n37349 , n37352 , n37353 );
and ( n37355 , n37193 , n37354 );
and ( n37356 , n37191 , n37354 );
or ( n37357 , n37194 , n37355 , n37356 );
xor ( n564643 , n36970 , n37172 );
xor ( n564644 , n564643 , n37175 );
and ( n564645 , n37357 , n564644 );
xor ( n37358 , n36972 , n37158 );
xor ( n37359 , n37358 , n37169 );
xor ( n37360 , n37161 , n37163 );
xor ( n37361 , n37360 , n37166 );
xor ( n37362 , n37082 , n37149 );
xor ( n37363 , n37362 , n37152 );
xor ( n37364 , n37127 , n37143 );
xor ( n37365 , n37364 , n37146 );
xor ( n37366 , n37130 , n37137 );
xor ( n37367 , n37366 , n37140 );
buf ( n564656 , n543260 );
buf ( n37369 , n564656 );
and ( n37370 , n32235 , n32508 );
and ( n37371 , n32525 , n32244 );
and ( n37372 , n37370 , n37371 );
and ( n37373 , n37369 , n37372 );
xor ( n37374 , n37209 , n37211 );
and ( n37375 , n37372 , n37374 );
and ( n37376 , n37369 , n37374 );
or ( n37377 , n37373 , n37375 , n37376 );
xor ( n37378 , n37131 , n37132 );
xor ( n37379 , n37378 , n37134 );
and ( n37380 , n37377 , n37379 );
xor ( n37381 , n37212 , n37213 );
and ( n37382 , n37379 , n37381 );
and ( n37383 , n37377 , n37381 );
or ( n37384 , n37380 , n37382 , n37383 );
and ( n37385 , n37367 , n37384 );
xor ( n37386 , n37218 , n37219 );
xor ( n37387 , n37230 , n37232 );
and ( n37388 , n32302 , n32850 );
and ( n37389 , n32868 , n32320 );
and ( n37390 , n37388 , n37389 );
buf ( n564679 , n543266 );
buf ( n37392 , n564679 );
and ( n37393 , n37390 , n37392 );
and ( n37394 , n37387 , n37393 );
and ( n37395 , n31783 , n33532 );
and ( n37396 , n33575 , n31766 );
and ( n37397 , n37395 , n37396 );
and ( n37398 , n37393 , n37397 );
and ( n37399 , n37387 , n37397 );
or ( n37400 , n37394 , n37398 , n37399 );
xor ( n37401 , n37300 , n37302 );
xor ( n37402 , n37305 , n37307 );
and ( n37403 , n37401 , n37402 );
and ( n37404 , n37400 , n37403 );
and ( n37405 , n37386 , n37404 );
and ( n37406 , n34480 , n31278 );
and ( n37407 , n33575 , n31871 );
and ( n37408 , n37406 , n37407 );
and ( n37409 , n32940 , n32244 );
and ( n37410 , n37407 , n37409 );
and ( n37411 , n37406 , n37409 );
or ( n37412 , n37408 , n37410 , n37411 );
and ( n37413 , n34315 , n31414 );
and ( n37414 , n34049 , n31453 );
and ( n37415 , n37413 , n37414 );
and ( n37416 , n33204 , n31997 );
and ( n37417 , n37414 , n37416 );
and ( n37418 , n37413 , n37416 );
or ( n37419 , n37415 , n37417 , n37418 );
and ( n37420 , n37412 , n37419 );
xor ( n37421 , n37241 , n37242 );
xor ( n37422 , n37421 , n37244 );
and ( n37423 , n37419 , n37422 );
and ( n37424 , n37412 , n37422 );
or ( n37425 , n37420 , n37423 , n37424 );
xor ( n37426 , n37277 , n37284 );
xor ( n37427 , n37426 , n37287 );
or ( n37428 , n37425 , n37427 );
and ( n37429 , n31269 , n34453 );
and ( n37430 , n31888 , n33532 );
and ( n37431 , n37429 , n37430 );
and ( n37432 , n32235 , n32922 );
and ( n37433 , n37430 , n37432 );
and ( n37434 , n37429 , n37432 );
or ( n37435 , n37431 , n37433 , n37434 );
and ( n37436 , n31405 , n34298 );
and ( n37437 , n31430 , n34032 );
and ( n37438 , n37436 , n37437 );
and ( n37439 , n32019 , n33213 );
and ( n37440 , n37437 , n37439 );
and ( n37441 , n37436 , n37439 );
or ( n37442 , n37438 , n37440 , n37441 );
and ( n37443 , n37435 , n37442 );
xor ( n37444 , n37234 , n37235 );
xor ( n37445 , n37444 , n37237 );
and ( n37446 , n37442 , n37445 );
and ( n37447 , n37435 , n37445 );
or ( n37448 , n37443 , n37446 , n37447 );
xor ( n37449 , n37257 , n37264 );
xor ( n37450 , n37449 , n37267 );
or ( n37451 , n37448 , n37450 );
and ( n37452 , n37428 , n37451 );
and ( n37453 , n37404 , n37452 );
and ( n37454 , n37386 , n37452 );
or ( n37455 , n37405 , n37453 , n37454 );
and ( n37456 , n37384 , n37455 );
and ( n37457 , n37367 , n37455 );
or ( n37458 , n37385 , n37456 , n37457 );
and ( n37459 , n37365 , n37458 );
xor ( n37460 , n37083 , n37084 );
xnor ( n37461 , n37233 , n37248 );
and ( n37462 , n37460 , n37461 );
xor ( n37463 , n37270 , n37290 );
and ( n37464 , n37461 , n37463 );
and ( n37465 , n37460 , n37463 );
or ( n37466 , n37462 , n37464 , n37465 );
xor ( n37467 , n37303 , n37308 );
xor ( n37468 , n37311 , n37313 );
and ( n37469 , n37467 , n37468 );
xor ( n37470 , n37316 , n37317 );
and ( n37471 , n37468 , n37470 );
and ( n37472 , n37467 , n37470 );
or ( n37473 , n37469 , n37471 , n37472 );
and ( n37474 , n37466 , n37473 );
xor ( n37475 , n37251 , n37252 );
xor ( n37476 , n37475 , n37254 );
xor ( n37477 , n37258 , n37259 );
xor ( n37478 , n37477 , n37261 );
or ( n37479 , n37476 , n37478 );
xor ( n37480 , n37271 , n37272 );
xor ( n37481 , n37480 , n37274 );
xor ( n37482 , n37278 , n37279 );
xor ( n37483 , n37482 , n37281 );
or ( n37484 , n37481 , n37483 );
and ( n37485 , n37479 , n37484 );
xor ( n37486 , n37370 , n37371 );
xor ( n37487 , n37240 , n37247 );
and ( n37488 , n37486 , n37487 );
and ( n37489 , n33894 , n31597 );
not ( n37490 , n37489 );
and ( n37491 , n33513 , n31766 );
and ( n37492 , n37490 , n37491 );
and ( n37493 , n31619 , n33914 );
not ( n37494 , n37493 );
and ( n37495 , n31783 , n33556 );
and ( n37496 , n37494 , n37495 );
and ( n37497 , n37492 , n37496 );
and ( n37498 , n37487 , n37497 );
and ( n37499 , n37486 , n37497 );
or ( n37500 , n37488 , n37498 , n37499 );
and ( n37501 , n37485 , n37500 );
xor ( n37502 , n37369 , n37372 );
xor ( n37503 , n37502 , n37374 );
and ( n37504 , n37500 , n37503 );
and ( n37505 , n37485 , n37503 );
or ( n37506 , n37501 , n37504 , n37505 );
and ( n37507 , n37473 , n37506 );
and ( n37508 , n37466 , n37506 );
or ( n37509 , n37474 , n37507 , n37508 );
xor ( n37510 , n37221 , n37222 );
xor ( n37511 , n37510 , n37224 );
xor ( n37512 , n37229 , n37249 );
xor ( n37513 , n37512 , n37291 );
and ( n37514 , n37511 , n37513 );
xor ( n37515 , n37309 , n37314 );
xor ( n37516 , n37515 , n37318 );
and ( n37517 , n37513 , n37516 );
and ( n37518 , n37511 , n37516 );
or ( n37519 , n37514 , n37517 , n37518 );
and ( n37520 , n37509 , n37519 );
xor ( n37521 , n37205 , n37206 );
xor ( n37522 , n37521 , n37214 );
and ( n37523 , n37519 , n37522 );
and ( n37524 , n37509 , n37522 );
or ( n37525 , n37520 , n37523 , n37524 );
and ( n37526 , n37458 , n37525 );
and ( n37527 , n37365 , n37525 );
or ( n37528 , n37459 , n37526 , n37527 );
and ( n37529 , n37363 , n37528 );
xor ( n37530 , n37196 , n37198 );
xor ( n37531 , n37530 , n37201 );
and ( n37532 , n37528 , n37531 );
and ( n37533 , n37363 , n37531 );
or ( n37534 , n37529 , n37532 , n37533 );
and ( n37535 , n37361 , n37534 );
xor ( n37536 , n37204 , n37348 );
xor ( n37537 , n37536 , n37351 );
and ( n37538 , n37534 , n37537 );
and ( n37539 , n37361 , n37537 );
or ( n37540 , n37535 , n37538 , n37539 );
and ( n37541 , n37359 , n37540 );
xor ( n37542 , n37191 , n37193 );
xor ( n37543 , n37542 , n37354 );
and ( n37544 , n37540 , n37543 );
and ( n37545 , n37359 , n37543 );
or ( n37546 , n37541 , n37544 , n37545 );
and ( n37547 , n564644 , n37546 );
and ( n37548 , n37357 , n37546 );
or ( n37549 , n564645 , n37547 , n37548 );
and ( n37550 , n37189 , n37549 );
xor ( n37551 , n37357 , n564644 );
xor ( n37552 , n37551 , n37546 );
xor ( n37553 , n37359 , n37540 );
xor ( n37554 , n37553 , n37543 );
xor ( n37555 , n37332 , n37342 );
xor ( n37556 , n37555 , n37345 );
xor ( n564845 , n37217 , n37297 );
xor ( n564846 , n564845 , n37329 );
xor ( n564847 , n37334 , n37336 );
xor ( n37557 , n564847 , n37339 );
and ( n37558 , n564846 , n37557 );
xor ( n37559 , n37220 , n37227 );
xor ( n37560 , n37559 , n37294 );
xor ( n37561 , n37321 , n37323 );
xor ( n37562 , n37561 , n37326 );
and ( n37563 , n37560 , n37562 );
xor ( n37564 , n37400 , n37403 );
xor ( n37565 , n37428 , n37451 );
and ( n37566 , n37564 , n37565 );
xor ( n37567 , n37390 , n37392 );
and ( n37568 , n33894 , n31766 );
and ( n37569 , n32940 , n32320 );
and ( n37570 , n37568 , n37569 );
and ( n37571 , n32868 , n32508 );
and ( n37572 , n37569 , n37571 );
and ( n37573 , n37568 , n37571 );
or ( n37574 , n37570 , n37572 , n37573 );
and ( n37575 , n31783 , n33914 );
and ( n37576 , n32302 , n32922 );
and ( n37577 , n37575 , n37576 );
and ( n37578 , n32525 , n32850 );
and ( n37579 , n37576 , n37578 );
and ( n37580 , n37575 , n37578 );
or ( n37581 , n37577 , n37579 , n37580 );
and ( n37582 , n37574 , n37581 );
and ( n37583 , n37567 , n37582 );
and ( n37584 , n34315 , n31453 );
and ( n37585 , n34049 , n31597 );
and ( n37586 , n37584 , n37585 );
and ( n37587 , n33204 , n32244 );
and ( n37588 , n37585 , n37587 );
and ( n37589 , n37584 , n37587 );
or ( n37590 , n37586 , n37588 , n37589 );
and ( n37591 , n31430 , n34298 );
and ( n37592 , n31619 , n34032 );
and ( n37593 , n37591 , n37592 );
and ( n37594 , n32235 , n33213 );
and ( n37595 , n37592 , n37594 );
and ( n37596 , n37591 , n37594 );
or ( n37597 , n37593 , n37595 , n37596 );
and ( n37598 , n37590 , n37597 );
and ( n37599 , n37582 , n37598 );
and ( n37600 , n37567 , n37598 );
or ( n37601 , n37583 , n37599 , n37600 );
xor ( n37602 , n37435 , n37442 );
xor ( n37603 , n37602 , n37445 );
xor ( n37604 , n37412 , n37419 );
xor ( n37605 , n37604 , n37422 );
and ( n37606 , n37603 , n37605 );
and ( n37607 , n37601 , n37606 );
xor ( n37608 , n37387 , n37393 );
xor ( n37609 , n37608 , n37397 );
and ( n37610 , n37606 , n37609 );
and ( n37611 , n37601 , n37609 );
or ( n37612 , n37607 , n37610 , n37611 );
and ( n37613 , n37565 , n37612 );
and ( n37614 , n37564 , n37612 );
or ( n37615 , n37566 , n37613 , n37614 );
xnor ( n37616 , n37425 , n37427 );
xnor ( n37617 , n37448 , n37450 );
and ( n37618 , n37616 , n37617 );
buf ( n564910 , n37489 );
buf ( n564911 , n37493 );
and ( n564912 , n564910 , n564911 );
xor ( n37619 , n37479 , n37484 );
and ( n37620 , n564912 , n37619 );
xor ( n37621 , n37401 , n37402 );
and ( n37622 , n37619 , n37621 );
and ( n37623 , n564912 , n37621 );
or ( n37624 , n37620 , n37622 , n37623 );
and ( n37625 , n37618 , n37624 );
buf ( n37626 , n32525 );
buf ( n564921 , n543269 );
buf ( n37628 , n564921 );
and ( n37629 , n37626 , n37628 );
xor ( n37630 , n37490 , n37491 );
xor ( n37631 , n37494 , n37495 );
and ( n37632 , n37630 , n37631 );
or ( n37633 , n37629 , n37632 );
and ( n37634 , n31405 , n34453 );
and ( n37635 , n31888 , n33556 );
and ( n37636 , n37634 , n37635 );
and ( n37637 , n32019 , n33532 );
and ( n37638 , n37635 , n37637 );
and ( n37639 , n37634 , n37637 );
or ( n37640 , n37636 , n37638 , n37639 );
xor ( n37641 , n37406 , n37407 );
xor ( n37642 , n37641 , n37409 );
and ( n37643 , n37640 , n37642 );
xor ( n37644 , n37413 , n37414 );
xor ( n37645 , n37644 , n37416 );
and ( n37646 , n37642 , n37645 );
and ( n37647 , n37640 , n37645 );
or ( n37648 , n37643 , n37646 , n37647 );
and ( n37649 , n34480 , n31414 );
and ( n37650 , n33513 , n31871 );
and ( n37651 , n37649 , n37650 );
and ( n37652 , n33575 , n31997 );
and ( n37653 , n37650 , n37652 );
and ( n37654 , n37649 , n37652 );
or ( n37655 , n37651 , n37653 , n37654 );
xor ( n37656 , n37429 , n37430 );
xor ( n37657 , n37656 , n37432 );
and ( n37658 , n37655 , n37657 );
xor ( n37659 , n37436 , n37437 );
xor ( n37660 , n37659 , n37439 );
and ( n37661 , n37657 , n37660 );
and ( n37662 , n37655 , n37660 );
or ( n37663 , n37658 , n37661 , n37662 );
and ( n37664 , n37648 , n37663 );
and ( n37665 , n37633 , n37664 );
xnor ( n37666 , n37476 , n37478 );
xnor ( n37667 , n37481 , n37483 );
and ( n37668 , n37666 , n37667 );
and ( n37669 , n37664 , n37668 );
and ( n37670 , n37633 , n37668 );
or ( n37671 , n37665 , n37669 , n37670 );
and ( n37672 , n37624 , n37671 );
and ( n37673 , n37618 , n37671 );
or ( n37674 , n37625 , n37672 , n37673 );
and ( n37675 , n37615 , n37674 );
xor ( n37676 , n37460 , n37461 );
xor ( n37677 , n37676 , n37463 );
xor ( n37678 , n37467 , n37468 );
xor ( n37679 , n37678 , n37470 );
and ( n37680 , n37677 , n37679 );
xor ( n37681 , n37485 , n37500 );
xor ( n37682 , n37681 , n37503 );
and ( n37683 , n37679 , n37682 );
and ( n37684 , n37677 , n37682 );
or ( n37685 , n37680 , n37683 , n37684 );
and ( n37686 , n37674 , n37685 );
and ( n37687 , n37615 , n37685 );
or ( n37688 , n37675 , n37686 , n37687 );
and ( n37689 , n37562 , n37688 );
and ( n37690 , n37560 , n37688 );
or ( n37691 , n37563 , n37689 , n37690 );
and ( n37692 , n37557 , n37691 );
and ( n37693 , n564846 , n37691 );
or ( n37694 , n37558 , n37692 , n37693 );
and ( n37695 , n37556 , n37694 );
xor ( n37696 , n37363 , n37528 );
xor ( n37697 , n37696 , n37531 );
and ( n37698 , n37694 , n37697 );
and ( n37699 , n37556 , n37697 );
or ( n37700 , n37695 , n37698 , n37699 );
xor ( n37701 , n37361 , n37534 );
xor ( n37702 , n37701 , n37537 );
and ( n37703 , n37700 , n37702 );
xor ( n37704 , n37377 , n37379 );
xor ( n37705 , n37704 , n37381 );
xor ( n37706 , n37386 , n37404 );
xor ( n37707 , n37706 , n37452 );
and ( n37708 , n37705 , n37707 );
xor ( n37709 , n37466 , n37473 );
xor ( n37710 , n37709 , n37506 );
and ( n37711 , n37707 , n37710 );
and ( n37712 , n37705 , n37710 );
or ( n37713 , n37708 , n37711 , n37712 );
xor ( n37714 , n37367 , n37384 );
xor ( n37715 , n37714 , n37455 );
and ( n37716 , n37713 , n37715 );
xor ( n37717 , n37509 , n37519 );
xor ( n37718 , n37717 , n37522 );
and ( n37719 , n37715 , n37718 );
and ( n37720 , n37713 , n37718 );
or ( n37721 , n37716 , n37719 , n37720 );
xor ( n37722 , n37365 , n37458 );
xor ( n37723 , n37722 , n37525 );
and ( n37724 , n37721 , n37723 );
xor ( n37725 , n37511 , n37513 );
xor ( n37726 , n37725 , n37516 );
xor ( n37727 , n37395 , n37396 );
xor ( n37728 , n37492 , n37496 );
and ( n37729 , n37727 , n37728 );
xor ( n37730 , n564910 , n564911 );
and ( n37731 , n37728 , n37730 );
and ( n37732 , n37727 , n37730 );
or ( n37733 , n37729 , n37731 , n37732 );
xor ( n37734 , n37486 , n37487 );
xor ( n37735 , n37734 , n37497 );
and ( n37736 , n37733 , n37735 );
xor ( n37737 , n37601 , n37606 );
xor ( n37738 , n37737 , n37609 );
and ( n37739 , n37735 , n37738 );
and ( n37740 , n37733 , n37738 );
or ( n37741 , n37736 , n37739 , n37740 );
xor ( n37742 , n37616 , n37617 );
xnor ( n37743 , n37629 , n37632 );
xor ( n37744 , n37626 , n37628 );
and ( n37745 , n32525 , n32922 );
and ( n37746 , n32940 , n32508 );
and ( n37747 , n37745 , n37746 );
buf ( n565042 , n543272 );
buf ( n37749 , n565042 );
and ( n37750 , n37747 , n37749 );
and ( n37751 , n37744 , n37750 );
and ( n37752 , n33894 , n31871 );
and ( n37753 , n33513 , n31997 );
and ( n37754 , n37752 , n37753 );
and ( n37755 , n33204 , n32320 );
and ( n37756 , n37753 , n37755 );
and ( n37757 , n37752 , n37755 );
or ( n37758 , n37754 , n37756 , n37757 );
and ( n37759 , n31888 , n33914 );
and ( n37760 , n32019 , n33556 );
and ( n37761 , n37759 , n37760 );
and ( n37762 , n32302 , n33213 );
and ( n37763 , n37760 , n37762 );
and ( n37764 , n37759 , n37762 );
or ( n37765 , n37761 , n37763 , n37764 );
and ( n37766 , n37758 , n37765 );
and ( n37767 , n37750 , n37766 );
and ( n37768 , n37744 , n37766 );
or ( n37769 , n37751 , n37767 , n37768 );
and ( n37770 , n37743 , n37769 );
xor ( n37771 , n37567 , n37582 );
xor ( n37772 , n37771 , n37598 );
and ( n37773 , n37769 , n37772 );
and ( n37774 , n37743 , n37772 );
or ( n37775 , n37770 , n37773 , n37774 );
and ( n37776 , n37742 , n37775 );
and ( n37777 , n34480 , n31453 );
and ( n37778 , n34315 , n31597 );
and ( n37779 , n37777 , n37778 );
and ( n37780 , n33575 , n32244 );
and ( n37781 , n37778 , n37780 );
and ( n37782 , n37777 , n37780 );
or ( n37783 , n37779 , n37781 , n37782 );
xor ( n37784 , n37634 , n37635 );
xor ( n37785 , n37784 , n37637 );
and ( n37786 , n37783 , n37785 );
xor ( n37787 , n37575 , n37576 );
xor ( n37788 , n37787 , n37578 );
and ( n37789 , n37785 , n37788 );
and ( n37790 , n37783 , n37788 );
or ( n37791 , n37786 , n37789 , n37790 );
xor ( n37792 , n37655 , n37657 );
xor ( n37793 , n37792 , n37660 );
and ( n37794 , n37791 , n37793 );
and ( n37795 , n31430 , n34453 );
and ( n37796 , n31619 , n34298 );
and ( n37797 , n37795 , n37796 );
and ( n37798 , n32235 , n33532 );
and ( n37799 , n37796 , n37798 );
and ( n37800 , n37795 , n37798 );
or ( n37801 , n37797 , n37799 , n37800 );
xor ( n37802 , n37649 , n37650 );
xor ( n37803 , n37802 , n37652 );
and ( n37804 , n37801 , n37803 );
xor ( n37805 , n37568 , n37569 );
xor ( n37806 , n37805 , n37571 );
and ( n37807 , n37803 , n37806 );
and ( n37808 , n37801 , n37806 );
or ( n37809 , n37804 , n37807 , n37808 );
xor ( n37810 , n37640 , n37642 );
xor ( n37811 , n37810 , n37645 );
and ( n37812 , n37809 , n37811 );
and ( n37813 , n37794 , n37812 );
and ( n37814 , n37775 , n37813 );
and ( n37815 , n37742 , n37813 );
or ( n37816 , n37776 , n37814 , n37815 );
and ( n37817 , n37741 , n37816 );
xor ( n37818 , n37648 , n37663 );
xor ( n37819 , n37603 , n37605 );
and ( n37820 , n37818 , n37819 );
xor ( n37821 , n37666 , n37667 );
and ( n37822 , n37819 , n37821 );
and ( n37823 , n37818 , n37821 );
or ( n37824 , n37820 , n37822 , n37823 );
xor ( n37825 , n564912 , n37619 );
xor ( n37826 , n37825 , n37621 );
and ( n37827 , n37824 , n37826 );
xor ( n37828 , n37633 , n37664 );
xor ( n37829 , n37828 , n37668 );
and ( n37830 , n37826 , n37829 );
and ( n37831 , n37824 , n37829 );
or ( n37832 , n37827 , n37830 , n37831 );
and ( n37833 , n37816 , n37832 );
and ( n37834 , n37741 , n37832 );
or ( n37835 , n37817 , n37833 , n37834 );
and ( n37836 , n37726 , n37835 );
xor ( n37837 , n37564 , n37565 );
xor ( n37838 , n37837 , n37612 );
xor ( n37839 , n37618 , n37624 );
xor ( n37840 , n37839 , n37671 );
and ( n37841 , n37838 , n37840 );
xor ( n37842 , n37677 , n37679 );
xor ( n37843 , n37842 , n37682 );
and ( n37844 , n37840 , n37843 );
and ( n37845 , n37838 , n37843 );
or ( n37846 , n37841 , n37844 , n37845 );
and ( n37847 , n37835 , n37846 );
and ( n37848 , n37726 , n37846 );
or ( n37849 , n37836 , n37847 , n37848 );
xor ( n37850 , n37560 , n37562 );
xor ( n37851 , n37850 , n37688 );
and ( n37852 , n37849 , n37851 );
xor ( n37853 , n37713 , n37715 );
xor ( n37854 , n37853 , n37718 );
and ( n37855 , n37851 , n37854 );
and ( n37856 , n37849 , n37854 );
or ( n37857 , n37852 , n37855 , n37856 );
and ( n37858 , n37723 , n37857 );
and ( n37859 , n37721 , n37857 );
or ( n37860 , n37724 , n37858 , n37859 );
xor ( n37861 , n37556 , n37694 );
xor ( n37862 , n37861 , n37697 );
and ( n37863 , n37860 , n37862 );
xor ( n37864 , n564846 , n37557 );
xor ( n37865 , n37864 , n37691 );
xor ( n37866 , n37721 , n37723 );
xor ( n37867 , n37866 , n37857 );
and ( n37868 , n37865 , n37867 );
xor ( n37869 , n37615 , n37674 );
xor ( n37870 , n37869 , n37685 );
xor ( n37871 , n37705 , n37707 );
xor ( n37872 , n37871 , n37710 );
and ( n37873 , n37870 , n37872 );
xor ( n37874 , n37747 , n37749 );
buf ( n37875 , n32868 );
buf ( n565170 , n543275 );
buf ( n37877 , n565170 );
and ( n37878 , n37875 , n37877 );
and ( n37879 , n37874 , n37878 );
and ( n37880 , n31783 , n34032 );
and ( n37881 , n34049 , n31766 );
and ( n37882 , n37880 , n37881 );
and ( n37883 , n37878 , n37882 );
and ( n37884 , n37874 , n37882 );
or ( n37885 , n37879 , n37883 , n37884 );
xor ( n37886 , n37584 , n37585 );
xor ( n37887 , n37886 , n37587 );
xor ( n37888 , n37591 , n37592 );
xor ( n37889 , n37888 , n37594 );
and ( n37890 , n37887 , n37889 );
and ( n37891 , n37885 , n37890 );
xor ( n37892 , n37744 , n37750 );
xor ( n37893 , n37892 , n37766 );
and ( n565188 , n37890 , n37893 );
and ( n565189 , n37885 , n37893 );
or ( n565190 , n37891 , n565188 , n565189 );
xor ( n37894 , n37791 , n37793 );
xor ( n37895 , n37809 , n37811 );
and ( n37896 , n37894 , n37895 );
and ( n37897 , n565190 , n37896 );
xor ( n37898 , n37388 , n37389 );
xor ( n37899 , n37574 , n37581 );
and ( n37900 , n37898 , n37899 );
xor ( n37901 , n37590 , n37597 );
and ( n37902 , n37899 , n37901 );
and ( n37903 , n37898 , n37901 );
or ( n37904 , n37900 , n37902 , n37903 );
xor ( n37905 , n37727 , n37728 );
xor ( n37906 , n37905 , n37730 );
and ( n37907 , n37904 , n37906 );
xor ( n37908 , n37743 , n37769 );
xor ( n37909 , n37908 , n37772 );
and ( n37910 , n37906 , n37909 );
and ( n37911 , n37904 , n37909 );
or ( n37912 , n37907 , n37910 , n37911 );
and ( n37913 , n37897 , n37912 );
xor ( n37914 , n37794 , n37812 );
and ( n37915 , n34049 , n31871 );
and ( n37916 , n33204 , n32508 );
and ( n37917 , n37915 , n37916 );
and ( n37918 , n32940 , n32850 );
and ( n37919 , n37916 , n37918 );
and ( n37920 , n37915 , n37918 );
or ( n37921 , n37917 , n37919 , n37920 );
and ( n37922 , n34480 , n31597 );
and ( n37923 , n34315 , n31766 );
and ( n37924 , n37922 , n37923 );
and ( n37925 , n33575 , n32320 );
and ( n37926 , n37923 , n37925 );
and ( n37927 , n37922 , n37925 );
or ( n37928 , n37924 , n37926 , n37927 );
and ( n37929 , n37921 , n37928 );
xor ( n565227 , n37759 , n37760 );
xor ( n565228 , n565227 , n37762 );
and ( n565229 , n37928 , n565228 );
and ( n37930 , n37921 , n565228 );
or ( n37931 , n37929 , n565229 , n37930 );
xor ( n37932 , n37783 , n37785 );
xor ( n37933 , n37932 , n37788 );
or ( n37934 , n37931 , n37933 );
and ( n37935 , n31888 , n34032 );
and ( n37936 , n32525 , n33213 );
and ( n37937 , n37935 , n37936 );
and ( n37938 , n32868 , n32922 );
and ( n37939 , n37936 , n37938 );
and ( n37940 , n37935 , n37938 );
or ( n37941 , n37937 , n37939 , n37940 );
and ( n37942 , n31619 , n34453 );
and ( n37943 , n31783 , n34298 );
and ( n37944 , n37942 , n37943 );
and ( n37945 , n32302 , n33532 );
and ( n37946 , n37943 , n37945 );
and ( n37947 , n37942 , n37945 );
or ( n37948 , n37944 , n37946 , n37947 );
and ( n37949 , n37941 , n37948 );
xor ( n37950 , n37752 , n37753 );
xor ( n37951 , n37950 , n37755 );
and ( n37952 , n37948 , n37951 );
and ( n37953 , n37941 , n37951 );
or ( n37954 , n37949 , n37952 , n37953 );
xor ( n37955 , n37801 , n37803 );
xor ( n37956 , n37955 , n37806 );
or ( n37957 , n37954 , n37956 );
and ( n37958 , n37934 , n37957 );
and ( n37959 , n37914 , n37958 );
xor ( n37960 , n37630 , n37631 );
xor ( n37961 , n37758 , n37765 );
xor ( n37962 , n37887 , n37889 );
and ( n37963 , n37961 , n37962 );
and ( n37964 , n33894 , n31997 );
and ( n37965 , n33513 , n32244 );
or ( n37966 , n37964 , n37965 );
and ( n37967 , n32019 , n33914 );
and ( n37968 , n32235 , n33556 );
or ( n37969 , n37967 , n37968 );
and ( n37970 , n37966 , n37969 );
and ( n37971 , n37962 , n37970 );
and ( n37972 , n37961 , n37970 );
or ( n37973 , n37963 , n37971 , n37972 );
and ( n37974 , n37960 , n37973 );
xor ( n37975 , n37898 , n37899 );
xor ( n37976 , n37975 , n37901 );
and ( n37977 , n37973 , n37976 );
and ( n37978 , n37960 , n37976 );
or ( n37979 , n37974 , n37977 , n37978 );
and ( n37980 , n37958 , n37979 );
and ( n37981 , n37914 , n37979 );
or ( n37982 , n37959 , n37980 , n37981 );
and ( n37983 , n37912 , n37982 );
and ( n37984 , n37897 , n37982 );
or ( n37985 , n37913 , n37983 , n37984 );
xor ( n37986 , n37733 , n37735 );
xor ( n37987 , n37986 , n37738 );
xor ( n37988 , n37742 , n37775 );
xor ( n37989 , n37988 , n37813 );
and ( n37990 , n37987 , n37989 );
xor ( n37991 , n37824 , n37826 );
xor ( n37992 , n37991 , n37829 );
and ( n37993 , n37989 , n37992 );
and ( n37994 , n37987 , n37992 );
or ( n37995 , n37990 , n37993 , n37994 );
and ( n37996 , n37985 , n37995 );
xor ( n37997 , n37741 , n37816 );
xor ( n37998 , n37997 , n37832 );
and ( n37999 , n37995 , n37998 );
and ( n38000 , n37985 , n37998 );
or ( n38001 , n37996 , n37999 , n38000 );
and ( n38002 , n37872 , n38001 );
and ( n38003 , n37870 , n38001 );
or ( n38004 , n37873 , n38002 , n38003 );
xor ( n38005 , n37849 , n37851 );
xor ( n38006 , n38005 , n37854 );
and ( n38007 , n38004 , n38006 );
xor ( n38008 , n37726 , n37835 );
xor ( n38009 , n38008 , n37846 );
xor ( n38010 , n37838 , n37840 );
xor ( n38011 , n38010 , n37843 );
xor ( n38012 , n37818 , n37819 );
xor ( n38013 , n38012 , n37821 );
xor ( n38014 , n565190 , n37896 );
and ( n38015 , n38013 , n38014 );
xor ( n38016 , n37885 , n37890 );
xor ( n38017 , n38016 , n37893 );
xor ( n38018 , n37934 , n37957 );
and ( n38019 , n38017 , n38018 );
xor ( n38020 , n37894 , n37895 );
and ( n38021 , n38018 , n38020 );
and ( n38022 , n38017 , n38020 );
or ( n38023 , n38019 , n38021 , n38022 );
and ( n38024 , n38014 , n38023 );
and ( n38025 , n38013 , n38023 );
or ( n38026 , n38015 , n38024 , n38025 );
and ( n38027 , n32868 , n33213 );
and ( n38028 , n33204 , n32850 );
and ( n38029 , n38027 , n38028 );
buf ( n565330 , n543278 );
buf ( n38031 , n565330 );
and ( n38032 , n38029 , n38031 );
and ( n38033 , n34315 , n31871 );
and ( n38034 , n34049 , n31997 );
and ( n38035 , n38033 , n38034 );
and ( n38036 , n33575 , n32508 );
and ( n38037 , n38034 , n38036 );
and ( n38038 , n38033 , n38036 );
or ( n38039 , n38035 , n38037 , n38038 );
and ( n38040 , n31888 , n34298 );
and ( n38041 , n32019 , n34032 );
and ( n38042 , n38040 , n38041 );
and ( n38043 , n32525 , n33532 );
and ( n38044 , n38041 , n38043 );
and ( n38045 , n38040 , n38043 );
or ( n38046 , n38042 , n38044 , n38045 );
and ( n38047 , n38039 , n38046 );
and ( n38048 , n38032 , n38047 );
and ( n38049 , n34480 , n31766 );
and ( n38050 , n33894 , n32244 );
and ( n38051 , n38049 , n38050 );
and ( n38052 , n33513 , n32320 );
and ( n38053 , n38050 , n38052 );
and ( n38054 , n38049 , n38052 );
or ( n38055 , n38051 , n38053 , n38054 );
and ( n38056 , n31783 , n34453 );
and ( n38057 , n32235 , n33914 );
and ( n38058 , n38056 , n38057 );
and ( n38059 , n32302 , n33556 );
and ( n38060 , n38057 , n38059 );
and ( n38061 , n38056 , n38059 );
or ( n38062 , n38058 , n38060 , n38061 );
and ( n38063 , n38055 , n38062 );
and ( n38064 , n38047 , n38063 );
and ( n38065 , n38032 , n38063 );
or ( n38066 , n38048 , n38064 , n38065 );
xor ( n38067 , n37941 , n37948 );
xor ( n38068 , n38067 , n37951 );
xor ( n38069 , n37921 , n37928 );
xor ( n38070 , n38069 , n565228 );
and ( n38071 , n38068 , n38070 );
or ( n38072 , n38066 , n38071 );
xnor ( n38073 , n37931 , n37933 );
xnor ( n38074 , n37954 , n37956 );
and ( n38075 , n38073 , n38074 );
and ( n38076 , n38072 , n38075 );
xor ( n38077 , n37777 , n37778 );
xor ( n38078 , n38077 , n37780 );
xor ( n38079 , n37795 , n37796 );
xor ( n38080 , n38079 , n37798 );
and ( n38081 , n38078 , n38080 );
xor ( n38082 , n37875 , n37877 );
xor ( n38083 , n37880 , n37881 );
and ( n38084 , n38082 , n38083 );
xor ( n38085 , n37745 , n37746 );
and ( n38086 , n38083 , n38085 );
and ( n38087 , n38082 , n38085 );
or ( n38088 , n38084 , n38086 , n38087 );
and ( n38089 , n38081 , n38088 );
xor ( n38090 , n37874 , n37878 );
xor ( n38091 , n38090 , n37882 );
and ( n38092 , n38088 , n38091 );
and ( n38093 , n38081 , n38091 );
or ( n38094 , n38089 , n38092 , n38093 );
and ( n38095 , n38075 , n38094 );
and ( n38096 , n38072 , n38094 );
or ( n38097 , n38076 , n38095 , n38096 );
xor ( n38098 , n37904 , n37906 );
xor ( n38099 , n38098 , n37909 );
and ( n38100 , n38097 , n38099 );
xor ( n38101 , n37914 , n37958 );
xor ( n38102 , n38101 , n37979 );
and ( n38103 , n38099 , n38102 );
and ( n38104 , n38097 , n38102 );
or ( n38105 , n38100 , n38103 , n38104 );
and ( n38106 , n38026 , n38105 );
xor ( n38107 , n37897 , n37912 );
xor ( n38108 , n38107 , n37982 );
and ( n38109 , n38105 , n38108 );
and ( n38110 , n38026 , n38108 );
or ( n38111 , n38106 , n38109 , n38110 );
and ( n565412 , n38011 , n38111 );
xor ( n38112 , n37985 , n37995 );
xor ( n38113 , n38112 , n37998 );
and ( n38114 , n38111 , n38113 );
and ( n38115 , n38011 , n38113 );
or ( n38116 , n565412 , n38114 , n38115 );
and ( n38117 , n38009 , n38116 );
xor ( n38118 , n37870 , n37872 );
xor ( n38119 , n38118 , n38001 );
and ( n38120 , n38116 , n38119 );
and ( n38121 , n38009 , n38119 );
or ( n38122 , n38117 , n38120 , n38121 );
and ( n38123 , n38006 , n38122 );
and ( n38124 , n38004 , n38122 );
or ( n38125 , n38007 , n38123 , n38124 );
and ( n38126 , n37867 , n38125 );
and ( n38127 , n37865 , n38125 );
or ( n38128 , n37868 , n38126 , n38127 );
and ( n38129 , n37862 , n38128 );
and ( n38130 , n37860 , n38128 );
or ( n38131 , n37863 , n38129 , n38130 );
and ( n38132 , n37702 , n38131 );
and ( n38133 , n37700 , n38131 );
or ( n38134 , n37703 , n38132 , n38133 );
or ( n38135 , n37554 , n38134 );
or ( n38136 , n37552 , n38135 );
and ( n38137 , n37549 , n38136 );
and ( n38138 , n37189 , n38136 );
or ( n38139 , n37550 , n38137 , n38138 );
and ( n38140 , n37186 , n38139 );
and ( n38141 , n37184 , n38139 );
or ( n38142 , n37187 , n38140 , n38141 );
and ( n38143 , n36966 , n38142 );
xor ( n38144 , n36966 , n38142 );
xor ( n38145 , n37184 , n37186 );
xor ( n38146 , n38145 , n38139 );
xor ( n38147 , n37189 , n37549 );
xor ( n38148 , n38147 , n38136 );
not ( n38149 , n38148 );
xnor ( n38150 , n37552 , n38135 );
xnor ( n38151 , n37554 , n38134 );
xor ( n38152 , n37700 , n37702 );
xor ( n38153 , n38152 , n38131 );
not ( n38154 , n38153 );
xor ( n38155 , n37860 , n37862 );
xor ( n38156 , n38155 , n38128 );
xor ( n38157 , n37865 , n37867 );
xor ( n38158 , n38157 , n38125 );
xor ( n38159 , n38004 , n38006 );
xor ( n38160 , n38159 , n38122 );
xor ( n38161 , n38009 , n38116 );
xor ( n38162 , n38161 , n38119 );
xor ( n38163 , n37987 , n37989 );
xor ( n38164 , n38163 , n37992 );
xor ( n38165 , n37966 , n37969 );
xor ( n38166 , n38078 , n38080 );
and ( n38167 , n38165 , n38166 );
xor ( n38168 , n37915 , n37916 );
xor ( n38169 , n38168 , n37918 );
xor ( n38170 , n37935 , n37936 );
xor ( n38171 , n38170 , n37938 );
and ( n38172 , n38169 , n38171 );
and ( n38173 , n38166 , n38172 );
and ( n38174 , n38165 , n38172 );
or ( n38175 , n38167 , n38173 , n38174 );
xor ( n38176 , n37922 , n37923 );
xor ( n38177 , n38176 , n37925 );
xor ( n38178 , n37942 , n37943 );
xor ( n38179 , n38178 , n37945 );
and ( n38180 , n38177 , n38179 );
xnor ( n38181 , n37964 , n37965 );
xnor ( n38182 , n37967 , n37968 );
and ( n38183 , n38181 , n38182 );
and ( n38184 , n38180 , n38183 );
xor ( n38185 , n38082 , n38083 );
xor ( n38186 , n38185 , n38085 );
and ( n38187 , n38183 , n38186 );
and ( n38188 , n38180 , n38186 );
or ( n38189 , n38184 , n38187 , n38188 );
and ( n38190 , n38175 , n38189 );
xor ( n38191 , n37961 , n37962 );
xor ( n38192 , n38191 , n37970 );
and ( n38193 , n38189 , n38192 );
and ( n38194 , n38175 , n38192 );
or ( n38195 , n38190 , n38193 , n38194 );
xor ( n38196 , n37960 , n37973 );
xor ( n38197 , n38196 , n37976 );
and ( n38198 , n38195 , n38197 );
xnor ( n38199 , n38066 , n38071 );
xor ( n38200 , n38073 , n38074 );
and ( n38201 , n38199 , n38200 );
xor ( n38202 , n38032 , n38047 );
xor ( n38203 , n38202 , n38063 );
xor ( n38204 , n38068 , n38070 );
and ( n38205 , n38203 , n38204 );
and ( n38206 , n31888 , n34453 );
and ( n38207 , n32302 , n33914 );
and ( n38208 , n38206 , n38207 );
and ( n38209 , n32525 , n33556 );
and ( n38210 , n38207 , n38209 );
and ( n38211 , n38206 , n38209 );
or ( n38212 , n38208 , n38210 , n38211 );
xor ( n38213 , n38033 , n38034 );
xor ( n38214 , n38213 , n38036 );
and ( n38215 , n38212 , n38214 );
xor ( n38216 , n38049 , n38050 );
xor ( n38217 , n38216 , n38052 );
and ( n38218 , n38214 , n38217 );
and ( n38219 , n38212 , n38217 );
or ( n38220 , n38215 , n38218 , n38219 );
and ( n38221 , n34480 , n31871 );
and ( n38222 , n33894 , n32320 );
and ( n38223 , n38221 , n38222 );
and ( n38224 , n33513 , n32508 );
and ( n38225 , n38222 , n38224 );
and ( n38226 , n38221 , n38224 );
or ( n38227 , n38223 , n38225 , n38226 );
xor ( n38228 , n38040 , n38041 );
xor ( n38229 , n38228 , n38043 );
and ( n38230 , n38227 , n38229 );
xor ( n38231 , n38056 , n38057 );
xor ( n38232 , n38231 , n38059 );
and ( n38233 , n38229 , n38232 );
and ( n38234 , n38227 , n38232 );
or ( n38235 , n38230 , n38233 , n38234 );
and ( n38236 , n38220 , n38235 );
and ( n38237 , n38204 , n38236 );
and ( n38238 , n38203 , n38236 );
or ( n38239 , n38205 , n38237 , n38238 );
and ( n38240 , n38200 , n38239 );
and ( n38241 , n38199 , n38239 );
or ( n38242 , n38201 , n38240 , n38241 );
and ( n38243 , n38197 , n38242 );
and ( n38244 , n38195 , n38242 );
or ( n38245 , n38198 , n38243 , n38244 );
xor ( n38246 , n38029 , n38031 );
xor ( n38247 , n38039 , n38046 );
and ( n38248 , n38246 , n38247 );
xor ( n38249 , n38055 , n38062 );
and ( n38250 , n38247 , n38249 );
and ( n38251 , n38246 , n38249 );
or ( n38252 , n38248 , n38250 , n38251 );
xor ( n38253 , n38169 , n38171 );
xor ( n38254 , n38177 , n38179 );
and ( n38255 , n38253 , n38254 );
xor ( n38256 , n38181 , n38182 );
and ( n38257 , n38254 , n38256 );
and ( n38258 , n38253 , n38256 );
or ( n38259 , n38255 , n38257 , n38258 );
and ( n38260 , n38252 , n38259 );
xor ( n38261 , n38165 , n38166 );
xor ( n38262 , n38261 , n38172 );
and ( n38263 , n38259 , n38262 );
and ( n38264 , n38252 , n38262 );
or ( n38265 , n38260 , n38263 , n38264 );
xor ( n38266 , n38081 , n38088 );
xor ( n38267 , n38266 , n38091 );
and ( n38268 , n38265 , n38267 );
xor ( n38269 , n38175 , n38189 );
xor ( n38270 , n38269 , n38192 );
and ( n38271 , n38267 , n38270 );
and ( n38272 , n38265 , n38270 );
or ( n38273 , n38268 , n38271 , n38272 );
xor ( n38274 , n38017 , n38018 );
xor ( n38275 , n38274 , n38020 );
and ( n38276 , n38273 , n38275 );
xor ( n38277 , n38072 , n38075 );
xor ( n38278 , n38277 , n38094 );
and ( n38279 , n38275 , n38278 );
and ( n38280 , n38273 , n38278 );
or ( n38281 , n38276 , n38279 , n38280 );
and ( n38282 , n38245 , n38281 );
xor ( n38283 , n38013 , n38014 );
xor ( n38284 , n38283 , n38023 );
and ( n38285 , n38281 , n38284 );
and ( n38286 , n38245 , n38284 );
or ( n38287 , n38282 , n38285 , n38286 );
and ( n38288 , n38164 , n38287 );
xor ( n38289 , n38026 , n38105 );
xor ( n38290 , n38289 , n38108 );
and ( n38291 , n38287 , n38290 );
and ( n38292 , n38164 , n38290 );
or ( n38293 , n38288 , n38291 , n38292 );
xor ( n38294 , n38011 , n38111 );
xor ( n38295 , n38294 , n38113 );
and ( n38296 , n38293 , n38295 );
xor ( n38297 , n38097 , n38099 );
xor ( n38298 , n38297 , n38102 );
xor ( n38299 , n38180 , n38183 );
xor ( n38300 , n38299 , n38186 );
and ( n38301 , n34315 , n31997 );
and ( n38302 , n33575 , n32850 );
and ( n38303 , n38301 , n38302 );
and ( n38304 , n33204 , n32922 );
and ( n38305 , n38302 , n38304 );
and ( n38306 , n38301 , n38304 );
or ( n38307 , n38303 , n38305 , n38306 );
and ( n38308 , n32019 , n34298 );
and ( n38309 , n32868 , n33532 );
and ( n38310 , n38308 , n38309 );
and ( n38311 , n32940 , n33213 );
and ( n38312 , n38309 , n38311 );
and ( n38313 , n38308 , n38311 );
or ( n38314 , n38310 , n38312 , n38313 );
and ( n38315 , n38307 , n38314 );
buf ( n38316 , n32940 );
buf ( n565618 , n543281 );
buf ( n38318 , n565618 );
and ( n38319 , n38316 , n38318 );
xor ( n38320 , n38027 , n38028 );
and ( n38321 , n38318 , n38320 );
and ( n38322 , n38316 , n38320 );
or ( n38323 , n38319 , n38321 , n38322 );
and ( n38324 , n38315 , n38323 );
xor ( n38325 , n38220 , n38235 );
and ( n38326 , n38323 , n38325 );
and ( n38327 , n38315 , n38325 );
or ( n38328 , n38324 , n38326 , n38327 );
and ( n38329 , n38300 , n38328 );
and ( n38330 , n32940 , n33532 );
and ( n38331 , n33575 , n32922 );
and ( n38332 , n38330 , n38331 );
buf ( n565634 , n543284 );
buf ( n38334 , n565634 );
and ( n38335 , n38332 , n38334 );
and ( n38336 , n32235 , n34032 );
and ( n38337 , n34049 , n32244 );
and ( n38338 , n38336 , n38337 );
or ( n38339 , n38335 , n38338 );
and ( n38340 , n32302 , n34032 );
and ( n38341 , n32525 , n33914 );
and ( n38342 , n38340 , n38341 );
and ( n38343 , n32868 , n33556 );
and ( n38344 , n38341 , n38343 );
and ( n38345 , n38340 , n38343 );
or ( n38346 , n38342 , n38344 , n38345 );
xor ( n38347 , n38221 , n38222 );
xor ( n38348 , n38347 , n38224 );
and ( n38349 , n38346 , n38348 );
xor ( n38350 , n38301 , n38302 );
xor ( n38351 , n38350 , n38304 );
and ( n38352 , n38348 , n38351 );
and ( n38353 , n38346 , n38351 );
or ( n38354 , n38349 , n38352 , n38353 );
and ( n38355 , n34049 , n32320 );
and ( n38356 , n33894 , n32508 );
and ( n38357 , n38355 , n38356 );
and ( n38358 , n33513 , n32850 );
and ( n38359 , n38356 , n38358 );
and ( n38360 , n38355 , n38358 );
or ( n38361 , n38357 , n38359 , n38360 );
xor ( n38362 , n38206 , n38207 );
xor ( n38363 , n38362 , n38209 );
and ( n38364 , n38361 , n38363 );
xor ( n38365 , n38308 , n38309 );
xor ( n38366 , n38365 , n38311 );
and ( n38367 , n38363 , n38366 );
and ( n38368 , n38361 , n38366 );
or ( n38369 , n38364 , n38367 , n38368 );
and ( n38370 , n38354 , n38369 );
and ( n38371 , n38339 , n38370 );
xor ( n38372 , n38212 , n38214 );
xor ( n38373 , n38372 , n38217 );
xor ( n38374 , n38227 , n38229 );
xor ( n38375 , n38374 , n38232 );
and ( n38376 , n38373 , n38375 );
and ( n38377 , n38370 , n38376 );
and ( n38378 , n38339 , n38376 );
or ( n38379 , n38371 , n38377 , n38378 );
and ( n38380 , n38328 , n38379 );
and ( n38381 , n38300 , n38379 );
or ( n38382 , n38329 , n38380 , n38381 );
xor ( n38383 , n38307 , n38314 );
and ( n38384 , n34480 , n31997 );
and ( n38385 , n34315 , n32244 );
or ( n38386 , n38384 , n38385 );
and ( n38387 , n32019 , n34453 );
and ( n38388 , n32235 , n34298 );
or ( n38389 , n38387 , n38388 );
and ( n38390 , n38386 , n38389 );
and ( n38391 , n38383 , n38390 );
xor ( n38392 , n38316 , n38318 );
xor ( n38393 , n38392 , n38320 );
and ( n38394 , n38390 , n38393 );
and ( n38395 , n38383 , n38393 );
or ( n38396 , n38391 , n38394 , n38395 );
xor ( n38397 , n38246 , n38247 );
xor ( n38398 , n38397 , n38249 );
and ( n38399 , n38396 , n38398 );
xor ( n38400 , n38253 , n38254 );
xor ( n38401 , n38400 , n38256 );
and ( n38402 , n38398 , n38401 );
and ( n38403 , n38396 , n38401 );
or ( n38404 , n38399 , n38402 , n38403 );
xor ( n38405 , n38203 , n38204 );
xor ( n38406 , n38405 , n38236 );
and ( n38407 , n38404 , n38406 );
xor ( n38408 , n38252 , n38259 );
xor ( n38409 , n38408 , n38262 );
and ( n38410 , n38406 , n38409 );
and ( n38411 , n38404 , n38409 );
or ( n38412 , n38407 , n38410 , n38411 );
and ( n38413 , n38382 , n38412 );
xor ( n38414 , n38199 , n38200 );
xor ( n38415 , n38414 , n38239 );
and ( n38416 , n38412 , n38415 );
and ( n38417 , n38382 , n38415 );
or ( n38418 , n38413 , n38416 , n38417 );
xor ( n38419 , n38195 , n38197 );
xor ( n38420 , n38419 , n38242 );
and ( n38421 , n38418 , n38420 );
xor ( n38422 , n38273 , n38275 );
xor ( n38423 , n38422 , n38278 );
and ( n38424 , n38420 , n38423 );
and ( n38425 , n38418 , n38423 );
or ( n38426 , n38421 , n38424 , n38425 );
and ( n38427 , n38298 , n38426 );
xor ( n38428 , n38245 , n38281 );
xor ( n38429 , n38428 , n38284 );
and ( n38430 , n38426 , n38429 );
and ( n38431 , n38298 , n38429 );
or ( n38432 , n38427 , n38430 , n38431 );
xor ( n38433 , n38164 , n38287 );
xor ( n38434 , n38433 , n38290 );
and ( n38435 , n38432 , n38434 );
xor ( n38436 , n38298 , n38426 );
xor ( n38437 , n38436 , n38429 );
xor ( n38438 , n38265 , n38267 );
xor ( n38439 , n38438 , n38270 );
xnor ( n38440 , n38335 , n38338 );
xor ( n38441 , n38354 , n38369 );
and ( n38442 , n38440 , n38441 );
xor ( n38443 , n38373 , n38375 );
and ( n38444 , n38441 , n38443 );
and ( n38445 , n38440 , n38443 );
or ( n38446 , n38442 , n38444 , n38445 );
buf ( n38447 , n33204 );
buf ( n565749 , n543287 );
buf ( n38449 , n565749 );
and ( n38450 , n38447 , n38449 );
xnor ( n38451 , n38384 , n38385 );
xnor ( n38452 , n38387 , n38388 );
and ( n38453 , n38451 , n38452 );
or ( n38454 , n38450 , n38453 );
and ( n38455 , n32302 , n34298 );
and ( n38456 , n32525 , n34032 );
and ( n38457 , n38455 , n38456 );
and ( n38458 , n32868 , n33914 );
and ( n38459 , n38456 , n38458 );
and ( n38460 , n38455 , n38458 );
or ( n38461 , n38457 , n38459 , n38460 );
and ( n38462 , n32235 , n34453 );
and ( n38463 , n32940 , n33556 );
and ( n38464 , n38462 , n38463 );
and ( n38465 , n33204 , n33532 );
and ( n38466 , n38463 , n38465 );
and ( n38467 , n38462 , n38465 );
or ( n38468 , n38464 , n38466 , n38467 );
and ( n38469 , n38461 , n38468 );
and ( n38470 , n34315 , n32320 );
and ( n38471 , n34049 , n32508 );
and ( n38472 , n38470 , n38471 );
and ( n38473 , n33894 , n32850 );
and ( n38474 , n38471 , n38473 );
and ( n38475 , n38470 , n38473 );
or ( n38476 , n38472 , n38474 , n38475 );
and ( n38477 , n34480 , n32244 );
and ( n38478 , n33513 , n32922 );
and ( n38479 , n38477 , n38478 );
and ( n38480 , n33575 , n33213 );
and ( n38481 , n38478 , n38480 );
and ( n38482 , n38477 , n38480 );
or ( n38483 , n38479 , n38481 , n38482 );
and ( n38484 , n38476 , n38483 );
and ( n38485 , n38469 , n38484 );
and ( n38486 , n38454 , n38485 );
xor ( n38487 , n38383 , n38390 );
xor ( n38488 , n38487 , n38393 );
and ( n38489 , n38485 , n38488 );
and ( n38490 , n38454 , n38488 );
or ( n38491 , n38486 , n38489 , n38490 );
and ( n38492 , n38446 , n38491 );
xor ( n38493 , n38315 , n38323 );
xor ( n38494 , n38493 , n38325 );
and ( n38495 , n38491 , n38494 );
and ( n38496 , n38446 , n38494 );
or ( n38497 , n38492 , n38495 , n38496 );
xor ( n38498 , n38300 , n38328 );
xor ( n38499 , n38498 , n38379 );
and ( n38500 , n38497 , n38499 );
xor ( n38501 , n38404 , n38406 );
xor ( n38502 , n38501 , n38409 );
and ( n38503 , n38499 , n38502 );
and ( n38504 , n38497 , n38502 );
or ( n38505 , n38500 , n38503 , n38504 );
and ( n38506 , n38439 , n38505 );
xor ( n38507 , n38382 , n38412 );
xor ( n38508 , n38507 , n38415 );
and ( n38509 , n38505 , n38508 );
and ( n38510 , n38439 , n38508 );
or ( n38511 , n38506 , n38509 , n38510 );
xor ( n38512 , n38418 , n38420 );
xor ( n38513 , n38512 , n38423 );
and ( n38514 , n38511 , n38513 );
xor ( n38515 , n38439 , n38505 );
xor ( n38516 , n38515 , n38508 );
xor ( n38517 , n38339 , n38370 );
xor ( n38518 , n38517 , n38376 );
xor ( n38519 , n38396 , n38398 );
xor ( n38520 , n38519 , n38401 );
and ( n38521 , n38518 , n38520 );
xnor ( n38522 , n38450 , n38453 );
xor ( n38523 , n38447 , n38449 );
and ( n38524 , n33204 , n33556 );
and ( n38525 , n33513 , n33213 );
and ( n38526 , n38524 , n38525 );
buf ( n565828 , n543290 );
buf ( n38528 , n565828 );
and ( n38529 , n38526 , n38528 );
and ( n38530 , n38523 , n38529 );
and ( n38531 , n34315 , n32508 );
and ( n38532 , n34049 , n32850 );
and ( n38533 , n38531 , n38532 );
and ( n38534 , n33894 , n32922 );
and ( n38535 , n38532 , n38534 );
and ( n38536 , n38531 , n38534 );
or ( n38537 , n38533 , n38535 , n38536 );
and ( n38538 , n32525 , n34298 );
and ( n38539 , n32868 , n34032 );
and ( n38540 , n38538 , n38539 );
and ( n38541 , n32940 , n33914 );
and ( n38542 , n38539 , n38541 );
and ( n38543 , n38538 , n38541 );
or ( n38544 , n38540 , n38542 , n38543 );
and ( n38545 , n38537 , n38544 );
and ( n38546 , n38529 , n38545 );
and ( n38547 , n38523 , n38545 );
or ( n38548 , n38530 , n38546 , n38547 );
and ( n38549 , n38522 , n38548 );
xor ( n38550 , n38355 , n38356 );
xor ( n38551 , n38550 , n38358 );
xor ( n38552 , n38340 , n38341 );
xor ( n38553 , n38552 , n38343 );
and ( n38554 , n38551 , n38553 );
and ( n38555 , n38548 , n38554 );
and ( n38556 , n38522 , n38554 );
or ( n38557 , n38549 , n38555 , n38556 );
xor ( n38558 , n38346 , n38348 );
xor ( n38559 , n38558 , n38351 );
xor ( n38560 , n38361 , n38363 );
xor ( n38561 , n38560 , n38366 );
and ( n38562 , n38559 , n38561 );
and ( n38563 , n38557 , n38562 );
and ( n38564 , n38520 , n38563 );
and ( n38565 , n38518 , n38563 );
or ( n38566 , n38521 , n38564 , n38565 );
xor ( n38567 , n38497 , n38499 );
xor ( n38568 , n38567 , n38502 );
and ( n38569 , n38566 , n38568 );
xor ( n38570 , n38461 , n38468 );
xor ( n38571 , n38476 , n38483 );
and ( n38572 , n38570 , n38571 );
xor ( n38573 , n38332 , n38334 );
and ( n38574 , n38572 , n38573 );
xor ( n38575 , n38336 , n38337 );
xor ( n38576 , n38386 , n38389 );
and ( n38577 , n38575 , n38576 );
xor ( n38578 , n38469 , n38484 );
and ( n38579 , n38576 , n38578 );
and ( n38580 , n38575 , n38578 );
or ( n38581 , n38577 , n38579 , n38580 );
and ( n38582 , n38574 , n38581 );
xor ( n38583 , n38559 , n38561 );
xor ( n38584 , n38455 , n38456 );
xor ( n38585 , n38584 , n38458 );
xor ( n38586 , n38462 , n38463 );
xor ( n38587 , n38586 , n38465 );
or ( n38588 , n38585 , n38587 );
xor ( n38589 , n38470 , n38471 );
xor ( n38590 , n38589 , n38473 );
xor ( n38591 , n38477 , n38478 );
xor ( n38592 , n38591 , n38480 );
or ( n38593 , n38590 , n38592 );
and ( n38594 , n38588 , n38593 );
and ( n38595 , n38583 , n38594 );
xor ( n38596 , n38330 , n38331 );
xor ( n38597 , n38551 , n38553 );
and ( n38598 , n38596 , n38597 );
xor ( n38599 , n38451 , n38452 );
and ( n38600 , n38597 , n38599 );
and ( n38601 , n38596 , n38599 );
or ( n38602 , n38598 , n38600 , n38601 );
and ( n38603 , n38594 , n38602 );
and ( n38604 , n38583 , n38602 );
or ( n38605 , n38595 , n38603 , n38604 );
and ( n38606 , n38581 , n38605 );
and ( n38607 , n38574 , n38605 );
or ( n38608 , n38582 , n38606 , n38607 );
xor ( n38609 , n38446 , n38491 );
xor ( n38610 , n38609 , n38494 );
and ( n38611 , n38608 , n38610 );
xor ( n38612 , n38440 , n38441 );
xor ( n38613 , n38612 , n38443 );
xor ( n38614 , n38454 , n38485 );
xor ( n38615 , n38614 , n38488 );
and ( n38616 , n38613 , n38615 );
xor ( n38617 , n38557 , n38562 );
and ( n38618 , n38615 , n38617 );
and ( n38619 , n38613 , n38617 );
or ( n38620 , n38616 , n38618 , n38619 );
and ( n38621 , n38610 , n38620 );
and ( n38622 , n38608 , n38620 );
or ( n38623 , n38611 , n38621 , n38622 );
and ( n38624 , n38568 , n38623 );
and ( n38625 , n38566 , n38623 );
or ( n38626 , n38569 , n38624 , n38625 );
and ( n38627 , n38516 , n38626 );
xor ( n38628 , n38522 , n38548 );
xor ( n38629 , n38628 , n38554 );
xor ( n38630 , n38572 , n38573 );
and ( n38631 , n38629 , n38630 );
xor ( n38632 , n38523 , n38529 );
xor ( n38633 , n38632 , n38545 );
xor ( n38634 , n38588 , n38593 );
and ( n38635 , n38633 , n38634 );
xor ( n38636 , n38570 , n38571 );
and ( n38637 , n38634 , n38636 );
and ( n38638 , n38633 , n38636 );
or ( n38639 , n38635 , n38637 , n38638 );
and ( n38640 , n38630 , n38639 );
and ( n38641 , n38629 , n38639 );
or ( n38642 , n38631 , n38640 , n38641 );
xor ( n38643 , n38526 , n38528 );
buf ( n38644 , n33575 );
buf ( n565946 , n543293 );
buf ( n38646 , n565946 );
and ( n38647 , n38644 , n38646 );
and ( n38648 , n38643 , n38647 );
and ( n38649 , n32302 , n34453 );
and ( n38650 , n34480 , n32320 );
and ( n38651 , n38649 , n38650 );
and ( n38652 , n38647 , n38651 );
and ( n38653 , n38643 , n38651 );
or ( n38654 , n38648 , n38652 , n38653 );
and ( n38655 , n32940 , n34032 );
and ( n38656 , n33204 , n33914 );
and ( n38657 , n38655 , n38656 );
and ( n38658 , n33575 , n33556 );
and ( n38659 , n38656 , n38658 );
and ( n38660 , n38655 , n38658 );
or ( n38661 , n38657 , n38659 , n38660 );
xor ( n38662 , n38538 , n38539 );
xor ( n38663 , n38662 , n38541 );
and ( n38664 , n38661 , n38663 );
and ( n38665 , n34049 , n32922 );
and ( n38666 , n33894 , n33213 );
and ( n38667 , n38665 , n38666 );
and ( n38668 , n33513 , n33532 );
and ( n38669 , n38666 , n38668 );
and ( n38670 , n38665 , n38668 );
or ( n38671 , n38667 , n38669 , n38670 );
xor ( n38672 , n38531 , n38532 );
xor ( n38673 , n38672 , n38534 );
and ( n38674 , n38671 , n38673 );
and ( n38675 , n38664 , n38674 );
and ( n38676 , n38654 , n38675 );
xnor ( n38677 , n38585 , n38587 );
xnor ( n38678 , n38590 , n38592 );
and ( n38679 , n38677 , n38678 );
and ( n38680 , n38675 , n38679 );
and ( n38681 , n38654 , n38679 );
or ( n38682 , n38676 , n38680 , n38681 );
xor ( n38683 , n38575 , n38576 );
xor ( n38684 , n38683 , n38578 );
and ( n38685 , n38682 , n38684 );
xor ( n38686 , n38583 , n38594 );
xor ( n38687 , n38686 , n38602 );
and ( n38688 , n38684 , n38687 );
and ( n38689 , n38682 , n38687 );
or ( n38690 , n38685 , n38688 , n38689 );
and ( n38691 , n38642 , n38690 );
xor ( n38692 , n38574 , n38581 );
xor ( n38693 , n38692 , n38605 );
and ( n38694 , n38690 , n38693 );
and ( n38695 , n38642 , n38693 );
or ( n38696 , n38691 , n38694 , n38695 );
xor ( n38697 , n38518 , n38520 );
xor ( n38698 , n38697 , n38563 );
and ( n38699 , n38696 , n38698 );
xor ( n38700 , n38596 , n38597 );
xor ( n38701 , n38700 , n38599 );
xor ( n38702 , n38537 , n38544 );
and ( n38703 , n34480 , n32508 );
and ( n38704 , n34315 , n32850 );
and ( n38705 , n38703 , n38704 );
and ( n38706 , n32525 , n34453 );
and ( n38707 , n32868 , n34298 );
and ( n38708 , n38706 , n38707 );
and ( n38709 , n38705 , n38708 );
and ( n38710 , n38702 , n38709 );
xor ( n38711 , n38664 , n38674 );
and ( n38712 , n38709 , n38711 );
and ( n38713 , n38702 , n38711 );
or ( n38714 , n38710 , n38712 , n38713 );
and ( n38715 , n38701 , n38714 );
xor ( n38716 , n38677 , n38678 );
xor ( n38717 , n38703 , n38704 );
xor ( n38718 , n38706 , n38707 );
and ( n38719 , n38717 , n38718 );
xor ( n38720 , n38644 , n38646 );
and ( n38721 , n38719 , n38720 );
and ( n38722 , n38716 , n38721 );
xor ( n38723 , n38661 , n38663 );
xor ( n38724 , n38671 , n38673 );
and ( n38725 , n38723 , n38724 );
and ( n38726 , n38721 , n38725 );
and ( n38727 , n38716 , n38725 );
or ( n38728 , n38722 , n38726 , n38727 );
and ( n38729 , n38714 , n38728 );
and ( n38730 , n38701 , n38728 );
or ( n38731 , n38715 , n38729 , n38730 );
xor ( n38732 , n38629 , n38630 );
xor ( n38733 , n38732 , n38639 );
and ( n38734 , n38731 , n38733 );
xor ( n38735 , n38682 , n38684 );
xor ( n38736 , n38735 , n38687 );
and ( n38737 , n38733 , n38736 );
and ( n38738 , n38731 , n38736 );
or ( n38739 , n38734 , n38737 , n38738 );
xor ( n38740 , n38613 , n38615 );
xor ( n38741 , n38740 , n38617 );
and ( n38742 , n38739 , n38741 );
xor ( n38743 , n38642 , n38690 );
xor ( n38744 , n38743 , n38693 );
and ( n38745 , n38741 , n38744 );
and ( n38746 , n38739 , n38744 );
or ( n38747 , n38742 , n38745 , n38746 );
and ( n38748 , n38698 , n38747 );
and ( n38749 , n38696 , n38747 );
or ( n38750 , n38699 , n38748 , n38749 );
xor ( n38751 , n38566 , n38568 );
xor ( n38752 , n38751 , n38623 );
and ( n38753 , n38750 , n38752 );
xor ( n38754 , n38608 , n38610 );
xor ( n38755 , n38754 , n38620 );
xor ( n38756 , n38696 , n38698 );
xor ( n38757 , n38756 , n38747 );
and ( n38758 , n38755 , n38757 );
xor ( n38759 , n38739 , n38741 );
xor ( n38760 , n38759 , n38744 );
xor ( n38761 , n38633 , n38634 );
xor ( n38762 , n38761 , n38636 );
xor ( n38763 , n38654 , n38675 );
xor ( n38764 , n38763 , n38679 );
and ( n38765 , n38762 , n38764 );
xor ( n38766 , n38719 , n38720 );
and ( n38767 , n33575 , n33914 );
and ( n38768 , n33894 , n33532 );
and ( n38769 , n38767 , n38768 );
buf ( n566071 , n543296 );
buf ( n38771 , n566071 );
and ( n38772 , n38769 , n38771 );
and ( n38773 , n38766 , n38772 );
and ( n38774 , n34480 , n32850 );
and ( n38775 , n34315 , n32922 );
and ( n38776 , n38774 , n38775 );
and ( n38777 , n34049 , n33213 );
and ( n38778 , n38775 , n38777 );
and ( n38779 , n38774 , n38777 );
or ( n38780 , n38776 , n38778 , n38779 );
and ( n38781 , n32868 , n34453 );
and ( n38782 , n32940 , n34298 );
and ( n38783 , n38781 , n38782 );
and ( n38784 , n33204 , n34032 );
and ( n38785 , n38782 , n38784 );
and ( n38786 , n38781 , n38784 );
or ( n38787 , n38783 , n38785 , n38786 );
and ( n38788 , n38780 , n38787 );
and ( n38789 , n38772 , n38788 );
and ( n38790 , n38766 , n38788 );
or ( n38791 , n38773 , n38789 , n38790 );
xor ( n38792 , n38643 , n38647 );
xor ( n38793 , n38792 , n38651 );
and ( n38794 , n38791 , n38793 );
and ( n38795 , n38764 , n38794 );
and ( n38796 , n38762 , n38794 );
or ( n38797 , n38765 , n38795 , n38796 );
xor ( n38798 , n38731 , n38733 );
xor ( n38799 , n38798 , n38736 );
and ( n38800 , n38797 , n38799 );
xor ( n38801 , n38649 , n38650 );
xor ( n38802 , n38524 , n38525 );
and ( n38803 , n38801 , n38802 );
xor ( n38804 , n38705 , n38708 );
and ( n38805 , n38802 , n38804 );
and ( n38806 , n38801 , n38804 );
or ( n38807 , n38803 , n38805 , n38806 );
xor ( n38808 , n38723 , n38724 );
xor ( n38809 , n38780 , n38787 );
xor ( n38810 , n38665 , n38666 );
xor ( n38811 , n38810 , n38668 );
xor ( n38812 , n38655 , n38656 );
xor ( n38813 , n38812 , n38658 );
xor ( n38814 , n38811 , n38813 );
and ( n38815 , n38809 , n38814 );
xor ( n38816 , n38717 , n38718 );
and ( n38817 , n38814 , n38816 );
and ( n38818 , n38809 , n38816 );
or ( n38819 , n38815 , n38817 , n38818 );
and ( n38820 , n38808 , n38819 );
xor ( n38821 , n38801 , n38802 );
xor ( n38822 , n38821 , n38804 );
and ( n38823 , n38819 , n38822 );
and ( n38824 , n38808 , n38822 );
or ( n38825 , n38820 , n38823 , n38824 );
and ( n38826 , n38807 , n38825 );
xor ( n38827 , n38702 , n38709 );
xor ( n38828 , n38827 , n38711 );
and ( n38829 , n38825 , n38828 );
and ( n38830 , n38807 , n38828 );
or ( n38831 , n38826 , n38829 , n38830 );
xor ( n38832 , n38701 , n38714 );
xor ( n38833 , n38832 , n38728 );
and ( n38834 , n38831 , n38833 );
xor ( n38835 , n38716 , n38721 );
xor ( n38836 , n38835 , n38725 );
xor ( n38837 , n38791 , n38793 );
and ( n38838 , n38836 , n38837 );
xor ( n38839 , n38769 , n38771 );
buf ( n38840 , n33513 );
buf ( n566142 , n543299 );
buf ( n38842 , n566142 );
and ( n38843 , n38840 , n38842 );
and ( n38844 , n38839 , n38843 );
and ( n38845 , n34315 , n33213 );
and ( n38846 , n34049 , n33532 );
and ( n38847 , n38845 , n38846 );
and ( n38848 , n33894 , n33556 );
and ( n38849 , n38846 , n38848 );
and ( n38850 , n38845 , n38848 );
or ( n38851 , n38847 , n38849 , n38850 );
and ( n38852 , n33204 , n34298 );
and ( n38853 , n33575 , n34032 );
and ( n38854 , n38852 , n38853 );
and ( n38855 , n33513 , n33914 );
and ( n38856 , n38853 , n38855 );
and ( n38857 , n38852 , n38855 );
or ( n38858 , n38854 , n38856 , n38857 );
and ( n38859 , n38851 , n38858 );
and ( n38860 , n38843 , n38859 );
and ( n38861 , n38839 , n38859 );
or ( n38862 , n38844 , n38860 , n38861 );
and ( n38863 , n38811 , n38813 );
and ( n38864 , n38862 , n38863 );
xor ( n38865 , n38766 , n38772 );
xor ( n38866 , n38865 , n38788 );
and ( n38867 , n38863 , n38866 );
and ( n38868 , n38862 , n38866 );
or ( n38869 , n38864 , n38867 , n38868 );
and ( n38870 , n38837 , n38869 );
and ( n38871 , n38836 , n38869 );
or ( n38872 , n38838 , n38870 , n38871 );
and ( n38873 , n38833 , n38872 );
and ( n38874 , n38831 , n38872 );
or ( n38875 , n38834 , n38873 , n38874 );
and ( n38876 , n38799 , n38875 );
and ( n38877 , n38797 , n38875 );
or ( n38878 , n38800 , n38876 , n38877 );
and ( n38879 , n38760 , n38878 );
xor ( n38880 , n38762 , n38764 );
xor ( n38881 , n38880 , n38794 );
xor ( n38882 , n38807 , n38825 );
xor ( n38883 , n38882 , n38828 );
xor ( n38884 , n38840 , n38842 );
and ( n38885 , n33513 , n34032 );
and ( n38886 , n34049 , n33556 );
and ( n38887 , n38885 , n38886 );
buf ( n566189 , n543302 );
buf ( n38889 , n566189 );
and ( n38890 , n38887 , n38889 );
and ( n38891 , n38884 , n38890 );
and ( n38892 , n32940 , n34453 );
and ( n38893 , n34480 , n32922 );
and ( n38894 , n38892 , n38893 );
and ( n38895 , n38890 , n38894 );
and ( n38896 , n38884 , n38894 );
or ( n38897 , n38891 , n38895 , n38896 );
xor ( n38898 , n38774 , n38775 );
xor ( n38899 , n38898 , n38777 );
xor ( n38900 , n38781 , n38782 );
xor ( n38901 , n38900 , n38784 );
and ( n38902 , n38899 , n38901 );
and ( n38903 , n38897 , n38902 );
xor ( n38904 , n38839 , n38843 );
xor ( n38905 , n38904 , n38859 );
and ( n38906 , n38902 , n38905 );
and ( n38907 , n38897 , n38905 );
or ( n38908 , n38903 , n38906 , n38907 );
xor ( n38909 , n38862 , n38863 );
xor ( n38910 , n38909 , n38866 );
or ( n38911 , n38908 , n38910 );
and ( n38912 , n38883 , n38911 );
xor ( n38913 , n38836 , n38837 );
xor ( n38914 , n38913 , n38869 );
and ( n38915 , n38911 , n38914 );
and ( n38916 , n38883 , n38914 );
or ( n38917 , n38912 , n38915 , n38916 );
and ( n38918 , n38881 , n38917 );
xor ( n38919 , n38831 , n38833 );
xor ( n38920 , n38919 , n38872 );
and ( n38921 , n38917 , n38920 );
and ( n38922 , n38881 , n38920 );
or ( n38923 , n38918 , n38921 , n38922 );
xor ( n38924 , n38797 , n38799 );
xor ( n38925 , n38924 , n38875 );
or ( n38926 , n38923 , n38925 );
and ( n38927 , n38878 , n38926 );
and ( n38928 , n38760 , n38926 );
or ( n38929 , n38879 , n38927 , n38928 );
and ( n38930 , n38757 , n38929 );
and ( n38931 , n38755 , n38929 );
or ( n38932 , n38758 , n38930 , n38931 );
and ( n38933 , n38752 , n38932 );
and ( n38934 , n38750 , n38932 );
or ( n38935 , n38753 , n38933 , n38934 );
and ( n38936 , n38626 , n38935 );
and ( n38937 , n38516 , n38935 );
or ( n38938 , n38627 , n38936 , n38937 );
and ( n38939 , n38513 , n38938 );
and ( n38940 , n38511 , n38938 );
or ( n38941 , n38514 , n38939 , n38940 );
or ( n38942 , n38437 , n38941 );
and ( n38943 , n38434 , n38942 );
and ( n38944 , n38432 , n38942 );
or ( n38945 , n38435 , n38943 , n38944 );
and ( n38946 , n38295 , n38945 );
and ( n38947 , n38293 , n38945 );
or ( n38948 , n38296 , n38946 , n38947 );
or ( n38949 , n38162 , n38948 );
or ( n38950 , n38160 , n38949 );
and ( n38951 , n38158 , n38950 );
xor ( n38952 , n38158 , n38950 );
xnor ( n38953 , n38160 , n38949 );
xnor ( n38954 , n38162 , n38948 );
xor ( n38955 , n38293 , n38295 );
xor ( n38956 , n38955 , n38945 );
xor ( n38957 , n38432 , n38434 );
xor ( n38958 , n38957 , n38942 );
not ( n38959 , n38958 );
xnor ( n38960 , n38437 , n38941 );
xor ( n38961 , n38511 , n38513 );
xor ( n38962 , n38961 , n38938 );
xor ( n38963 , n38516 , n38626 );
xor ( n38964 , n38963 , n38935 );
xor ( n38965 , n38750 , n38752 );
xor ( n38966 , n38965 , n38932 );
xor ( n38967 , n38755 , n38757 );
xor ( n38968 , n38967 , n38929 );
xor ( n38969 , n38760 , n38878 );
xor ( n38970 , n38969 , n38926 );
not ( n38971 , n38970 );
xnor ( n38972 , n38923 , n38925 );
xor ( n38973 , n38881 , n38917 );
xor ( n38974 , n38973 , n38920 );
xor ( n38975 , n38808 , n38819 );
xor ( n38976 , n38975 , n38822 );
xor ( n38977 , n38767 , n38768 );
xor ( n38978 , n38851 , n38858 );
and ( n38979 , n38977 , n38978 );
xor ( n38980 , n38899 , n38901 );
and ( n38981 , n38978 , n38980 );
and ( n38982 , n38977 , n38980 );
or ( n38983 , n38979 , n38981 , n38982 );
xor ( n38984 , n38809 , n38814 );
xor ( n38985 , n38984 , n38816 );
and ( n38986 , n38983 , n38985 );
xor ( n38987 , n38897 , n38902 );
xor ( n38988 , n38987 , n38905 );
and ( n38989 , n38985 , n38988 );
and ( n38990 , n38983 , n38988 );
or ( n38991 , n38986 , n38989 , n38990 );
and ( n38992 , n38976 , n38991 );
xnor ( n38993 , n38908 , n38910 );
and ( n38994 , n38991 , n38993 );
and ( n38995 , n38976 , n38993 );
or ( n38996 , n38992 , n38994 , n38995 );
xor ( n38997 , n38883 , n38911 );
xor ( n38998 , n38997 , n38914 );
and ( n38999 , n38996 , n38998 );
and ( n39000 , n34480 , n33213 );
and ( n39001 , n34315 , n33532 );
or ( n39002 , n39000 , n39001 );
and ( n39003 , n33204 , n34453 );
and ( n39004 , n33575 , n34298 );
or ( n39005 , n39003 , n39004 );
and ( n39006 , n39002 , n39005 );
xor ( n39007 , n38845 , n38846 );
xor ( n39008 , n39007 , n38848 );
xor ( n39009 , n38852 , n38853 );
xor ( n39010 , n39009 , n38855 );
and ( n39011 , n39008 , n39010 );
and ( n39012 , n39006 , n39011 );
xor ( n39013 , n38884 , n38890 );
xor ( n39014 , n39013 , n38894 );
and ( n39015 , n39011 , n39014 );
and ( n39016 , n39006 , n39014 );
or ( n39017 , n39012 , n39015 , n39016 );
buf ( n39018 , n33894 );
buf ( n566320 , n543305 );
buf ( n39020 , n566320 );
and ( n39021 , n39018 , n39020 );
xnor ( n39022 , n39000 , n39001 );
xnor ( n39023 , n39003 , n39004 );
and ( n39024 , n39022 , n39023 );
or ( n39025 , n39021 , n39024 );
xor ( n39026 , n38892 , n38893 );
xor ( n39027 , n39002 , n39005 );
and ( n39028 , n39026 , n39027 );
xor ( n39029 , n39008 , n39010 );
and ( n39030 , n39027 , n39029 );
and ( n39031 , n39026 , n39029 );
or ( n39032 , n39028 , n39030 , n39031 );
and ( n39033 , n39025 , n39032 );
xor ( n39034 , n38977 , n38978 );
xor ( n39035 , n39034 , n38980 );
and ( n39036 , n39032 , n39035 );
and ( n39037 , n39025 , n39035 );
or ( n39038 , n39033 , n39036 , n39037 );
and ( n39039 , n39017 , n39038 );
xor ( n39040 , n38887 , n38889 );
and ( n39041 , n34480 , n33532 );
and ( n39042 , n34315 , n33556 );
and ( n39043 , n39041 , n39042 );
and ( n39044 , n34049 , n33914 );
and ( n39045 , n39042 , n39044 );
and ( n39046 , n39041 , n39044 );
or ( n39047 , n39043 , n39045 , n39046 );
and ( n39048 , n33575 , n34453 );
and ( n39049 , n33513 , n34298 );
and ( n39050 , n39048 , n39049 );
and ( n39051 , n33894 , n34032 );
and ( n39052 , n39049 , n39051 );
and ( n39053 , n39048 , n39051 );
or ( n39054 , n39050 , n39052 , n39053 );
and ( n39055 , n39047 , n39054 );
and ( n39056 , n39040 , n39055 );
xnor ( n39057 , n39021 , n39024 );
and ( n39058 , n39055 , n39057 );
and ( n39059 , n39040 , n39057 );
or ( n39060 , n39056 , n39058 , n39059 );
xor ( n39061 , n39006 , n39011 );
xor ( n39062 , n39061 , n39014 );
and ( n39063 , n39060 , n39062 );
xor ( n39064 , n39025 , n39032 );
xor ( n39065 , n39064 , n39035 );
and ( n39066 , n39062 , n39065 );
and ( n39067 , n39060 , n39065 );
or ( n39068 , n39063 , n39066 , n39067 );
and ( n39069 , n39038 , n39068 );
and ( n39070 , n39017 , n39068 );
or ( n39071 , n39039 , n39069 , n39070 );
xor ( n39072 , n38983 , n38985 );
xor ( n39073 , n39072 , n38988 );
xor ( n39074 , n39018 , n39020 );
and ( n39075 , n33894 , n34298 );
and ( n39076 , n34315 , n33914 );
and ( n39077 , n39075 , n39076 );
buf ( n566379 , n543308 );
buf ( n39079 , n566379 );
and ( n39080 , n39077 , n39079 );
and ( n39081 , n39074 , n39080 );
xor ( n39082 , n39041 , n39042 );
xor ( n39083 , n39082 , n39044 );
xor ( n39084 , n39048 , n39049 );
xor ( n39085 , n39084 , n39051 );
and ( n39086 , n39083 , n39085 );
and ( n39087 , n39080 , n39086 );
and ( n39088 , n39074 , n39086 );
or ( n39089 , n39081 , n39087 , n39088 );
xor ( n39090 , n39040 , n39055 );
xor ( n39091 , n39090 , n39057 );
or ( n39092 , n39089 , n39091 );
xor ( n39093 , n38885 , n38886 );
xor ( n39094 , n39047 , n39054 );
and ( n39095 , n39093 , n39094 );
xor ( n39096 , n39022 , n39023 );
and ( n39097 , n39094 , n39096 );
and ( n39098 , n39093 , n39096 );
or ( n39099 , n39095 , n39097 , n39098 );
xor ( n39100 , n39026 , n39027 );
xor ( n39101 , n39100 , n39029 );
and ( n39102 , n39099 , n39101 );
xor ( n39103 , n39077 , n39079 );
buf ( n39104 , n34049 );
buf ( n566406 , n543311 );
buf ( n39106 , n566406 );
and ( n39107 , n39104 , n39106 );
and ( n39108 , n39103 , n39107 );
and ( n39109 , n33513 , n34453 );
and ( n39110 , n34480 , n33556 );
and ( n39111 , n39109 , n39110 );
and ( n39112 , n39107 , n39111 );
and ( n39113 , n39103 , n39111 );
or ( n39114 , n39108 , n39112 , n39113 );
xor ( n39115 , n39074 , n39080 );
xor ( n39116 , n39115 , n39086 );
or ( n39117 , n39114 , n39116 );
and ( n39118 , n39101 , n39117 );
and ( n39119 , n39099 , n39117 );
or ( n39120 , n39102 , n39118 , n39119 );
and ( n39121 , n39092 , n39120 );
xor ( n39122 , n39060 , n39062 );
xor ( n39123 , n39122 , n39065 );
and ( n39124 , n39120 , n39123 );
and ( n39125 , n39092 , n39123 );
or ( n39126 , n39121 , n39124 , n39125 );
or ( n39127 , n39073 , n39126 );
and ( n39128 , n39071 , n39127 );
xor ( n39129 , n38976 , n38991 );
xor ( n39130 , n39129 , n38993 );
and ( n39131 , n39127 , n39130 );
and ( n39132 , n39071 , n39130 );
or ( n39133 , n39128 , n39131 , n39132 );
and ( n39134 , n38998 , n39133 );
and ( n39135 , n38996 , n39133 );
or ( n39136 , n38999 , n39134 , n39135 );
and ( n39137 , n38974 , n39136 );
xor ( n39138 , n38974 , n39136 );
xor ( n39139 , n38996 , n38998 );
xor ( n39140 , n39139 , n39133 );
not ( n39141 , n39140 );
xor ( n39142 , n39071 , n39127 );
xor ( n39143 , n39142 , n39130 );
xor ( n39144 , n39017 , n39038 );
xor ( n39145 , n39144 , n39068 );
xnor ( n39146 , n39073 , n39126 );
and ( n39147 , n39145 , n39146 );
xor ( n39148 , n39145 , n39146 );
xnor ( n39149 , n39089 , n39091 );
xor ( n39150 , n39093 , n39094 );
xor ( n39151 , n39150 , n39096 );
xnor ( n39152 , n39114 , n39116 );
and ( n39153 , n39151 , n39152 );
xor ( n39154 , n39083 , n39085 );
and ( n39155 , n34480 , n33914 );
and ( n39156 , n34315 , n34032 );
or ( n39157 , n39155 , n39156 );
and ( n39158 , n33894 , n34453 );
and ( n39159 , n34049 , n34298 );
or ( n39160 , n39158 , n39159 );
and ( n39161 , n39157 , n39160 );
and ( n39162 , n39154 , n39161 );
xor ( n39163 , n39103 , n39107 );
xor ( n39164 , n39163 , n39111 );
and ( n39165 , n39161 , n39164 );
and ( n39166 , n39154 , n39164 );
or ( n39167 , n39162 , n39165 , n39166 );
and ( n39168 , n39152 , n39167 );
and ( n39169 , n39151 , n39167 );
or ( n39170 , n39153 , n39168 , n39169 );
and ( n39171 , n39149 , n39170 );
xor ( n39172 , n39099 , n39101 );
xor ( n39173 , n39172 , n39117 );
and ( n39174 , n39170 , n39173 );
and ( n39175 , n39149 , n39173 );
or ( n39176 , n39171 , n39174 , n39175 );
xor ( n39177 , n39092 , n39120 );
xor ( n39178 , n39177 , n39123 );
and ( n39179 , n39176 , n39178 );
xor ( n39180 , n39176 , n39178 );
xor ( n39181 , n39149 , n39170 );
xor ( n39182 , n39181 , n39173 );
xnor ( n39183 , n39155 , n39156 );
xnor ( n39184 , n39158 , n39159 );
and ( n39185 , n39183 , n39184 );
xor ( n39186 , n39104 , n39106 );
or ( n39187 , n39185 , n39186 );
xor ( n39188 , n39109 , n39110 );
xor ( n39189 , n39075 , n39076 );
and ( n39190 , n39188 , n39189 );
xor ( n39191 , n39157 , n39160 );
and ( n39192 , n39189 , n39191 );
and ( n39193 , n39188 , n39191 );
or ( n39194 , n39190 , n39192 , n39193 );
and ( n39195 , n39187 , n39194 );
and ( n39196 , n34049 , n34453 );
and ( n39197 , n34480 , n34032 );
and ( n39198 , n39196 , n39197 );
buf ( n566500 , n543314 );
buf ( n39200 , n566500 );
and ( n39201 , n39198 , n39200 );
xnor ( n39202 , n39185 , n39186 );
or ( n39203 , n39201 , n39202 );
and ( n39204 , n39194 , n39203 );
and ( n39205 , n39187 , n39203 );
or ( n39206 , n39195 , n39204 , n39205 );
xor ( n39207 , n39151 , n39152 );
xor ( n39208 , n39207 , n39167 );
and ( n39209 , n39206 , n39208 );
xor ( n39210 , n39154 , n39161 );
xor ( n39211 , n39210 , n39164 );
buf ( n39212 , n34315 );
buf ( n566514 , n543317 );
buf ( n39214 , n566514 );
and ( n39215 , n39212 , n39214 );
xor ( n39216 , n39198 , n39200 );
and ( n39217 , n39215 , n39216 );
xor ( n39218 , n39183 , n39184 );
and ( n39219 , n39216 , n39218 );
and ( n39220 , n39215 , n39218 );
or ( n39221 , n39217 , n39219 , n39220 );
xor ( n39222 , n39188 , n39189 );
xor ( n39223 , n39222 , n39191 );
and ( n39224 , n39221 , n39223 );
xnor ( n39225 , n39201 , n39202 );
and ( n39226 , n39223 , n39225 );
and ( n39227 , n39221 , n39225 );
or ( n39228 , n39224 , n39226 , n39227 );
and ( n39229 , n39211 , n39228 );
xor ( n39230 , n39187 , n39194 );
xor ( n39231 , n39230 , n39203 );
and ( n39232 , n39228 , n39231 );
and ( n39233 , n39211 , n39231 );
or ( n39234 , n39229 , n39232 , n39233 );
and ( n39235 , n39208 , n39234 );
and ( n39236 , n39206 , n39234 );
or ( n39237 , n39209 , n39235 , n39236 );
and ( n39238 , n39182 , n39237 );
xor ( n39239 , n39182 , n39237 );
xor ( n39240 , n39206 , n39208 );
xor ( n39241 , n39240 , n39234 );
xor ( n39242 , n39211 , n39228 );
xor ( n39243 , n39242 , n39231 );
and ( n39244 , n34315 , n34453 );
and ( n39245 , n34480 , n34298 );
and ( n39246 , n39244 , n39245 );
xor ( n39247 , n39212 , n39214 );
or ( n39248 , n39246 , n39247 );
xor ( n39249 , n39196 , n39197 );
xnor ( n39250 , n39246 , n39247 );
or ( n39251 , n39249 , n39250 );
or ( n39252 , n39248 , n39251 );
xor ( n39253 , n39221 , n39223 );
xor ( n39254 , n39253 , n39225 );
and ( n39255 , n39252 , n39254 );
xor ( n39256 , n39252 , n39254 );
xor ( n39257 , n39215 , n39216 );
xor ( n39258 , n39257 , n39218 );
xnor ( n39259 , n39248 , n39251 );
and ( n39260 , n39258 , n39259 );
xor ( n39261 , n39258 , n39259 );
xnor ( n39262 , n39249 , n39250 );
buf ( n566564 , n543320 );
buf ( n39264 , n566564 );
xor ( n39265 , n39244 , n39245 );
and ( n39266 , n39264 , n39265 );
xor ( n39267 , n39264 , n39265 );
buf ( n39268 , n34480 );
buf ( n566570 , n543323 );
buf ( n39270 , n566570 );
and ( n39271 , n39268 , n39270 );
and ( n39272 , n39267 , n39271 );
or ( n39273 , n39266 , n39272 );
and ( n39274 , n39262 , n39273 );
and ( n39275 , n39261 , n39274 );
or ( n39276 , n39260 , n39275 );
and ( n39277 , n39256 , n39276 );
or ( n39278 , n39255 , n39277 );
and ( n39279 , n39243 , n39278 );
and ( n39280 , n39241 , n39279 );
and ( n39281 , n39239 , n39280 );
or ( n39282 , n39238 , n39281 );
and ( n39283 , n39180 , n39282 );
or ( n39284 , n39179 , n39283 );
and ( n39285 , n39148 , n39284 );
or ( n39286 , n39147 , n39285 );
and ( n39287 , n39143 , n39286 );
and ( n39288 , n39141 , n39287 );
or ( n39289 , n39140 , n39288 );
and ( n39290 , n39138 , n39289 );
or ( n39291 , n39137 , n39290 );
and ( n39292 , n38972 , n39291 );
and ( n39293 , n38971 , n39292 );
or ( n39294 , n38970 , n39293 );
and ( n39295 , n38968 , n39294 );
and ( n39296 , n38966 , n39295 );
and ( n39297 , n38964 , n39296 );
and ( n39298 , n38962 , n39297 );
and ( n39299 , n38960 , n39298 );
and ( n39300 , n38959 , n39299 );
or ( n39301 , n38958 , n39300 );
and ( n39302 , n38956 , n39301 );
and ( n39303 , n38954 , n39302 );
and ( n39304 , n38953 , n39303 );
and ( n39305 , n38952 , n39304 );
or ( n39306 , n38951 , n39305 );
and ( n39307 , n38156 , n39306 );
and ( n39308 , n38154 , n39307 );
or ( n39309 , n38153 , n39308 );
and ( n39310 , n38151 , n39309 );
and ( n39311 , n38150 , n39310 );
and ( n39312 , n38149 , n39311 );
or ( n39313 , n38148 , n39312 );
and ( n39314 , n38146 , n39313 );
and ( n39315 , n38144 , n39314 );
or ( n39316 , n38143 , n39315 );
and ( n39317 , n36964 , n39316 );
or ( n39318 , n36963 , n39317 );
and ( n39319 , n36961 , n39318 );
and ( n39320 , n36959 , n39319 );
and ( n39321 , n36958 , n39320 );
and ( n39322 , n36956 , n39321 );
and ( n39323 , n36954 , n39322 );
and ( n39324 , n36952 , n39323 );
or ( n39325 , n36951 , n39324 );
and ( n39326 , n36949 , n39325 );
and ( n39327 , n36947 , n39326 );
or ( n39328 , n36946 , n39327 );
and ( n39329 , n34956 , n39328 );
and ( n39330 , n34954 , n39329 );
or ( n39331 , n34953 , n39330 );
and ( n39332 , n34951 , n39331 );
and ( n39333 , n34950 , n39332 );
and ( n39334 , n34949 , n39333 );
and ( n39335 , n34947 , n39334 );
or ( n39336 , n34946 , n39335 );
and ( n39337 , n34944 , n39336 );
or ( n39338 , n34943 , n39337 );
and ( n39339 , n34941 , n39338 );
and ( n39340 , n34939 , n39339 );
and ( n39341 , n34937 , n39340 );
or ( n39342 , n34936 , n39341 );
and ( n39343 , n34934 , n39342 );
or ( n39344 , n34933 , n39343 );
and ( n39345 , n32137 , n39344 );
and ( n39346 , n32135 , n39345 );
and ( n39347 , n32134 , n39346 );
or ( n39348 , n32133 , n39347 );
and ( n39349 , n32131 , n39348 );
and ( n39350 , n32129 , n39349 );
or ( n39351 , n32128 , n39350 );
and ( n39352 , n31389 , n39351 );
and ( n39353 , n31388 , n39352 );
or ( n39354 , n31387 , n39353 );
and ( n39355 , n31385 , n39354 );
or ( n39356 , n31384 , n39355 );
and ( n39357 , n31382 , n39356 );
and ( n39358 , n31380 , n39357 );
and ( n39359 , n31379 , n39358 );
or ( n39360 , n31378 , n39359 );
and ( n39361 , n31376 , n39360 );
xor ( n39362 , n31375 , n39361 );
buf ( n566664 , n39362 );
buf ( n566665 , n566664 );
buf ( n39365 , n566665 );
buf ( n566667 , n1154 );
buf ( n39367 , n566667 );
buf ( n566669 , n1155 );
buf ( n39369 , n566669 );
xor ( n39370 , n39367 , n39369 );
buf ( n566672 , n1156 );
buf ( n39372 , n566672 );
xor ( n39373 , n39369 , n39372 );
not ( n39374 , n39373 );
and ( n39375 , n39370 , n39374 );
and ( n39376 , n39365 , n39375 );
not ( n39377 , n39376 );
and ( n39378 , n39369 , n39372 );
not ( n39379 , n39378 );
and ( n39380 , n39367 , n39379 );
xnor ( n39381 , n39377 , n39380 );
buf ( n39382 , n39381 );
not ( n39383 , n39380 );
and ( n39384 , n39382 , n39383 );
and ( n39385 , n39365 , n39367 );
and ( n39386 , n39383 , n39385 );
and ( n39387 , n39382 , n39385 );
or ( n39388 , n39384 , n39386 , n39387 );
buf ( n566690 , n1157 );
buf ( n39390 , n566690 );
xor ( n39391 , n39372 , n39390 );
buf ( n566693 , n1158 );
buf ( n39393 , n566693 );
xor ( n39394 , n39390 , n39393 );
not ( n39395 , n39394 );
and ( n39396 , n39391 , n39395 );
and ( n39397 , n39365 , n39396 );
not ( n39398 , n39397 );
and ( n39399 , n39390 , n39393 );
not ( n39400 , n39399 );
and ( n39401 , n39372 , n39400 );
xnor ( n39402 , n39398 , n39401 );
buf ( n39403 , n39402 );
not ( n39404 , n39401 );
and ( n39405 , n39403 , n39404 );
xor ( n39406 , n31376 , n39360 );
buf ( n566708 , n39406 );
buf ( n566709 , n566708 );
buf ( n39409 , n566709 );
and ( n39410 , n39409 , n39375 );
and ( n39411 , n39365 , n39373 );
nor ( n39412 , n39410 , n39411 );
xnor ( n39413 , n39412 , n39380 );
and ( n39414 , n39404 , n39413 );
and ( n39415 , n39403 , n39413 );
or ( n39416 , n39405 , n39414 , n39415 );
not ( n39417 , n39381 );
and ( n39418 , n39416 , n39417 );
and ( n39419 , n39409 , n39367 );
and ( n39420 , n39417 , n39419 );
and ( n39421 , n39416 , n39419 );
or ( n39422 , n39418 , n39420 , n39421 );
xor ( n39423 , n39382 , n39383 );
xor ( n39424 , n39423 , n39385 );
and ( n39425 , n39422 , n39424 );
xor ( n39426 , n39416 , n39417 );
xor ( n39427 , n39426 , n39419 );
not ( n39428 , n39402 );
xor ( n39429 , n31379 , n39358 );
buf ( n566731 , n39429 );
buf ( n566732 , n566731 );
buf ( n39432 , n566732 );
and ( n39433 , n39432 , n39375 );
and ( n39434 , n39409 , n39373 );
nor ( n39435 , n39433 , n39434 );
xnor ( n39436 , n39435 , n39380 );
and ( n39437 , n39428 , n39436 );
xor ( n39438 , n31380 , n39357 );
buf ( n566740 , n39438 );
buf ( n566741 , n566740 );
buf ( n39441 , n566741 );
and ( n39442 , n39441 , n39367 );
and ( n39443 , n39436 , n39442 );
and ( n39444 , n39428 , n39442 );
or ( n39445 , n39437 , n39443 , n39444 );
and ( n39446 , n39432 , n39367 );
and ( n39447 , n39445 , n39446 );
xor ( n39448 , n39403 , n39404 );
xor ( n39449 , n39448 , n39413 );
and ( n39450 , n39446 , n39449 );
and ( n39451 , n39445 , n39449 );
or ( n39452 , n39447 , n39450 , n39451 );
and ( n39453 , n39427 , n39452 );
xor ( n39454 , n39445 , n39446 );
xor ( n39455 , n39454 , n39449 );
buf ( n566757 , n1159 );
buf ( n39457 , n566757 );
buf ( n566759 , n1160 );
buf ( n39459 , n566759 );
and ( n39460 , n39457 , n39459 );
not ( n39461 , n39460 );
and ( n39462 , n39393 , n39461 );
not ( n39463 , n39462 );
and ( n39464 , n39409 , n39396 );
and ( n39465 , n39365 , n39394 );
nor ( n39466 , n39464 , n39465 );
xnor ( n39467 , n39466 , n39401 );
and ( n39468 , n39463 , n39467 );
xor ( n39469 , n31382 , n39356 );
buf ( n566771 , n39469 );
buf ( n566772 , n566771 );
buf ( n39472 , n566772 );
and ( n39473 , n39472 , n39367 );
and ( n39474 , n39467 , n39473 );
and ( n39475 , n39463 , n39473 );
or ( n39476 , n39468 , n39474 , n39475 );
xor ( n39477 , n39393 , n39457 );
xor ( n39478 , n39457 , n39459 );
not ( n39479 , n39478 );
and ( n39480 , n39477 , n39479 );
and ( n39481 , n39365 , n39480 );
not ( n39482 , n39481 );
xnor ( n39483 , n39482 , n39462 );
not ( n39484 , n39483 );
and ( n39485 , n39432 , n39396 );
and ( n39486 , n39409 , n39394 );
nor ( n39487 , n39485 , n39486 );
xnor ( n39488 , n39487 , n39401 );
and ( n39489 , n39484 , n39488 );
xor ( n39490 , n31385 , n39354 );
buf ( n566792 , n39490 );
buf ( n566793 , n566792 );
buf ( n39493 , n566793 );
and ( n39494 , n39493 , n39367 );
and ( n39495 , n39488 , n39494 );
and ( n39496 , n39484 , n39494 );
or ( n39497 , n39489 , n39495 , n39496 );
buf ( n39498 , n39483 );
and ( n39499 , n39497 , n39498 );
and ( n39500 , n39441 , n39375 );
and ( n39501 , n39432 , n39373 );
nor ( n39502 , n39500 , n39501 );
xnor ( n39503 , n39502 , n39380 );
and ( n39504 , n39498 , n39503 );
and ( n39505 , n39497 , n39503 );
or ( n39506 , n39499 , n39504 , n39505 );
and ( n39507 , n39476 , n39506 );
xor ( n39508 , n39428 , n39436 );
xor ( n39509 , n39508 , n39442 );
and ( n39510 , n39506 , n39509 );
and ( n39511 , n39476 , n39509 );
or ( n39512 , n39507 , n39510 , n39511 );
and ( n39513 , n39455 , n39512 );
xor ( n39514 , n39476 , n39506 );
xor ( n39515 , n39514 , n39509 );
buf ( n566817 , n1161 );
buf ( n39517 , n566817 );
buf ( n566819 , n1162 );
buf ( n39519 , n566819 );
and ( n39520 , n39517 , n39519 );
not ( n39521 , n39520 );
and ( n39522 , n39459 , n39521 );
not ( n39523 , n39522 );
and ( n39524 , n39409 , n39480 );
and ( n39525 , n39365 , n39478 );
nor ( n39526 , n39524 , n39525 );
xnor ( n39527 , n39526 , n39462 );
and ( n39528 , n39523 , n39527 );
and ( n39529 , n39493 , n39375 );
and ( n39530 , n39472 , n39373 );
nor ( n39531 , n39529 , n39530 );
xnor ( n39532 , n39531 , n39380 );
and ( n39533 , n39527 , n39532 );
and ( n39534 , n39523 , n39532 );
or ( n39535 , n39528 , n39533 , n39534 );
xor ( n39536 , n39459 , n39517 );
xor ( n39537 , n39517 , n39519 );
not ( n39538 , n39537 );
and ( n39539 , n39536 , n39538 );
and ( n39540 , n39365 , n39539 );
not ( n39541 , n39540 );
xnor ( n39542 , n39541 , n39522 );
buf ( n39543 , n39542 );
and ( n39544 , n39441 , n39396 );
and ( n39545 , n39432 , n39394 );
nor ( n39546 , n39544 , n39545 );
xnor ( n39547 , n39546 , n39401 );
and ( n39548 , n39543 , n39547 );
xor ( n39549 , n31388 , n39352 );
buf ( n566851 , n39549 );
buf ( n566852 , n566851 );
buf ( n39552 , n566852 );
and ( n39553 , n39552 , n39367 );
and ( n39554 , n39547 , n39553 );
and ( n39555 , n39543 , n39553 );
or ( n39556 , n39548 , n39554 , n39555 );
and ( n39557 , n39535 , n39556 );
and ( n39558 , n39472 , n39375 );
and ( n39559 , n39441 , n39373 );
nor ( n39560 , n39558 , n39559 );
xnor ( n39561 , n39560 , n39380 );
and ( n39562 , n39556 , n39561 );
and ( n39563 , n39535 , n39561 );
or ( n39564 , n39557 , n39562 , n39563 );
xor ( n39565 , n39463 , n39467 );
xor ( n39566 , n39565 , n39473 );
and ( n39567 , n39564 , n39566 );
xor ( n39568 , n39497 , n39498 );
xor ( n39569 , n39568 , n39503 );
and ( n39570 , n39566 , n39569 );
and ( n39571 , n39564 , n39569 );
or ( n39572 , n39567 , n39570 , n39571 );
and ( n39573 , n39515 , n39572 );
xor ( n39574 , n39564 , n39566 );
xor ( n39575 , n39574 , n39569 );
not ( n39576 , n39542 );
and ( n39577 , n39432 , n39480 );
and ( n39578 , n39409 , n39478 );
nor ( n39579 , n39577 , n39578 );
xnor ( n39580 , n39579 , n39462 );
and ( n39581 , n39576 , n39580 );
and ( n39582 , n39552 , n39375 );
and ( n39583 , n39493 , n39373 );
nor ( n39584 , n39582 , n39583 );
xnor ( n39585 , n39584 , n39380 );
and ( n39586 , n39580 , n39585 );
and ( n39587 , n39576 , n39585 );
or ( n39588 , n39581 , n39586 , n39587 );
xor ( n39589 , n39523 , n39527 );
xor ( n39590 , n39589 , n39532 );
and ( n39591 , n39588 , n39590 );
xor ( n39592 , n39543 , n39547 );
xor ( n39593 , n39592 , n39553 );
and ( n39594 , n39590 , n39593 );
and ( n39595 , n39588 , n39593 );
or ( n39596 , n39591 , n39594 , n39595 );
xor ( n39597 , n39535 , n39556 );
xor ( n39598 , n39597 , n39561 );
and ( n39599 , n39596 , n39598 );
xor ( n39600 , n39484 , n39488 );
xor ( n39601 , n39600 , n39494 );
and ( n39602 , n39598 , n39601 );
and ( n39603 , n39596 , n39601 );
or ( n39604 , n39599 , n39602 , n39603 );
and ( n39605 , n39575 , n39604 );
xor ( n39606 , n39596 , n39598 );
xor ( n39607 , n39606 , n39601 );
and ( n39608 , n39441 , n39480 );
and ( n39609 , n39432 , n39478 );
nor ( n39610 , n39608 , n39609 );
xnor ( n39611 , n39610 , n39462 );
and ( n39612 , n39493 , n39396 );
and ( n39613 , n39472 , n39394 );
nor ( n39614 , n39612 , n39613 );
xnor ( n39615 , n39614 , n39401 );
and ( n39616 , n39611 , n39615 );
xor ( n39617 , n31389 , n39351 );
buf ( n566919 , n39617 );
buf ( n566920 , n566919 );
buf ( n39620 , n566920 );
and ( n39621 , n39620 , n39375 );
and ( n39622 , n39552 , n39373 );
nor ( n39623 , n39621 , n39622 );
xnor ( n39624 , n39623 , n39380 );
and ( n39625 , n39615 , n39624 );
and ( n39626 , n39611 , n39624 );
or ( n39627 , n39616 , n39625 , n39626 );
and ( n39628 , n39472 , n39396 );
and ( n39629 , n39441 , n39394 );
nor ( n39630 , n39628 , n39629 );
xnor ( n39631 , n39630 , n39401 );
and ( n39632 , n39627 , n39631 );
and ( n39633 , n39620 , n39367 );
and ( n39634 , n39631 , n39633 );
and ( n39635 , n39627 , n39633 );
or ( n39636 , n39632 , n39634 , n39635 );
buf ( n566938 , n1163 );
buf ( n39638 , n566938 );
buf ( n566940 , n1164 );
buf ( n39640 , n566940 );
and ( n39641 , n39638 , n39640 );
not ( n39642 , n39641 );
and ( n39643 , n39519 , n39642 );
not ( n39644 , n39643 );
and ( n39645 , n39409 , n39539 );
and ( n39646 , n39365 , n39537 );
nor ( n39647 , n39645 , n39646 );
xnor ( n39648 , n39647 , n39522 );
and ( n39649 , n39644 , n39648 );
xor ( n39650 , n32129 , n39349 );
buf ( n566952 , n39650 );
buf ( n566953 , n566952 );
buf ( n39653 , n566953 );
and ( n39654 , n39653 , n39367 );
and ( n39655 , n39648 , n39654 );
and ( n39656 , n39644 , n39654 );
or ( n39657 , n39649 , n39655 , n39656 );
and ( n39658 , n39432 , n39539 );
and ( n39659 , n39409 , n39537 );
nor ( n39660 , n39658 , n39659 );
xnor ( n39661 , n39660 , n39522 );
and ( n39662 , n39552 , n39396 );
and ( n39663 , n39493 , n39394 );
nor ( n39664 , n39662 , n39663 );
xnor ( n39665 , n39664 , n39401 );
and ( n39666 , n39661 , n39665 );
xor ( n39667 , n32131 , n39348 );
buf ( n566969 , n39667 );
buf ( n566970 , n566969 );
buf ( n39670 , n566970 );
and ( n39671 , n39670 , n39367 );
and ( n39672 , n39665 , n39671 );
and ( n39673 , n39661 , n39671 );
or ( n39674 , n39666 , n39672 , n39673 );
xor ( n39675 , n39519 , n39638 );
xor ( n39676 , n39638 , n39640 );
not ( n39677 , n39676 );
and ( n39678 , n39675 , n39677 );
and ( n39679 , n39365 , n39678 );
not ( n39680 , n39679 );
xnor ( n39681 , n39680 , n39643 );
not ( n39682 , n39681 );
and ( n39683 , n39472 , n39480 );
and ( n39684 , n39441 , n39478 );
nor ( n39685 , n39683 , n39684 );
xnor ( n39686 , n39685 , n39462 );
and ( n39687 , n39682 , n39686 );
and ( n39688 , n39653 , n39375 );
and ( n39689 , n39620 , n39373 );
nor ( n39690 , n39688 , n39689 );
xnor ( n39691 , n39690 , n39380 );
and ( n39692 , n39686 , n39691 );
and ( n39693 , n39682 , n39691 );
or ( n39694 , n39687 , n39692 , n39693 );
and ( n39695 , n39674 , n39694 );
buf ( n39696 , n39681 );
and ( n39697 , n39694 , n39696 );
and ( n39698 , n39674 , n39696 );
or ( n39699 , n39695 , n39697 , n39698 );
and ( n39700 , n39657 , n39699 );
xor ( n39701 , n39576 , n39580 );
xor ( n39702 , n39701 , n39585 );
and ( n39703 , n39699 , n39702 );
and ( n39704 , n39657 , n39702 );
or ( n39705 , n39700 , n39703 , n39704 );
and ( n39706 , n39636 , n39705 );
xor ( n39707 , n39588 , n39590 );
xor ( n39708 , n39707 , n39593 );
and ( n39709 , n39705 , n39708 );
and ( n39710 , n39636 , n39708 );
or ( n39711 , n39706 , n39709 , n39710 );
and ( n39712 , n39607 , n39711 );
xor ( n39713 , n39636 , n39705 );
xor ( n39714 , n39713 , n39708 );
xor ( n39715 , n39644 , n39648 );
xor ( n39716 , n39715 , n39654 );
xor ( n39717 , n39611 , n39615 );
xor ( n39718 , n39717 , n39624 );
and ( n39719 , n39716 , n39718 );
xor ( n39720 , n39674 , n39694 );
xor ( n39721 , n39720 , n39696 );
and ( n39722 , n39718 , n39721 );
and ( n39723 , n39716 , n39721 );
or ( n39724 , n39719 , n39722 , n39723 );
xor ( n39725 , n39627 , n39631 );
xor ( n39726 , n39725 , n39633 );
and ( n39727 , n39724 , n39726 );
xor ( n39728 , n39657 , n39699 );
xor ( n39729 , n39728 , n39702 );
and ( n39730 , n39726 , n39729 );
and ( n39731 , n39724 , n39729 );
or ( n39732 , n39727 , n39730 , n39731 );
and ( n39733 , n39714 , n39732 );
xor ( n39734 , n39724 , n39726 );
xor ( n39735 , n39734 , n39729 );
buf ( n567037 , n1165 );
buf ( n39737 , n567037 );
buf ( n567039 , n1166 );
buf ( n39739 , n567039 );
and ( n39740 , n39737 , n39739 );
not ( n39741 , n39740 );
and ( n39742 , n39640 , n39741 );
not ( n39743 , n39742 );
and ( n39744 , n39670 , n39375 );
and ( n39745 , n39653 , n39373 );
nor ( n39746 , n39744 , n39745 );
xnor ( n39747 , n39746 , n39380 );
and ( n39748 , n39743 , n39747 );
xor ( n39749 , n32134 , n39346 );
buf ( n567051 , n39749 );
buf ( n567052 , n567051 );
buf ( n39752 , n567052 );
and ( n39753 , n39752 , n39367 );
and ( n39754 , n39747 , n39753 );
and ( n39755 , n39743 , n39753 );
or ( n39756 , n39748 , n39754 , n39755 );
xor ( n39757 , n39640 , n39737 );
xor ( n39758 , n39737 , n39739 );
not ( n39759 , n39758 );
and ( n39760 , n39757 , n39759 );
and ( n39761 , n39365 , n39760 );
not ( n39762 , n39761 );
xnor ( n39763 , n39762 , n39742 );
buf ( n39764 , n39763 );
and ( n39765 , n39409 , n39678 );
and ( n39766 , n39365 , n39676 );
nor ( n39767 , n39765 , n39766 );
xnor ( n39768 , n39767 , n39643 );
and ( n39769 , n39764 , n39768 );
and ( n39770 , n39493 , n39480 );
and ( n39771 , n39472 , n39478 );
nor ( n39772 , n39770 , n39771 );
xnor ( n39773 , n39772 , n39462 );
and ( n39774 , n39768 , n39773 );
and ( n39775 , n39764 , n39773 );
or ( n39776 , n39769 , n39774 , n39775 );
and ( n39777 , n39756 , n39776 );
xor ( n39778 , n39682 , n39686 );
xor ( n39779 , n39778 , n39691 );
and ( n39780 , n39776 , n39779 );
and ( n39781 , n39756 , n39779 );
or ( n39782 , n39777 , n39780 , n39781 );
and ( n39783 , n39432 , n39678 );
and ( n39784 , n39409 , n39676 );
nor ( n39785 , n39783 , n39784 );
xnor ( n39786 , n39785 , n39643 );
and ( n39787 , n39752 , n39375 );
and ( n39788 , n39670 , n39373 );
nor ( n39789 , n39787 , n39788 );
xnor ( n39790 , n39789 , n39380 );
and ( n39791 , n39786 , n39790 );
xor ( n39792 , n32135 , n39345 );
buf ( n567094 , n39792 );
buf ( n567095 , n567094 );
buf ( n39795 , n567095 );
and ( n39796 , n39795 , n39367 );
and ( n39797 , n39790 , n39796 );
and ( n39798 , n39786 , n39796 );
or ( n39799 , n39791 , n39797 , n39798 );
and ( n39800 , n39441 , n39539 );
and ( n39801 , n39432 , n39537 );
nor ( n39802 , n39800 , n39801 );
xnor ( n39803 , n39802 , n39522 );
and ( n39804 , n39799 , n39803 );
and ( n39805 , n39620 , n39396 );
and ( n39806 , n39552 , n39394 );
nor ( n39807 , n39805 , n39806 );
xnor ( n39808 , n39807 , n39401 );
and ( n39809 , n39803 , n39808 );
and ( n39810 , n39799 , n39808 );
or ( n39811 , n39804 , n39809 , n39810 );
and ( n39812 , n39472 , n39539 );
and ( n39813 , n39441 , n39537 );
nor ( n39814 , n39812 , n39813 );
xnor ( n39815 , n39814 , n39522 );
and ( n39816 , n39552 , n39480 );
and ( n39817 , n39493 , n39478 );
nor ( n39818 , n39816 , n39817 );
xnor ( n39819 , n39818 , n39462 );
and ( n39820 , n39815 , n39819 );
and ( n39821 , n39653 , n39396 );
and ( n39822 , n39620 , n39394 );
nor ( n39823 , n39821 , n39822 );
xnor ( n39824 , n39823 , n39401 );
and ( n39825 , n39819 , n39824 );
and ( n39826 , n39815 , n39824 );
or ( n39827 , n39820 , n39825 , n39826 );
xor ( n39828 , n39743 , n39747 );
xor ( n39829 , n39828 , n39753 );
and ( n39830 , n39827 , n39829 );
xor ( n39831 , n39764 , n39768 );
xor ( n39832 , n39831 , n39773 );
and ( n39833 , n39829 , n39832 );
and ( n39834 , n39827 , n39832 );
or ( n39835 , n39830 , n39833 , n39834 );
and ( n39836 , n39811 , n39835 );
xor ( n39837 , n39661 , n39665 );
xor ( n39838 , n39837 , n39671 );
and ( n39839 , n39835 , n39838 );
and ( n39840 , n39811 , n39838 );
or ( n39841 , n39836 , n39839 , n39840 );
and ( n39842 , n39782 , n39841 );
xor ( n39843 , n39716 , n39718 );
xor ( n39844 , n39843 , n39721 );
and ( n39845 , n39841 , n39844 );
and ( n39846 , n39782 , n39844 );
or ( n39847 , n39842 , n39845 , n39846 );
and ( n39848 , n39735 , n39847 );
xor ( n39849 , n39782 , n39841 );
xor ( n39850 , n39849 , n39844 );
buf ( n567152 , n1167 );
buf ( n39852 , n567152 );
buf ( n567154 , n1168 );
buf ( n39854 , n567154 );
and ( n39855 , n39852 , n39854 );
not ( n39856 , n39855 );
and ( n39857 , n39739 , n39856 );
not ( n39858 , n39857 );
and ( n39859 , n39670 , n39396 );
and ( n39860 , n39653 , n39394 );
nor ( n39861 , n39859 , n39860 );
xnor ( n39862 , n39861 , n39401 );
and ( n39863 , n39858 , n39862 );
xor ( n39864 , n32137 , n39344 );
buf ( n567166 , n39864 );
buf ( n567167 , n567166 );
buf ( n39867 , n567167 );
and ( n39868 , n39867 , n39367 );
and ( n39869 , n39862 , n39868 );
and ( n39870 , n39858 , n39868 );
or ( n39871 , n39863 , n39869 , n39870 );
and ( n39872 , n39409 , n39760 );
and ( n39873 , n39365 , n39758 );
nor ( n39874 , n39872 , n39873 );
xnor ( n39875 , n39874 , n39742 );
and ( n39876 , n39493 , n39539 );
and ( n39877 , n39472 , n39537 );
nor ( n39878 , n39876 , n39877 );
xnor ( n39879 , n39878 , n39522 );
and ( n39880 , n39875 , n39879 );
and ( n39881 , n39795 , n39375 );
and ( n39882 , n39752 , n39373 );
nor ( n39883 , n39881 , n39882 );
xnor ( n39884 , n39883 , n39380 );
and ( n39885 , n39879 , n39884 );
and ( n39886 , n39875 , n39884 );
or ( n39887 , n39880 , n39885 , n39886 );
and ( n39888 , n39871 , n39887 );
not ( n39889 , n39763 );
and ( n39890 , n39887 , n39889 );
and ( n39891 , n39871 , n39889 );
or ( n39892 , n39888 , n39890 , n39891 );
xor ( n39893 , n39739 , n39852 );
xor ( n39894 , n39852 , n39854 );
not ( n39895 , n39894 );
and ( n39896 , n39893 , n39895 );
and ( n39897 , n39365 , n39896 );
not ( n39898 , n39897 );
xnor ( n39899 , n39898 , n39857 );
buf ( n39900 , n39899 );
and ( n39901 , n39441 , n39678 );
and ( n39902 , n39432 , n39676 );
nor ( n39903 , n39901 , n39902 );
xnor ( n39904 , n39903 , n39643 );
and ( n39905 , n39900 , n39904 );
and ( n39906 , n39620 , n39480 );
and ( n39907 , n39552 , n39478 );
nor ( n39908 , n39906 , n39907 );
xnor ( n39909 , n39908 , n39462 );
and ( n39910 , n39904 , n39909 );
and ( n39911 , n39900 , n39909 );
or ( n39912 , n39905 , n39910 , n39911 );
xor ( n39913 , n39786 , n39790 );
xor ( n39914 , n39913 , n39796 );
and ( n39915 , n39912 , n39914 );
xor ( n39916 , n39815 , n39819 );
xor ( n39917 , n39916 , n39824 );
and ( n39918 , n39914 , n39917 );
and ( n39919 , n39912 , n39917 );
or ( n39920 , n39915 , n39918 , n39919 );
and ( n39921 , n39892 , n39920 );
xor ( n39922 , n39799 , n39803 );
xor ( n39923 , n39922 , n39808 );
and ( n39924 , n39920 , n39923 );
and ( n39925 , n39892 , n39923 );
or ( n39926 , n39921 , n39924 , n39925 );
xor ( n39927 , n39756 , n39776 );
xor ( n39928 , n39927 , n39779 );
and ( n39929 , n39926 , n39928 );
xor ( n39930 , n39811 , n39835 );
xor ( n39931 , n39930 , n39838 );
and ( n39932 , n39928 , n39931 );
and ( n39933 , n39926 , n39931 );
or ( n39934 , n39929 , n39932 , n39933 );
and ( n39935 , n39850 , n39934 );
and ( n39936 , n39752 , n39396 );
and ( n39937 , n39670 , n39394 );
nor ( n39938 , n39936 , n39937 );
xnor ( n39939 , n39938 , n39401 );
and ( n39940 , n39867 , n39375 );
and ( n39941 , n39795 , n39373 );
nor ( n39942 , n39940 , n39941 );
xnor ( n39943 , n39942 , n39380 );
and ( n39944 , n39939 , n39943 );
xor ( n39945 , n34934 , n39342 );
buf ( n567247 , n39945 );
buf ( n567248 , n567247 );
buf ( n39948 , n567248 );
and ( n39949 , n39948 , n39367 );
and ( n39950 , n39943 , n39949 );
and ( n39951 , n39939 , n39949 );
or ( n39952 , n39944 , n39950 , n39951 );
not ( n39953 , n39899 );
and ( n39954 , n39432 , n39760 );
and ( n39955 , n39409 , n39758 );
nor ( n39956 , n39954 , n39955 );
xnor ( n39957 , n39956 , n39742 );
and ( n39958 , n39953 , n39957 );
and ( n39959 , n39552 , n39539 );
and ( n39960 , n39493 , n39537 );
nor ( n39961 , n39959 , n39960 );
xnor ( n39962 , n39961 , n39522 );
and ( n39963 , n39957 , n39962 );
and ( n39964 , n39953 , n39962 );
or ( n39965 , n39958 , n39963 , n39964 );
and ( n39966 , n39952 , n39965 );
xor ( n39967 , n39858 , n39862 );
xor ( n39968 , n39967 , n39868 );
and ( n39969 , n39965 , n39968 );
and ( n39970 , n39952 , n39968 );
or ( n39971 , n39966 , n39969 , n39970 );
xor ( n39972 , n39871 , n39887 );
xor ( n39973 , n39972 , n39889 );
and ( n39974 , n39971 , n39973 );
xor ( n39975 , n39912 , n39914 );
xor ( n39976 , n39975 , n39917 );
and ( n39977 , n39973 , n39976 );
and ( n39978 , n39971 , n39976 );
or ( n39979 , n39974 , n39977 , n39978 );
xor ( n39980 , n39827 , n39829 );
xor ( n39981 , n39980 , n39832 );
and ( n39982 , n39979 , n39981 );
xor ( n39983 , n39892 , n39920 );
xor ( n39984 , n39983 , n39923 );
and ( n39985 , n39981 , n39984 );
and ( n39986 , n39979 , n39984 );
or ( n39987 , n39982 , n39985 , n39986 );
xor ( n39988 , n39926 , n39928 );
xor ( n39989 , n39988 , n39931 );
and ( n39990 , n39987 , n39989 );
xor ( n39991 , n39979 , n39981 );
xor ( n39992 , n39991 , n39984 );
buf ( n567294 , n1169 );
buf ( n39994 , n567294 );
buf ( n567296 , n1170 );
buf ( n39996 , n567296 );
and ( n39997 , n39994 , n39996 );
not ( n39998 , n39997 );
and ( n39999 , n39854 , n39998 );
not ( n40000 , n39999 );
and ( n40001 , n39948 , n39375 );
and ( n40002 , n39867 , n39373 );
nor ( n40003 , n40001 , n40002 );
xnor ( n40004 , n40003 , n39380 );
and ( n40005 , n40000 , n40004 );
xor ( n40006 , n34937 , n39340 );
buf ( n567308 , n40006 );
buf ( n567309 , n567308 );
buf ( n40009 , n567309 );
and ( n40010 , n40009 , n39367 );
and ( n40011 , n40004 , n40010 );
and ( n40012 , n40000 , n40010 );
or ( n40013 , n40005 , n40011 , n40012 );
and ( n40014 , n39472 , n39678 );
and ( n40015 , n39441 , n39676 );
nor ( n40016 , n40014 , n40015 );
xnor ( n40017 , n40016 , n39643 );
and ( n40018 , n40013 , n40017 );
and ( n40019 , n39653 , n39480 );
and ( n40020 , n39620 , n39478 );
nor ( n40021 , n40019 , n40020 );
xnor ( n40022 , n40021 , n39462 );
and ( n40023 , n40017 , n40022 );
and ( n40024 , n40013 , n40022 );
or ( n40025 , n40018 , n40023 , n40024 );
xor ( n40026 , n39875 , n39879 );
xor ( n40027 , n40026 , n39884 );
and ( n40028 , n40025 , n40027 );
xor ( n40029 , n39900 , n39904 );
xor ( n40030 , n40029 , n39909 );
and ( n40031 , n40027 , n40030 );
and ( n40032 , n40025 , n40030 );
or ( n40033 , n40028 , n40031 , n40032 );
and ( n40034 , n39493 , n39678 );
and ( n40035 , n39472 , n39676 );
nor ( n40036 , n40034 , n40035 );
xnor ( n40037 , n40036 , n39643 );
and ( n40038 , n39670 , n39480 );
and ( n40039 , n39653 , n39478 );
nor ( n40040 , n40038 , n40039 );
xnor ( n40041 , n40040 , n39462 );
and ( n40042 , n40037 , n40041 );
and ( n40043 , n39795 , n39396 );
and ( n40044 , n39752 , n39394 );
nor ( n40045 , n40043 , n40044 );
xnor ( n40046 , n40045 , n39401 );
and ( n40047 , n40041 , n40046 );
and ( n40048 , n40037 , n40046 );
or ( n40049 , n40042 , n40047 , n40048 );
xor ( n40050 , n39854 , n39994 );
xor ( n40051 , n39994 , n39996 );
not ( n40052 , n40051 );
and ( n40053 , n40050 , n40052 );
and ( n40054 , n39365 , n40053 );
not ( n40055 , n40054 );
xnor ( n40056 , n40055 , n39999 );
buf ( n40057 , n40056 );
and ( n40058 , n39409 , n39896 );
and ( n40059 , n39365 , n39894 );
nor ( n40060 , n40058 , n40059 );
xnor ( n40061 , n40060 , n39857 );
and ( n40062 , n40057 , n40061 );
and ( n40063 , n39620 , n39539 );
and ( n40064 , n39552 , n39537 );
nor ( n40065 , n40063 , n40064 );
xnor ( n40066 , n40065 , n39522 );
and ( n40067 , n40061 , n40066 );
and ( n40068 , n40057 , n40066 );
or ( n40069 , n40062 , n40067 , n40068 );
and ( n40070 , n40049 , n40069 );
xor ( n40071 , n39939 , n39943 );
xor ( n40072 , n40071 , n39949 );
and ( n40073 , n40069 , n40072 );
and ( n40074 , n40049 , n40072 );
or ( n40075 , n40070 , n40073 , n40074 );
xor ( n40076 , n39952 , n39965 );
xor ( n40077 , n40076 , n39968 );
and ( n40078 , n40075 , n40077 );
xor ( n40079 , n40025 , n40027 );
xor ( n40080 , n40079 , n40030 );
and ( n40081 , n40077 , n40080 );
and ( n40082 , n40075 , n40080 );
or ( n40083 , n40078 , n40081 , n40082 );
and ( n40084 , n40033 , n40083 );
xor ( n40085 , n39971 , n39973 );
xor ( n40086 , n40085 , n39976 );
and ( n40087 , n40083 , n40086 );
and ( n40088 , n40033 , n40086 );
or ( n40089 , n40084 , n40087 , n40088 );
and ( n40090 , n39992 , n40089 );
xor ( n40091 , n40033 , n40083 );
xor ( n40092 , n40091 , n40086 );
and ( n40093 , n39432 , n39896 );
and ( n40094 , n39409 , n39894 );
nor ( n40095 , n40093 , n40094 );
xnor ( n40096 , n40095 , n39857 );
and ( n40097 , n39472 , n39760 );
and ( n40098 , n39441 , n39758 );
nor ( n40099 , n40097 , n40098 );
xnor ( n40100 , n40099 , n39742 );
and ( n40101 , n40096 , n40100 );
and ( n40102 , n39653 , n39539 );
and ( n40103 , n39620 , n39537 );
nor ( n40104 , n40102 , n40103 );
xnor ( n40105 , n40104 , n39522 );
and ( n40106 , n40100 , n40105 );
and ( n40107 , n40096 , n40105 );
or ( n40108 , n40101 , n40106 , n40107 );
not ( n40109 , n40056 );
and ( n40110 , n39552 , n39678 );
and ( n40111 , n39493 , n39676 );
nor ( n40112 , n40110 , n40111 );
xnor ( n40113 , n40112 , n39643 );
and ( n40114 , n40109 , n40113 );
and ( n40115 , n39867 , n39396 );
and ( n40116 , n39795 , n39394 );
nor ( n40117 , n40115 , n40116 );
xnor ( n40118 , n40117 , n39401 );
and ( n40119 , n40113 , n40118 );
and ( n40120 , n40109 , n40118 );
or ( n40121 , n40114 , n40119 , n40120 );
and ( n40122 , n40108 , n40121 );
xor ( n40123 , n40037 , n40041 );
xor ( n40124 , n40123 , n40046 );
and ( n40125 , n40121 , n40124 );
and ( n40126 , n40108 , n40124 );
or ( n40127 , n40122 , n40125 , n40126 );
xor ( n40128 , n40013 , n40017 );
xor ( n40129 , n40128 , n40022 );
and ( n40130 , n40127 , n40129 );
xor ( n40131 , n39953 , n39957 );
xor ( n40132 , n40131 , n39962 );
and ( n40133 , n40129 , n40132 );
and ( n40134 , n40127 , n40132 );
or ( n40135 , n40130 , n40133 , n40134 );
and ( n40136 , n39752 , n39480 );
and ( n40137 , n39670 , n39478 );
nor ( n40138 , n40136 , n40137 );
xnor ( n40139 , n40138 , n39462 );
and ( n40140 , n40009 , n39375 );
and ( n40141 , n39948 , n39373 );
nor ( n40142 , n40140 , n40141 );
xnor ( n40143 , n40142 , n39380 );
and ( n40144 , n40139 , n40143 );
xor ( n40145 , n34939 , n39339 );
buf ( n567447 , n40145 );
buf ( n567448 , n567447 );
buf ( n40148 , n567448 );
and ( n40149 , n40148 , n39367 );
and ( n40150 , n40143 , n40149 );
and ( n40151 , n40139 , n40149 );
or ( n40152 , n40144 , n40150 , n40151 );
and ( n40153 , n39441 , n39760 );
and ( n40154 , n39432 , n39758 );
nor ( n40155 , n40153 , n40154 );
xnor ( n40156 , n40155 , n39742 );
and ( n40157 , n40152 , n40156 );
xor ( n40158 , n40000 , n40004 );
xor ( n40159 , n40158 , n40010 );
and ( n40160 , n40156 , n40159 );
and ( n40161 , n40152 , n40159 );
or ( n40162 , n40157 , n40160 , n40161 );
buf ( n567464 , n1171 );
buf ( n40164 , n567464 );
buf ( n567466 , n1172 );
buf ( n40166 , n567466 );
and ( n40167 , n40164 , n40166 );
not ( n40168 , n40167 );
and ( n40169 , n39996 , n40168 );
not ( n40170 , n40169 );
and ( n40171 , n39948 , n39396 );
and ( n40172 , n39867 , n39394 );
nor ( n40173 , n40171 , n40172 );
xnor ( n40174 , n40173 , n39401 );
and ( n40175 , n40170 , n40174 );
and ( n40176 , n40148 , n39375 );
and ( n40177 , n40009 , n39373 );
nor ( n40178 , n40176 , n40177 );
xnor ( n40179 , n40178 , n39380 );
and ( n40180 , n40174 , n40179 );
and ( n40181 , n40170 , n40179 );
or ( n40182 , n40175 , n40180 , n40181 );
xor ( n40183 , n34944 , n39336 );
buf ( n567485 , n40183 );
buf ( n567486 , n567485 );
buf ( n40186 , n567486 );
and ( n40187 , n40186 , n39367 );
buf ( n40188 , n40187 );
and ( n40189 , n39670 , n39539 );
and ( n40190 , n39653 , n39537 );
nor ( n40191 , n40189 , n40190 );
xnor ( n40192 , n40191 , n39522 );
and ( n40193 , n40188 , n40192 );
xor ( n40194 , n34941 , n39338 );
buf ( n567496 , n40194 );
buf ( n567497 , n567496 );
buf ( n40197 , n567497 );
and ( n40198 , n40197 , n39367 );
and ( n40199 , n40192 , n40198 );
and ( n40200 , n40188 , n40198 );
or ( n40201 , n40193 , n40199 , n40200 );
and ( n40202 , n40182 , n40201 );
xor ( n40203 , n40139 , n40143 );
xor ( n40204 , n40203 , n40149 );
and ( n40205 , n40201 , n40204 );
and ( n40206 , n40182 , n40204 );
or ( n40207 , n40202 , n40205 , n40206 );
xor ( n40208 , n40057 , n40061 );
xor ( n40209 , n40208 , n40066 );
and ( n40210 , n40207 , n40209 );
xor ( n40211 , n40152 , n40156 );
xor ( n40212 , n40211 , n40159 );
and ( n40213 , n40209 , n40212 );
and ( n40214 , n40207 , n40212 );
or ( n40215 , n40210 , n40213 , n40214 );
and ( n40216 , n40162 , n40215 );
xor ( n40217 , n40049 , n40069 );
xor ( n40218 , n40217 , n40072 );
and ( n40219 , n40215 , n40218 );
and ( n40220 , n40162 , n40218 );
or ( n40221 , n40216 , n40219 , n40220 );
and ( n40222 , n40135 , n40221 );
xor ( n40223 , n40075 , n40077 );
xor ( n40224 , n40223 , n40080 );
and ( n40225 , n40221 , n40224 );
and ( n40226 , n40135 , n40224 );
or ( n40227 , n40222 , n40225 , n40226 );
and ( n40228 , n40092 , n40227 );
xor ( n40229 , n40135 , n40221 );
xor ( n40230 , n40229 , n40224 );
and ( n40231 , n39409 , n40053 );
and ( n40232 , n39365 , n40051 );
nor ( n40233 , n40231 , n40232 );
xnor ( n40234 , n40233 , n39999 );
and ( n40235 , n39493 , n39760 );
and ( n40236 , n39472 , n39758 );
nor ( n40237 , n40235 , n40236 );
xnor ( n40238 , n40237 , n39742 );
and ( n40239 , n40234 , n40238 );
and ( n40240 , n39795 , n39480 );
and ( n40241 , n39752 , n39478 );
nor ( n40242 , n40240 , n40241 );
xnor ( n40243 , n40242 , n39462 );
and ( n40244 , n40238 , n40243 );
and ( n40245 , n40234 , n40243 );
or ( n40246 , n40239 , n40244 , n40245 );
xor ( n40247 , n40096 , n40100 );
xor ( n40248 , n40247 , n40105 );
and ( n40249 , n40246 , n40248 );
xor ( n40250 , n40109 , n40113 );
xor ( n40251 , n40250 , n40118 );
and ( n40252 , n40248 , n40251 );
and ( n40253 , n40246 , n40251 );
or ( n40254 , n40249 , n40252 , n40253 );
xor ( n40255 , n39996 , n40164 );
xor ( n40256 , n40164 , n40166 );
not ( n40257 , n40256 );
and ( n40258 , n40255 , n40257 );
and ( n40259 , n39365 , n40258 );
not ( n40260 , n40259 );
xnor ( n40261 , n40260 , n40169 );
and ( n40262 , n40009 , n39396 );
and ( n40263 , n39948 , n39394 );
nor ( n40264 , n40262 , n40263 );
xnor ( n40265 , n40264 , n39401 );
and ( n40266 , n40261 , n40265 );
and ( n40267 , n40197 , n39375 );
and ( n40268 , n40148 , n39373 );
nor ( n40269 , n40267 , n40268 );
xnor ( n40270 , n40269 , n39380 );
and ( n40271 , n40265 , n40270 );
and ( n40272 , n40261 , n40270 );
or ( n40273 , n40266 , n40271 , n40272 );
and ( n40274 , n39441 , n39896 );
and ( n40275 , n39432 , n39894 );
nor ( n40276 , n40274 , n40275 );
xnor ( n40277 , n40276 , n39857 );
and ( n40278 , n40273 , n40277 );
and ( n40279 , n39620 , n39678 );
and ( n40280 , n39552 , n39676 );
nor ( n40281 , n40279 , n40280 );
xnor ( n40282 , n40281 , n39643 );
and ( n40283 , n40277 , n40282 );
and ( n40284 , n40273 , n40282 );
or ( n40285 , n40278 , n40283 , n40284 );
and ( n40286 , n39752 , n39539 );
and ( n40287 , n39670 , n39537 );
nor ( n40288 , n40286 , n40287 );
xnor ( n40289 , n40288 , n39522 );
and ( n40290 , n39867 , n39480 );
and ( n40291 , n39795 , n39478 );
nor ( n40292 , n40290 , n40291 );
xnor ( n40293 , n40292 , n39462 );
and ( n40294 , n40289 , n40293 );
not ( n40295 , n40187 );
and ( n40296 , n40293 , n40295 );
and ( n40297 , n40289 , n40295 );
or ( n40298 , n40294 , n40296 , n40297 );
xor ( n40299 , n40170 , n40174 );
xor ( n40300 , n40299 , n40179 );
and ( n40301 , n40298 , n40300 );
xor ( n40302 , n40188 , n40192 );
xor ( n40303 , n40302 , n40198 );
and ( n40304 , n40300 , n40303 );
and ( n40305 , n40298 , n40303 );
or ( n40306 , n40301 , n40304 , n40305 );
and ( n40307 , n40285 , n40306 );
xor ( n40308 , n40182 , n40201 );
xor ( n40309 , n40308 , n40204 );
and ( n40310 , n40306 , n40309 );
and ( n40311 , n40285 , n40309 );
or ( n40312 , n40307 , n40310 , n40311 );
and ( n40313 , n40254 , n40312 );
xor ( n40314 , n40108 , n40121 );
xor ( n40315 , n40314 , n40124 );
and ( n40316 , n40312 , n40315 );
and ( n40317 , n40254 , n40315 );
or ( n40318 , n40313 , n40316 , n40317 );
xor ( n40319 , n40127 , n40129 );
xor ( n40320 , n40319 , n40132 );
and ( n40321 , n40318 , n40320 );
xor ( n40322 , n40162 , n40215 );
xor ( n40323 , n40322 , n40218 );
and ( n40324 , n40320 , n40323 );
and ( n40325 , n40318 , n40323 );
or ( n40326 , n40321 , n40324 , n40325 );
and ( n40327 , n40230 , n40326 );
xor ( n40328 , n40318 , n40320 );
xor ( n40329 , n40328 , n40323 );
and ( n40330 , n39432 , n40053 );
and ( n40331 , n39409 , n40051 );
nor ( n40332 , n40330 , n40331 );
xnor ( n40333 , n40332 , n39999 );
and ( n40334 , n39552 , n39760 );
and ( n40335 , n39493 , n39758 );
nor ( n40336 , n40334 , n40335 );
xnor ( n40337 , n40336 , n39742 );
and ( n40338 , n40333 , n40337 );
and ( n40339 , n39653 , n39678 );
and ( n40340 , n39620 , n39676 );
nor ( n40341 , n40339 , n40340 );
xnor ( n40342 , n40341 , n39643 );
and ( n40343 , n40337 , n40342 );
and ( n40344 , n40333 , n40342 );
or ( n40345 , n40338 , n40343 , n40344 );
xor ( n40346 , n40234 , n40238 );
xor ( n40347 , n40346 , n40243 );
and ( n40348 , n40345 , n40347 );
xor ( n40349 , n40273 , n40277 );
xor ( n40350 , n40349 , n40282 );
and ( n40351 , n40347 , n40350 );
and ( n40352 , n40345 , n40350 );
or ( n40353 , n40348 , n40351 , n40352 );
and ( n40354 , n39948 , n39480 );
and ( n40355 , n39867 , n39478 );
nor ( n40356 , n40354 , n40355 );
xnor ( n40357 , n40356 , n39462 );
and ( n40358 , n40148 , n39396 );
and ( n40359 , n40009 , n39394 );
nor ( n40360 , n40358 , n40359 );
xnor ( n40361 , n40360 , n39401 );
and ( n40362 , n40357 , n40361 );
and ( n40363 , n40186 , n39375 );
and ( n40364 , n40197 , n39373 );
nor ( n40365 , n40363 , n40364 );
xnor ( n40366 , n40365 , n39380 );
and ( n40367 , n40361 , n40366 );
and ( n40368 , n40357 , n40366 );
or ( n40369 , n40362 , n40367 , n40368 );
xor ( n40370 , n34949 , n39333 );
buf ( n567672 , n40370 );
buf ( n567673 , n567672 );
buf ( n40373 , n567673 );
and ( n40374 , n40373 , n39367 );
buf ( n40375 , n40374 );
buf ( n567677 , n1173 );
buf ( n40377 , n567677 );
buf ( n567679 , n1174 );
buf ( n40379 , n567679 );
and ( n40380 , n40377 , n40379 );
not ( n40381 , n40380 );
and ( n40382 , n40166 , n40381 );
not ( n40383 , n40382 );
and ( n40384 , n40375 , n40383 );
xor ( n40385 , n34947 , n39334 );
buf ( n567687 , n40385 );
buf ( n567688 , n567687 );
buf ( n40388 , n567688 );
and ( n40389 , n40388 , n39367 );
and ( n40390 , n40383 , n40389 );
and ( n40391 , n40375 , n40389 );
or ( n40392 , n40384 , n40390 , n40391 );
and ( n40393 , n40369 , n40392 );
and ( n40394 , n39472 , n39896 );
and ( n40395 , n39441 , n39894 );
nor ( n40396 , n40394 , n40395 );
xnor ( n40397 , n40396 , n39857 );
and ( n40398 , n40392 , n40397 );
and ( n40399 , n40369 , n40397 );
or ( n40400 , n40393 , n40398 , n40399 );
and ( n40401 , n39409 , n40258 );
and ( n40402 , n39365 , n40256 );
nor ( n40403 , n40401 , n40402 );
xnor ( n40404 , n40403 , n40169 );
and ( n40405 , n39620 , n39760 );
and ( n40406 , n39552 , n39758 );
nor ( n40407 , n40405 , n40406 );
xnor ( n40408 , n40407 , n39742 );
and ( n40409 , n40404 , n40408 );
xor ( n40410 , n40375 , n40383 );
xor ( n40411 , n40410 , n40389 );
and ( n40412 , n40408 , n40411 );
and ( n40413 , n40404 , n40411 );
or ( n40414 , n40409 , n40412 , n40413 );
xor ( n40415 , n40261 , n40265 );
xor ( n40416 , n40415 , n40270 );
and ( n40417 , n40414 , n40416 );
xor ( n40418 , n40289 , n40293 );
xor ( n40419 , n40418 , n40295 );
and ( n40420 , n40416 , n40419 );
and ( n40421 , n40414 , n40419 );
or ( n40422 , n40417 , n40420 , n40421 );
and ( n40423 , n40400 , n40422 );
xor ( n40424 , n40298 , n40300 );
xor ( n40425 , n40424 , n40303 );
and ( n40426 , n40422 , n40425 );
and ( n40427 , n40400 , n40425 );
or ( n40428 , n40423 , n40426 , n40427 );
and ( n40429 , n40353 , n40428 );
xor ( n40430 , n40246 , n40248 );
xor ( n40431 , n40430 , n40251 );
and ( n40432 , n40428 , n40431 );
and ( n40433 , n40353 , n40431 );
or ( n40434 , n40429 , n40432 , n40433 );
xor ( n40435 , n40207 , n40209 );
xor ( n40436 , n40435 , n40212 );
and ( n40437 , n40434 , n40436 );
xor ( n40438 , n40254 , n40312 );
xor ( n40439 , n40438 , n40315 );
and ( n40440 , n40436 , n40439 );
and ( n40441 , n40434 , n40439 );
or ( n40442 , n40437 , n40440 , n40441 );
and ( n40443 , n40329 , n40442 );
xor ( n40444 , n40434 , n40436 );
xor ( n40445 , n40444 , n40439 );
and ( n40446 , n39493 , n39896 );
and ( n40447 , n39472 , n39894 );
nor ( n40448 , n40446 , n40447 );
xnor ( n40449 , n40448 , n39857 );
and ( n40450 , n39670 , n39678 );
and ( n40451 , n39653 , n39676 );
nor ( n40452 , n40450 , n40451 );
xnor ( n40453 , n40452 , n39643 );
and ( n40454 , n40449 , n40453 );
and ( n40455 , n39795 , n39539 );
and ( n40456 , n39752 , n39537 );
nor ( n40457 , n40455 , n40456 );
xnor ( n40458 , n40457 , n39522 );
and ( n40459 , n40453 , n40458 );
and ( n40460 , n40449 , n40458 );
or ( n40461 , n40454 , n40459 , n40460 );
xor ( n40462 , n40333 , n40337 );
xor ( n40463 , n40462 , n40342 );
and ( n40464 , n40461 , n40463 );
xor ( n40465 , n40369 , n40392 );
xor ( n40466 , n40465 , n40397 );
and ( n40467 , n40463 , n40466 );
and ( n40468 , n40461 , n40466 );
or ( n40469 , n40464 , n40467 , n40468 );
xor ( n40470 , n40345 , n40347 );
xor ( n40471 , n40470 , n40350 );
and ( n40472 , n40469 , n40471 );
xor ( n40473 , n40400 , n40422 );
xor ( n40474 , n40473 , n40425 );
and ( n40475 , n40471 , n40474 );
and ( n40476 , n40469 , n40474 );
or ( n40477 , n40472 , n40475 , n40476 );
xor ( n40478 , n40285 , n40306 );
xor ( n40479 , n40478 , n40309 );
and ( n40480 , n40477 , n40479 );
xor ( n40481 , n40353 , n40428 );
xor ( n40482 , n40481 , n40431 );
and ( n40483 , n40479 , n40482 );
and ( n40484 , n40477 , n40482 );
or ( n40485 , n40480 , n40483 , n40484 );
and ( n40486 , n40445 , n40485 );
xor ( n40487 , n40477 , n40479 );
xor ( n40488 , n40487 , n40482 );
xor ( n40489 , n34951 , n39331 );
buf ( n567791 , n40489 );
buf ( n567792 , n567791 );
buf ( n40492 , n567792 );
and ( n40493 , n40492 , n39367 );
buf ( n40494 , n40493 );
buf ( n567796 , n1175 );
buf ( n40496 , n567796 );
buf ( n567798 , n1176 );
buf ( n40498 , n567798 );
and ( n40499 , n40496 , n40498 );
not ( n40500 , n40499 );
and ( n40501 , n40379 , n40500 );
not ( n40502 , n40501 );
and ( n40503 , n40494 , n40502 );
xor ( n40504 , n34950 , n39332 );
buf ( n567806 , n40504 );
buf ( n567807 , n567806 );
buf ( n40507 , n567807 );
and ( n40508 , n40507 , n39367 );
and ( n40509 , n40502 , n40508 );
and ( n40510 , n40494 , n40508 );
or ( n40511 , n40503 , n40509 , n40510 );
and ( n40512 , n40009 , n39480 );
and ( n40513 , n39948 , n39478 );
nor ( n40514 , n40512 , n40513 );
xnor ( n40515 , n40514 , n39462 );
and ( n40516 , n40511 , n40515 );
and ( n40517 , n40197 , n39396 );
and ( n40518 , n40148 , n39394 );
nor ( n40519 , n40517 , n40518 );
xnor ( n40520 , n40519 , n39401 );
and ( n40521 , n40515 , n40520 );
and ( n40522 , n40511 , n40520 );
or ( n40523 , n40516 , n40521 , n40522 );
xor ( n40524 , n40166 , n40377 );
xor ( n40525 , n40377 , n40379 );
not ( n40526 , n40525 );
and ( n40527 , n40524 , n40526 );
and ( n40528 , n39365 , n40527 );
not ( n40529 , n40528 );
xnor ( n40530 , n40529 , n40382 );
and ( n40531 , n40388 , n39375 );
and ( n40532 , n40186 , n39373 );
nor ( n40533 , n40531 , n40532 );
xnor ( n40534 , n40533 , n39380 );
and ( n40535 , n40530 , n40534 );
not ( n40536 , n40374 );
and ( n40537 , n40534 , n40536 );
and ( n40538 , n40530 , n40536 );
or ( n40539 , n40535 , n40537 , n40538 );
and ( n40540 , n40523 , n40539 );
and ( n40541 , n39441 , n40053 );
and ( n40542 , n39432 , n40051 );
nor ( n40543 , n40541 , n40542 );
xnor ( n40544 , n40543 , n39999 );
and ( n40545 , n40539 , n40544 );
and ( n40546 , n40523 , n40544 );
or ( n40547 , n40540 , n40545 , n40546 );
and ( n40548 , n39552 , n39896 );
and ( n40549 , n39493 , n39894 );
nor ( n40550 , n40548 , n40549 );
xnor ( n40551 , n40550 , n39857 );
and ( n40552 , n39752 , n39678 );
and ( n40553 , n39670 , n39676 );
nor ( n40554 , n40552 , n40553 );
xnor ( n40555 , n40554 , n39643 );
and ( n40556 , n40551 , n40555 );
and ( n40557 , n39867 , n39539 );
and ( n40558 , n39795 , n39537 );
nor ( n40559 , n40557 , n40558 );
xnor ( n40560 , n40559 , n39522 );
and ( n40561 , n40555 , n40560 );
and ( n40562 , n40551 , n40560 );
or ( n40563 , n40556 , n40561 , n40562 );
and ( n40564 , n39432 , n40258 );
and ( n40565 , n39409 , n40256 );
nor ( n40566 , n40564 , n40565 );
xnor ( n40567 , n40566 , n40169 );
and ( n40568 , n39472 , n40053 );
and ( n40569 , n39441 , n40051 );
nor ( n40570 , n40568 , n40569 );
xnor ( n40571 , n40570 , n39999 );
and ( n40572 , n40567 , n40571 );
and ( n40573 , n39653 , n39760 );
and ( n40574 , n39620 , n39758 );
nor ( n40575 , n40573 , n40574 );
xnor ( n40576 , n40575 , n39742 );
and ( n40577 , n40571 , n40576 );
and ( n40578 , n40567 , n40576 );
or ( n40579 , n40572 , n40577 , n40578 );
and ( n40580 , n40563 , n40579 );
xor ( n40581 , n40449 , n40453 );
xor ( n40582 , n40581 , n40458 );
and ( n40583 , n40579 , n40582 );
and ( n40584 , n40563 , n40582 );
or ( n40585 , n40580 , n40583 , n40584 );
and ( n40586 , n40547 , n40585 );
xor ( n40587 , n40414 , n40416 );
xor ( n40588 , n40587 , n40419 );
and ( n40589 , n40585 , n40588 );
and ( n40590 , n40547 , n40588 );
or ( n40591 , n40586 , n40589 , n40590 );
and ( n40592 , n39670 , n39760 );
and ( n40593 , n39653 , n39758 );
nor ( n40594 , n40592 , n40593 );
xnor ( n40595 , n40594 , n39742 );
and ( n40596 , n39948 , n39539 );
and ( n40597 , n39867 , n39537 );
nor ( n40598 , n40596 , n40597 );
xnor ( n40599 , n40598 , n39522 );
and ( n40600 , n40595 , n40599 );
and ( n40601 , n40148 , n39480 );
and ( n40602 , n40009 , n39478 );
nor ( n40603 , n40601 , n40602 );
xnor ( n40604 , n40603 , n39462 );
and ( n40605 , n40599 , n40604 );
and ( n40606 , n40595 , n40604 );
or ( n40607 , n40600 , n40605 , n40606 );
and ( n40608 , n40186 , n39396 );
and ( n40609 , n40197 , n39394 );
nor ( n40610 , n40608 , n40609 );
xnor ( n40611 , n40610 , n39401 );
and ( n40612 , n40373 , n39375 );
and ( n40613 , n40388 , n39373 );
nor ( n40614 , n40612 , n40613 );
xnor ( n40615 , n40614 , n39380 );
and ( n40616 , n40611 , n40615 );
xor ( n40617 , n40494 , n40502 );
xor ( n40618 , n40617 , n40508 );
and ( n40619 , n40615 , n40618 );
and ( n40620 , n40611 , n40618 );
or ( n40621 , n40616 , n40619 , n40620 );
and ( n40622 , n40607 , n40621 );
xor ( n40623 , n40530 , n40534 );
xor ( n40624 , n40623 , n40536 );
and ( n40625 , n40621 , n40624 );
and ( n40626 , n40607 , n40624 );
or ( n40627 , n40622 , n40625 , n40626 );
xor ( n40628 , n40357 , n40361 );
xor ( n40629 , n40628 , n40366 );
and ( n40630 , n40627 , n40629 );
xor ( n40631 , n40404 , n40408 );
xor ( n40632 , n40631 , n40411 );
and ( n40633 , n40629 , n40632 );
and ( n40634 , n40627 , n40632 );
or ( n40635 , n40630 , n40633 , n40634 );
and ( n40636 , n39409 , n40527 );
and ( n40637 , n39365 , n40525 );
nor ( n40638 , n40636 , n40637 );
xnor ( n40639 , n40638 , n40382 );
and ( n40640 , n39493 , n40053 );
and ( n40641 , n39472 , n40051 );
nor ( n40642 , n40640 , n40641 );
xnor ( n40643 , n40642 , n39999 );
and ( n40644 , n40639 , n40643 );
and ( n40645 , n39795 , n39678 );
and ( n40646 , n39752 , n39676 );
nor ( n40647 , n40645 , n40646 );
xnor ( n40648 , n40647 , n39643 );
and ( n40649 , n40643 , n40648 );
and ( n40650 , n40639 , n40648 );
or ( n40651 , n40644 , n40649 , n40650 );
and ( n40652 , n40388 , n39396 );
and ( n40653 , n40186 , n39394 );
nor ( n40654 , n40652 , n40653 );
xnor ( n40655 , n40654 , n39401 );
and ( n40656 , n40507 , n39375 );
and ( n40657 , n40373 , n39373 );
nor ( n40658 , n40656 , n40657 );
xnor ( n40659 , n40658 , n39380 );
and ( n40660 , n40655 , n40659 );
not ( n40661 , n40493 );
and ( n40662 , n40659 , n40661 );
and ( n40663 , n40655 , n40661 );
or ( n40664 , n40660 , n40662 , n40663 );
and ( n40665 , n39441 , n40258 );
and ( n40666 , n39432 , n40256 );
nor ( n40667 , n40665 , n40666 );
xnor ( n40668 , n40667 , n40169 );
and ( n40669 , n40664 , n40668 );
and ( n40670 , n39620 , n39896 );
and ( n40671 , n39552 , n39894 );
nor ( n40672 , n40670 , n40671 );
xnor ( n40673 , n40672 , n39857 );
and ( n40674 , n40668 , n40673 );
and ( n40675 , n40664 , n40673 );
or ( n40676 , n40669 , n40674 , n40675 );
and ( n40677 , n40651 , n40676 );
xor ( n40678 , n40511 , n40515 );
xor ( n40679 , n40678 , n40520 );
and ( n40680 , n40676 , n40679 );
and ( n40681 , n40651 , n40679 );
or ( n40682 , n40677 , n40680 , n40681 );
xor ( n40683 , n40523 , n40539 );
xor ( n40684 , n40683 , n40544 );
and ( n40685 , n40682 , n40684 );
xor ( n40686 , n40563 , n40579 );
xor ( n40687 , n40686 , n40582 );
and ( n40688 , n40684 , n40687 );
and ( n40689 , n40682 , n40687 );
or ( n40690 , n40685 , n40688 , n40689 );
and ( n40691 , n40635 , n40690 );
xor ( n40692 , n40461 , n40463 );
xor ( n40693 , n40692 , n40466 );
and ( n40694 , n40690 , n40693 );
and ( n40695 , n40635 , n40693 );
or ( n40696 , n40691 , n40694 , n40695 );
and ( n40697 , n40591 , n40696 );
xor ( n40698 , n40469 , n40471 );
xor ( n40699 , n40698 , n40474 );
and ( n40700 , n40696 , n40699 );
and ( n40701 , n40591 , n40699 );
or ( n40702 , n40697 , n40700 , n40701 );
and ( n40703 , n40488 , n40702 );
xor ( n40704 , n40591 , n40696 );
xor ( n40705 , n40704 , n40699 );
and ( n40706 , n39752 , n39760 );
and ( n40707 , n39670 , n39758 );
nor ( n40708 , n40706 , n40707 );
xnor ( n40709 , n40708 , n39742 );
and ( n40710 , n39867 , n39678 );
and ( n40711 , n39795 , n39676 );
nor ( n40712 , n40710 , n40711 );
xnor ( n40713 , n40712 , n39643 );
and ( n40714 , n40709 , n40713 );
and ( n40715 , n40009 , n39539 );
and ( n40716 , n39948 , n39537 );
nor ( n40717 , n40715 , n40716 );
xnor ( n40718 , n40717 , n39522 );
and ( n40719 , n40713 , n40718 );
and ( n40720 , n40709 , n40718 );
or ( n40721 , n40714 , n40719 , n40720 );
buf ( n568023 , n1177 );
buf ( n40723 , n568023 );
buf ( n568025 , n1178 );
buf ( n40725 , n568025 );
and ( n40726 , n40723 , n40725 );
not ( n40727 , n40726 );
and ( n40728 , n40498 , n40727 );
not ( n40729 , n40728 );
and ( n40730 , n40492 , n39375 );
and ( n40731 , n40507 , n39373 );
nor ( n40732 , n40730 , n40731 );
xnor ( n40733 , n40732 , n39380 );
and ( n40734 , n40729 , n40733 );
xor ( n40735 , n34954 , n39329 );
buf ( n568037 , n40735 );
buf ( n568038 , n568037 );
buf ( n40738 , n568038 );
and ( n40739 , n40738 , n39367 );
and ( n40740 , n40733 , n40739 );
and ( n40741 , n40729 , n40739 );
or ( n40742 , n40734 , n40740 , n40741 );
xor ( n40743 , n40379 , n40496 );
xor ( n40744 , n40496 , n40498 );
not ( n40745 , n40744 );
and ( n40746 , n40743 , n40745 );
and ( n40747 , n39365 , n40746 );
not ( n40748 , n40747 );
xnor ( n40749 , n40748 , n40501 );
and ( n40750 , n40742 , n40749 );
and ( n40751 , n40197 , n39480 );
and ( n40752 , n40148 , n39478 );
nor ( n40753 , n40751 , n40752 );
xnor ( n40754 , n40753 , n39462 );
and ( n40755 , n40749 , n40754 );
and ( n40756 , n40742 , n40754 );
or ( n40757 , n40750 , n40755 , n40756 );
and ( n40758 , n40721 , n40757 );
xor ( n40759 , n40611 , n40615 );
xor ( n40760 , n40759 , n40618 );
and ( n40761 , n40757 , n40760 );
and ( n40762 , n40721 , n40760 );
or ( n40763 , n40758 , n40761 , n40762 );
xor ( n40764 , n40551 , n40555 );
xor ( n40765 , n40764 , n40560 );
and ( n40766 , n40763 , n40765 );
xor ( n40767 , n40567 , n40571 );
xor ( n40768 , n40767 , n40576 );
and ( n40769 , n40765 , n40768 );
and ( n40770 , n40763 , n40768 );
or ( n40771 , n40766 , n40769 , n40770 );
and ( n40772 , n39432 , n40527 );
and ( n40773 , n39409 , n40525 );
nor ( n40774 , n40772 , n40773 );
xnor ( n40775 , n40774 , n40382 );
and ( n40776 , n39552 , n40053 );
and ( n40777 , n39493 , n40051 );
nor ( n40778 , n40776 , n40777 );
xnor ( n40779 , n40778 , n39999 );
and ( n40780 , n40775 , n40779 );
and ( n40781 , n39653 , n39896 );
and ( n40782 , n39620 , n39894 );
nor ( n40783 , n40781 , n40782 );
xnor ( n40784 , n40783 , n39857 );
and ( n40785 , n40779 , n40784 );
and ( n40786 , n40775 , n40784 );
or ( n40787 , n40780 , n40785 , n40786 );
and ( n40788 , n40738 , n39375 );
and ( n40789 , n40492 , n39373 );
nor ( n40790 , n40788 , n40789 );
xnor ( n40791 , n40790 , n39380 );
buf ( n40792 , n40791 );
and ( n40793 , n40373 , n39396 );
and ( n40794 , n40388 , n39394 );
nor ( n40795 , n40793 , n40794 );
xnor ( n40796 , n40795 , n39401 );
and ( n40797 , n40792 , n40796 );
xor ( n40798 , n40729 , n40733 );
xor ( n40799 , n40798 , n40739 );
and ( n40800 , n40796 , n40799 );
and ( n40801 , n40792 , n40799 );
or ( n40802 , n40797 , n40800 , n40801 );
and ( n40803 , n39472 , n40258 );
and ( n40804 , n39441 , n40256 );
nor ( n40805 , n40803 , n40804 );
xnor ( n40806 , n40805 , n40169 );
and ( n40807 , n40802 , n40806 );
xor ( n40808 , n40655 , n40659 );
xor ( n40809 , n40808 , n40661 );
and ( n40810 , n40806 , n40809 );
and ( n40811 , n40802 , n40809 );
or ( n40812 , n40807 , n40810 , n40811 );
and ( n40813 , n40787 , n40812 );
xor ( n40814 , n40595 , n40599 );
xor ( n40815 , n40814 , n40604 );
and ( n40816 , n40812 , n40815 );
and ( n40817 , n40787 , n40815 );
or ( n40818 , n40813 , n40816 , n40817 );
xor ( n40819 , n40607 , n40621 );
xor ( n40820 , n40819 , n40624 );
and ( n40821 , n40818 , n40820 );
xor ( n40822 , n40651 , n40676 );
xor ( n40823 , n40822 , n40679 );
and ( n40824 , n40820 , n40823 );
and ( n40825 , n40818 , n40823 );
or ( n40826 , n40821 , n40824 , n40825 );
and ( n40827 , n40771 , n40826 );
xor ( n40828 , n40627 , n40629 );
xor ( n40829 , n40828 , n40632 );
and ( n40830 , n40826 , n40829 );
and ( n40831 , n40771 , n40829 );
or ( n40832 , n40827 , n40830 , n40831 );
xor ( n40833 , n40547 , n40585 );
xor ( n40834 , n40833 , n40588 );
and ( n40835 , n40832 , n40834 );
xor ( n40836 , n40635 , n40690 );
xor ( n40837 , n40836 , n40693 );
and ( n40838 , n40834 , n40837 );
and ( n40839 , n40832 , n40837 );
or ( n40840 , n40835 , n40838 , n40839 );
and ( n40841 , n40705 , n40840 );
xor ( n40842 , n40832 , n40834 );
xor ( n40843 , n40842 , n40837 );
and ( n40844 , n39670 , n39896 );
and ( n40845 , n39653 , n39894 );
nor ( n40846 , n40844 , n40845 );
xnor ( n40847 , n40846 , n39857 );
and ( n40848 , n39795 , n39760 );
and ( n40849 , n39752 , n39758 );
nor ( n40850 , n40848 , n40849 );
xnor ( n40851 , n40850 , n39742 );
and ( n40852 , n40847 , n40851 );
and ( n40853 , n40186 , n39480 );
and ( n40854 , n40197 , n39478 );
nor ( n40855 , n40853 , n40854 );
xnor ( n40856 , n40855 , n39462 );
and ( n40857 , n40851 , n40856 );
and ( n40858 , n40847 , n40856 );
or ( n40859 , n40852 , n40857 , n40858 );
and ( n40860 , n40507 , n39396 );
and ( n40861 , n40373 , n39394 );
nor ( n40862 , n40860 , n40861 );
xnor ( n40863 , n40862 , n39401 );
not ( n40864 , n40791 );
and ( n40865 , n40863 , n40864 );
xor ( n40866 , n34956 , n39328 );
buf ( n568168 , n40866 );
buf ( n568169 , n568168 );
buf ( n40869 , n568169 );
and ( n40870 , n40869 , n39367 );
and ( n40871 , n40864 , n40870 );
and ( n40872 , n40863 , n40870 );
or ( n40873 , n40865 , n40871 , n40872 );
and ( n40874 , n39948 , n39678 );
and ( n40875 , n39867 , n39676 );
nor ( n40876 , n40874 , n40875 );
xnor ( n40877 , n40876 , n39643 );
and ( n40878 , n40873 , n40877 );
and ( n40879 , n40148 , n39539 );
and ( n40880 , n40009 , n39537 );
nor ( n40881 , n40879 , n40880 );
xnor ( n40882 , n40881 , n39522 );
and ( n40883 , n40877 , n40882 );
and ( n40884 , n40873 , n40882 );
or ( n40885 , n40878 , n40883 , n40884 );
and ( n40886 , n40859 , n40885 );
xor ( n40887 , n40742 , n40749 );
xor ( n40888 , n40887 , n40754 );
and ( n40889 , n40885 , n40888 );
and ( n40890 , n40859 , n40888 );
or ( n40891 , n40886 , n40889 , n40890 );
xor ( n40892 , n40639 , n40643 );
xor ( n40893 , n40892 , n40648 );
and ( n40894 , n40891 , n40893 );
xor ( n40895 , n40664 , n40668 );
xor ( n40896 , n40895 , n40673 );
and ( n40897 , n40893 , n40896 );
and ( n40898 , n40891 , n40896 );
or ( n40899 , n40894 , n40897 , n40898 );
and ( n40900 , n39409 , n40746 );
and ( n40901 , n39365 , n40744 );
nor ( n40902 , n40900 , n40901 );
xnor ( n40903 , n40902 , n40501 );
and ( n40904 , n39441 , n40527 );
and ( n40905 , n39432 , n40525 );
nor ( n40906 , n40904 , n40905 );
xnor ( n40907 , n40906 , n40382 );
and ( n40908 , n40903 , n40907 );
and ( n40909 , n39493 , n40258 );
and ( n40910 , n39472 , n40256 );
nor ( n40911 , n40909 , n40910 );
xnor ( n40912 , n40911 , n40169 );
and ( n40913 , n40907 , n40912 );
and ( n40914 , n40903 , n40912 );
or ( n40915 , n40908 , n40913 , n40914 );
xor ( n40916 , n40709 , n40713 );
xor ( n40917 , n40916 , n40718 );
and ( n40918 , n40915 , n40917 );
xor ( n40919 , n40775 , n40779 );
xor ( n40920 , n40919 , n40784 );
and ( n40921 , n40917 , n40920 );
and ( n40922 , n40915 , n40920 );
or ( n40923 , n40918 , n40921 , n40922 );
xor ( n40924 , n40787 , n40812 );
xor ( n40925 , n40924 , n40815 );
and ( n40926 , n40923 , n40925 );
xor ( n40927 , n40721 , n40757 );
xor ( n40928 , n40927 , n40760 );
and ( n40929 , n40925 , n40928 );
and ( n40930 , n40923 , n40928 );
or ( n40931 , n40926 , n40929 , n40930 );
and ( n40932 , n40899 , n40931 );
xor ( n40933 , n40763 , n40765 );
xor ( n40934 , n40933 , n40768 );
and ( n40935 , n40931 , n40934 );
and ( n40936 , n40899 , n40934 );
or ( n40937 , n40932 , n40935 , n40936 );
xor ( n40938 , n40682 , n40684 );
xor ( n40939 , n40938 , n40687 );
and ( n40940 , n40937 , n40939 );
xor ( n40941 , n40771 , n40826 );
xor ( n40942 , n40941 , n40829 );
and ( n40943 , n40939 , n40942 );
and ( n40944 , n40937 , n40942 );
or ( n40945 , n40940 , n40943 , n40944 );
and ( n40946 , n40843 , n40945 );
xor ( n40947 , n40937 , n40939 );
xor ( n40948 , n40947 , n40942 );
and ( n40949 , n39432 , n40746 );
and ( n40950 , n39409 , n40744 );
nor ( n40951 , n40949 , n40950 );
xnor ( n40952 , n40951 , n40501 );
and ( n40953 , n39552 , n40258 );
and ( n40954 , n39493 , n40256 );
nor ( n40955 , n40953 , n40954 );
xnor ( n40956 , n40955 , n40169 );
and ( n40957 , n40952 , n40956 );
and ( n40958 , n39653 , n40053 );
and ( n40959 , n39620 , n40051 );
nor ( n40960 , n40958 , n40959 );
xnor ( n40961 , n40960 , n39999 );
and ( n40962 , n40956 , n40961 );
and ( n40963 , n40952 , n40961 );
or ( n40964 , n40957 , n40962 , n40963 );
xor ( n40965 , n40847 , n40851 );
xor ( n40966 , n40965 , n40856 );
and ( n40967 , n40964 , n40966 );
xor ( n40968 , n40903 , n40907 );
xor ( n40969 , n40968 , n40912 );
and ( n40970 , n40966 , n40969 );
and ( n40971 , n40964 , n40969 );
or ( n40972 , n40967 , n40970 , n40971 );
xor ( n40973 , n40915 , n40917 );
xor ( n40974 , n40973 , n40920 );
and ( n40975 , n40972 , n40974 );
xor ( n40976 , n40859 , n40885 );
xor ( n40977 , n40976 , n40888 );
and ( n40978 , n40974 , n40977 );
and ( n40979 , n40972 , n40977 );
or ( n40980 , n40975 , n40978 , n40979 );
and ( n40981 , n40373 , n39480 );
and ( n40982 , n40388 , n39478 );
nor ( n40983 , n40981 , n40982 );
xnor ( n40984 , n40983 , n39462 );
and ( n40985 , n40492 , n39396 );
and ( n40986 , n40507 , n39394 );
nor ( n40987 , n40985 , n40986 );
xnor ( n40988 , n40987 , n39401 );
and ( n40989 , n40984 , n40988 );
and ( n40990 , n40869 , n39375 );
and ( n40991 , n40738 , n39373 );
nor ( n40992 , n40990 , n40991 );
xnor ( n40993 , n40992 , n39380 );
and ( n40994 , n40988 , n40993 );
and ( n40995 , n40984 , n40993 );
or ( n40996 , n40989 , n40994 , n40995 );
and ( n40997 , n40009 , n39678 );
and ( n40998 , n39948 , n39676 );
nor ( n40999 , n40997 , n40998 );
xnor ( n41000 , n40999 , n39643 );
and ( n41001 , n40996 , n41000 );
and ( n41002 , n40197 , n39539 );
and ( n41003 , n40148 , n39537 );
nor ( n41004 , n41002 , n41003 );
xnor ( n41005 , n41004 , n39522 );
and ( n41006 , n41000 , n41005 );
and ( n41007 , n40996 , n41005 );
or ( n41008 , n41001 , n41006 , n41007 );
and ( n41009 , n39752 , n39896 );
and ( n41010 , n39670 , n39894 );
nor ( n41011 , n41009 , n41010 );
xnor ( n41012 , n41011 , n39857 );
and ( n41013 , n39867 , n39760 );
and ( n41014 , n39795 , n39758 );
nor ( n41015 , n41013 , n41014 );
xnor ( n41016 , n41015 , n39742 );
and ( n41017 , n41012 , n41016 );
xor ( n41018 , n40863 , n40864 );
xor ( n41019 , n41018 , n40870 );
and ( n41020 , n41016 , n41019 );
and ( n41021 , n41012 , n41019 );
or ( n41022 , n41017 , n41020 , n41021 );
and ( n41023 , n41008 , n41022 );
xor ( n41024 , n40873 , n40877 );
xor ( n41025 , n41024 , n40882 );
and ( n41026 , n41022 , n41025 );
and ( n41027 , n41008 , n41025 );
or ( n41028 , n41023 , n41026 , n41027 );
xor ( n41029 , n36949 , n39325 );
buf ( n568331 , n41029 );
buf ( n568332 , n568331 );
buf ( n41032 , n568332 );
and ( n41033 , n41032 , n39367 );
buf ( n41034 , n41033 );
buf ( n568336 , n1179 );
buf ( n41036 , n568336 );
buf ( n568338 , n1180 );
buf ( n41038 , n568338 );
and ( n41039 , n41036 , n41038 );
not ( n41040 , n41039 );
and ( n41041 , n40725 , n41040 );
not ( n41042 , n41041 );
and ( n41043 , n41034 , n41042 );
xor ( n41044 , n36947 , n39326 );
buf ( n568346 , n41044 );
buf ( n568347 , n568346 );
buf ( n41047 , n568347 );
and ( n41048 , n41047 , n39367 );
and ( n41049 , n41042 , n41048 );
and ( n41050 , n41034 , n41048 );
or ( n41051 , n41043 , n41049 , n41050 );
xor ( n41052 , n40498 , n40723 );
xor ( n41053 , n40723 , n40725 );
not ( n41054 , n41053 );
and ( n41055 , n41052 , n41054 );
and ( n41056 , n39365 , n41055 );
not ( n41057 , n41056 );
xnor ( n41058 , n41057 , n40728 );
and ( n41059 , n41051 , n41058 );
and ( n41060 , n40388 , n39480 );
and ( n41061 , n40186 , n39478 );
nor ( n41062 , n41060 , n41061 );
xnor ( n41063 , n41062 , n39462 );
and ( n41064 , n41058 , n41063 );
and ( n41065 , n41051 , n41063 );
or ( n41066 , n41059 , n41064 , n41065 );
and ( n41067 , n39620 , n40053 );
and ( n41068 , n39552 , n40051 );
nor ( n41069 , n41067 , n41068 );
xnor ( n41070 , n41069 , n39999 );
and ( n41071 , n41066 , n41070 );
xor ( n41072 , n40792 , n40796 );
xor ( n41073 , n41072 , n40799 );
and ( n41074 , n41070 , n41073 );
and ( n41075 , n41066 , n41073 );
or ( n41076 , n41071 , n41074 , n41075 );
and ( n41077 , n41028 , n41076 );
xor ( n41078 , n40802 , n40806 );
xor ( n41079 , n41078 , n40809 );
and ( n41080 , n41076 , n41079 );
and ( n41081 , n41028 , n41079 );
or ( n41082 , n41077 , n41080 , n41081 );
and ( n41083 , n40980 , n41082 );
xor ( n41084 , n40891 , n40893 );
xor ( n41085 , n41084 , n40896 );
and ( n41086 , n41082 , n41085 );
and ( n41087 , n40980 , n41085 );
or ( n41088 , n41083 , n41086 , n41087 );
xor ( n41089 , n40818 , n40820 );
xor ( n41090 , n41089 , n40823 );
and ( n41091 , n41088 , n41090 );
xor ( n41092 , n40899 , n40931 );
xor ( n41093 , n41092 , n40934 );
and ( n41094 , n41090 , n41093 );
and ( n41095 , n41088 , n41093 );
or ( n41096 , n41091 , n41094 , n41095 );
and ( n41097 , n40948 , n41096 );
xor ( n41098 , n41088 , n41090 );
xor ( n41099 , n41098 , n41093 );
and ( n41100 , n39493 , n40527 );
and ( n41101 , n39472 , n40525 );
nor ( n41102 , n41100 , n41101 );
xnor ( n41103 , n41102 , n40382 );
and ( n41104 , n39795 , n39896 );
and ( n41105 , n39752 , n39894 );
nor ( n41106 , n41104 , n41105 );
xnor ( n41107 , n41106 , n39857 );
and ( n41108 , n41103 , n41107 );
xor ( n41109 , n40984 , n40988 );
xor ( n41110 , n41109 , n40993 );
and ( n41111 , n41107 , n41110 );
and ( n41112 , n41103 , n41110 );
or ( n41113 , n41108 , n41111 , n41112 );
xor ( n41114 , n40952 , n40956 );
xor ( n41115 , n41114 , n40961 );
and ( n41116 , n41113 , n41115 );
xor ( n41117 , n40996 , n41000 );
xor ( n41118 , n41117 , n41005 );
and ( n41119 , n41115 , n41118 );
and ( n41120 , n41113 , n41118 );
or ( n41121 , n41116 , n41119 , n41120 );
xor ( n41122 , n40964 , n40966 );
xor ( n41123 , n41122 , n40969 );
and ( n41124 , n41121 , n41123 );
xor ( n41125 , n41008 , n41022 );
xor ( n41126 , n41125 , n41025 );
and ( n41127 , n41123 , n41126 );
and ( n41128 , n41121 , n41126 );
or ( n41129 , n41124 , n41127 , n41128 );
and ( n41130 , n40738 , n39396 );
and ( n41131 , n40492 , n39394 );
nor ( n41132 , n41130 , n41131 );
xnor ( n41133 , n41132 , n39401 );
and ( n41134 , n41047 , n39375 );
and ( n41135 , n40869 , n39373 );
nor ( n41136 , n41134 , n41135 );
xnor ( n41137 , n41136 , n39380 );
and ( n41138 , n41133 , n41137 );
not ( n41139 , n41033 );
and ( n41140 , n41137 , n41139 );
and ( n41141 , n41133 , n41139 );
or ( n41142 , n41138 , n41140 , n41141 );
and ( n41143 , n40148 , n39678 );
and ( n41144 , n40009 , n39676 );
nor ( n41145 , n41143 , n41144 );
xnor ( n41146 , n41145 , n39643 );
and ( n41147 , n41142 , n41146 );
xor ( n41148 , n41034 , n41042 );
xor ( n41149 , n41148 , n41048 );
and ( n41150 , n41146 , n41149 );
and ( n41151 , n41142 , n41149 );
or ( n41152 , n41147 , n41150 , n41151 );
and ( n41153 , n39472 , n40527 );
and ( n41154 , n39441 , n40525 );
nor ( n41155 , n41153 , n41154 );
xnor ( n41156 , n41155 , n40382 );
and ( n41157 , n41152 , n41156 );
xor ( n41158 , n41051 , n41058 );
xor ( n41159 , n41158 , n41063 );
and ( n41160 , n41156 , n41159 );
and ( n41161 , n41152 , n41159 );
or ( n41162 , n41157 , n41160 , n41161 );
and ( n41163 , n39670 , n40053 );
and ( n41164 , n39653 , n40051 );
nor ( n41165 , n41163 , n41164 );
xnor ( n41166 , n41165 , n39999 );
and ( n41167 , n39948 , n39760 );
and ( n41168 , n39867 , n39758 );
nor ( n41169 , n41167 , n41168 );
xnor ( n41170 , n41169 , n39742 );
and ( n41171 , n41166 , n41170 );
and ( n41172 , n40186 , n39539 );
and ( n41173 , n40197 , n39537 );
nor ( n41174 , n41172 , n41173 );
xnor ( n41175 , n41174 , n39522 );
and ( n41176 , n41170 , n41175 );
and ( n41177 , n41166 , n41175 );
or ( n41178 , n41171 , n41176 , n41177 );
xor ( n41179 , n36952 , n39323 );
buf ( n568481 , n41179 );
buf ( n568482 , n568481 );
buf ( n41182 , n568482 );
and ( n41183 , n41182 , n39375 );
and ( n41184 , n41032 , n39373 );
nor ( n41185 , n41183 , n41184 );
xnor ( n41186 , n41185 , n39380 );
buf ( n41187 , n41186 );
buf ( n568489 , n1181 );
buf ( n41189 , n568489 );
buf ( n568491 , n1182 );
buf ( n41191 , n568491 );
and ( n41192 , n41189 , n41191 );
not ( n41193 , n41192 );
and ( n41194 , n41038 , n41193 );
not ( n41195 , n41194 );
and ( n41196 , n41187 , n41195 );
and ( n41197 , n41182 , n39367 );
and ( n41198 , n41195 , n41197 );
and ( n41199 , n41187 , n41197 );
or ( n41200 , n41196 , n41198 , n41199 );
and ( n41201 , n40388 , n39539 );
and ( n41202 , n40186 , n39537 );
nor ( n41203 , n41201 , n41202 );
xnor ( n41204 , n41203 , n39522 );
and ( n41205 , n41200 , n41204 );
and ( n41206 , n40507 , n39480 );
and ( n41207 , n40373 , n39478 );
nor ( n41208 , n41206 , n41207 );
xnor ( n41209 , n41208 , n39462 );
and ( n41210 , n41204 , n41209 );
and ( n41211 , n41200 , n41209 );
or ( n41212 , n41205 , n41210 , n41211 );
and ( n41213 , n39409 , n41055 );
and ( n41214 , n39365 , n41053 );
nor ( n41215 , n41213 , n41214 );
xnor ( n41216 , n41215 , n40728 );
and ( n41217 , n41212 , n41216 );
and ( n41218 , n39620 , n40258 );
and ( n41219 , n39552 , n40256 );
nor ( n41220 , n41218 , n41219 );
xnor ( n41221 , n41220 , n40169 );
and ( n41222 , n41216 , n41221 );
and ( n41223 , n41212 , n41221 );
or ( n41224 , n41217 , n41222 , n41223 );
and ( n41225 , n41178 , n41224 );
xor ( n41226 , n41012 , n41016 );
xor ( n41227 , n41226 , n41019 );
and ( n41228 , n41224 , n41227 );
and ( n41229 , n41178 , n41227 );
or ( n41230 , n41225 , n41228 , n41229 );
and ( n41231 , n41162 , n41230 );
xor ( n41232 , n41066 , n41070 );
xor ( n41233 , n41232 , n41073 );
and ( n41234 , n41230 , n41233 );
and ( n41235 , n41162 , n41233 );
or ( n41236 , n41231 , n41234 , n41235 );
and ( n41237 , n41129 , n41236 );
xor ( n41238 , n41028 , n41076 );
xor ( n41239 , n41238 , n41079 );
and ( n41240 , n41236 , n41239 );
and ( n41241 , n41129 , n41239 );
or ( n41242 , n41237 , n41240 , n41241 );
xor ( n41243 , n40980 , n41082 );
xor ( n41244 , n41243 , n41085 );
and ( n41245 , n41242 , n41244 );
xor ( n41246 , n40923 , n40925 );
xor ( n41247 , n41246 , n40928 );
and ( n41248 , n41244 , n41247 );
and ( n41249 , n41242 , n41247 );
or ( n41250 , n41245 , n41248 , n41249 );
and ( n41251 , n41099 , n41250 );
xor ( n41252 , n41242 , n41244 );
xor ( n41253 , n41252 , n41247 );
xor ( n41254 , n40972 , n40974 );
xor ( n41255 , n41254 , n40977 );
xor ( n41256 , n41129 , n41236 );
xor ( n41257 , n41256 , n41239 );
and ( n41258 , n41255 , n41257 );
and ( n41259 , n41253 , n41258 );
and ( n41260 , n40197 , n39678 );
and ( n41261 , n40148 , n39676 );
nor ( n41262 , n41260 , n41261 );
xnor ( n41263 , n41262 , n39643 );
buf ( n41264 , n41263 );
buf ( n41265 , n41264 );
buf ( n41266 , n41265 );
buf ( n41267 , n41266 );
xor ( n41268 , n41121 , n41123 );
xor ( n41269 , n41268 , n41126 );
not ( n41270 , n41266 );
and ( n41271 , n41269 , n41270 );
not ( n41272 , n41265 );
and ( n41273 , n40492 , n39480 );
and ( n41274 , n40507 , n39478 );
nor ( n41275 , n41273 , n41274 );
xnor ( n41276 , n41275 , n39462 );
and ( n41277 , n40869 , n39396 );
and ( n41278 , n40738 , n39394 );
nor ( n41279 , n41277 , n41278 );
xnor ( n41280 , n41279 , n39401 );
and ( n41281 , n41276 , n41280 );
and ( n41282 , n41032 , n39375 );
and ( n41283 , n41047 , n39373 );
nor ( n41284 , n41282 , n41283 );
xnor ( n41285 , n41284 , n39380 );
and ( n41286 , n41280 , n41285 );
and ( n41287 , n41276 , n41285 );
or ( n41288 , n41281 , n41286 , n41287 );
xor ( n41289 , n40725 , n41036 );
xor ( n41290 , n41036 , n41038 );
not ( n41291 , n41290 );
and ( n41292 , n41289 , n41291 );
and ( n41293 , n39365 , n41292 );
not ( n41294 , n41293 );
xnor ( n41295 , n41294 , n41041 );
and ( n41296 , n41288 , n41295 );
xor ( n41297 , n41133 , n41137 );
xor ( n41298 , n41297 , n41139 );
and ( n41299 , n41295 , n41298 );
and ( n41300 , n41288 , n41298 );
or ( n41301 , n41296 , n41299 , n41300 );
and ( n41302 , n39441 , n40746 );
and ( n41303 , n39432 , n40744 );
nor ( n41304 , n41302 , n41303 );
xnor ( n41305 , n41304 , n40501 );
and ( n41306 , n41301 , n41305 );
and ( n41307 , n41272 , n41306 );
xor ( n41308 , n41152 , n41156 );
xor ( n41309 , n41308 , n41159 );
and ( n41310 , n41306 , n41309 );
and ( n41311 , n41272 , n41309 );
or ( n41312 , n41307 , n41310 , n41311 );
and ( n41313 , n41270 , n41312 );
and ( n41314 , n41269 , n41312 );
or ( n41315 , n41271 , n41313 , n41314 );
and ( n41316 , n41267 , n41315 );
xor ( n41317 , n41162 , n41230 );
xor ( n41318 , n41317 , n41233 );
and ( n41319 , n39432 , n41055 );
and ( n41320 , n39409 , n41053 );
nor ( n41321 , n41319 , n41320 );
xnor ( n41322 , n41321 , n40728 );
and ( n41323 , n39653 , n40258 );
and ( n41324 , n39620 , n40256 );
nor ( n41325 , n41323 , n41324 );
xnor ( n41326 , n41325 , n40169 );
and ( n41327 , n41322 , n41326 );
xor ( n41328 , n41200 , n41204 );
xor ( n41329 , n41328 , n41209 );
and ( n41330 , n41326 , n41329 );
and ( n41331 , n41322 , n41329 );
or ( n41332 , n41327 , n41330 , n41331 );
xor ( n41333 , n41166 , n41170 );
xor ( n41334 , n41333 , n41175 );
and ( n41335 , n41332 , n41334 );
xor ( n41336 , n41212 , n41216 );
xor ( n41337 , n41336 , n41221 );
and ( n41338 , n41334 , n41337 );
and ( n41339 , n41332 , n41337 );
or ( n41340 , n41335 , n41338 , n41339 );
xor ( n41341 , n41113 , n41115 );
xor ( n41342 , n41341 , n41118 );
and ( n41343 , n41340 , n41342 );
xor ( n41344 , n41178 , n41224 );
xor ( n41345 , n41344 , n41227 );
and ( n41346 , n41342 , n41345 );
and ( n41347 , n41340 , n41345 );
or ( n41348 , n41343 , n41346 , n41347 );
and ( n41349 , n41318 , n41348 );
and ( n41350 , n39552 , n40527 );
and ( n41351 , n39493 , n40525 );
nor ( n41352 , n41350 , n41351 );
xnor ( n41353 , n41352 , n40382 );
and ( n41354 , n39752 , n40053 );
and ( n41355 , n39670 , n40051 );
nor ( n41356 , n41354 , n41355 );
xnor ( n41357 , n41356 , n39999 );
and ( n41358 , n41353 , n41357 );
and ( n41359 , n39867 , n39896 );
and ( n41360 , n39795 , n39894 );
nor ( n41361 , n41359 , n41360 );
xnor ( n41362 , n41361 , n39857 );
and ( n41363 , n41357 , n41362 );
and ( n41364 , n41353 , n41362 );
or ( n41365 , n41358 , n41363 , n41364 );
xor ( n41366 , n41103 , n41107 );
xor ( n41367 , n41366 , n41110 );
and ( n41368 , n41365 , n41367 );
xor ( n41369 , n41142 , n41146 );
xor ( n41370 , n41369 , n41149 );
and ( n41371 , n41367 , n41370 );
and ( n41372 , n41365 , n41370 );
or ( n41373 , n41368 , n41371 , n41372 );
not ( n41374 , n41264 );
and ( n41375 , n39670 , n40258 );
and ( n41376 , n39653 , n40256 );
nor ( n41377 , n41375 , n41376 );
xnor ( n41378 , n41377 , n40169 );
and ( n41379 , n39948 , n39896 );
and ( n41380 , n39867 , n39894 );
nor ( n41381 , n41379 , n41380 );
xnor ( n41382 , n41381 , n39857 );
and ( n41383 , n41378 , n41382 );
and ( n41384 , n40186 , n39678 );
and ( n41385 , n40197 , n39676 );
nor ( n41386 , n41384 , n41385 );
xnor ( n41387 , n41386 , n39643 );
and ( n41388 , n41382 , n41387 );
and ( n41389 , n41378 , n41387 );
or ( n41390 , n41383 , n41388 , n41389 );
and ( n41391 , n39409 , n41292 );
and ( n41392 , n39365 , n41290 );
nor ( n41393 , n41391 , n41392 );
xnor ( n41394 , n41393 , n41041 );
and ( n41395 , n39493 , n40746 );
and ( n41396 , n39472 , n40744 );
nor ( n41397 , n41395 , n41396 );
xnor ( n41398 , n41397 , n40501 );
and ( n41399 , n41394 , n41398 );
and ( n41400 , n39795 , n40053 );
and ( n41401 , n39752 , n40051 );
nor ( n41402 , n41400 , n41401 );
xnor ( n41403 , n41402 , n39999 );
and ( n41404 , n41398 , n41403 );
and ( n41405 , n41394 , n41403 );
or ( n41406 , n41399 , n41404 , n41405 );
and ( n41407 , n41390 , n41406 );
xor ( n41408 , n41353 , n41357 );
xor ( n41409 , n41408 , n41362 );
and ( n41410 , n41406 , n41409 );
and ( n41411 , n41390 , n41409 );
or ( n41412 , n41407 , n41410 , n41411 );
and ( n41413 , n41374 , n41412 );
xor ( n41414 , n41301 , n41305 );
and ( n41415 , n41412 , n41414 );
and ( n41416 , n41374 , n41414 );
or ( n41417 , n41413 , n41415 , n41416 );
and ( n41418 , n41373 , n41417 );
and ( n41419 , n40507 , n39539 );
and ( n41420 , n40373 , n39537 );
nor ( n41421 , n41419 , n41420 );
xnor ( n41422 , n41421 , n39522 );
and ( n41423 , n40738 , n39480 );
and ( n41424 , n40492 , n39478 );
nor ( n41425 , n41423 , n41424 );
xnor ( n41426 , n41425 , n39462 );
and ( n41427 , n41422 , n41426 );
and ( n41428 , n41047 , n39396 );
and ( n41429 , n40869 , n39394 );
nor ( n41430 , n41428 , n41429 );
xnor ( n41431 , n41430 , n39401 );
and ( n41432 , n41426 , n41431 );
and ( n41433 , n41422 , n41431 );
or ( n41434 , n41427 , n41432 , n41433 );
and ( n41435 , n40148 , n39760 );
and ( n41436 , n40009 , n39758 );
nor ( n41437 , n41435 , n41436 );
xnor ( n41438 , n41437 , n39742 );
and ( n41439 , n41434 , n41438 );
xor ( n41440 , n41276 , n41280 );
xor ( n41441 , n41440 , n41285 );
and ( n41442 , n41438 , n41441 );
and ( n41443 , n41434 , n41441 );
or ( n41444 , n41439 , n41442 , n41443 );
and ( n41445 , n39472 , n40746 );
and ( n41446 , n39441 , n40744 );
nor ( n41447 , n41445 , n41446 );
xnor ( n41448 , n41447 , n40501 );
and ( n41449 , n41444 , n41448 );
xor ( n41450 , n41288 , n41295 );
xor ( n41451 , n41450 , n41298 );
and ( n41452 , n41448 , n41451 );
and ( n41453 , n41444 , n41451 );
or ( n41454 , n41449 , n41452 , n41453 );
and ( n41455 , n40009 , n39760 );
and ( n41456 , n39948 , n39758 );
nor ( n41457 , n41455 , n41456 );
xnor ( n41458 , n41457 , n39742 );
not ( n41459 , n41263 );
and ( n41460 , n41458 , n41459 );
xor ( n41461 , n41390 , n41406 );
xor ( n41462 , n41461 , n41409 );
and ( n41463 , n41459 , n41462 );
and ( n41464 , n41458 , n41462 );
or ( n41465 , n41460 , n41463 , n41464 );
and ( n41466 , n41454 , n41465 );
xor ( n41467 , n41365 , n41367 );
xor ( n41468 , n41467 , n41370 );
and ( n41469 , n41465 , n41468 );
and ( n41470 , n41454 , n41468 );
or ( n41471 , n41466 , n41469 , n41470 );
and ( n41472 , n41417 , n41471 );
and ( n41473 , n41373 , n41471 );
or ( n41474 , n41418 , n41472 , n41473 );
and ( n41475 , n41348 , n41474 );
and ( n41476 , n41318 , n41474 );
or ( n41477 , n41349 , n41475 , n41476 );
and ( n41478 , n41315 , n41477 );
and ( n41479 , n41267 , n41477 );
or ( n41480 , n41316 , n41478 , n41479 );
and ( n41481 , n41258 , n41480 );
and ( n41482 , n41253 , n41480 );
or ( n41483 , n41259 , n41481 , n41482 );
and ( n41484 , n41250 , n41483 );
and ( n41485 , n41099 , n41483 );
or ( n41486 , n41251 , n41484 , n41485 );
and ( n41487 , n41096 , n41486 );
and ( n41488 , n40948 , n41486 );
or ( n41489 , n41097 , n41487 , n41488 );
and ( n41490 , n40945 , n41489 );
and ( n41491 , n40843 , n41489 );
or ( n41492 , n40946 , n41490 , n41491 );
and ( n41493 , n40840 , n41492 );
and ( n41494 , n40705 , n41492 );
or ( n41495 , n40841 , n41493 , n41494 );
and ( n41496 , n40702 , n41495 );
and ( n41497 , n40488 , n41495 );
or ( n41498 , n40703 , n41496 , n41497 );
and ( n41499 , n40485 , n41498 );
and ( n41500 , n40445 , n41498 );
or ( n41501 , n40486 , n41499 , n41500 );
and ( n41502 , n40442 , n41501 );
and ( n41503 , n40329 , n41501 );
or ( n41504 , n40443 , n41502 , n41503 );
and ( n41505 , n40326 , n41504 );
and ( n41506 , n40230 , n41504 );
or ( n41507 , n40327 , n41505 , n41506 );
and ( n41508 , n40227 , n41507 );
and ( n41509 , n40092 , n41507 );
or ( n41510 , n40228 , n41508 , n41509 );
and ( n41511 , n40089 , n41510 );
and ( n41512 , n39992 , n41510 );
or ( n41513 , n40090 , n41511 , n41512 );
and ( n41514 , n39989 , n41513 );
and ( n41515 , n39987 , n41513 );
or ( n41516 , n39990 , n41514 , n41515 );
and ( n41517 , n39934 , n41516 );
and ( n41518 , n39850 , n41516 );
or ( n41519 , n39935 , n41517 , n41518 );
and ( n41520 , n39847 , n41519 );
and ( n41521 , n39735 , n41519 );
or ( n41522 , n39848 , n41520 , n41521 );
and ( n41523 , n39732 , n41522 );
and ( n41524 , n39714 , n41522 );
or ( n41525 , n39733 , n41523 , n41524 );
and ( n41526 , n39711 , n41525 );
and ( n41527 , n39607 , n41525 );
or ( n41528 , n39712 , n41526 , n41527 );
and ( n41529 , n39604 , n41528 );
and ( n41530 , n39575 , n41528 );
or ( n41531 , n39605 , n41529 , n41530 );
and ( n41532 , n39572 , n41531 );
and ( n41533 , n39515 , n41531 );
or ( n41534 , n39573 , n41532 , n41533 );
and ( n41535 , n39512 , n41534 );
and ( n41536 , n39455 , n41534 );
or ( n41537 , n39513 , n41535 , n41536 );
and ( n41538 , n39452 , n41537 );
and ( n41539 , n39427 , n41537 );
or ( n41540 , n39453 , n41538 , n41539 );
and ( n41541 , n39424 , n41540 );
and ( n41542 , n39422 , n41540 );
or ( n41543 , n39425 , n41541 , n41542 );
and ( n41544 , n39388 , n41543 );
xor ( n41545 , n39422 , n39424 );
xor ( n41546 , n41545 , n41540 );
xor ( n41547 , n39427 , n39452 );
xor ( n41548 , n41547 , n41537 );
xor ( n41549 , n39455 , n39512 );
xor ( n41550 , n41549 , n41534 );
xor ( n41551 , n39515 , n39572 );
xor ( n41552 , n41551 , n41531 );
xor ( n41553 , n39575 , n39604 );
xor ( n41554 , n41553 , n41528 );
xor ( n41555 , n39607 , n39711 );
xor ( n41556 , n41555 , n41525 );
xor ( n41557 , n39714 , n39732 );
xor ( n41558 , n41557 , n41522 );
xor ( n41559 , n39735 , n39847 );
xor ( n41560 , n41559 , n41519 );
xor ( n41561 , n39850 , n39934 );
xor ( n41562 , n41561 , n41516 );
xor ( n41563 , n39987 , n39989 );
xor ( n41564 , n41563 , n41513 );
xor ( n41565 , n39992 , n40089 );
xor ( n41566 , n41565 , n41510 );
xor ( n41567 , n40092 , n40227 );
xor ( n41568 , n41567 , n41507 );
xor ( n41569 , n40230 , n40326 );
xor ( n41570 , n41569 , n41504 );
xor ( n41571 , n40329 , n40442 );
xor ( n41572 , n41571 , n41501 );
xor ( n41573 , n40445 , n40485 );
xor ( n41574 , n41573 , n41498 );
xor ( n41575 , n40488 , n40702 );
xor ( n41576 , n41575 , n41495 );
xor ( n41577 , n40705 , n40840 );
xor ( n41578 , n41577 , n41492 );
xor ( n41579 , n40843 , n40945 );
xor ( n41580 , n41579 , n41489 );
xor ( n41581 , n40948 , n41096 );
xor ( n41582 , n41581 , n41486 );
xor ( n41583 , n41099 , n41250 );
xor ( n41584 , n41583 , n41483 );
xor ( n41585 , n41255 , n41257 );
xor ( n41586 , n41269 , n41270 );
xor ( n41587 , n41586 , n41312 );
and ( n41588 , n39441 , n41055 );
and ( n41589 , n39432 , n41053 );
nor ( n41590 , n41588 , n41589 );
xnor ( n41591 , n41590 , n40728 );
and ( n41592 , n39620 , n40527 );
and ( n41593 , n39552 , n40525 );
nor ( n41594 , n41592 , n41593 );
xnor ( n41595 , n41594 , n40382 );
and ( n41596 , n41591 , n41595 );
xor ( n41597 , n41394 , n41398 );
xor ( n41598 , n41597 , n41403 );
and ( n41599 , n41595 , n41598 );
and ( n41600 , n41591 , n41598 );
or ( n41601 , n41596 , n41599 , n41600 );
and ( n41602 , n39752 , n40258 );
and ( n41603 , n39670 , n40256 );
nor ( n41604 , n41602 , n41603 );
xnor ( n41605 , n41604 , n40169 );
and ( n41606 , n39867 , n40053 );
and ( n41607 , n39795 , n40051 );
nor ( n41608 , n41606 , n41607 );
xnor ( n41609 , n41608 , n39999 );
and ( n41610 , n41605 , n41609 );
not ( n41611 , n41186 );
xor ( n41612 , n36954 , n39322 );
buf ( n568914 , n41612 );
buf ( n568915 , n568914 );
buf ( n41615 , n568915 );
and ( n41616 , n41615 , n39367 );
and ( n41617 , n41611 , n41616 );
and ( n41618 , n41610 , n41617 );
xor ( n41619 , n41038 , n41189 );
xor ( n41620 , n41189 , n41191 );
not ( n41621 , n41620 );
and ( n41622 , n41619 , n41621 );
and ( n41623 , n39365 , n41622 );
not ( n41624 , n41623 );
xnor ( n41625 , n41624 , n41194 );
and ( n41626 , n39472 , n41055 );
and ( n41627 , n39441 , n41053 );
nor ( n41628 , n41626 , n41627 );
xnor ( n41629 , n41628 , n40728 );
and ( n41630 , n41625 , n41629 );
and ( n41631 , n40388 , n39678 );
and ( n41632 , n40186 , n39676 );
nor ( n41633 , n41631 , n41632 );
xnor ( n41634 , n41633 , n39643 );
and ( n41635 , n41629 , n41634 );
and ( n41636 , n41625 , n41634 );
or ( n41637 , n41630 , n41635 , n41636 );
and ( n41638 , n41617 , n41637 );
and ( n41639 , n41610 , n41637 );
or ( n41640 , n41618 , n41638 , n41639 );
and ( n41641 , n41601 , n41640 );
xor ( n41642 , n41444 , n41448 );
xor ( n41643 , n41642 , n41451 );
and ( n41644 , n41640 , n41643 );
and ( n41645 , n41601 , n41643 );
or ( n41646 , n41641 , n41644 , n41645 );
and ( n41647 , n40373 , n39539 );
and ( n41648 , n40388 , n39537 );
nor ( n41649 , n41647 , n41648 );
xnor ( n41650 , n41649 , n39522 );
xor ( n41651 , n41187 , n41195 );
xor ( n41652 , n41651 , n41197 );
and ( n41653 , n41650 , n41652 );
xor ( n41654 , n41434 , n41438 );
xor ( n41655 , n41654 , n41441 );
xor ( n41656 , n41422 , n41426 );
xor ( n41657 , n41656 , n41431 );
xor ( n41658 , n41605 , n41609 );
and ( n41659 , n41657 , n41658 );
xor ( n41660 , n41611 , n41616 );
and ( n41661 , n41658 , n41660 );
and ( n41662 , n41657 , n41660 );
or ( n41663 , n41659 , n41661 , n41662 );
and ( n41664 , n41655 , n41663 );
and ( n41665 , n39670 , n40527 );
and ( n41666 , n39653 , n40525 );
nor ( n41667 , n41665 , n41666 );
xnor ( n41668 , n41667 , n40382 );
and ( n41669 , n39948 , n40053 );
and ( n41670 , n39867 , n40051 );
nor ( n41671 , n41669 , n41670 );
xnor ( n41672 , n41671 , n39999 );
and ( n41673 , n41668 , n41672 );
and ( n41674 , n40186 , n39760 );
and ( n41675 , n40197 , n39758 );
nor ( n41676 , n41674 , n41675 );
xnor ( n41677 , n41676 , n39742 );
and ( n41678 , n41672 , n41677 );
and ( n41679 , n41668 , n41677 );
or ( n41680 , n41673 , n41678 , n41679 );
buf ( n568982 , n1183 );
buf ( n41682 , n568982 );
buf ( n568984 , n1184 );
buf ( n41684 , n568984 );
and ( n41685 , n41682 , n41684 );
not ( n41686 , n41685 );
and ( n41687 , n41191 , n41686 );
not ( n41688 , n41687 );
xor ( n41689 , n36956 , n39321 );
buf ( n568991 , n41689 );
buf ( n568992 , n568991 );
buf ( n41692 , n568992 );
and ( n41693 , n41692 , n39367 );
and ( n41694 , n41688 , n41693 );
and ( n41695 , n41680 , n41694 );
and ( n41696 , n39441 , n41292 );
and ( n41697 , n39432 , n41290 );
nor ( n41698 , n41696 , n41697 );
xnor ( n41699 , n41698 , n41041 );
and ( n41700 , n40148 , n39896 );
and ( n41701 , n40009 , n39894 );
nor ( n41702 , n41700 , n41701 );
xnor ( n41703 , n41702 , n39857 );
and ( n41704 , n41699 , n41703 );
and ( n41705 , n40492 , n39539 );
and ( n41706 , n40507 , n39537 );
nor ( n41707 , n41705 , n41706 );
xnor ( n41708 , n41707 , n39522 );
and ( n41709 , n41703 , n41708 );
and ( n41710 , n41699 , n41708 );
or ( n41711 , n41704 , n41709 , n41710 );
and ( n41712 , n41694 , n41711 );
and ( n41713 , n41680 , n41711 );
or ( n41714 , n41695 , n41712 , n41713 );
and ( n41715 , n41663 , n41714 );
and ( n41716 , n41655 , n41714 );
or ( n41717 , n41664 , n41715 , n41716 );
and ( n41718 , n41653 , n41717 );
xor ( n41719 , n41458 , n41459 );
xor ( n41720 , n41719 , n41462 );
and ( n41721 , n41717 , n41720 );
and ( n41722 , n41653 , n41720 );
or ( n41723 , n41718 , n41721 , n41722 );
and ( n41724 , n41646 , n41723 );
xor ( n41725 , n41374 , n41412 );
xor ( n41726 , n41725 , n41414 );
and ( n41727 , n41723 , n41726 );
and ( n41728 , n41646 , n41726 );
or ( n41729 , n41724 , n41727 , n41728 );
xor ( n41730 , n41272 , n41306 );
xor ( n41731 , n41730 , n41309 );
and ( n41732 , n41729 , n41731 );
xor ( n41733 , n41340 , n41342 );
xor ( n41734 , n41733 , n41345 );
and ( n41735 , n41731 , n41734 );
and ( n41736 , n41729 , n41734 );
or ( n41737 , n41732 , n41735 , n41736 );
and ( n41738 , n41587 , n41737 );
xor ( n41739 , n41318 , n41348 );
xor ( n41740 , n41739 , n41474 );
and ( n41741 , n41737 , n41740 );
and ( n41742 , n41587 , n41740 );
or ( n41743 , n41738 , n41741 , n41742 );
and ( n41744 , n41585 , n41743 );
xor ( n41745 , n41267 , n41315 );
xor ( n41746 , n41745 , n41477 );
and ( n41747 , n41743 , n41746 );
and ( n41748 , n41585 , n41746 );
or ( n41749 , n41744 , n41747 , n41748 );
xor ( n41750 , n41253 , n41258 );
xor ( n41751 , n41750 , n41480 );
and ( n41752 , n41749 , n41751 );
xor ( n41753 , n41585 , n41743 );
xor ( n41754 , n41753 , n41746 );
xor ( n41755 , n41332 , n41334 );
xor ( n41756 , n41755 , n41337 );
xor ( n41757 , n41322 , n41326 );
xor ( n41758 , n41757 , n41329 );
xor ( n41759 , n41591 , n41595 );
xor ( n41760 , n41759 , n41598 );
xor ( n41761 , n41610 , n41617 );
xor ( n41762 , n41761 , n41637 );
and ( n41763 , n41760 , n41762 );
xor ( n41764 , n41650 , n41652 );
and ( n41765 , n41762 , n41764 );
and ( n41766 , n41760 , n41764 );
or ( n41767 , n41763 , n41765 , n41766 );
and ( n41768 , n41758 , n41767 );
xor ( n41769 , n41601 , n41640 );
xor ( n41770 , n41769 , n41643 );
and ( n41771 , n41767 , n41770 );
and ( n41772 , n41758 , n41770 );
or ( n41773 , n41768 , n41771 , n41772 );
and ( n41774 , n41756 , n41773 );
xor ( n41775 , n41454 , n41465 );
xor ( n41776 , n41775 , n41468 );
and ( n41777 , n41773 , n41776 );
and ( n41778 , n41756 , n41776 );
or ( n41779 , n41774 , n41777 , n41778 );
xor ( n41780 , n41373 , n41417 );
xor ( n41781 , n41780 , n41471 );
and ( n41782 , n41779 , n41781 );
xor ( n41783 , n41646 , n41723 );
xor ( n41784 , n41783 , n41726 );
xor ( n41785 , n41653 , n41717 );
xor ( n41786 , n41785 , n41720 );
and ( n41787 , n39432 , n41292 );
and ( n41788 , n39409 , n41290 );
nor ( n41789 , n41787 , n41788 );
xnor ( n41790 , n41789 , n41041 );
and ( n41791 , n39552 , n40746 );
and ( n41792 , n39493 , n40744 );
nor ( n41793 , n41791 , n41792 );
xnor ( n41794 , n41793 , n40501 );
and ( n41795 , n41790 , n41794 );
and ( n41796 , n39653 , n40527 );
and ( n41797 , n39620 , n40525 );
nor ( n41798 , n41796 , n41797 );
xnor ( n41799 , n41798 , n40382 );
and ( n41800 , n41794 , n41799 );
and ( n41801 , n41790 , n41799 );
or ( n41802 , n41795 , n41800 , n41801 );
not ( n41803 , n41684 );
xor ( n41804 , n36958 , n39320 );
buf ( n569106 , n41804 );
buf ( n569107 , n569106 );
buf ( n41807 , n569107 );
and ( n41808 , n41807 , n39375 );
and ( n41809 , n41692 , n39373 );
nor ( n41810 , n41808 , n41809 );
xnor ( n41811 , n41810 , n39380 );
and ( n41812 , n41803 , n41811 );
xor ( n41813 , n36959 , n39319 );
buf ( n569115 , n41813 );
buf ( n569116 , n569115 );
buf ( n41816 , n569116 );
and ( n41817 , n41816 , n39367 );
and ( n41818 , n41811 , n41817 );
and ( n41819 , n41803 , n41817 );
or ( n41820 , n41812 , n41818 , n41819 );
and ( n41821 , n40738 , n39539 );
and ( n41822 , n40492 , n39537 );
nor ( n41823 , n41821 , n41822 );
xnor ( n41824 , n41823 , n39522 );
and ( n41825 , n41820 , n41824 );
and ( n41826 , n41047 , n39480 );
and ( n41827 , n40869 , n39478 );
nor ( n41828 , n41826 , n41827 );
xnor ( n41829 , n41828 , n39462 );
and ( n41830 , n41824 , n41829 );
and ( n41831 , n41820 , n41829 );
or ( n41832 , n41825 , n41830 , n41831 );
and ( n41833 , n40373 , n39678 );
and ( n41834 , n40388 , n39676 );
nor ( n41835 , n41833 , n41834 );
xnor ( n41836 , n41835 , n39643 );
and ( n41837 , n41832 , n41836 );
and ( n41838 , n41807 , n39367 );
buf ( n41839 , n41838 );
and ( n41840 , n40869 , n39480 );
and ( n41841 , n40738 , n39478 );
nor ( n41842 , n41840 , n41841 );
xnor ( n41843 , n41842 , n39462 );
xor ( n41844 , n41839 , n41843 );
and ( n41845 , n41032 , n39396 );
and ( n41846 , n41047 , n39394 );
nor ( n41847 , n41845 , n41846 );
xnor ( n41848 , n41847 , n39401 );
xor ( n41849 , n41844 , n41848 );
and ( n41850 , n41836 , n41849 );
and ( n41851 , n41832 , n41849 );
or ( n41852 , n41837 , n41850 , n41851 );
and ( n41853 , n40009 , n39896 );
and ( n41854 , n39948 , n39894 );
nor ( n41855 , n41853 , n41854 );
xnor ( n41856 , n41855 , n39857 );
and ( n41857 , n41852 , n41856 );
and ( n41858 , n40197 , n39760 );
and ( n41859 , n40148 , n39758 );
nor ( n41860 , n41858 , n41859 );
xnor ( n41861 , n41860 , n39742 );
and ( n41862 , n41856 , n41861 );
and ( n41863 , n41852 , n41861 );
or ( n41864 , n41857 , n41862 , n41863 );
and ( n41865 , n41802 , n41864 );
xor ( n41866 , n41378 , n41382 );
xor ( n41867 , n41866 , n41387 );
and ( n41868 , n41864 , n41867 );
and ( n41869 , n41802 , n41867 );
or ( n41870 , n41865 , n41868 , n41869 );
and ( n41871 , n41786 , n41870 );
xor ( n41872 , n41625 , n41629 );
xor ( n41873 , n41872 , n41634 );
and ( n41874 , n41839 , n41843 );
and ( n41875 , n41843 , n41848 );
and ( n41876 , n41839 , n41848 );
or ( n41877 , n41874 , n41875 , n41876 );
and ( n41878 , n41873 , n41877 );
and ( n41879 , n41615 , n39375 );
and ( n41880 , n41182 , n39373 );
nor ( n41881 , n41879 , n41880 );
xnor ( n41882 , n41881 , n39380 );
xor ( n41883 , n41688 , n41693 );
and ( n41884 , n41882 , n41883 );
and ( n41885 , n39752 , n40527 );
and ( n41886 , n39670 , n40525 );
nor ( n41887 , n41885 , n41886 );
xnor ( n41888 , n41887 , n40382 );
and ( n41889 , n40009 , n40053 );
and ( n41890 , n39948 , n40051 );
nor ( n41891 , n41889 , n41890 );
xnor ( n41892 , n41891 , n39999 );
and ( n41893 , n41888 , n41892 );
and ( n41894 , n41883 , n41893 );
and ( n41895 , n41882 , n41893 );
or ( n41896 , n41884 , n41894 , n41895 );
and ( n41897 , n41877 , n41896 );
and ( n41898 , n41873 , n41896 );
or ( n41899 , n41878 , n41897 , n41898 );
xor ( n41900 , n41655 , n41663 );
xor ( n41901 , n41900 , n41714 );
and ( n41902 , n41899 , n41901 );
xor ( n41903 , n41657 , n41658 );
xor ( n41904 , n41903 , n41660 );
xor ( n41905 , n41680 , n41694 );
xor ( n41906 , n41905 , n41711 );
and ( n41907 , n41904 , n41906 );
and ( n41908 , n41182 , n39396 );
and ( n41909 , n41032 , n39394 );
nor ( n41910 , n41908 , n41909 );
xnor ( n41911 , n41910 , n39401 );
buf ( n41912 , n41911 );
xor ( n41913 , n41699 , n41703 );
xor ( n41914 , n41913 , n41708 );
and ( n41915 , n41912 , n41914 );
and ( n41916 , n40507 , n39678 );
and ( n41917 , n40373 , n39676 );
nor ( n41918 , n41916 , n41917 );
xnor ( n41919 , n41918 , n39643 );
and ( n41920 , n41692 , n39375 );
and ( n41921 , n41615 , n39373 );
nor ( n41922 , n41920 , n41921 );
xnor ( n41923 , n41922 , n39380 );
and ( n41924 , n41919 , n41923 );
xor ( n41925 , n41888 , n41892 );
and ( n41926 , n41923 , n41925 );
and ( n41927 , n41919 , n41925 );
or ( n41928 , n41924 , n41926 , n41927 );
and ( n41929 , n41914 , n41928 );
and ( n41930 , n41912 , n41928 );
or ( n41931 , n41915 , n41929 , n41930 );
and ( n41932 , n41906 , n41931 );
and ( n41933 , n41904 , n41931 );
or ( n41934 , n41907 , n41932 , n41933 );
and ( n41935 , n41901 , n41934 );
and ( n41936 , n41899 , n41934 );
or ( n41937 , n41902 , n41935 , n41936 );
and ( n41938 , n41870 , n41937 );
and ( n41939 , n41786 , n41937 );
or ( n41940 , n41871 , n41938 , n41939 );
and ( n41941 , n41784 , n41940 );
xor ( n41942 , n41756 , n41773 );
xor ( n41943 , n41942 , n41776 );
and ( n41944 , n41940 , n41943 );
and ( n41945 , n41784 , n41943 );
or ( n41946 , n41941 , n41944 , n41945 );
and ( n41947 , n41781 , n41946 );
and ( n41948 , n41779 , n41946 );
or ( n41949 , n41782 , n41947 , n41948 );
xor ( n41950 , n41587 , n41737 );
xor ( n41951 , n41950 , n41740 );
and ( n41952 , n41949 , n41951 );
xor ( n41953 , n41729 , n41731 );
xor ( n41954 , n41953 , n41734 );
xor ( n41955 , n41779 , n41781 );
xor ( n41956 , n41955 , n41946 );
and ( n41957 , n41954 , n41956 );
xor ( n41958 , n41758 , n41767 );
xor ( n41959 , n41958 , n41770 );
xor ( n41960 , n41760 , n41762 );
xor ( n41961 , n41960 , n41764 );
xor ( n41962 , n41873 , n41877 );
xor ( n41963 , n41962 , n41896 );
xor ( n41964 , n41852 , n41856 );
xor ( n41965 , n41964 , n41861 );
and ( n41966 , n41963 , n41965 );
xor ( n41967 , n41882 , n41883 );
xor ( n41968 , n41967 , n41893 );
not ( n41969 , n41911 );
not ( n41970 , n41838 );
and ( n41971 , n41969 , n41970 );
and ( n41972 , n39948 , n40258 );
and ( n41973 , n39867 , n40256 );
nor ( n41974 , n41972 , n41973 );
xnor ( n41975 , n41974 , n40169 );
and ( n41976 , n40148 , n40053 );
and ( n41977 , n40009 , n40051 );
nor ( n41978 , n41976 , n41977 );
xnor ( n41979 , n41978 , n39999 );
and ( n41980 , n41975 , n41979 );
xor ( n41981 , n41191 , n41682 );
xor ( n41982 , n41682 , n41684 );
not ( n41983 , n41982 );
and ( n41984 , n41981 , n41983 );
and ( n41985 , n39409 , n41984 );
and ( n41986 , n39365 , n41982 );
nor ( n41987 , n41985 , n41986 );
xnor ( n41988 , n41987 , n41687 );
and ( n41989 , n39493 , n41292 );
and ( n41990 , n39472 , n41290 );
nor ( n41991 , n41989 , n41990 );
xnor ( n41992 , n41991 , n41041 );
xor ( n41993 , n41988 , n41992 );
and ( n41994 , n39795 , n40527 );
and ( n41995 , n39752 , n40525 );
nor ( n41996 , n41994 , n41995 );
xnor ( n41997 , n41996 , n40382 );
xor ( n41998 , n41993 , n41997 );
and ( n41999 , n41979 , n41998 );
and ( n42000 , n41975 , n41998 );
or ( n42001 , n41980 , n41999 , n42000 );
and ( n42002 , n41970 , n42001 );
and ( n42003 , n41969 , n42001 );
or ( n42004 , n41971 , n42002 , n42003 );
and ( n42005 , n41968 , n42004 );
xor ( n42006 , n41912 , n41914 );
xor ( n42007 , n42006 , n41928 );
and ( n42008 , n42004 , n42007 );
and ( n42009 , n41968 , n42007 );
or ( n42010 , n42005 , n42008 , n42009 );
and ( n42011 , n41965 , n42010 );
and ( n42012 , n41963 , n42010 );
or ( n42013 , n41966 , n42011 , n42012 );
and ( n42014 , n41961 , n42013 );
xor ( n42015 , n41899 , n41901 );
xor ( n42016 , n42015 , n41934 );
and ( n42017 , n42013 , n42016 );
and ( n42018 , n41961 , n42016 );
or ( n42019 , n42014 , n42017 , n42018 );
and ( n42020 , n41959 , n42019 );
xor ( n42021 , n41786 , n41870 );
xor ( n42022 , n42021 , n41937 );
and ( n42023 , n42019 , n42022 );
and ( n42024 , n41959 , n42022 );
or ( n42025 , n42020 , n42023 , n42024 );
xor ( n42026 , n41784 , n41940 );
xor ( n42027 , n42026 , n41943 );
and ( n42028 , n42025 , n42027 );
and ( n42029 , n39409 , n41622 );
and ( n42030 , n39365 , n41620 );
nor ( n42031 , n42029 , n42030 );
xnor ( n42032 , n42031 , n41194 );
and ( n42033 , n39493 , n41055 );
and ( n42034 , n39472 , n41053 );
nor ( n42035 , n42033 , n42034 );
xnor ( n42036 , n42035 , n40728 );
and ( n42037 , n42032 , n42036 );
and ( n42038 , n39795 , n40258 );
and ( n42039 , n39752 , n40256 );
nor ( n42040 , n42038 , n42039 );
xnor ( n42041 , n42040 , n40169 );
and ( n42042 , n42036 , n42041 );
and ( n42043 , n42032 , n42041 );
or ( n42044 , n42037 , n42042 , n42043 );
xor ( n42045 , n36964 , n39316 );
buf ( n569347 , n42045 );
buf ( n569348 , n569347 );
buf ( n42048 , n569348 );
and ( n42049 , n42048 , n39367 );
buf ( n42050 , n557768 );
not ( n42051 , n42050 );
and ( n42052 , n42049 , n42051 );
and ( n42053 , n41182 , n39480 );
and ( n42054 , n41032 , n39478 );
nor ( n42055 , n42053 , n42054 );
xnor ( n42056 , n42055 , n39462 );
and ( n42057 , n42052 , n42056 );
xor ( n42058 , n36961 , n39318 );
buf ( n569360 , n42058 );
buf ( n569361 , n569360 );
buf ( n42061 , n569361 );
and ( n42062 , n42061 , n39367 );
and ( n42063 , n42056 , n42062 );
and ( n42064 , n42052 , n42062 );
or ( n42065 , n42057 , n42063 , n42064 );
and ( n42066 , n40869 , n39539 );
and ( n42067 , n40738 , n39537 );
nor ( n42068 , n42066 , n42067 );
xnor ( n42069 , n42068 , n39522 );
and ( n42070 , n42065 , n42069 );
xor ( n42071 , n41803 , n41811 );
xor ( n42072 , n42071 , n41817 );
and ( n42073 , n42069 , n42072 );
and ( n42074 , n42065 , n42072 );
or ( n42075 , n42070 , n42073 , n42074 );
and ( n42076 , n40388 , n39760 );
and ( n42077 , n40186 , n39758 );
nor ( n42078 , n42076 , n42077 );
xnor ( n42079 , n42078 , n39742 );
and ( n42080 , n42075 , n42079 );
xor ( n42081 , n41820 , n41824 );
xor ( n42082 , n42081 , n41829 );
and ( n42083 , n42079 , n42082 );
and ( n42084 , n42075 , n42082 );
or ( n42085 , n42080 , n42083 , n42084 );
and ( n42086 , n39620 , n40746 );
and ( n42087 , n39552 , n40744 );
nor ( n42088 , n42086 , n42087 );
xnor ( n42089 , n42088 , n40501 );
and ( n42090 , n42085 , n42089 );
xor ( n42091 , n41832 , n41836 );
xor ( n42092 , n42091 , n41849 );
and ( n42093 , n42089 , n42092 );
and ( n42094 , n42085 , n42092 );
or ( n42095 , n42090 , n42093 , n42094 );
and ( n42096 , n42044 , n42095 );
xor ( n42097 , n41790 , n41794 );
xor ( n42098 , n42097 , n41799 );
and ( n42099 , n42095 , n42098 );
and ( n42100 , n42044 , n42098 );
or ( n42101 , n42096 , n42099 , n42100 );
xor ( n42102 , n41802 , n41864 );
xor ( n42103 , n42102 , n41867 );
and ( n42104 , n42101 , n42103 );
xor ( n42105 , n41959 , n42019 );
xor ( n42106 , n42105 , n42022 );
and ( n42107 , n42104 , n42106 );
xor ( n42108 , n41961 , n42013 );
xor ( n42109 , n42108 , n42016 );
xor ( n42110 , n42101 , n42103 );
and ( n42111 , n42109 , n42110 );
and ( n42112 , n40738 , n39678 );
and ( n42113 , n40492 , n39676 );
nor ( n42114 , n42112 , n42113 );
xnor ( n42115 , n42114 , n39643 );
and ( n42116 , n41047 , n39539 );
and ( n42117 , n40869 , n39537 );
nor ( n42118 , n42116 , n42117 );
xnor ( n42119 , n42118 , n39522 );
and ( n42120 , n42115 , n42119 );
xor ( n42121 , n42052 , n42056 );
xor ( n42122 , n42121 , n42062 );
and ( n42123 , n42119 , n42122 );
and ( n42124 , n42115 , n42122 );
or ( n42125 , n42120 , n42123 , n42124 );
and ( n42126 , n40373 , n39760 );
and ( n42127 , n40388 , n39758 );
nor ( n42128 , n42126 , n42127 );
xnor ( n42129 , n42128 , n39742 );
and ( n42130 , n42125 , n42129 );
xor ( n42131 , n42065 , n42069 );
xor ( n42132 , n42131 , n42072 );
and ( n42133 , n42129 , n42132 );
and ( n42134 , n42125 , n42132 );
or ( n42135 , n42130 , n42133 , n42134 );
and ( n42136 , n39472 , n41292 );
and ( n42137 , n39441 , n41290 );
nor ( n42138 , n42136 , n42137 );
xnor ( n42139 , n42138 , n41041 );
and ( n42140 , n42135 , n42139 );
and ( n42141 , n39552 , n41055 );
and ( n42142 , n39493 , n41053 );
nor ( n42143 , n42141 , n42142 );
xnor ( n42144 , n42143 , n40728 );
and ( n42145 , n42139 , n42144 );
and ( n42146 , n42135 , n42144 );
or ( n42147 , n42140 , n42145 , n42146 );
xor ( n42148 , n42032 , n42036 );
xor ( n42149 , n42148 , n42041 );
and ( n42150 , n42147 , n42149 );
xor ( n42151 , n42085 , n42089 );
xor ( n42152 , n42151 , n42092 );
and ( n42153 , n42149 , n42152 );
and ( n42154 , n42147 , n42152 );
or ( n42155 , n42150 , n42153 , n42154 );
xor ( n42156 , n42044 , n42095 );
xor ( n42157 , n42156 , n42098 );
and ( n42158 , n42155 , n42157 );
and ( n42159 , n42110 , n42158 );
and ( n42160 , n42109 , n42158 );
or ( n42161 , n42111 , n42159 , n42160 );
and ( n42162 , n42106 , n42161 );
and ( n42163 , n42104 , n42161 );
or ( n42164 , n42107 , n42162 , n42163 );
and ( n42165 , n42027 , n42164 );
and ( n42166 , n42025 , n42164 );
or ( n42167 , n42028 , n42165 , n42166 );
and ( n42168 , n41956 , n42167 );
and ( n42169 , n41954 , n42167 );
or ( n42170 , n41957 , n42168 , n42169 );
and ( n42171 , n41951 , n42170 );
and ( n42172 , n41949 , n42170 );
or ( n42173 , n41952 , n42171 , n42172 );
or ( n42174 , n41754 , n42173 );
and ( n42175 , n41751 , n42174 );
and ( n42176 , n41749 , n42174 );
or ( n42177 , n41752 , n42175 , n42176 );
or ( n42178 , n41584 , n42177 );
or ( n42179 , n41582 , n42178 );
or ( n42180 , n41580 , n42179 );
or ( n42181 , n41578 , n42180 );
or ( n42182 , n41576 , n42181 );
or ( n42183 , n41574 , n42182 );
or ( n42184 , n41572 , n42183 );
or ( n42185 , n41570 , n42184 );
or ( n42186 , n41568 , n42185 );
or ( n42187 , n41566 , n42186 );
or ( n42188 , n41564 , n42187 );
or ( n42189 , n41562 , n42188 );
or ( n42190 , n41560 , n42189 );
or ( n42191 , n41558 , n42190 );
or ( n42192 , n41556 , n42191 );
or ( n42193 , n41554 , n42192 );
or ( n42194 , n41552 , n42193 );
or ( n42195 , n41550 , n42194 );
or ( n42196 , n41548 , n42195 );
or ( n42197 , n41546 , n42196 );
and ( n42198 , n41543 , n42197 );
and ( n42199 , n39388 , n42197 );
or ( n42200 , n41544 , n42198 , n42199 );
not ( n42201 , n42200 );
xor ( n42202 , n39388 , n41543 );
xor ( n42203 , n42202 , n42197 );
xnor ( n42204 , n41546 , n42196 );
xnor ( n42205 , n41548 , n42195 );
xnor ( n42206 , n41550 , n42194 );
xnor ( n42207 , n41552 , n42193 );
xnor ( n42208 , n41554 , n42192 );
xnor ( n42209 , n41556 , n42191 );
xnor ( n42210 , n41558 , n42190 );
xnor ( n42211 , n41560 , n42189 );
xnor ( n42212 , n41562 , n42188 );
xnor ( n42213 , n41564 , n42187 );
xnor ( n42214 , n41566 , n42186 );
xnor ( n42215 , n41568 , n42185 );
xnor ( n42216 , n41570 , n42184 );
xnor ( n42217 , n41572 , n42183 );
xnor ( n42218 , n41574 , n42182 );
xnor ( n42219 , n41576 , n42181 );
xnor ( n42220 , n41578 , n42180 );
xnor ( n42221 , n41580 , n42179 );
xnor ( n42222 , n41582 , n42178 );
xnor ( n42223 , n41584 , n42177 );
xor ( n42224 , n41749 , n41751 );
xor ( n42225 , n42224 , n42174 );
not ( n42226 , n42225 );
xnor ( n42227 , n41754 , n42173 );
xor ( n42228 , n41949 , n41951 );
xor ( n42229 , n42228 , n42170 );
xor ( n42230 , n41954 , n41956 );
xor ( n42231 , n42230 , n42167 );
xor ( n42232 , n42025 , n42027 );
xor ( n42233 , n42232 , n42164 );
xor ( n42234 , n41904 , n41906 );
xor ( n42235 , n42234 , n41931 );
xor ( n42236 , n41963 , n41965 );
xor ( n42237 , n42236 , n42010 );
and ( n42238 , n42235 , n42237 );
and ( n42239 , n39432 , n41984 );
and ( n42240 , n39409 , n41982 );
nor ( n42241 , n42239 , n42240 );
xnor ( n42242 , n42241 , n41687 );
and ( n42243 , n39653 , n41055 );
and ( n42244 , n39620 , n41053 );
nor ( n42245 , n42243 , n42244 );
xnor ( n42246 , n42245 , n40728 );
and ( n42247 , n42242 , n42246 );
and ( n42248 , n39867 , n40527 );
and ( n42249 , n39795 , n40525 );
nor ( n42250 , n42248 , n42249 );
xnor ( n42251 , n42250 , n40382 );
and ( n42252 , n42246 , n42251 );
and ( n42253 , n42242 , n42251 );
or ( n42254 , n42247 , n42252 , n42253 );
and ( n42255 , n39752 , n40746 );
and ( n42256 , n39670 , n40744 );
nor ( n42257 , n42255 , n42256 );
xnor ( n42258 , n42257 , n40501 );
and ( n42259 , n40009 , n40258 );
and ( n42260 , n39948 , n40256 );
nor ( n42261 , n42259 , n42260 );
xnor ( n42262 , n42261 , n40169 );
and ( n42263 , n42258 , n42262 );
and ( n42264 , n42254 , n42263 );
buf ( n569566 , n1185 );
buf ( n42266 , n569566 );
xor ( n42267 , n41684 , n42266 );
not ( n42268 , n42266 );
and ( n42269 , n42267 , n42268 );
and ( n42270 , n39365 , n42269 );
not ( n42271 , n42270 );
xnor ( n42272 , n42271 , n41684 );
and ( n42273 , n39472 , n41622 );
and ( n42274 , n39441 , n41620 );
nor ( n42275 , n42273 , n42274 );
xnor ( n42276 , n42275 , n41194 );
and ( n42277 , n42272 , n42276 );
and ( n42278 , n39552 , n41292 );
and ( n42279 , n39493 , n41290 );
nor ( n42280 , n42278 , n42279 );
xnor ( n42281 , n42280 , n41041 );
and ( n42282 , n42276 , n42281 );
and ( n42283 , n42272 , n42281 );
or ( n42284 , n42277 , n42282 , n42283 );
and ( n42285 , n42263 , n42284 );
and ( n42286 , n42254 , n42284 );
or ( n42287 , n42264 , n42285 , n42286 );
xor ( n42288 , n41919 , n41923 );
xor ( n42289 , n42288 , n41925 );
and ( n42290 , n42287 , n42289 );
and ( n42291 , n39409 , n42269 );
and ( n42292 , n39365 , n42266 );
nor ( n42293 , n42291 , n42292 );
xnor ( n42294 , n42293 , n41684 );
and ( n42295 , n39493 , n41622 );
and ( n42296 , n39472 , n41620 );
nor ( n42297 , n42295 , n42296 );
xnor ( n42298 , n42297 , n41194 );
and ( n42299 , n42294 , n42298 );
and ( n42300 , n39620 , n41292 );
and ( n42301 , n39552 , n41290 );
nor ( n42302 , n42300 , n42301 );
xnor ( n42303 , n42302 , n41041 );
and ( n42304 , n42298 , n42303 );
and ( n42305 , n42294 , n42303 );
or ( n42306 , n42299 , n42304 , n42305 );
xor ( n42307 , n42242 , n42246 );
xor ( n42308 , n42307 , n42251 );
and ( n42309 , n42306 , n42308 );
and ( n42310 , n40197 , n40053 );
and ( n42311 , n40148 , n40051 );
nor ( n42312 , n42310 , n42311 );
xnor ( n42313 , n42312 , n39999 );
and ( n42314 , n40507 , n39760 );
and ( n42315 , n40373 , n39758 );
nor ( n42316 , n42314 , n42315 );
xnor ( n42317 , n42316 , n39742 );
and ( n42318 , n42313 , n42317 );
xor ( n42319 , n42258 , n42262 );
and ( n42320 , n42317 , n42319 );
and ( n42321 , n42313 , n42319 );
or ( n42322 , n42318 , n42320 , n42321 );
and ( n42323 , n42309 , n42322 );
and ( n42324 , n40492 , n39760 );
and ( n42325 , n40507 , n39758 );
nor ( n42326 , n42324 , n42325 );
xnor ( n42327 , n42326 , n39742 );
and ( n42328 , n40869 , n39678 );
and ( n42329 , n40738 , n39676 );
nor ( n42330 , n42328 , n42329 );
xnor ( n42331 , n42330 , n39643 );
and ( n42332 , n42327 , n42331 );
and ( n42333 , n39441 , n41984 );
and ( n42334 , n39432 , n41982 );
nor ( n42335 , n42333 , n42334 );
xnor ( n42336 , n42335 , n41687 );
and ( n42337 , n39795 , n40746 );
and ( n42338 , n39752 , n40744 );
nor ( n42339 , n42337 , n42338 );
xnor ( n42340 , n42339 , n40501 );
and ( n42341 , n42336 , n42340 );
and ( n42342 , n40148 , n40258 );
and ( n42343 , n40009 , n40256 );
nor ( n42344 , n42342 , n42343 );
xnor ( n42345 , n42344 , n40169 );
and ( n42346 , n42340 , n42345 );
and ( n42347 , n42336 , n42345 );
or ( n42348 , n42341 , n42346 , n42347 );
and ( n42349 , n42332 , n42348 );
xor ( n42350 , n42272 , n42276 );
xor ( n42351 , n42350 , n42281 );
and ( n42352 , n42348 , n42351 );
and ( n42353 , n42332 , n42351 );
or ( n42354 , n42349 , n42352 , n42353 );
and ( n42355 , n42322 , n42354 );
and ( n42356 , n42309 , n42354 );
or ( n42357 , n42323 , n42355 , n42356 );
and ( n42358 , n42289 , n42357 );
and ( n42359 , n42287 , n42357 );
or ( n42360 , n42290 , n42358 , n42359 );
xor ( n42361 , n41968 , n42004 );
xor ( n42362 , n42361 , n42007 );
and ( n42363 , n42360 , n42362 );
xor ( n42364 , n41969 , n41970 );
xor ( n42365 , n42364 , n42001 );
and ( n42366 , n41816 , n39375 );
and ( n42367 , n41807 , n39373 );
nor ( n42368 , n42366 , n42367 );
xnor ( n42369 , n42368 , n39380 );
buf ( n42370 , n42369 );
and ( n42371 , n41032 , n39480 );
and ( n42372 , n41047 , n39478 );
nor ( n42373 , n42371 , n42372 );
xnor ( n42374 , n42373 , n39462 );
and ( n42375 , n42370 , n42374 );
and ( n42376 , n41615 , n39396 );
and ( n42377 , n41182 , n39394 );
nor ( n42378 , n42376 , n42377 );
xnor ( n42379 , n42378 , n39401 );
and ( n42380 , n42374 , n42379 );
and ( n42381 , n42370 , n42379 );
or ( n42382 , n42375 , n42380 , n42381 );
and ( n42383 , n42365 , n42382 );
xor ( n42384 , n41975 , n41979 );
xor ( n42385 , n42384 , n41998 );
xor ( n42386 , n42254 , n42263 );
xor ( n42387 , n42386 , n42284 );
and ( n42388 , n42385 , n42387 );
xor ( n42389 , n42306 , n42308 );
and ( n42390 , n41615 , n39480 );
and ( n42391 , n41182 , n39478 );
nor ( n42392 , n42390 , n42391 );
xnor ( n42393 , n42392 , n39462 );
xor ( n42394 , n42049 , n42051 );
and ( n42395 , n42393 , n42394 );
and ( n42396 , n42389 , n42395 );
and ( n42397 , n40373 , n39896 );
and ( n42398 , n40388 , n39894 );
nor ( n42399 , n42397 , n42398 );
xnor ( n42400 , n42399 , n39857 );
and ( n42401 , n39670 , n41055 );
and ( n42402 , n39653 , n41053 );
nor ( n42403 , n42401 , n42402 );
xnor ( n42404 , n42403 , n40728 );
and ( n42405 , n39948 , n40527 );
and ( n42406 , n39867 , n40525 );
nor ( n42407 , n42405 , n42406 );
xnor ( n42408 , n42407 , n40382 );
xor ( n42409 , n42404 , n42408 );
and ( n42410 , n40186 , n40053 );
and ( n42411 , n40197 , n40051 );
nor ( n42412 , n42410 , n42411 );
xnor ( n42413 , n42412 , n39999 );
xor ( n42414 , n42409 , n42413 );
and ( n42415 , n42400 , n42414 );
xor ( n42416 , n42294 , n42298 );
xor ( n42417 , n42416 , n42303 );
and ( n42418 , n42414 , n42417 );
and ( n42419 , n42400 , n42417 );
or ( n42420 , n42415 , n42418 , n42419 );
and ( n42421 , n42395 , n42420 );
and ( n42422 , n42389 , n42420 );
or ( n42423 , n42396 , n42421 , n42422 );
and ( n42424 , n42387 , n42423 );
and ( n42425 , n42385 , n42423 );
or ( n42426 , n42388 , n42424 , n42425 );
and ( n42427 , n42382 , n42426 );
and ( n42428 , n42365 , n42426 );
or ( n42429 , n42383 , n42427 , n42428 );
and ( n42430 , n42362 , n42429 );
and ( n42431 , n42360 , n42429 );
or ( n42432 , n42363 , n42430 , n42431 );
and ( n42433 , n42237 , n42432 );
and ( n42434 , n42235 , n42432 );
or ( n42435 , n42238 , n42433 , n42434 );
xor ( n42436 , n42155 , n42157 );
and ( n42437 , n39432 , n41622 );
and ( n42438 , n39409 , n41620 );
nor ( n42439 , n42437 , n42438 );
xnor ( n42440 , n42439 , n41194 );
and ( n42441 , n39653 , n40746 );
and ( n42442 , n39620 , n40744 );
nor ( n42443 , n42441 , n42442 );
xnor ( n42444 , n42443 , n40501 );
and ( n42445 , n42440 , n42444 );
and ( n42446 , n39867 , n40258 );
and ( n42447 , n39795 , n40256 );
nor ( n42448 , n42446 , n42447 );
xnor ( n42449 , n42448 , n40169 );
and ( n42450 , n42444 , n42449 );
and ( n42451 , n42440 , n42449 );
or ( n42452 , n42445 , n42450 , n42451 );
xor ( n42453 , n38144 , n39314 );
buf ( n569755 , n42453 );
buf ( n569756 , n569755 );
buf ( n42456 , n569756 );
and ( n42457 , n42456 , n39367 );
buf ( n42458 , n557769 );
not ( n42459 , n42458 );
and ( n42460 , n42457 , n42459 );
and ( n42461 , n41807 , n39396 );
and ( n42462 , n41692 , n39394 );
nor ( n42463 , n42461 , n42462 );
xnor ( n42464 , n42463 , n39401 );
and ( n42465 , n42460 , n42464 );
and ( n42466 , n42061 , n39375 );
and ( n42467 , n41816 , n39373 );
nor ( n42468 , n42466 , n42467 );
xnor ( n42469 , n42468 , n39380 );
and ( n42470 , n42464 , n42469 );
and ( n42471 , n42460 , n42469 );
or ( n42472 , n42465 , n42470 , n42471 );
and ( n42473 , n41692 , n39396 );
and ( n42474 , n41615 , n39394 );
nor ( n42475 , n42473 , n42474 );
xnor ( n42476 , n42475 , n39401 );
and ( n42477 , n42472 , n42476 );
not ( n42478 , n42369 );
and ( n42479 , n42476 , n42478 );
and ( n42480 , n42472 , n42478 );
or ( n42481 , n42477 , n42479 , n42480 );
and ( n42482 , n40492 , n39678 );
and ( n42483 , n40507 , n39676 );
nor ( n42484 , n42482 , n42483 );
xnor ( n42485 , n42484 , n39643 );
and ( n42486 , n42481 , n42485 );
xor ( n42487 , n42370 , n42374 );
xor ( n42488 , n42487 , n42379 );
and ( n42489 , n42485 , n42488 );
and ( n42490 , n42481 , n42488 );
or ( n42491 , n42486 , n42489 , n42490 );
and ( n42492 , n39365 , n41984 );
not ( n42493 , n42492 );
xnor ( n42494 , n42493 , n41687 );
and ( n42495 , n42491 , n42494 );
and ( n42496 , n40197 , n39896 );
and ( n42497 , n40148 , n39894 );
nor ( n42498 , n42496 , n42497 );
xnor ( n42499 , n42498 , n39857 );
and ( n42500 , n42494 , n42499 );
and ( n42501 , n42491 , n42499 );
or ( n42502 , n42495 , n42500 , n42501 );
and ( n42503 , n42452 , n42502 );
xor ( n42504 , n41668 , n41672 );
xor ( n42505 , n42504 , n41677 );
and ( n42506 , n42502 , n42505 );
and ( n42507 , n42452 , n42505 );
or ( n42508 , n42503 , n42506 , n42507 );
and ( n42509 , n42436 , n42508 );
xor ( n42510 , n42235 , n42237 );
xor ( n42511 , n42510 , n42432 );
and ( n42512 , n42508 , n42511 );
and ( n42513 , n42436 , n42511 );
or ( n42514 , n42509 , n42512 , n42513 );
and ( n42515 , n42435 , n42514 );
xor ( n42516 , n42109 , n42110 );
xor ( n42517 , n42516 , n42158 );
and ( n42518 , n42514 , n42517 );
and ( n42519 , n42435 , n42517 );
or ( n42520 , n42515 , n42518 , n42519 );
xor ( n42521 , n42104 , n42106 );
xor ( n42522 , n42521 , n42161 );
and ( n42523 , n42520 , n42522 );
and ( n42524 , n41988 , n41992 );
and ( n42525 , n41992 , n41997 );
and ( n42526 , n41988 , n41997 );
or ( n42527 , n42524 , n42525 , n42526 );
xor ( n42528 , n42440 , n42444 );
xor ( n42529 , n42528 , n42449 );
and ( n42530 , n42527 , n42529 );
xor ( n42531 , n42135 , n42139 );
xor ( n42532 , n42531 , n42144 );
and ( n42533 , n42529 , n42532 );
and ( n42534 , n42527 , n42532 );
or ( n42535 , n42530 , n42533 , n42534 );
xor ( n42536 , n42452 , n42502 );
xor ( n42537 , n42536 , n42505 );
and ( n42538 , n42535 , n42537 );
xor ( n42539 , n42147 , n42149 );
xor ( n42540 , n42539 , n42152 );
and ( n42541 , n42537 , n42540 );
and ( n42542 , n42535 , n42540 );
or ( n42543 , n42538 , n42541 , n42542 );
xor ( n42544 , n42287 , n42289 );
xor ( n42545 , n42544 , n42357 );
xor ( n42546 , n42457 , n42459 );
and ( n42547 , n41182 , n39539 );
and ( n42548 , n41032 , n39537 );
nor ( n42549 , n42547 , n42548 );
xnor ( n42550 , n42549 , n39522 );
and ( n42551 , n42546 , n42550 );
and ( n42552 , n41692 , n39480 );
and ( n42553 , n41615 , n39478 );
nor ( n42554 , n42552 , n42553 );
xnor ( n42555 , n42554 , n39462 );
and ( n42556 , n42550 , n42555 );
and ( n42557 , n42546 , n42555 );
or ( n42558 , n42551 , n42556 , n42557 );
and ( n42559 , n41032 , n39539 );
and ( n42560 , n41047 , n39537 );
nor ( n42561 , n42559 , n42560 );
xnor ( n42562 , n42561 , n39522 );
and ( n42563 , n42558 , n42562 );
xor ( n42564 , n42460 , n42464 );
xor ( n42565 , n42564 , n42469 );
and ( n42566 , n42562 , n42565 );
and ( n42567 , n42558 , n42565 );
or ( n42568 , n42563 , n42566 , n42567 );
and ( n42569 , n40388 , n39896 );
and ( n42570 , n40186 , n39894 );
nor ( n42571 , n42569 , n42570 );
xnor ( n42572 , n42571 , n39857 );
and ( n42573 , n42568 , n42572 );
xor ( n42574 , n42115 , n42119 );
xor ( n42575 , n42574 , n42122 );
and ( n42576 , n42572 , n42575 );
and ( n42577 , n42568 , n42575 );
or ( n42578 , n42573 , n42576 , n42577 );
and ( n42579 , n39441 , n41622 );
and ( n42580 , n39432 , n41620 );
nor ( n42581 , n42579 , n42580 );
xnor ( n42582 , n42581 , n41194 );
and ( n42583 , n42578 , n42582 );
and ( n42584 , n39620 , n41055 );
and ( n42585 , n39552 , n41053 );
nor ( n42586 , n42584 , n42585 );
xnor ( n42587 , n42586 , n40728 );
and ( n42588 , n42582 , n42587 );
and ( n42589 , n42578 , n42587 );
or ( n42590 , n42583 , n42588 , n42589 );
and ( n42591 , n42545 , n42590 );
xor ( n42592 , n42327 , n42331 );
and ( n42593 , n39752 , n41055 );
and ( n42594 , n39670 , n41053 );
nor ( n42595 , n42593 , n42594 );
xnor ( n42596 , n42595 , n40728 );
and ( n42597 , n40009 , n40527 );
and ( n42598 , n39948 , n40525 );
nor ( n42599 , n42597 , n42598 );
xnor ( n42600 , n42599 , n40382 );
and ( n42601 , n42596 , n42600 );
and ( n42602 , n40197 , n40258 );
and ( n42603 , n40148 , n40256 );
nor ( n42604 , n42602 , n42603 );
xnor ( n42605 , n42604 , n40169 );
and ( n42606 , n42600 , n42605 );
and ( n42607 , n42596 , n42605 );
or ( n42608 , n42601 , n42606 , n42607 );
and ( n42609 , n42592 , n42608 );
and ( n42610 , n39472 , n41984 );
and ( n42611 , n39441 , n41982 );
nor ( n42612 , n42610 , n42611 );
xnor ( n42613 , n42612 , n41687 );
and ( n42614 , n39552 , n41622 );
and ( n42615 , n39493 , n41620 );
nor ( n42616 , n42614 , n42615 );
xnor ( n42617 , n42616 , n41194 );
and ( n42618 , n42613 , n42617 );
and ( n42619 , n42608 , n42618 );
and ( n42620 , n42592 , n42618 );
or ( n42621 , n42609 , n42619 , n42620 );
and ( n42622 , n39432 , n42269 );
and ( n42623 , n39409 , n42266 );
nor ( n42624 , n42622 , n42623 );
xnor ( n42625 , n42624 , n41684 );
and ( n42626 , n39653 , n41292 );
and ( n42627 , n39620 , n41290 );
nor ( n42628 , n42626 , n42627 );
xnor ( n42629 , n42628 , n41041 );
and ( n42630 , n42625 , n42629 );
and ( n42631 , n39867 , n40746 );
and ( n42632 , n39795 , n40744 );
nor ( n42633 , n42631 , n42632 );
xnor ( n42634 , n42633 , n40501 );
and ( n42635 , n42629 , n42634 );
and ( n42636 , n42625 , n42634 );
or ( n42637 , n42630 , n42635 , n42636 );
and ( n42638 , n40388 , n40053 );
and ( n42639 , n40186 , n40051 );
nor ( n42640 , n42638 , n42639 );
xnor ( n42641 , n42640 , n39999 );
and ( n42642 , n40507 , n39896 );
and ( n42643 , n40373 , n39894 );
nor ( n42644 , n42642 , n42643 );
xnor ( n42645 , n42644 , n39857 );
and ( n42646 , n42641 , n42645 );
and ( n42647 , n41816 , n39396 );
and ( n42648 , n41807 , n39394 );
nor ( n42649 , n42647 , n42648 );
xnor ( n42650 , n42649 , n39401 );
and ( n42651 , n42645 , n42650 );
and ( n42652 , n42641 , n42650 );
or ( n42653 , n42646 , n42651 , n42652 );
and ( n42654 , n42637 , n42653 );
xor ( n42655 , n42336 , n42340 );
xor ( n42656 , n42655 , n42345 );
and ( n42657 , n42653 , n42656 );
and ( n42658 , n42637 , n42656 );
or ( n42659 , n42654 , n42657 , n42658 );
and ( n42660 , n42621 , n42659 );
xor ( n42661 , n42313 , n42317 );
xor ( n42662 , n42661 , n42319 );
and ( n42663 , n42659 , n42662 );
and ( n42664 , n42621 , n42662 );
or ( n42665 , n42660 , n42663 , n42664 );
xor ( n42666 , n42309 , n42322 );
xor ( n42667 , n42666 , n42354 );
and ( n42668 , n42665 , n42667 );
xor ( n42669 , n42125 , n42129 );
xor ( n42670 , n42669 , n42132 );
and ( n42671 , n42667 , n42670 );
and ( n42672 , n42665 , n42670 );
or ( n42673 , n42668 , n42671 , n42672 );
and ( n42674 , n42590 , n42673 );
and ( n42675 , n42545 , n42673 );
or ( n42676 , n42591 , n42674 , n42675 );
xor ( n42677 , n42360 , n42362 );
xor ( n42678 , n42677 , n42429 );
and ( n42679 , n42676 , n42678 );
and ( n42680 , n39670 , n40746 );
and ( n42681 , n39653 , n40744 );
nor ( n42682 , n42680 , n42681 );
xnor ( n42683 , n42682 , n40501 );
and ( n42684 , n40186 , n39896 );
and ( n42685 , n40197 , n39894 );
nor ( n42686 , n42684 , n42685 );
xnor ( n42687 , n42686 , n39857 );
and ( n42688 , n42683 , n42687 );
xor ( n42689 , n42481 , n42485 );
xor ( n42690 , n42689 , n42488 );
and ( n42691 , n42687 , n42690 );
and ( n42692 , n42683 , n42690 );
or ( n42693 , n42688 , n42691 , n42692 );
xor ( n42694 , n42075 , n42079 );
xor ( n42695 , n42694 , n42082 );
and ( n42696 , n42693 , n42695 );
and ( n42697 , n42678 , n42696 );
and ( n42698 , n42676 , n42696 );
or ( n42699 , n42679 , n42697 , n42698 );
and ( n42700 , n42543 , n42699 );
xor ( n42701 , n42436 , n42508 );
xor ( n42702 , n42701 , n42511 );
and ( n42703 , n42699 , n42702 );
and ( n42704 , n42543 , n42702 );
or ( n42705 , n42700 , n42703 , n42704 );
xor ( n42706 , n42435 , n42514 );
xor ( n42707 , n42706 , n42517 );
and ( n42708 , n42705 , n42707 );
xor ( n42709 , n42332 , n42348 );
xor ( n42710 , n42709 , n42351 );
xor ( n42711 , n42472 , n42476 );
xor ( n42712 , n42711 , n42478 );
and ( n42713 , n42710 , n42712 );
xor ( n42714 , n42393 , n42394 );
and ( n42715 , n42048 , n39375 );
and ( n42716 , n42061 , n39373 );
nor ( n42717 , n42715 , n42716 );
xnor ( n42718 , n42717 , n39380 );
xor ( n42719 , n42596 , n42600 );
xor ( n42720 , n42719 , n42605 );
and ( n42721 , n42718 , n42720 );
xor ( n42722 , n42613 , n42617 );
and ( n42723 , n42720 , n42722 );
and ( n42724 , n42718 , n42722 );
or ( n42725 , n42721 , n42723 , n42724 );
and ( n42726 , n42714 , n42725 );
and ( n42727 , n41807 , n39480 );
and ( n42728 , n41692 , n39478 );
nor ( n42729 , n42727 , n42728 );
xnor ( n42730 , n42729 , n39462 );
and ( n42731 , n42061 , n39396 );
and ( n42732 , n41816 , n39394 );
nor ( n42733 , n42731 , n42732 );
xnor ( n42734 , n42733 , n39401 );
and ( n42735 , n42730 , n42734 );
and ( n42736 , n39670 , n41292 );
and ( n42737 , n39653 , n41290 );
nor ( n42738 , n42736 , n42737 );
xnor ( n42739 , n42738 , n41041 );
and ( n42740 , n39795 , n41055 );
and ( n42741 , n39752 , n41053 );
nor ( n42742 , n42740 , n42741 );
xnor ( n42743 , n42742 , n40728 );
and ( n42744 , n42739 , n42743 );
and ( n42745 , n42735 , n42744 );
and ( n42746 , n39441 , n42269 );
and ( n42747 , n39432 , n42266 );
nor ( n42748 , n42746 , n42747 );
xnor ( n42749 , n42748 , n41684 );
and ( n42750 , n39948 , n40746 );
and ( n42751 , n39867 , n40744 );
nor ( n42752 , n42750 , n42751 );
xnor ( n42753 , n42752 , n40501 );
and ( n42754 , n42749 , n42753 );
and ( n42755 , n40148 , n40527 );
and ( n42756 , n40009 , n40525 );
nor ( n42757 , n42755 , n42756 );
xnor ( n42758 , n42757 , n40382 );
and ( n42759 , n42753 , n42758 );
and ( n42760 , n42749 , n42758 );
or ( n42761 , n42754 , n42759 , n42760 );
and ( n42762 , n42744 , n42761 );
and ( n42763 , n42735 , n42761 );
or ( n42764 , n42745 , n42762 , n42763 );
and ( n42765 , n42725 , n42764 );
and ( n42766 , n42714 , n42764 );
or ( n42767 , n42726 , n42765 , n42766 );
and ( n42768 , n42712 , n42767 );
and ( n42769 , n42710 , n42767 );
or ( n42770 , n42713 , n42768 , n42769 );
and ( n42771 , n40186 , n40258 );
and ( n42772 , n40197 , n40256 );
nor ( n42773 , n42771 , n42772 );
xnor ( n42774 , n42773 , n40169 );
and ( n42775 , n40373 , n40053 );
and ( n42776 , n40388 , n40051 );
nor ( n42777 , n42775 , n42776 );
xnor ( n42778 , n42777 , n39999 );
and ( n42779 , n42774 , n42778 );
and ( n42780 , n40492 , n39896 );
and ( n42781 , n40507 , n39894 );
nor ( n42782 , n42780 , n42781 );
xnor ( n42783 , n42782 , n39857 );
and ( n42784 , n42778 , n42783 );
and ( n42785 , n42774 , n42783 );
or ( n42786 , n42779 , n42784 , n42785 );
and ( n42787 , n40869 , n39760 );
and ( n42788 , n40738 , n39758 );
nor ( n42789 , n42787 , n42788 );
xnor ( n42790 , n42789 , n39742 );
and ( n42791 , n41032 , n39678 );
and ( n42792 , n41047 , n39676 );
nor ( n42793 , n42791 , n42792 );
xnor ( n42794 , n42793 , n39643 );
and ( n42795 , n42790 , n42794 );
and ( n42796 , n41615 , n39539 );
and ( n42797 , n41182 , n39537 );
nor ( n42798 , n42796 , n42797 );
xnor ( n42799 , n42798 , n39522 );
and ( n42800 , n42794 , n42799 );
and ( n42801 , n42790 , n42799 );
or ( n42802 , n42795 , n42800 , n42801 );
and ( n42803 , n42786 , n42802 );
and ( n42804 , n42456 , n39375 );
and ( n42805 , n42048 , n39373 );
nor ( n42806 , n42804 , n42805 );
xnor ( n42807 , n42806 , n39380 );
xor ( n42808 , n38146 , n39313 );
buf ( n570110 , n42808 );
buf ( n570111 , n570110 );
buf ( n42811 , n570111 );
and ( n42812 , n42811 , n39367 );
and ( n42813 , n42807 , n42812 );
buf ( n42814 , n557770 );
not ( n42815 , n42814 );
and ( n42816 , n42812 , n42815 );
and ( n42817 , n42807 , n42815 );
or ( n42818 , n42813 , n42816 , n42817 );
and ( n42819 , n42802 , n42818 );
and ( n42820 , n42786 , n42818 );
or ( n42821 , n42803 , n42819 , n42820 );
xor ( n42822 , n42400 , n42414 );
xor ( n42823 , n42822 , n42417 );
and ( n42824 , n42821 , n42823 );
xor ( n42825 , n42592 , n42608 );
xor ( n42826 , n42825 , n42618 );
and ( n42827 , n42823 , n42826 );
and ( n42828 , n42821 , n42826 );
or ( n42829 , n42824 , n42827 , n42828 );
xor ( n42830 , n42389 , n42395 );
xor ( n42831 , n42830 , n42420 );
and ( n42832 , n42829 , n42831 );
xor ( n42833 , n42621 , n42659 );
xor ( n42834 , n42833 , n42662 );
and ( n42835 , n42831 , n42834 );
and ( n42836 , n42829 , n42834 );
or ( n42837 , n42832 , n42835 , n42836 );
and ( n42838 , n42770 , n42837 );
xor ( n42839 , n42385 , n42387 );
xor ( n42840 , n42839 , n42423 );
and ( n42841 , n42837 , n42840 );
and ( n42842 , n42770 , n42840 );
or ( n42843 , n42838 , n42841 , n42842 );
xor ( n42844 , n42365 , n42382 );
xor ( n42845 , n42844 , n42426 );
and ( n42846 , n42843 , n42845 );
xor ( n42847 , n42491 , n42494 );
xor ( n42848 , n42847 , n42499 );
and ( n42849 , n42845 , n42848 );
and ( n42850 , n42843 , n42848 );
or ( n42851 , n42846 , n42849 , n42850 );
xor ( n42852 , n42527 , n42529 );
xor ( n42853 , n42852 , n42532 );
xor ( n42854 , n42578 , n42582 );
xor ( n42855 , n42854 , n42587 );
and ( n42856 , n42404 , n42408 );
and ( n42857 , n42408 , n42413 );
and ( n42858 , n42404 , n42413 );
or ( n42859 , n42856 , n42857 , n42858 );
xor ( n42860 , n42568 , n42572 );
xor ( n42861 , n42860 , n42575 );
and ( n42862 , n42859 , n42861 );
and ( n42863 , n42855 , n42862 );
xor ( n42864 , n42637 , n42653 );
xor ( n42865 , n42864 , n42656 );
xor ( n42866 , n42558 , n42562 );
xor ( n42867 , n42866 , n42565 );
and ( n42868 , n42865 , n42867 );
and ( n42869 , n40738 , n39760 );
and ( n42870 , n40492 , n39758 );
nor ( n42871 , n42869 , n42870 );
xnor ( n42872 , n42871 , n39742 );
and ( n42873 , n41047 , n39678 );
and ( n42874 , n40869 , n39676 );
nor ( n42875 , n42873 , n42874 );
xnor ( n42876 , n42875 , n39643 );
and ( n42877 , n42872 , n42876 );
xor ( n42878 , n42546 , n42550 );
xor ( n42879 , n42878 , n42555 );
and ( n42880 , n42876 , n42879 );
and ( n42881 , n42872 , n42879 );
or ( n42882 , n42877 , n42880 , n42881 );
and ( n42883 , n42867 , n42882 );
and ( n42884 , n42865 , n42882 );
or ( n42885 , n42868 , n42883 , n42884 );
xor ( n42886 , n42625 , n42629 );
xor ( n42887 , n42886 , n42634 );
xor ( n42888 , n42641 , n42645 );
xor ( n42889 , n42888 , n42650 );
and ( n42890 , n42887 , n42889 );
xor ( n42891 , n42730 , n42734 );
xor ( n42892 , n42739 , n42743 );
and ( n42893 , n42891 , n42892 );
and ( n42894 , n39472 , n42269 );
and ( n42895 , n39441 , n42266 );
nor ( n42896 , n42894 , n42895 );
xnor ( n42897 , n42896 , n41684 );
and ( n42898 , n39867 , n41055 );
and ( n42899 , n39795 , n41053 );
nor ( n42900 , n42898 , n42899 );
xnor ( n42901 , n42900 , n40728 );
and ( n42902 , n42897 , n42901 );
and ( n42903 , n40009 , n40746 );
and ( n42904 , n39948 , n40744 );
nor ( n42905 , n42903 , n42904 );
xnor ( n42906 , n42905 , n40501 );
and ( n42907 , n42901 , n42906 );
and ( n42908 , n42897 , n42906 );
or ( n42909 , n42902 , n42907 , n42908 );
and ( n42910 , n42892 , n42909 );
and ( n42911 , n42891 , n42909 );
or ( n42912 , n42893 , n42910 , n42911 );
and ( n42913 , n42889 , n42912 );
and ( n42914 , n42887 , n42912 );
or ( n42915 , n42890 , n42913 , n42914 );
and ( n42916 , n41182 , n39678 );
and ( n42917 , n41032 , n39676 );
nor ( n42918 , n42916 , n42917 );
xnor ( n42919 , n42918 , n39643 );
and ( n42920 , n41692 , n39539 );
and ( n42921 , n41615 , n39537 );
nor ( n42922 , n42920 , n42921 );
xnor ( n42923 , n42922 , n39522 );
and ( n42924 , n42919 , n42923 );
and ( n42925 , n42811 , n39375 );
and ( n42926 , n42456 , n39373 );
nor ( n42927 , n42925 , n42926 );
xnor ( n42928 , n42927 , n39380 );
and ( n42929 , n42923 , n42928 );
and ( n42930 , n42919 , n42928 );
or ( n42931 , n42924 , n42929 , n42930 );
xor ( n42932 , n42749 , n42753 );
xor ( n42933 , n42932 , n42758 );
and ( n42934 , n42931 , n42933 );
xor ( n42935 , n42774 , n42778 );
xor ( n42936 , n42935 , n42783 );
and ( n42937 , n42933 , n42936 );
and ( n42938 , n42931 , n42936 );
or ( n42939 , n42934 , n42937 , n42938 );
xor ( n42940 , n42718 , n42720 );
xor ( n42941 , n42940 , n42722 );
and ( n42942 , n42939 , n42941 );
xor ( n42943 , n42735 , n42744 );
xor ( n42944 , n42943 , n42761 );
and ( n42945 , n42941 , n42944 );
and ( n42946 , n42939 , n42944 );
or ( n42947 , n42942 , n42945 , n42946 );
and ( n42948 , n42915 , n42947 );
xor ( n42949 , n42714 , n42725 );
xor ( n42950 , n42949 , n42764 );
and ( n42951 , n42947 , n42950 );
and ( n42952 , n42915 , n42950 );
or ( n42953 , n42948 , n42951 , n42952 );
and ( n42954 , n42885 , n42953 );
xor ( n42955 , n42710 , n42712 );
xor ( n42956 , n42955 , n42767 );
and ( n42957 , n42953 , n42956 );
and ( n42958 , n42885 , n42956 );
or ( n42959 , n42954 , n42957 , n42958 );
and ( n42960 , n42862 , n42959 );
and ( n42961 , n42855 , n42959 );
or ( n42962 , n42863 , n42960 , n42961 );
and ( n42963 , n42853 , n42962 );
xor ( n42964 , n42545 , n42590 );
xor ( n42965 , n42964 , n42673 );
and ( n42966 , n42962 , n42965 );
and ( n42967 , n42853 , n42965 );
or ( n42968 , n42963 , n42966 , n42967 );
and ( n42969 , n42851 , n42968 );
xor ( n42970 , n42535 , n42537 );
xor ( n42971 , n42970 , n42540 );
and ( n42972 , n42968 , n42971 );
and ( n42973 , n42851 , n42971 );
or ( n42974 , n42969 , n42972 , n42973 );
xor ( n42975 , n42543 , n42699 );
xor ( n42976 , n42975 , n42702 );
and ( n42977 , n42974 , n42976 );
xor ( n42978 , n42693 , n42695 );
xor ( n42979 , n42665 , n42667 );
xor ( n42980 , n42979 , n42670 );
xor ( n42981 , n42770 , n42837 );
xor ( n42982 , n42981 , n42840 );
and ( n42983 , n42980 , n42982 );
xor ( n42984 , n42683 , n42687 );
xor ( n42985 , n42984 , n42690 );
and ( n42986 , n42982 , n42985 );
and ( n42987 , n42980 , n42985 );
or ( n42988 , n42983 , n42986 , n42987 );
and ( n42989 , n42978 , n42988 );
xor ( n42990 , n42843 , n42845 );
xor ( n42991 , n42990 , n42848 );
and ( n42992 , n42988 , n42991 );
and ( n42993 , n42978 , n42991 );
or ( n42994 , n42989 , n42992 , n42993 );
xor ( n42995 , n42676 , n42678 );
xor ( n42996 , n42995 , n42696 );
and ( n42997 , n42994 , n42996 );
xor ( n42998 , n42853 , n42962 );
xor ( n42999 , n42998 , n42965 );
xor ( n43000 , n42829 , n42831 );
xor ( n43001 , n43000 , n42834 );
xor ( n43002 , n42859 , n42861 );
and ( n43003 , n43001 , n43002 );
xor ( n43004 , n42821 , n42823 );
xor ( n43005 , n43004 , n42826 );
xor ( n43006 , n42786 , n42802 );
xor ( n43007 , n43006 , n42818 );
xor ( n43008 , n42872 , n42876 );
xor ( n43009 , n43008 , n42879 );
and ( n43010 , n43007 , n43009 );
xor ( n43011 , n42790 , n42794 );
xor ( n43012 , n43011 , n42799 );
xor ( n43013 , n42807 , n42812 );
xor ( n43014 , n43013 , n42815 );
and ( n43015 , n43012 , n43014 );
xor ( n43016 , n38149 , n39311 );
buf ( n570318 , n43016 );
buf ( n570319 , n570318 );
buf ( n43019 , n570319 );
and ( n43020 , n43019 , n39375 );
and ( n43021 , n42811 , n39373 );
nor ( n43022 , n43020 , n43021 );
xnor ( n43023 , n43022 , n39380 );
xor ( n43024 , n38150 , n39310 );
buf ( n570326 , n43024 );
buf ( n570327 , n570326 );
buf ( n43027 , n570327 );
and ( n43028 , n43027 , n39367 );
and ( n43029 , n43023 , n43028 );
buf ( n43030 , n557771 );
not ( n43031 , n43030 );
and ( n43032 , n43029 , n43031 );
and ( n43033 , n43014 , n43032 );
and ( n43034 , n43012 , n43032 );
or ( n43035 , n43015 , n43033 , n43034 );
and ( n43036 , n43009 , n43035 );
and ( n43037 , n43007 , n43035 );
or ( n43038 , n43010 , n43036 , n43037 );
and ( n43039 , n43005 , n43038 );
xor ( n43040 , n42865 , n42867 );
xor ( n43041 , n43040 , n42882 );
and ( n43042 , n43038 , n43041 );
and ( n43043 , n43005 , n43041 );
or ( n43044 , n43039 , n43042 , n43043 );
and ( n43045 , n43002 , n43044 );
and ( n43046 , n43001 , n43044 );
or ( n43047 , n43003 , n43045 , n43046 );
xor ( n43048 , n42855 , n42862 );
xor ( n43049 , n43048 , n42959 );
and ( n43050 , n43047 , n43049 );
xor ( n43051 , n42885 , n42953 );
xor ( n43052 , n43051 , n42956 );
xor ( n43053 , n42915 , n42947 );
xor ( n43054 , n43053 , n42950 );
xor ( n43055 , n42887 , n42889 );
xor ( n43056 , n43055 , n42912 );
xor ( n43057 , n42939 , n42941 );
xor ( n43058 , n43057 , n42944 );
and ( n43059 , n43056 , n43058 );
xor ( n43060 , n42891 , n42892 );
xor ( n43061 , n43060 , n42909 );
xor ( n43062 , n42931 , n42933 );
xor ( n43063 , n43062 , n42936 );
and ( n43064 , n43061 , n43063 );
xor ( n43065 , n43023 , n43028 );
and ( n43066 , n43027 , n39375 );
and ( n43067 , n43019 , n39373 );
nor ( n43068 , n43066 , n43067 );
xnor ( n43069 , n43068 , n39380 );
xor ( n43070 , n38151 , n39309 );
buf ( n570372 , n43070 );
buf ( n570373 , n570372 );
buf ( n43073 , n570373 );
and ( n43074 , n43073 , n39367 );
and ( n43075 , n43069 , n43074 );
and ( n43076 , n43065 , n43075 );
buf ( n43077 , n557772 );
not ( n43078 , n43077 );
and ( n43079 , n43075 , n43078 );
and ( n43080 , n43065 , n43078 );
or ( n43081 , n43076 , n43079 , n43080 );
and ( n43082 , n41816 , n39480 );
and ( n43083 , n41807 , n39478 );
nor ( n43084 , n43082 , n43083 );
xnor ( n43085 , n43084 , n39462 );
and ( n43086 , n43081 , n43085 );
and ( n43087 , n42048 , n39396 );
and ( n43088 , n42061 , n39394 );
nor ( n43089 , n43087 , n43088 );
xnor ( n43090 , n43089 , n39401 );
and ( n43091 , n43085 , n43090 );
and ( n43092 , n43081 , n43090 );
or ( n43093 , n43086 , n43091 , n43092 );
and ( n43094 , n43063 , n43093 );
and ( n43095 , n43061 , n43093 );
or ( n43096 , n43064 , n43094 , n43095 );
and ( n43097 , n43058 , n43096 );
and ( n43098 , n43056 , n43096 );
or ( n43099 , n43059 , n43097 , n43098 );
and ( n43100 , n43054 , n43099 );
xor ( n43101 , n43005 , n43038 );
xor ( n43102 , n43101 , n43041 );
and ( n43103 , n43099 , n43102 );
and ( n43104 , n43054 , n43102 );
or ( n43105 , n43100 , n43103 , n43104 );
and ( n43106 , n43052 , n43105 );
xor ( n43107 , n43001 , n43002 );
xor ( n43108 , n43107 , n43044 );
and ( n43109 , n43105 , n43108 );
and ( n43110 , n43052 , n43108 );
or ( n43111 , n43106 , n43109 , n43110 );
and ( n43112 , n43049 , n43111 );
and ( n43113 , n43047 , n43111 );
or ( n43114 , n43050 , n43112 , n43113 );
and ( n43115 , n42999 , n43114 );
xor ( n43116 , n42978 , n42988 );
xor ( n43117 , n43116 , n42991 );
and ( n43118 , n43114 , n43117 );
and ( n43119 , n42999 , n43117 );
or ( n43120 , n43115 , n43118 , n43119 );
and ( n43121 , n42996 , n43120 );
and ( n43122 , n42994 , n43120 );
or ( n43123 , n42997 , n43121 , n43122 );
and ( n43124 , n42976 , n43123 );
and ( n43125 , n42974 , n43123 );
or ( n43126 , n42977 , n43124 , n43125 );
and ( n43127 , n42707 , n43126 );
and ( n43128 , n42705 , n43126 );
or ( n43129 , n42708 , n43127 , n43128 );
and ( n43130 , n42522 , n43129 );
and ( n43131 , n42520 , n43129 );
or ( n43132 , n42523 , n43130 , n43131 );
and ( n43133 , n42233 , n43132 );
xor ( n43134 , n42233 , n43132 );
xor ( n43135 , n42520 , n42522 );
xor ( n43136 , n43135 , n43129 );
xor ( n43137 , n42705 , n42707 );
xor ( n43138 , n43137 , n43126 );
xor ( n43139 , n42974 , n42976 );
xor ( n43140 , n43139 , n43123 );
xor ( n43141 , n42851 , n42968 );
xor ( n43142 , n43141 , n42971 );
xor ( n43143 , n42994 , n42996 );
xor ( n43144 , n43143 , n43120 );
and ( n43145 , n43142 , n43144 );
xor ( n43146 , n42999 , n43114 );
xor ( n43147 , n43146 , n43117 );
xor ( n43148 , n42980 , n42982 );
xor ( n43149 , n43148 , n42985 );
xor ( n43150 , n43047 , n43049 );
xor ( n43151 , n43150 , n43111 );
and ( n43152 , n43149 , n43151 );
xor ( n43153 , n43052 , n43105 );
xor ( n43154 , n43153 , n43108 );
xor ( n43155 , n43007 , n43009 );
xor ( n43156 , n43155 , n43035 );
and ( n43157 , n43019 , n39367 );
xor ( n43158 , n42919 , n42923 );
xor ( n43159 , n43158 , n42928 );
and ( n43160 , n43157 , n43159 );
xor ( n43161 , n43029 , n43031 );
and ( n43162 , n43159 , n43161 );
and ( n43163 , n43157 , n43161 );
or ( n43164 , n43160 , n43162 , n43163 );
xor ( n43165 , n43012 , n43014 );
xor ( n43166 , n43165 , n43032 );
and ( n43167 , n43164 , n43166 );
and ( n43168 , n41047 , n39760 );
and ( n43169 , n40869 , n39758 );
nor ( n43170 , n43168 , n43169 );
xnor ( n43171 , n43170 , n39742 );
xor ( n43172 , n43081 , n43085 );
xor ( n43173 , n43172 , n43090 );
and ( n43174 , n43171 , n43173 );
and ( n43175 , n43166 , n43174 );
and ( n43176 , n43164 , n43174 );
or ( n43177 , n43167 , n43175 , n43176 );
and ( n43178 , n43156 , n43177 );
xor ( n43179 , n43056 , n43058 );
xor ( n43180 , n43179 , n43096 );
and ( n43181 , n43177 , n43180 );
and ( n43182 , n43156 , n43180 );
or ( n43183 , n43178 , n43181 , n43182 );
xor ( n43184 , n43054 , n43099 );
xor ( n43185 , n43184 , n43102 );
and ( n43186 , n43183 , n43185 );
xor ( n43187 , n43061 , n43063 );
xor ( n43188 , n43187 , n43093 );
xor ( n43189 , n38154 , n39307 );
buf ( n570491 , n43189 );
buf ( n570492 , n570491 );
buf ( n43192 , n570492 );
and ( n43193 , n43192 , n39375 );
and ( n43194 , n43073 , n39373 );
nor ( n43195 , n43193 , n43194 );
xnor ( n43196 , n43195 , n39380 );
xor ( n43197 , n38156 , n39306 );
buf ( n570499 , n43197 );
buf ( n570500 , n570499 );
buf ( n43200 , n570500 );
and ( n43201 , n43200 , n39367 );
and ( n43202 , n43196 , n43201 );
and ( n43203 , n43192 , n39367 );
and ( n43204 , n43202 , n43203 );
and ( n43205 , n42811 , n39396 );
and ( n43206 , n42456 , n39394 );
nor ( n43207 , n43205 , n43206 );
xnor ( n43208 , n43207 , n39401 );
and ( n43209 , n43204 , n43208 );
buf ( n43210 , n557773 );
not ( n43211 , n43210 );
and ( n43212 , n43208 , n43211 );
and ( n43213 , n43204 , n43211 );
or ( n43214 , n43209 , n43212 , n43213 );
and ( n43215 , n41807 , n39539 );
and ( n43216 , n41692 , n39537 );
nor ( n43217 , n43215 , n43216 );
xnor ( n43218 , n43217 , n39522 );
and ( n43219 , n43214 , n43218 );
and ( n43220 , n42456 , n39396 );
and ( n43221 , n42048 , n39394 );
nor ( n43222 , n43220 , n43221 );
xnor ( n43223 , n43222 , n39401 );
and ( n43224 , n43218 , n43223 );
and ( n43225 , n43214 , n43223 );
or ( n43226 , n43219 , n43224 , n43225 );
and ( n43227 , n41615 , n39678 );
and ( n43228 , n41182 , n39676 );
nor ( n43229 , n43227 , n43228 );
xnor ( n43230 , n43229 , n39643 );
and ( n43231 , n42061 , n39480 );
and ( n43232 , n41816 , n39478 );
nor ( n43233 , n43231 , n43232 );
xnor ( n43234 , n43233 , n39462 );
and ( n43235 , n43230 , n43234 );
xor ( n43236 , n43065 , n43075 );
xor ( n43237 , n43236 , n43078 );
and ( n43238 , n43234 , n43237 );
and ( n43239 , n43230 , n43237 );
or ( n43240 , n43235 , n43238 , n43239 );
and ( n43241 , n43226 , n43240 );
and ( n43242 , n40738 , n39896 );
and ( n43243 , n40492 , n39894 );
nor ( n43244 , n43242 , n43243 );
xnor ( n43245 , n43244 , n39857 );
and ( n43246 , n43240 , n43245 );
and ( n43247 , n43226 , n43245 );
or ( n43248 , n43241 , n43246 , n43247 );
and ( n43249 , n43188 , n43248 );
and ( n43250 , n39620 , n41984 );
and ( n43251 , n39552 , n41982 );
nor ( n43252 , n43250 , n43251 );
xnor ( n43253 , n43252 , n41687 );
and ( n43254 , n39552 , n42269 );
and ( n43255 , n39493 , n42266 );
nor ( n43256 , n43254 , n43255 );
xnor ( n43257 , n43256 , n41684 );
and ( n43258 , n39653 , n41984 );
and ( n43259 , n39620 , n41982 );
nor ( n43260 , n43258 , n43259 );
xnor ( n43261 , n43260 , n41687 );
and ( n43262 , n43257 , n43261 );
and ( n43263 , n40197 , n40746 );
and ( n43264 , n40148 , n40744 );
nor ( n43265 , n43263 , n43264 );
xnor ( n43266 , n43265 , n40501 );
and ( n43267 , n43261 , n43266 );
and ( n43268 , n43257 , n43266 );
or ( n43269 , n43262 , n43267 , n43268 );
and ( n43270 , n43253 , n43269 );
and ( n43271 , n40388 , n40527 );
and ( n43272 , n40186 , n40525 );
nor ( n43273 , n43271 , n43272 );
xnor ( n43274 , n43273 , n40382 );
and ( n43275 , n39752 , n41622 );
and ( n43276 , n39670 , n41620 );
nor ( n43277 , n43275 , n43276 );
xnor ( n43278 , n43277 , n41194 );
and ( n43279 , n39867 , n41292 );
and ( n43280 , n39795 , n41290 );
nor ( n43281 , n43279 , n43280 );
xnor ( n43282 , n43281 , n41041 );
xor ( n43283 , n43278 , n43282 );
and ( n43284 , n40009 , n41055 );
and ( n43285 , n39948 , n41053 );
nor ( n43286 , n43284 , n43285 );
xnor ( n43287 , n43286 , n40728 );
xor ( n43288 , n43283 , n43287 );
and ( n43289 , n43274 , n43288 );
and ( n43290 , n39620 , n42269 );
and ( n43291 , n39552 , n42266 );
nor ( n43292 , n43290 , n43291 );
xnor ( n43293 , n43292 , n41684 );
and ( n43294 , n40186 , n40746 );
and ( n43295 , n40197 , n40744 );
nor ( n43296 , n43294 , n43295 );
xnor ( n43297 , n43296 , n40501 );
and ( n43298 , n43293 , n43297 );
and ( n43299 , n43288 , n43298 );
and ( n43300 , n43274 , n43298 );
or ( n43301 , n43289 , n43299 , n43300 );
and ( n43302 , n43269 , n43301 );
and ( n43303 , n43253 , n43301 );
or ( n43304 , n43270 , n43302 , n43303 );
xor ( n43305 , n43157 , n43159 );
xor ( n43306 , n43305 , n43161 );
and ( n43307 , n43304 , n43306 );
xor ( n43308 , n43171 , n43173 );
and ( n43309 , n43306 , n43308 );
and ( n43310 , n43304 , n43308 );
or ( n43311 , n43307 , n43309 , n43310 );
and ( n43312 , n43248 , n43311 );
and ( n43313 , n43188 , n43311 );
or ( n43314 , n43249 , n43312 , n43313 );
xor ( n43315 , n43156 , n43177 );
xor ( n43316 , n43315 , n43180 );
and ( n43317 , n43314 , n43316 );
xor ( n43318 , n43069 , n43074 );
and ( n43319 , n43019 , n39396 );
and ( n43320 , n42811 , n39394 );
nor ( n43321 , n43319 , n43320 );
xnor ( n43322 , n43321 , n39401 );
and ( n43323 , n43073 , n39375 );
and ( n43324 , n43027 , n39373 );
nor ( n43325 , n43323 , n43324 );
xnor ( n43326 , n43325 , n39380 );
and ( n43327 , n43322 , n43326 );
buf ( n43328 , n557774 );
not ( n43329 , n43328 );
and ( n43330 , n43326 , n43329 );
and ( n43331 , n43322 , n43329 );
or ( n43332 , n43327 , n43330 , n43331 );
and ( n43333 , n43318 , n43332 );
xor ( n43334 , n43204 , n43208 );
xor ( n43335 , n43334 , n43211 );
and ( n43336 , n43332 , n43335 );
and ( n43337 , n43318 , n43335 );
or ( n43338 , n43333 , n43336 , n43337 );
and ( n43339 , n41032 , n39760 );
and ( n43340 , n41047 , n39758 );
nor ( n43341 , n43339 , n43340 );
xnor ( n43342 , n43341 , n39742 );
and ( n43343 , n43338 , n43342 );
xor ( n43344 , n43214 , n43218 );
xor ( n43345 , n43344 , n43223 );
and ( n43346 , n43342 , n43345 );
and ( n43347 , n43338 , n43345 );
or ( n43348 , n43343 , n43346 , n43347 );
and ( n43349 , n40388 , n40258 );
and ( n43350 , n40186 , n40256 );
nor ( n43351 , n43349 , n43350 );
xnor ( n43352 , n43351 , n40169 );
and ( n43353 , n43348 , n43352 );
and ( n43354 , n40507 , n40053 );
and ( n43355 , n40373 , n40051 );
nor ( n43356 , n43354 , n43355 );
xnor ( n43357 , n43356 , n39999 );
and ( n43358 , n43352 , n43357 );
and ( n43359 , n43348 , n43357 );
or ( n43360 , n43353 , n43358 , n43359 );
and ( n43361 , n39493 , n41984 );
and ( n43362 , n39472 , n41982 );
nor ( n43363 , n43361 , n43362 );
xnor ( n43364 , n43363 , n41687 );
and ( n43365 , n43360 , n43364 );
and ( n43366 , n39620 , n41622 );
and ( n43367 , n39552 , n41620 );
nor ( n43368 , n43366 , n43367 );
xnor ( n43369 , n43368 , n41194 );
and ( n43370 , n43364 , n43369 );
and ( n43371 , n43360 , n43369 );
or ( n43372 , n43365 , n43370 , n43371 );
and ( n43373 , n43316 , n43372 );
and ( n43374 , n43314 , n43372 );
or ( n43375 , n43317 , n43373 , n43374 );
and ( n43376 , n43185 , n43375 );
and ( n43377 , n43183 , n43375 );
or ( n43378 , n43186 , n43376 , n43377 );
and ( n43379 , n43154 , n43378 );
xor ( n43380 , n43164 , n43166 );
xor ( n43381 , n43380 , n43174 );
and ( n43382 , n41692 , n39678 );
and ( n43383 , n41615 , n39676 );
nor ( n43384 , n43382 , n43383 );
xnor ( n43385 , n43384 , n39643 );
and ( n43386 , n41816 , n39539 );
and ( n43387 , n41807 , n39537 );
nor ( n43388 , n43386 , n43387 );
xnor ( n43389 , n43388 , n39522 );
and ( n43390 , n43385 , n43389 );
and ( n43391 , n42048 , n39480 );
and ( n43392 , n42061 , n39478 );
nor ( n43393 , n43391 , n43392 );
xnor ( n43394 , n43393 , n39462 );
and ( n43395 , n43389 , n43394 );
and ( n43396 , n43385 , n43394 );
or ( n43397 , n43390 , n43395 , n43396 );
and ( n43398 , n40492 , n40053 );
and ( n43399 , n40507 , n40051 );
nor ( n43400 , n43398 , n43399 );
xnor ( n43401 , n43400 , n39999 );
and ( n43402 , n43397 , n43401 );
and ( n43403 , n40869 , n39896 );
and ( n43404 , n40738 , n39894 );
nor ( n43405 , n43403 , n43404 );
xnor ( n43406 , n43405 , n39857 );
and ( n43407 , n43401 , n43406 );
and ( n43408 , n43397 , n43406 );
or ( n43409 , n43402 , n43407 , n43408 );
xor ( n43410 , n43226 , n43240 );
xor ( n43411 , n43410 , n43245 );
and ( n43412 , n43409 , n43411 );
and ( n43413 , n43381 , n43412 );
xor ( n43414 , n43188 , n43248 );
xor ( n43415 , n43414 , n43311 );
and ( n43416 , n43412 , n43415 );
and ( n43417 , n43381 , n43415 );
or ( n43418 , n43413 , n43416 , n43417 );
xor ( n43419 , n43360 , n43364 );
xor ( n43420 , n43419 , n43369 );
and ( n43421 , n43200 , n39375 );
and ( n43422 , n43192 , n39373 );
nor ( n43423 , n43421 , n43422 );
xnor ( n43424 , n43423 , n39380 );
xor ( n43425 , n38952 , n39304 );
buf ( n570727 , n43425 );
buf ( n570728 , n570727 );
buf ( n43428 , n570728 );
and ( n43429 , n43428 , n39367 );
xor ( n43430 , n43424 , n43429 );
and ( n570732 , n43428 , n39375 );
and ( n43431 , n43200 , n39373 );
nor ( n43432 , n570732 , n43431 );
xnor ( n43433 , n43432 , n39380 );
xor ( n43434 , n38953 , n39303 );
buf ( n570737 , n43434 );
buf ( n570738 , n570737 );
buf ( n43437 , n570738 );
and ( n43438 , n43437 , n39367 );
and ( n43439 , n43433 , n43438 );
and ( n43440 , n43430 , n43439 );
and ( n43441 , n43073 , n39396 );
and ( n43442 , n43027 , n39394 );
nor ( n43443 , n43441 , n43442 );
xnor ( n43444 , n43443 , n39401 );
and ( n43445 , n43439 , n43444 );
and ( n43446 , n43430 , n43444 );
or ( n43447 , n43440 , n43445 , n43446 );
and ( n43448 , n42811 , n39480 );
and ( n43449 , n42456 , n39478 );
nor ( n43450 , n43448 , n43449 );
xnor ( n43451 , n43450 , n39462 );
and ( n43452 , n43447 , n43451 );
and ( n43453 , n43027 , n39396 );
and ( n43454 , n43019 , n39394 );
nor ( n43455 , n43453 , n43454 );
xnor ( n43456 , n43455 , n39401 );
and ( n43457 , n43451 , n43456 );
and ( n43458 , n43447 , n43456 );
or ( n43459 , n43452 , n43457 , n43458 );
and ( n43460 , n41807 , n39678 );
and ( n43461 , n41692 , n39676 );
nor ( n43462 , n43460 , n43461 );
xnor ( n43463 , n43462 , n39643 );
and ( n43464 , n43459 , n43463 );
and ( n43465 , n42456 , n39480 );
and ( n43466 , n42048 , n39478 );
nor ( n43467 , n43465 , n43466 );
xnor ( n43468 , n43467 , n39462 );
and ( n43469 , n43463 , n43468 );
and ( n43470 , n43459 , n43468 );
or ( n43471 , n43464 , n43469 , n43470 );
xor ( n43472 , n43202 , n43203 );
xor ( n43473 , n43196 , n43201 );
and ( n43474 , n43424 , n43429 );
and ( n43475 , n43473 , n43474 );
buf ( n43476 , n557775 );
not ( n43477 , n43476 );
and ( n43478 , n43474 , n43477 );
and ( n43479 , n43473 , n43477 );
or ( n43480 , n43475 , n43478 , n43479 );
and ( n43481 , n43472 , n43480 );
xor ( n43482 , n43322 , n43326 );
xor ( n43483 , n43482 , n43329 );
and ( n43484 , n43480 , n43483 );
and ( n43485 , n43472 , n43483 );
or ( n43486 , n43481 , n43484 , n43485 );
and ( n43487 , n43471 , n43486 );
and ( n43488 , n41182 , n39760 );
and ( n43489 , n41032 , n39758 );
nor ( n43490 , n43488 , n43489 );
xnor ( n43491 , n43490 , n39742 );
and ( n43492 , n43486 , n43491 );
and ( n43493 , n43471 , n43491 );
or ( n43494 , n43487 , n43492 , n43493 );
and ( n43495 , n40373 , n40258 );
and ( n43496 , n40388 , n40256 );
nor ( n43497 , n43495 , n43496 );
xnor ( n43498 , n43497 , n40169 );
and ( n43499 , n43494 , n43498 );
xor ( n43500 , n43230 , n43234 );
xor ( n43501 , n43500 , n43237 );
and ( n43502 , n43498 , n43501 );
and ( n43503 , n43494 , n43501 );
or ( n43504 , n43499 , n43502 , n43503 );
and ( n43505 , n39752 , n41292 );
and ( n43506 , n39670 , n41290 );
nor ( n43507 , n43505 , n43506 );
xnor ( n43508 , n43507 , n41041 );
and ( n43509 , n43504 , n43508 );
and ( n43510 , n40197 , n40527 );
and ( n43511 , n40148 , n40525 );
nor ( n43512 , n43510 , n43511 );
xnor ( n43513 , n43512 , n40382 );
and ( n43514 , n43508 , n43513 );
and ( n43515 , n43504 , n43513 );
or ( n43516 , n43509 , n43514 , n43515 );
and ( n43517 , n43420 , n43516 );
and ( n43518 , n39552 , n41984 );
and ( n43519 , n39493 , n41982 );
nor ( n43520 , n43518 , n43519 );
xnor ( n43521 , n43520 , n41687 );
and ( n43522 , n39653 , n41622 );
and ( n43523 , n39620 , n41620 );
nor ( n43524 , n43522 , n43523 );
xnor ( n43525 , n43524 , n41194 );
and ( n43526 , n43521 , n43525 );
xor ( n43527 , n43348 , n43352 );
xor ( n43528 , n43527 , n43357 );
and ( n43529 , n43525 , n43528 );
and ( n43530 , n43521 , n43528 );
or ( n43531 , n43526 , n43529 , n43530 );
and ( n43532 , n43516 , n43531 );
and ( n43533 , n43420 , n43531 );
or ( n43534 , n43517 , n43532 , n43533 );
and ( n43535 , n43418 , n43534 );
xor ( n43536 , n43314 , n43316 );
xor ( n43537 , n43536 , n43372 );
and ( n43538 , n43534 , n43537 );
and ( n43539 , n43418 , n43537 );
or ( n43540 , n43535 , n43538 , n43539 );
xor ( n43541 , n43183 , n43185 );
xor ( n43542 , n43541 , n43375 );
and ( n43543 , n43540 , n43542 );
and ( n43544 , n39670 , n41984 );
and ( n43545 , n39653 , n41982 );
nor ( n43546 , n43544 , n43545 );
xnor ( n43547 , n43546 , n41687 );
and ( n43548 , n39795 , n41622 );
and ( n43549 , n39752 , n41620 );
nor ( n43550 , n43548 , n43549 );
xnor ( n43551 , n43550 , n41194 );
and ( n43552 , n43547 , n43551 );
and ( n43553 , n39948 , n41292 );
and ( n43554 , n39867 , n41290 );
nor ( n43555 , n43553 , n43554 );
xnor ( n43556 , n43555 , n41041 );
and ( n43557 , n43551 , n43556 );
and ( n43558 , n43547 , n43556 );
or ( n43559 , n43552 , n43557 , n43558 );
and ( n43560 , n40148 , n41055 );
and ( n43561 , n40009 , n41053 );
nor ( n43562 , n43560 , n43561 );
xnor ( n43563 , n43562 , n40728 );
and ( n43564 , n40373 , n40527 );
and ( n43565 , n40388 , n40525 );
nor ( n43566 , n43564 , n43565 );
xnor ( n43567 , n43566 , n40382 );
and ( n43568 , n43563 , n43567 );
and ( n43569 , n40869 , n40053 );
and ( n43570 , n40738 , n40051 );
nor ( n43571 , n43569 , n43570 );
xnor ( n43572 , n43571 , n39999 );
and ( n43573 , n43567 , n43572 );
and ( n43574 , n43563 , n43572 );
or ( n43575 , n43568 , n43573 , n43574 );
and ( n43576 , n43559 , n43575 );
xor ( n43577 , n43257 , n43261 );
xor ( n43578 , n43577 , n43266 );
and ( n43579 , n43575 , n43578 );
and ( n43580 , n43559 , n43578 );
or ( n43581 , n43576 , n43579 , n43580 );
and ( n43582 , n41032 , n39896 );
and ( n43583 , n41047 , n39894 );
nor ( n43584 , n43582 , n43583 );
xnor ( n43585 , n43584 , n39857 );
xor ( n43586 , n43293 , n43297 );
and ( n43587 , n43585 , n43586 );
and ( n43588 , n39653 , n42269 );
and ( n43589 , n39620 , n42266 );
nor ( n43590 , n43588 , n43589 );
xnor ( n43591 , n43590 , n41684 );
and ( n43592 , n39752 , n41984 );
and ( n43593 , n39670 , n41982 );
nor ( n43594 , n43592 , n43593 );
xnor ( n43595 , n43594 , n41687 );
and ( n43596 , n43591 , n43595 );
and ( n43597 , n40197 , n41055 );
and ( n43598 , n40148 , n41053 );
nor ( n43599 , n43597 , n43598 );
xnor ( n43600 , n43599 , n40728 );
and ( n43601 , n43595 , n43600 );
and ( n43602 , n43591 , n43600 );
or ( n43603 , n43596 , n43601 , n43602 );
and ( n43604 , n43586 , n43603 );
and ( n43605 , n43585 , n43603 );
or ( n43606 , n43587 , n43604 , n43605 );
and ( n43607 , n39867 , n41622 );
and ( n43608 , n39795 , n41620 );
nor ( n43609 , n43607 , n43608 );
xnor ( n43610 , n43609 , n41194 );
and ( n43611 , n40009 , n41292 );
and ( n43612 , n39948 , n41290 );
nor ( n43613 , n43611 , n43612 );
xnor ( n43614 , n43613 , n41041 );
and ( n43615 , n43610 , n43614 );
and ( n43616 , n40388 , n40746 );
and ( n43617 , n40186 , n40744 );
nor ( n43618 , n43616 , n43617 );
xnor ( n43619 , n43618 , n40501 );
and ( n43620 , n40507 , n40527 );
and ( n43621 , n40373 , n40525 );
nor ( n43622 , n43620 , n43621 );
xnor ( n43623 , n43622 , n40382 );
and ( n43624 , n43619 , n43623 );
and ( n43625 , n40738 , n40258 );
and ( n43626 , n40492 , n40256 );
nor ( n43627 , n43625 , n43626 );
xnor ( n43628 , n43627 , n40169 );
and ( n43629 , n43623 , n43628 );
and ( n43630 , n43619 , n43628 );
or ( n43631 , n43624 , n43629 , n43630 );
and ( n43632 , n43615 , n43631 );
and ( n43633 , n41047 , n40053 );
and ( n43634 , n40869 , n40051 );
nor ( n43635 , n43633 , n43634 );
xnor ( n43636 , n43635 , n39999 );
and ( n43637 , n41692 , n39760 );
and ( n43638 , n41615 , n39758 );
nor ( n43639 , n43637 , n43638 );
xnor ( n43640 , n43639 , n39742 );
and ( n43641 , n43636 , n43640 );
and ( n43642 , n41816 , n39678 );
and ( n43643 , n41807 , n39676 );
nor ( n43644 , n43642 , n43643 );
xnor ( n43645 , n43644 , n39643 );
and ( n43646 , n43640 , n43645 );
and ( n43647 , n43636 , n43645 );
or ( n43648 , n43641 , n43646 , n43647 );
and ( n43649 , n43631 , n43648 );
and ( n43650 , n43615 , n43648 );
or ( n43651 , n43632 , n43649 , n43650 );
and ( n43652 , n43606 , n43651 );
xor ( n43653 , n43274 , n43288 );
xor ( n43654 , n43653 , n43298 );
and ( n43655 , n43651 , n43654 );
and ( n43656 , n43606 , n43654 );
or ( n43657 , n43652 , n43655 , n43656 );
and ( n43658 , n43581 , n43657 );
xor ( n43659 , n43253 , n43269 );
xor ( n43660 , n43659 , n43301 );
and ( n43661 , n43657 , n43660 );
and ( n43662 , n43581 , n43660 );
or ( n43663 , n43658 , n43661 , n43662 );
xor ( n43664 , n43304 , n43306 );
xor ( n43665 , n43664 , n43308 );
and ( n43666 , n43663 , n43665 );
xor ( n43667 , n43409 , n43411 );
and ( n43668 , n43665 , n43667 );
and ( n43669 , n43663 , n43667 );
or ( n43670 , n43666 , n43668 , n43669 );
xor ( n570973 , n43381 , n43412 );
xor ( n43671 , n570973 , n43415 );
and ( n43672 , n43670 , n43671 );
and ( n43673 , n41615 , n39760 );
and ( n43674 , n41182 , n39758 );
nor ( n43675 , n43673 , n43674 );
xnor ( n43676 , n43675 , n39742 );
and ( n43677 , n42061 , n39539 );
and ( n43678 , n41816 , n39537 );
nor ( n43679 , n43677 , n43678 );
xnor ( n43680 , n43679 , n39522 );
and ( n43681 , n43676 , n43680 );
xor ( n43682 , n43472 , n43480 );
xor ( n43683 , n43682 , n43483 );
and ( n43684 , n43680 , n43683 );
and ( n43685 , n43676 , n43683 );
or ( n43686 , n43681 , n43684 , n43685 );
and ( n43687 , n40507 , n40258 );
and ( n43688 , n40373 , n40256 );
nor ( n43689 , n43687 , n43688 );
xnor ( n43690 , n43689 , n40169 );
and ( n43691 , n43686 , n43690 );
xor ( n43692 , n43385 , n43389 );
xor ( n43693 , n43692 , n43394 );
and ( n43694 , n43690 , n43693 );
and ( n43695 , n43686 , n43693 );
or ( n43696 , n43691 , n43694 , n43695 );
and ( n43697 , n39670 , n41622 );
and ( n43698 , n39653 , n41620 );
nor ( n43699 , n43697 , n43698 );
xnor ( n43700 , n43699 , n41194 );
and ( n43701 , n43696 , n43700 );
and ( n43702 , n40186 , n40527 );
and ( n43703 , n40197 , n40525 );
nor ( n43704 , n43702 , n43703 );
xnor ( n43705 , n43704 , n40382 );
and ( n43706 , n43700 , n43705 );
and ( n43707 , n43696 , n43705 );
or ( n43708 , n43701 , n43706 , n43707 );
xor ( n43709 , n42897 , n42901 );
xor ( n43710 , n43709 , n42906 );
and ( n43711 , n43708 , n43710 );
xor ( n43712 , n43504 , n43508 );
xor ( n43713 , n43712 , n43513 );
and ( n43714 , n43710 , n43713 );
and ( n43715 , n43708 , n43713 );
or ( n43716 , n43711 , n43714 , n43715 );
and ( n43717 , n43671 , n43716 );
and ( n43718 , n43670 , n43716 );
or ( n43719 , n43672 , n43717 , n43718 );
and ( n43720 , n39493 , n42269 );
and ( n43721 , n39472 , n42266 );
nor ( n43722 , n43720 , n43721 );
xnor ( n43723 , n43722 , n41684 );
and ( n43724 , n40148 , n40746 );
and ( n43725 , n40009 , n40744 );
nor ( n43726 , n43724 , n43725 );
xnor ( n43727 , n43726 , n40501 );
and ( n43728 , n43723 , n43727 );
and ( n43729 , n40738 , n40053 );
and ( n43730 , n40492 , n40051 );
nor ( n43731 , n43729 , n43730 );
xnor ( n43732 , n43731 , n39999 );
and ( n43733 , n41047 , n39896 );
and ( n43734 , n40869 , n39894 );
nor ( n43735 , n43733 , n43734 );
xnor ( n43736 , n43735 , n39857 );
and ( n43737 , n43732 , n43736 );
xor ( n43738 , n43318 , n43332 );
xor ( n43739 , n43738 , n43335 );
and ( n43740 , n43736 , n43739 );
and ( n43741 , n43732 , n43739 );
or ( n43742 , n43737 , n43740 , n43741 );
xor ( n43743 , n43397 , n43401 );
xor ( n43744 , n43743 , n43406 );
xor ( n43745 , n43742 , n43744 );
xor ( n43746 , n43338 , n43342 );
xor ( n43747 , n43746 , n43345 );
xor ( n43748 , n43745 , n43747 );
and ( n43749 , n43727 , n43748 );
and ( n43750 , n43723 , n43748 );
or ( n43751 , n43728 , n43749 , n43750 );
xor ( n43752 , n43521 , n43525 );
xor ( n43753 , n43752 , n43528 );
and ( n43754 , n43751 , n43753 );
and ( n43755 , n43742 , n43744 );
and ( n43756 , n43744 , n43747 );
and ( n43757 , n43742 , n43747 );
or ( n43758 , n43755 , n43756 , n43757 );
xor ( n43759 , n43559 , n43575 );
xor ( n43760 , n43759 , n43578 );
xor ( n43761 , n43547 , n43551 );
xor ( n43762 , n43761 , n43556 );
xor ( n43763 , n43563 , n43567 );
xor ( n43764 , n43763 , n43572 );
and ( n43765 , n43762 , n43764 );
xor ( n43766 , n43591 , n43595 );
xor ( n43767 , n43766 , n43600 );
xor ( n43768 , n43610 , n43614 );
and ( n43769 , n43767 , n43768 );
and ( n43770 , n39670 , n42269 );
and ( n43771 , n39653 , n42266 );
nor ( n43772 , n43770 , n43771 );
xnor ( n43773 , n43772 , n41684 );
and ( n43774 , n40148 , n41292 );
and ( n43775 , n40009 , n41290 );
nor ( n43776 , n43774 , n43775 );
xnor ( n43777 , n43776 , n41041 );
and ( n43778 , n43773 , n43777 );
and ( n43779 , n40186 , n41055 );
and ( n43780 , n40197 , n41053 );
nor ( n43781 , n43779 , n43780 );
xnor ( n43782 , n43781 , n40728 );
and ( n43783 , n43777 , n43782 );
and ( n43784 , n43773 , n43782 );
or ( n43785 , n43778 , n43783 , n43784 );
and ( n43786 , n43768 , n43785 );
and ( n43787 , n43767 , n43785 );
or ( n43788 , n43769 , n43786 , n43787 );
and ( n43789 , n43764 , n43788 );
and ( n43790 , n43762 , n43788 );
or ( n43791 , n43765 , n43789 , n43790 );
and ( n43792 , n43760 , n43791 );
and ( n43793 , n41615 , n39896 );
and ( n43794 , n41182 , n39894 );
nor ( n43795 , n43793 , n43794 );
xnor ( n43796 , n43795 , n39857 );
and ( n43797 , n41807 , n39760 );
and ( n43798 , n41692 , n39758 );
nor ( n43799 , n43797 , n43798 );
xnor ( n43800 , n43799 , n39742 );
and ( n43801 , n43796 , n43800 );
and ( n43802 , n39795 , n41984 );
and ( n43803 , n39752 , n41982 );
nor ( n43804 , n43802 , n43803 );
xnor ( n43805 , n43804 , n41687 );
and ( n43806 , n39948 , n41622 );
and ( n43807 , n39867 , n41620 );
nor ( n43808 , n43806 , n43807 );
xnor ( n43809 , n43808 , n41194 );
and ( n43810 , n43805 , n43809 );
and ( n43811 , n40373 , n40746 );
and ( n43812 , n40388 , n40744 );
nor ( n43813 , n43811 , n43812 );
xnor ( n43814 , n43813 , n40501 );
and ( n43815 , n43809 , n43814 );
and ( n43816 , n43805 , n43814 );
or ( n43817 , n43810 , n43815 , n43816 );
and ( n43818 , n43801 , n43817 );
and ( n43819 , n40492 , n40527 );
and ( n43820 , n40507 , n40525 );
nor ( n43821 , n43819 , n43820 );
xnor ( n43822 , n43821 , n40382 );
and ( n43823 , n40869 , n40258 );
and ( n43824 , n40738 , n40256 );
nor ( n43825 , n43823 , n43824 );
xnor ( n43826 , n43825 , n40169 );
and ( n43827 , n43822 , n43826 );
and ( n43828 , n41032 , n40053 );
and ( n43829 , n41047 , n40051 );
nor ( n43830 , n43828 , n43829 );
xnor ( n43831 , n43830 , n39999 );
and ( n43832 , n43826 , n43831 );
and ( n43833 , n43822 , n43831 );
or ( n43834 , n43827 , n43832 , n43833 );
and ( n43835 , n43817 , n43834 );
and ( n43836 , n43801 , n43834 );
or ( n43837 , n43818 , n43835 , n43836 );
and ( n43838 , n42061 , n39678 );
and ( n43839 , n41816 , n39676 );
nor ( n43840 , n43838 , n43839 );
xnor ( n43841 , n43840 , n39643 );
and ( n43842 , n42456 , n39539 );
and ( n43843 , n42048 , n39537 );
nor ( n43844 , n43842 , n43843 );
xnor ( n43845 , n43844 , n39522 );
and ( n43846 , n43841 , n43845 );
and ( n43847 , n43019 , n39480 );
and ( n43848 , n42811 , n39478 );
nor ( n43849 , n43847 , n43848 );
xnor ( n43850 , n43849 , n39462 );
and ( n43851 , n43845 , n43850 );
and ( n43852 , n43841 , n43850 );
or ( n43853 , n43846 , n43851 , n43852 );
xor ( n43854 , n43619 , n43623 );
xor ( n43855 , n43854 , n43628 );
and ( n43856 , n43853 , n43855 );
xor ( n43857 , n43636 , n43640 );
xor ( n43858 , n43857 , n43645 );
and ( n43859 , n43855 , n43858 );
and ( n43860 , n43853 , n43858 );
or ( n43861 , n43856 , n43859 , n43860 );
and ( n43862 , n43837 , n43861 );
xor ( n43863 , n43585 , n43586 );
xor ( n43864 , n43863 , n43603 );
and ( n43865 , n43861 , n43864 );
and ( n43866 , n43837 , n43864 );
or ( n43867 , n43862 , n43865 , n43866 );
and ( n43868 , n43791 , n43867 );
and ( n43869 , n43760 , n43867 );
or ( n43870 , n43792 , n43868 , n43869 );
xor ( n43871 , n43581 , n43657 );
xor ( n43872 , n43871 , n43660 );
and ( n43873 , n43870 , n43872 );
xor ( n43874 , n43606 , n43651 );
xor ( n43875 , n43874 , n43654 );
xor ( n43876 , n43615 , n43631 );
xor ( n43877 , n43876 , n43648 );
xor ( n43878 , n43473 , n43474 );
xor ( n43879 , n43878 , n43477 );
buf ( n43880 , n557776 );
not ( n43881 , n43880 );
xor ( n43882 , n43773 , n43777 );
xor ( n43883 , n43882 , n43782 );
and ( n43884 , n43881 , n43883 );
xor ( n43885 , n43796 , n43800 );
and ( n43886 , n43883 , n43885 );
and ( n43887 , n43881 , n43885 );
or ( n43888 , n43884 , n43886 , n43887 );
and ( n43889 , n43879 , n43888 );
and ( n43890 , n39752 , n42269 );
and ( n43891 , n39670 , n42266 );
nor ( n43892 , n43890 , n43891 );
xnor ( n43893 , n43892 , n41684 );
and ( n43894 , n39867 , n41984 );
and ( n43895 , n39795 , n41982 );
nor ( n43896 , n43894 , n43895 );
xnor ( n43897 , n43896 , n41687 );
and ( n43898 , n43893 , n43897 );
and ( n43899 , n40197 , n41292 );
and ( n43900 , n40148 , n41290 );
nor ( n43901 , n43899 , n43900 );
xnor ( n43902 , n43901 , n41041 );
and ( n43903 , n43897 , n43902 );
and ( n43904 , n43893 , n43902 );
or ( n43905 , n43898 , n43903 , n43904 );
and ( n43906 , n42811 , n39539 );
and ( n43907 , n42456 , n39537 );
nor ( n43908 , n43906 , n43907 );
xnor ( n43909 , n43908 , n39522 );
and ( n43910 , n43027 , n39480 );
and ( n43911 , n43019 , n39478 );
nor ( n43912 , n43910 , n43911 );
xnor ( n43913 , n43912 , n39462 );
and ( n43914 , n43909 , n43913 );
and ( n43915 , n43905 , n43914 );
and ( n43916 , n40009 , n41622 );
and ( n43917 , n39948 , n41620 );
nor ( n43918 , n43916 , n43917 );
xnor ( n43919 , n43918 , n41194 );
and ( n43920 , n40388 , n41055 );
and ( n43921 , n40186 , n41053 );
nor ( n43922 , n43920 , n43921 );
xnor ( n43923 , n43922 , n40728 );
and ( n43924 , n43919 , n43923 );
and ( n43925 , n40507 , n40746 );
and ( n43926 , n40373 , n40744 );
nor ( n43927 , n43925 , n43926 );
xnor ( n43928 , n43927 , n40501 );
and ( n43929 , n43923 , n43928 );
and ( n43930 , n43919 , n43928 );
or ( n43931 , n43924 , n43929 , n43930 );
and ( n43932 , n43914 , n43931 );
and ( n43933 , n43905 , n43931 );
or ( n43934 , n43915 , n43932 , n43933 );
and ( n43935 , n43888 , n43934 );
and ( n43936 , n43879 , n43934 );
or ( n43937 , n43889 , n43935 , n43936 );
and ( n43938 , n43877 , n43937 );
and ( n43939 , n40738 , n40527 );
and ( n43940 , n40492 , n40525 );
nor ( n43941 , n43939 , n43940 );
xnor ( n43942 , n43941 , n40382 );
and ( n43943 , n41047 , n40258 );
and ( n43944 , n40869 , n40256 );
nor ( n43945 , n43943 , n43944 );
xnor ( n43946 , n43945 , n40169 );
and ( n43947 , n43942 , n43946 );
and ( n43948 , n41182 , n40053 );
and ( n43949 , n41032 , n40051 );
nor ( n43950 , n43948 , n43949 );
xnor ( n43951 , n43950 , n39999 );
and ( n43952 , n43946 , n43951 );
and ( n43953 , n43942 , n43951 );
or ( n43954 , n43947 , n43952 , n43953 );
and ( n43955 , n41692 , n39896 );
and ( n43956 , n41615 , n39894 );
nor ( n43957 , n43955 , n43956 );
xnor ( n43958 , n43957 , n39857 );
and ( n43959 , n41816 , n39760 );
and ( n43960 , n41807 , n39758 );
nor ( n43961 , n43959 , n43960 );
xnor ( n43962 , n43961 , n39742 );
and ( n43963 , n43958 , n43962 );
and ( n43964 , n42048 , n39678 );
and ( n43965 , n42061 , n39676 );
nor ( n43966 , n43964 , n43965 );
xnor ( n43967 , n43966 , n39643 );
and ( n43968 , n43962 , n43967 );
and ( n43969 , n43958 , n43967 );
or ( n43970 , n43963 , n43968 , n43969 );
and ( n43971 , n43954 , n43970 );
xor ( n43972 , n43805 , n43809 );
xor ( n43973 , n43972 , n43814 );
and ( n43974 , n43970 , n43973 );
and ( n43975 , n43954 , n43973 );
or ( n43976 , n43971 , n43974 , n43975 );
xor ( n43977 , n43767 , n43768 );
xor ( n43978 , n43977 , n43785 );
and ( n43979 , n43976 , n43978 );
xor ( n43980 , n43801 , n43817 );
xor ( n43981 , n43980 , n43834 );
and ( n43982 , n43978 , n43981 );
and ( n43983 , n43976 , n43981 );
or ( n43984 , n43979 , n43982 , n43983 );
and ( n43985 , n43937 , n43984 );
and ( n43986 , n43877 , n43984 );
or ( n43987 , n43938 , n43985 , n43986 );
and ( n43988 , n43875 , n43987 );
xor ( n43989 , n43760 , n43791 );
xor ( n43990 , n43989 , n43867 );
and ( n43991 , n43987 , n43990 );
and ( n43992 , n43875 , n43990 );
or ( n43993 , n43988 , n43991 , n43992 );
and ( n43994 , n43872 , n43993 );
and ( n43995 , n43870 , n43993 );
or ( n43996 , n43873 , n43994 , n43995 );
and ( n43997 , n43758 , n43996 );
and ( n43998 , n39795 , n41292 );
and ( n43999 , n39752 , n41290 );
nor ( n44000 , n43998 , n43999 );
xnor ( n44001 , n44000 , n41041 );
and ( n44002 , n39948 , n41055 );
and ( n44003 , n39867 , n41053 );
nor ( n44004 , n44002 , n44003 );
xnor ( n44005 , n44004 , n40728 );
and ( n44006 , n44001 , n44005 );
xor ( n44007 , n43494 , n43498 );
xor ( n44008 , n44007 , n43501 );
and ( n44009 , n44005 , n44008 );
and ( n44010 , n44001 , n44008 );
or ( n44011 , n44006 , n44009 , n44010 );
and ( n44012 , n43996 , n44011 );
and ( n44013 , n43758 , n44011 );
or ( n44014 , n43997 , n44012 , n44013 );
and ( n44015 , n43754 , n44014 );
xor ( n44016 , n43420 , n43516 );
xor ( n44017 , n44016 , n43531 );
and ( n44018 , n44014 , n44017 );
and ( n44019 , n43754 , n44017 );
or ( n44020 , n44015 , n44018 , n44019 );
and ( n44021 , n43719 , n44020 );
xor ( n44022 , n43418 , n43534 );
xor ( n44023 , n44022 , n43537 );
and ( n44024 , n44020 , n44023 );
and ( n44025 , n43719 , n44023 );
or ( n44026 , n44021 , n44024 , n44025 );
and ( n44027 , n43542 , n44026 );
and ( n44028 , n43540 , n44026 );
or ( n44029 , n43543 , n44027 , n44028 );
and ( n44030 , n43378 , n44029 );
and ( n44031 , n43154 , n44029 );
or ( n44032 , n43379 , n44030 , n44031 );
and ( n44033 , n43151 , n44032 );
and ( n44034 , n43149 , n44032 );
or ( n44035 , n43152 , n44033 , n44034 );
or ( n44036 , n43147 , n44035 );
and ( n44037 , n43144 , n44036 );
and ( n44038 , n43142 , n44036 );
or ( n44039 , n43145 , n44037 , n44038 );
or ( n44040 , n43140 , n44039 );
or ( n44041 , n43138 , n44040 );
and ( n44042 , n43136 , n44041 );
xor ( n44043 , n43136 , n44041 );
xnor ( n44044 , n43138 , n44040 );
xnor ( n44045 , n43140 , n44039 );
xor ( n44046 , n43142 , n43144 );
xor ( n44047 , n44046 , n44036 );
not ( n44048 , n44047 );
xnor ( n44049 , n43147 , n44035 );
xor ( n44050 , n43149 , n43151 );
xor ( n44051 , n44050 , n44032 );
xor ( n44052 , n43154 , n43378 );
xor ( n44053 , n44052 , n44029 );
xor ( n44054 , n43540 , n43542 );
xor ( n44055 , n44054 , n44026 );
and ( n44056 , n41182 , n39896 );
and ( n44057 , n41032 , n39894 );
nor ( n44058 , n44056 , n44057 );
xnor ( n44059 , n44058 , n39857 );
and ( n44060 , n42048 , n39539 );
and ( n44061 , n42061 , n39537 );
nor ( n44062 , n44060 , n44061 );
xnor ( n44063 , n44062 , n39522 );
and ( n44064 , n44059 , n44063 );
xor ( n44065 , n43447 , n43451 );
xor ( n44066 , n44065 , n43456 );
and ( n44067 , n44063 , n44066 );
and ( n44068 , n44059 , n44066 );
or ( n44069 , n44064 , n44067 , n44068 );
and ( n44070 , n40492 , n40258 );
and ( n44071 , n40507 , n40256 );
nor ( n44072 , n44070 , n44071 );
xnor ( n44073 , n44072 , n40169 );
and ( n44074 , n44069 , n44073 );
xor ( n44075 , n43459 , n43463 );
xor ( n44076 , n44075 , n43468 );
and ( n44077 , n44073 , n44076 );
and ( n44078 , n44069 , n44076 );
or ( n44079 , n44074 , n44077 , n44078 );
xor ( n44080 , n43686 , n43690 );
xor ( n44081 , n44080 , n43693 );
and ( n44082 , n44079 , n44081 );
xor ( n44083 , n43732 , n43736 );
xor ( n44084 , n44083 , n43739 );
and ( n44085 , n44081 , n44084 );
and ( n44086 , n44079 , n44084 );
or ( n44087 , n44082 , n44085 , n44086 );
xor ( n44088 , n43471 , n43486 );
xor ( n44089 , n44088 , n43491 );
xor ( n44090 , n43762 , n43764 );
xor ( n44091 , n44090 , n43788 );
xor ( n44092 , n43837 , n43861 );
xor ( n44093 , n44092 , n43864 );
and ( n44094 , n44091 , n44093 );
xor ( n44095 , n43676 , n43680 );
xor ( n44096 , n44095 , n43683 );
and ( n44097 , n44093 , n44096 );
and ( n44098 , n44091 , n44096 );
or ( n44099 , n44094 , n44097 , n44098 );
and ( n44100 , n44089 , n44099 );
xor ( n44101 , n43853 , n43855 );
xor ( n44102 , n44101 , n43858 );
xor ( n44103 , n43822 , n43826 );
xor ( n44104 , n44103 , n43831 );
xor ( n44105 , n43841 , n43845 );
xor ( n44106 , n44105 , n43850 );
and ( n44107 , n44104 , n44106 );
xor ( n44108 , n43430 , n43439 );
xor ( n44109 , n44108 , n43444 );
and ( n44110 , n44106 , n44109 );
and ( n44111 , n44104 , n44109 );
or ( n44112 , n44107 , n44110 , n44111 );
and ( n44113 , n44102 , n44112 );
and ( n44114 , n43192 , n39396 );
and ( n44115 , n43073 , n39394 );
nor ( n44116 , n44114 , n44115 );
xnor ( n44117 , n44116 , n39401 );
buf ( n44118 , n557777 );
not ( n44119 , n44118 );
and ( n44120 , n44117 , n44119 );
xor ( n44121 , n43893 , n43897 );
xor ( n44122 , n44121 , n43902 );
and ( n44123 , n44119 , n44122 );
and ( n44124 , n44117 , n44122 );
or ( n44125 , n44120 , n44123 , n44124 );
xor ( n44126 , n43433 , n43438 );
xor ( n44127 , n43909 , n43913 );
and ( n44128 , n44126 , n44127 );
and ( n44129 , n41032 , n40258 );
and ( n44130 , n41047 , n40256 );
nor ( n44131 , n44129 , n44130 );
xnor ( n44132 , n44131 , n40169 );
and ( n44133 , n41615 , n40053 );
and ( n44134 , n41182 , n40051 );
nor ( n44135 , n44133 , n44134 );
xnor ( n44136 , n44135 , n39999 );
and ( n44137 , n44132 , n44136 );
and ( n44138 , n42061 , n39760 );
and ( n44139 , n41816 , n39758 );
nor ( n44140 , n44138 , n44139 );
xnor ( n44141 , n44140 , n39742 );
and ( n44142 , n44136 , n44141 );
and ( n44143 , n44132 , n44141 );
or ( n44144 , n44137 , n44142 , n44143 );
and ( n44145 , n44127 , n44144 );
and ( n44146 , n44126 , n44144 );
or ( n44147 , n44128 , n44145 , n44146 );
and ( n44148 , n44125 , n44147 );
and ( n44149 , n43200 , n39396 );
and ( n44150 , n43192 , n39394 );
nor ( n44151 , n44149 , n44150 );
xnor ( n44152 , n44151 , n39401 );
and ( n44153 , n43437 , n39375 );
and ( n44154 , n43428 , n39373 );
nor ( n44155 , n44153 , n44154 );
xnor ( n44156 , n44155 , n39380 );
and ( n44157 , n44152 , n44156 );
and ( n44158 , n39795 , n42269 );
and ( n44159 , n39752 , n42266 );
nor ( n44160 , n44158 , n44159 );
xnor ( n44161 , n44160 , n41684 );
and ( n44162 , n40186 , n41292 );
and ( n44163 , n40197 , n41290 );
nor ( n44164 , n44162 , n44163 );
xnor ( n44165 , n44164 , n41041 );
and ( n44166 , n44161 , n44165 );
and ( n44167 , n40869 , n40527 );
and ( n44168 , n40738 , n40525 );
nor ( n44169 , n44167 , n44168 );
xnor ( n44170 , n44169 , n40382 );
and ( n44171 , n44165 , n44170 );
and ( n44172 , n44161 , n44170 );
or ( n44173 , n44166 , n44171 , n44172 );
and ( n44174 , n44157 , n44173 );
xor ( n44175 , n43919 , n43923 );
xor ( n44176 , n44175 , n43928 );
and ( n44177 , n44173 , n44176 );
and ( n44178 , n44157 , n44176 );
or ( n44179 , n44174 , n44177 , n44178 );
and ( n44180 , n44147 , n44179 );
and ( n44181 , n44125 , n44179 );
or ( n44182 , n44148 , n44180 , n44181 );
and ( n44183 , n44112 , n44182 );
and ( n44184 , n44102 , n44182 );
or ( n44185 , n44113 , n44183 , n44184 );
xor ( n44186 , n43881 , n43883 );
xor ( n44187 , n44186 , n43885 );
xor ( n44188 , n43905 , n43914 );
xor ( n44189 , n44188 , n43931 );
and ( n44190 , n44187 , n44189 );
xor ( n44191 , n43954 , n43970 );
xor ( n44192 , n44191 , n43973 );
and ( n44193 , n44189 , n44192 );
and ( n44194 , n44187 , n44192 );
or ( n44195 , n44190 , n44193 , n44194 );
xor ( n44196 , n43879 , n43888 );
xor ( n44197 , n44196 , n43934 );
and ( n44198 , n44195 , n44197 );
xor ( n44199 , n43976 , n43978 );
xor ( n44200 , n44199 , n43981 );
and ( n44201 , n44197 , n44200 );
and ( n44202 , n44195 , n44200 );
or ( n44203 , n44198 , n44201 , n44202 );
and ( n44204 , n44185 , n44203 );
xor ( n44205 , n43877 , n43937 );
xor ( n44206 , n44205 , n43984 );
and ( n44207 , n44203 , n44206 );
and ( n44208 , n44185 , n44206 );
or ( n44209 , n44204 , n44207 , n44208 );
and ( n44210 , n44099 , n44209 );
and ( n44211 , n44089 , n44209 );
or ( n44212 , n44100 , n44210 , n44211 );
and ( n44213 , n44087 , n44212 );
xor ( n44214 , n43870 , n43872 );
xor ( n44215 , n44214 , n43993 );
and ( n44216 , n44212 , n44215 );
and ( n44217 , n44087 , n44215 );
or ( n44218 , n44213 , n44216 , n44217 );
xor ( n44219 , n43663 , n43665 );
xor ( n44220 , n44219 , n43667 );
and ( n44221 , n44218 , n44220 );
xor ( n44222 , n43708 , n43710 );
xor ( n44223 , n44222 , n43713 );
and ( n44224 , n44220 , n44223 );
and ( n44225 , n44218 , n44223 );
or ( n44226 , n44221 , n44224 , n44225 );
xor ( n44227 , n43751 , n43753 );
and ( n44228 , n43278 , n43282 );
and ( n44229 , n43282 , n43287 );
and ( n44230 , n43278 , n43287 );
or ( n44231 , n44228 , n44229 , n44230 );
xor ( n44232 , n43696 , n43700 );
xor ( n44233 , n44232 , n43705 );
and ( n44234 , n44231 , n44233 );
xor ( n44235 , n44001 , n44005 );
xor ( n44236 , n44235 , n44008 );
and ( n44237 , n44233 , n44236 );
and ( n44238 , n44231 , n44236 );
or ( n44239 , n44234 , n44237 , n44238 );
and ( n44240 , n44227 , n44239 );
xor ( n44241 , n43723 , n43727 );
xor ( n44242 , n44241 , n43748 );
xor ( n44243 , n43875 , n43987 );
xor ( n44244 , n44243 , n43990 );
xor ( n44245 , n44079 , n44081 );
xor ( n44246 , n44245 , n44084 );
and ( n44247 , n44244 , n44246 );
xor ( n44248 , n44069 , n44073 );
xor ( n44249 , n44248 , n44076 );
xor ( n44250 , n44059 , n44063 );
xor ( n44251 , n44250 , n44066 );
xor ( n44252 , n43942 , n43946 );
xor ( n44253 , n44252 , n43951 );
xor ( n44254 , n43958 , n43962 );
xor ( n44255 , n44254 , n43967 );
and ( n44256 , n44253 , n44255 );
and ( n44257 , n42456 , n39678 );
and ( n44258 , n42048 , n39676 );
nor ( n44259 , n44257 , n44258 );
xnor ( n44260 , n44259 , n39643 );
xor ( n44261 , n38954 , n39302 );
buf ( n571565 , n44261 );
buf ( n571566 , n571565 );
buf ( n44264 , n571566 );
and ( n44265 , n44264 , n39367 );
and ( n44266 , n44260 , n44265 );
xor ( n44267 , n44152 , n44156 );
and ( n44268 , n44265 , n44267 );
and ( n44269 , n44260 , n44267 );
or ( n44270 , n44266 , n44268 , n44269 );
and ( n44271 , n44255 , n44270 );
and ( n44272 , n44253 , n44270 );
or ( n44273 , n44256 , n44271 , n44272 );
xor ( n44274 , n44117 , n44119 );
xor ( n44275 , n44274 , n44122 );
xor ( n44276 , n44126 , n44127 );
xor ( n44277 , n44276 , n44144 );
and ( n44278 , n44275 , n44277 );
xor ( n44279 , n44157 , n44173 );
xor ( n44280 , n44279 , n44176 );
and ( n44281 , n44277 , n44280 );
and ( n44282 , n44275 , n44280 );
or ( n44283 , n44278 , n44281 , n44282 );
and ( n44284 , n44273 , n44283 );
xor ( n44285 , n44104 , n44106 );
xor ( n44286 , n44285 , n44109 );
and ( n44287 , n44283 , n44286 );
and ( n44288 , n44273 , n44286 );
or ( n44289 , n44284 , n44287 , n44288 );
and ( n44290 , n44251 , n44289 );
xor ( n44291 , n44102 , n44112 );
xor ( n44292 , n44291 , n44182 );
and ( n44293 , n44289 , n44292 );
and ( n44294 , n44251 , n44292 );
or ( n44295 , n44290 , n44293 , n44294 );
and ( n44296 , n44249 , n44295 );
xor ( n44297 , n44091 , n44093 );
xor ( n44298 , n44297 , n44096 );
and ( n44299 , n44295 , n44298 );
and ( n44300 , n44249 , n44298 );
or ( n44301 , n44296 , n44299 , n44300 );
and ( n44302 , n44246 , n44301 );
and ( n44303 , n44244 , n44301 );
or ( n44304 , n44247 , n44302 , n44303 );
and ( n44305 , n44242 , n44304 );
xor ( n44306 , n44087 , n44212 );
xor ( n44307 , n44306 , n44215 );
and ( n44308 , n44304 , n44307 );
and ( n44309 , n44242 , n44307 );
or ( n44310 , n44305 , n44308 , n44309 );
and ( n44311 , n44239 , n44310 );
and ( n44312 , n44227 , n44310 );
or ( n44313 , n44240 , n44311 , n44312 );
and ( n44314 , n44226 , n44313 );
xor ( n44315 , n43670 , n43671 );
xor ( n44316 , n44315 , n43716 );
and ( n44317 , n44313 , n44316 );
and ( n44318 , n44226 , n44316 );
or ( n44319 , n44314 , n44317 , n44318 );
xor ( n44320 , n43719 , n44020 );
xor ( n44321 , n44320 , n44023 );
and ( n44322 , n44319 , n44321 );
xor ( n44323 , n43754 , n44014 );
xor ( n44324 , n44323 , n44017 );
xor ( n44325 , n43758 , n43996 );
xor ( n44326 , n44325 , n44011 );
xor ( n44327 , n44231 , n44233 );
xor ( n44328 , n44327 , n44236 );
xor ( n44329 , n44089 , n44099 );
xor ( n44330 , n44329 , n44209 );
xor ( n44331 , n44185 , n44203 );
xor ( n44332 , n44331 , n44206 );
xor ( n44333 , n44195 , n44197 );
xor ( n44334 , n44333 , n44200 );
xor ( n44335 , n44125 , n44147 );
xor ( n44336 , n44335 , n44179 );
xor ( n44337 , n44187 , n44189 );
xor ( n44338 , n44337 , n44192 );
and ( n44339 , n44336 , n44338 );
and ( n44340 , n44264 , n39375 );
and ( n44341 , n43437 , n39373 );
nor ( n44342 , n44340 , n44341 );
xnor ( n44343 , n44342 , n39380 );
xor ( n44344 , n38956 , n39301 );
buf ( n571648 , n44344 );
buf ( n571649 , n571648 );
buf ( n44347 , n571649 );
and ( n44348 , n44347 , n39367 );
xor ( n44349 , n44343 , n44348 );
and ( n44350 , n44347 , n39375 );
and ( n44351 , n44264 , n39373 );
nor ( n44352 , n44350 , n44351 );
xnor ( n44353 , n44352 , n39380 );
xor ( n44354 , n38959 , n39299 );
buf ( n571658 , n44354 );
buf ( n571659 , n571658 );
buf ( n44357 , n571659 );
and ( n44358 , n44357 , n39367 );
and ( n44359 , n44353 , n44358 );
and ( n44360 , n44349 , n44359 );
and ( n44361 , n43428 , n39396 );
and ( n44362 , n43200 , n39394 );
nor ( n44363 , n44361 , n44362 );
xnor ( n44364 , n44363 , n39401 );
and ( n44365 , n44359 , n44364 );
and ( n44366 , n44349 , n44364 );
or ( n44367 , n44360 , n44365 , n44366 );
buf ( n44368 , n557778 );
not ( n44369 , n44368 );
and ( n44370 , n44367 , n44369 );
and ( n44371 , n44343 , n44348 );
xor ( n44372 , n44161 , n44165 );
xor ( n44373 , n44372 , n44170 );
and ( n44374 , n44371 , n44373 );
xor ( n44375 , n44260 , n44265 );
xor ( n44376 , n44375 , n44267 );
and ( n44377 , n44373 , n44376 );
and ( n44378 , n44371 , n44376 );
or ( n44379 , n44374 , n44377 , n44378 );
and ( n44380 , n44370 , n44379 );
xor ( n44381 , n44253 , n44255 );
xor ( n44382 , n44381 , n44270 );
and ( n44383 , n44379 , n44382 );
and ( n44384 , n44370 , n44382 );
or ( n44385 , n44380 , n44383 , n44384 );
and ( n44386 , n44338 , n44385 );
and ( n44387 , n44336 , n44385 );
or ( n44388 , n44339 , n44386 , n44387 );
and ( n44389 , n44334 , n44388 );
xor ( n44390 , n44251 , n44289 );
xor ( n44391 , n44390 , n44292 );
and ( n44392 , n44388 , n44391 );
and ( n44393 , n44334 , n44391 );
or ( n44394 , n44389 , n44392 , n44393 );
and ( n44395 , n44332 , n44394 );
xor ( n44396 , n44249 , n44295 );
xor ( n44397 , n44396 , n44298 );
and ( n44398 , n44394 , n44397 );
and ( n44399 , n44332 , n44397 );
or ( n44400 , n44395 , n44398 , n44399 );
and ( n44401 , n44330 , n44400 );
xor ( n44402 , n44244 , n44246 );
xor ( n44403 , n44402 , n44301 );
and ( n44404 , n44400 , n44403 );
and ( n44405 , n44330 , n44403 );
or ( n44406 , n44401 , n44404 , n44405 );
and ( n44407 , n44328 , n44406 );
xor ( n44408 , n44242 , n44304 );
xor ( n44409 , n44408 , n44307 );
and ( n44410 , n44406 , n44409 );
and ( n44411 , n44328 , n44409 );
or ( n44412 , n44407 , n44410 , n44411 );
and ( n44413 , n44326 , n44412 );
xor ( n44414 , n44218 , n44220 );
xor ( n44415 , n44414 , n44223 );
and ( n44416 , n44412 , n44415 );
and ( n44417 , n44326 , n44415 );
or ( n44418 , n44413 , n44416 , n44417 );
and ( n44419 , n44324 , n44418 );
xor ( n44420 , n44226 , n44313 );
xor ( n44421 , n44420 , n44316 );
and ( n44422 , n44418 , n44421 );
and ( n44423 , n44324 , n44421 );
or ( n44424 , n44419 , n44422 , n44423 );
and ( n44425 , n44321 , n44424 );
and ( n44426 , n44319 , n44424 );
or ( n44427 , n44322 , n44425 , n44426 );
and ( n44428 , n44055 , n44427 );
xor ( n44429 , n44055 , n44427 );
xor ( n44430 , n44319 , n44321 );
xor ( n44431 , n44430 , n44424 );
xor ( n44432 , n44324 , n44418 );
xor ( n44433 , n44432 , n44421 );
xor ( n44434 , n44227 , n44239 );
xor ( n44435 , n44434 , n44310 );
xor ( n44436 , n44326 , n44412 );
xor ( n44437 , n44436 , n44415 );
and ( n44438 , n44435 , n44437 );
xor ( n44439 , n44435 , n44437 );
xor ( n44440 , n44328 , n44406 );
xor ( n44441 , n44440 , n44409 );
xor ( n44442 , n44330 , n44400 );
xor ( n44443 , n44442 , n44403 );
xor ( n44444 , n44332 , n44394 );
xor ( n44445 , n44444 , n44397 );
xor ( n44446 , n44273 , n44283 );
xor ( n44447 , n44446 , n44286 );
xor ( n44448 , n44275 , n44277 );
xor ( n44449 , n44448 , n44280 );
xor ( n44450 , n44353 , n44358 );
and ( n44451 , n44357 , n39375 );
and ( n44452 , n44347 , n39373 );
nor ( n44453 , n44451 , n44452 );
xnor ( n44454 , n44453 , n39380 );
xor ( n44455 , n38960 , n39298 );
buf ( n571759 , n44455 );
buf ( n571760 , n571759 );
buf ( n44458 , n571760 );
and ( n44459 , n44458 , n39367 );
and ( n44460 , n44454 , n44459 );
and ( n44461 , n44450 , n44460 );
and ( n44462 , n43200 , n39480 );
and ( n44463 , n43192 , n39478 );
nor ( n44464 , n44462 , n44463 );
xnor ( n44465 , n44464 , n39462 );
and ( n44466 , n44460 , n44465 );
and ( n44467 , n44450 , n44465 );
or ( n44468 , n44461 , n44466 , n44467 );
and ( n44469 , n43192 , n39480 );
and ( n44470 , n43073 , n39478 );
nor ( n44471 , n44469 , n44470 );
xnor ( n44472 , n44471 , n39462 );
and ( n44473 , n44468 , n44472 );
xor ( n44474 , n44349 , n44359 );
xor ( n44475 , n44474 , n44364 );
and ( n44476 , n44472 , n44475 );
and ( n44477 , n44468 , n44475 );
or ( n44478 , n44473 , n44476 , n44477 );
and ( n44479 , n43019 , n39539 );
and ( n44480 , n42811 , n39537 );
nor ( n44481 , n44479 , n44480 );
xnor ( n44482 , n44481 , n39522 );
and ( n44483 , n44478 , n44482 );
and ( n44484 , n43073 , n39480 );
and ( n44485 , n43027 , n39478 );
nor ( n44486 , n44484 , n44485 );
xnor ( n44487 , n44486 , n39462 );
and ( n44488 , n44482 , n44487 );
and ( n44489 , n44478 , n44487 );
or ( n44490 , n44483 , n44488 , n44489 );
and ( n44491 , n44449 , n44490 );
xor ( n44492 , n44370 , n44379 );
xor ( n44493 , n44492 , n44382 );
and ( n44494 , n44490 , n44493 );
and ( n44495 , n44449 , n44493 );
or ( n44496 , n44491 , n44494 , n44495 );
and ( n44497 , n44447 , n44496 );
xor ( n44498 , n44336 , n44338 );
xor ( n44499 , n44498 , n44385 );
and ( n44500 , n44496 , n44499 );
and ( n44501 , n44447 , n44499 );
or ( n44502 , n44497 , n44500 , n44501 );
xor ( n44503 , n44334 , n44388 );
xor ( n44504 , n44503 , n44391 );
and ( n44505 , n44502 , n44504 );
xor ( n44506 , n44447 , n44496 );
xor ( n44507 , n44506 , n44499 );
xor ( n44508 , n44367 , n44369 );
xor ( n44509 , n44371 , n44373 );
xor ( n44510 , n44509 , n44376 );
and ( n44511 , n44508 , n44510 );
xor ( n44512 , n44454 , n44459 );
and ( n44513 , n44458 , n39375 );
and ( n44514 , n44357 , n39373 );
nor ( n44515 , n44513 , n44514 );
xnor ( n44516 , n44515 , n39380 );
xor ( n44517 , n38962 , n39297 );
buf ( n571821 , n44517 );
buf ( n571822 , n571821 );
buf ( n44520 , n571822 );
and ( n44521 , n44520 , n39367 );
and ( n44522 , n44516 , n44521 );
and ( n44523 , n44512 , n44522 );
and ( n44524 , n44264 , n39396 );
and ( n44525 , n43437 , n39394 );
nor ( n44526 , n44524 , n44525 );
xnor ( n44527 , n44526 , n39401 );
and ( n44528 , n44522 , n44527 );
and ( n44529 , n44512 , n44527 );
or ( n44530 , n44523 , n44528 , n44529 );
and ( n44531 , n43437 , n39396 );
and ( n44532 , n43428 , n39394 );
nor ( n44533 , n44531 , n44532 );
xnor ( n44534 , n44533 , n39401 );
and ( n44535 , n44530 , n44534 );
xor ( n44536 , n44450 , n44460 );
xor ( n44537 , n44536 , n44465 );
and ( n44538 , n44534 , n44537 );
and ( n44539 , n44530 , n44537 );
or ( n44540 , n44535 , n44538 , n44539 );
and ( n44541 , n43027 , n39539 );
and ( n44542 , n43019 , n39537 );
nor ( n44543 , n44541 , n44542 );
xnor ( n44544 , n44543 , n39522 );
and ( n44545 , n44540 , n44544 );
buf ( n44546 , n557779 );
not ( n44547 , n44546 );
and ( n44548 , n44544 , n44547 );
and ( n44549 , n44540 , n44547 );
or ( n44550 , n44545 , n44548 , n44549 );
and ( n44551 , n44510 , n44550 );
and ( n44552 , n44508 , n44550 );
or ( n44553 , n44511 , n44551 , n44552 );
xor ( n44554 , n44449 , n44490 );
xor ( n44555 , n44554 , n44493 );
and ( n44556 , n44553 , n44555 );
xor ( n44557 , n44516 , n44521 );
and ( n44558 , n44520 , n39375 );
and ( n44559 , n44458 , n39373 );
nor ( n44560 , n44558 , n44559 );
xnor ( n44561 , n44560 , n39380 );
xor ( n44562 , n38964 , n39296 );
buf ( n571866 , n44562 );
buf ( n571867 , n571866 );
buf ( n44565 , n571867 );
and ( n44566 , n44565 , n39367 );
and ( n44567 , n44561 , n44566 );
and ( n44568 , n44557 , n44567 );
and ( n44569 , n44347 , n39396 );
and ( n44570 , n44264 , n39394 );
nor ( n44571 , n44569 , n44570 );
xnor ( n44572 , n44571 , n39401 );
and ( n44573 , n44567 , n44572 );
and ( n44574 , n44557 , n44572 );
or ( n44575 , n44568 , n44573 , n44574 );
and ( n44576 , n43428 , n39480 );
and ( n44577 , n43200 , n39478 );
nor ( n44578 , n44576 , n44577 );
xnor ( n44579 , n44578 , n39462 );
and ( n44580 , n44575 , n44579 );
xor ( n44581 , n44512 , n44522 );
xor ( n44582 , n44581 , n44527 );
and ( n44583 , n44579 , n44582 );
and ( n44584 , n44575 , n44582 );
or ( n44585 , n44580 , n44583 , n44584 );
and ( n44586 , n43073 , n39539 );
and ( n44587 , n43027 , n39537 );
nor ( n44588 , n44586 , n44587 );
xnor ( n44589 , n44588 , n39522 );
and ( n44590 , n44585 , n44589 );
buf ( n44591 , n557780 );
not ( n44592 , n44591 );
and ( n44593 , n44589 , n44592 );
and ( n44594 , n44585 , n44592 );
or ( n44595 , n44590 , n44593 , n44594 );
and ( n44596 , n42811 , n39678 );
and ( n44597 , n42456 , n39676 );
nor ( n44598 , n44596 , n44597 );
xnor ( n44599 , n44598 , n39643 );
and ( n44600 , n44595 , n44599 );
xor ( n44601 , n44468 , n44472 );
xor ( n44602 , n44601 , n44475 );
and ( n44603 , n44599 , n44602 );
and ( n44604 , n44595 , n44602 );
or ( n44605 , n44600 , n44603 , n44604 );
and ( n44606 , n41807 , n39896 );
and ( n44607 , n41692 , n39894 );
nor ( n44608 , n44606 , n44607 );
xnor ( n44609 , n44608 , n39857 );
and ( n44610 , n44605 , n44609 );
xor ( n44611 , n44478 , n44482 );
xor ( n44612 , n44611 , n44487 );
and ( n44613 , n44609 , n44612 );
and ( n44614 , n44605 , n44612 );
or ( n44615 , n44610 , n44613 , n44614 );
and ( n44616 , n44555 , n44615 );
and ( n44617 , n44553 , n44615 );
or ( n44618 , n44556 , n44616 , n44617 );
and ( n44619 , n44507 , n44618 );
and ( n44620 , n41182 , n40258 );
and ( n44621 , n41032 , n40256 );
nor ( n44622 , n44620 , n44621 );
xnor ( n44623 , n44622 , n40169 );
and ( n44624 , n41692 , n40053 );
and ( n44625 , n41615 , n40051 );
nor ( n44626 , n44624 , n44625 );
xnor ( n44627 , n44626 , n39999 );
and ( n44628 , n44623 , n44627 );
and ( n44629 , n42048 , n39760 );
and ( n44630 , n42061 , n39758 );
nor ( n44631 , n44629 , n44630 );
xnor ( n44632 , n44631 , n39742 );
and ( n44633 , n44627 , n44632 );
and ( n44634 , n44623 , n44632 );
or ( n44635 , n44628 , n44633 , n44634 );
and ( n44636 , n40492 , n40746 );
and ( n44637 , n40507 , n40744 );
nor ( n44638 , n44636 , n44637 );
xnor ( n44639 , n44638 , n40501 );
and ( n44640 , n44635 , n44639 );
xor ( n44641 , n44605 , n44609 );
xor ( n44642 , n44641 , n44612 );
and ( n44643 , n44639 , n44642 );
and ( n44644 , n44635 , n44642 );
or ( n44645 , n44640 , n44643 , n44644 );
xor ( n44646 , n44553 , n44555 );
xor ( n44647 , n44646 , n44615 );
and ( n44648 , n44645 , n44647 );
and ( n44649 , n44520 , n39396 );
and ( n44650 , n44458 , n39394 );
nor ( n44651 , n44649 , n44650 );
xnor ( n44652 , n44651 , n39401 );
xor ( n44653 , n38966 , n39295 );
buf ( n571957 , n44653 );
buf ( n571958 , n571957 );
buf ( n44656 , n571958 );
and ( n44657 , n44656 , n39375 );
and ( n44658 , n44565 , n39373 );
nor ( n44659 , n44657 , n44658 );
xnor ( n44660 , n44659 , n39380 );
and ( n44661 , n44652 , n44660 );
xor ( n44662 , n38968 , n39294 );
buf ( n571966 , n44662 );
buf ( n571967 , n571966 );
buf ( n44665 , n571967 );
and ( n44666 , n44665 , n39367 );
and ( n44667 , n44660 , n44666 );
and ( n44668 , n44652 , n44666 );
or ( n44669 , n44661 , n44667 , n44668 );
and ( n44670 , n44347 , n39480 );
and ( n44671 , n44264 , n39478 );
nor ( n44672 , n44670 , n44671 );
xnor ( n44673 , n44672 , n39462 );
and ( n44674 , n44669 , n44673 );
and ( n44675 , n44458 , n39396 );
and ( n44676 , n44357 , n39394 );
nor ( n44677 , n44675 , n44676 );
xnor ( n44678 , n44677 , n39401 );
and ( n44679 , n44565 , n39375 );
and ( n44680 , n44520 , n39373 );
nor ( n44681 , n44679 , n44680 );
xnor ( n44682 , n44681 , n39380 );
xor ( n44683 , n44678 , n44682 );
and ( n44684 , n44656 , n39367 );
xor ( n44685 , n44683 , n44684 );
and ( n44686 , n44673 , n44685 );
and ( n44687 , n44669 , n44685 );
or ( n44688 , n44674 , n44686 , n44687 );
and ( n44689 , n43192 , n39678 );
and ( n44690 , n43073 , n39676 );
nor ( n44691 , n44689 , n44690 );
xnor ( n44692 , n44691 , n39643 );
and ( n44693 , n44688 , n44692 );
and ( n44694 , n43428 , n39539 );
and ( n44695 , n43200 , n39537 );
nor ( n44696 , n44694 , n44695 );
xnor ( n44697 , n44696 , n39522 );
and ( n44698 , n44692 , n44697 );
and ( n44699 , n44688 , n44697 );
or ( n44700 , n44693 , n44698 , n44699 );
and ( n44701 , n43073 , n39678 );
and ( n44702 , n43027 , n39676 );
nor ( n44703 , n44701 , n44702 );
xnor ( n44704 , n44703 , n39643 );
and ( n44705 , n44700 , n44704 );
buf ( n44706 , n557782 );
not ( n44707 , n44706 );
and ( n44708 , n44704 , n44707 );
and ( n44709 , n44700 , n44707 );
or ( n44710 , n44705 , n44708 , n44709 );
and ( n44711 , n42811 , n39760 );
and ( n44712 , n42456 , n39758 );
nor ( n44713 , n44711 , n44712 );
xnor ( n44714 , n44713 , n39742 );
and ( n44715 , n44710 , n44714 );
and ( n44716 , n44357 , n39396 );
and ( n44717 , n44347 , n39394 );
nor ( n44718 , n44716 , n44717 );
xnor ( n44719 , n44718 , n39401 );
xor ( n44720 , n44561 , n44566 );
and ( n44721 , n44719 , n44720 );
and ( n44722 , n43200 , n39539 );
and ( n44723 , n43192 , n39537 );
nor ( n44724 , n44722 , n44723 );
xnor ( n44725 , n44724 , n39522 );
and ( n44726 , n44721 , n44725 );
xor ( n44727 , n44557 , n44567 );
xor ( n44728 , n44727 , n44572 );
and ( n44729 , n44725 , n44728 );
and ( n44730 , n44721 , n44728 );
or ( n44731 , n44726 , n44729 , n44730 );
and ( n44732 , n43192 , n39539 );
and ( n44733 , n43073 , n39537 );
nor ( n44734 , n44732 , n44733 );
xnor ( n44735 , n44734 , n39522 );
xor ( n44736 , n44731 , n44735 );
buf ( n44737 , n557781 );
not ( n44738 , n44737 );
xor ( n44739 , n44736 , n44738 );
and ( n44740 , n44714 , n44739 );
and ( n44741 , n44710 , n44739 );
or ( n44742 , n44715 , n44740 , n44741 );
and ( n44743 , n41807 , n40053 );
and ( n44744 , n41692 , n40051 );
nor ( n44745 , n44743 , n44744 );
xnor ( n44746 , n44745 , n39999 );
and ( n44747 , n44742 , n44746 );
and ( n44748 , n42061 , n39896 );
and ( n44749 , n41816 , n39894 );
nor ( n44750 , n44748 , n44749 );
xnor ( n44751 , n44750 , n39857 );
and ( n44752 , n44746 , n44751 );
and ( n44753 , n44742 , n44751 );
or ( n44754 , n44747 , n44752 , n44753 );
xor ( n44755 , n44719 , n44720 );
and ( n44756 , n44678 , n44682 );
and ( n44757 , n44682 , n44684 );
and ( n44758 , n44678 , n44684 );
or ( n44759 , n44756 , n44757 , n44758 );
and ( n44760 , n44755 , n44759 );
and ( n44761 , n44264 , n39480 );
and ( n44762 , n43437 , n39478 );
nor ( n44763 , n44761 , n44762 );
xnor ( n44764 , n44763 , n39462 );
and ( n44765 , n44759 , n44764 );
and ( n44766 , n44755 , n44764 );
or ( n44767 , n44760 , n44765 , n44766 );
and ( n44768 , n43437 , n39480 );
and ( n44769 , n43428 , n39478 );
nor ( n44770 , n44768 , n44769 );
xnor ( n44771 , n44770 , n39462 );
and ( n44772 , n44767 , n44771 );
xor ( n44773 , n44721 , n44725 );
xor ( n44774 , n44773 , n44728 );
and ( n44775 , n44771 , n44774 );
and ( n44776 , n44767 , n44774 );
or ( n44777 , n44772 , n44775 , n44776 );
and ( n44778 , n43027 , n39678 );
and ( n44779 , n43019 , n39676 );
nor ( n44780 , n44778 , n44779 );
xnor ( n44781 , n44780 , n39643 );
and ( n44782 , n44777 , n44781 );
xor ( n44783 , n44575 , n44579 );
xor ( n44784 , n44783 , n44582 );
and ( n44785 , n44781 , n44784 );
and ( n44786 , n44777 , n44784 );
or ( n44787 , n44782 , n44785 , n44786 );
and ( n44788 , n42456 , n39760 );
and ( n44789 , n42048 , n39758 );
nor ( n44790 , n44788 , n44789 );
xnor ( n44791 , n44790 , n39742 );
and ( n44792 , n44787 , n44791 );
xor ( n44793 , n44585 , n44589 );
xor ( n44794 , n44793 , n44592 );
and ( n44795 , n44791 , n44794 );
and ( n44796 , n44787 , n44794 );
or ( n44797 , n44792 , n44795 , n44796 );
and ( n44798 , n44754 , n44797 );
xor ( n44799 , n44595 , n44599 );
xor ( n44800 , n44799 , n44602 );
and ( n44801 , n44797 , n44800 );
and ( n44802 , n44754 , n44800 );
or ( n44803 , n44798 , n44801 , n44802 );
xor ( n44804 , n44132 , n44136 );
xor ( n44805 , n44804 , n44141 );
and ( n44806 , n44803 , n44805 );
and ( n44807 , n44647 , n44806 );
and ( n44808 , n44645 , n44806 );
or ( n44809 , n44648 , n44807 , n44808 );
and ( n44810 , n44618 , n44809 );
and ( n44811 , n44507 , n44809 );
or ( n44812 , n44619 , n44810 , n44811 );
and ( n44813 , n44504 , n44812 );
and ( n44814 , n44502 , n44812 );
or ( n44815 , n44505 , n44813 , n44814 );
and ( n44816 , n44445 , n44815 );
xor ( n44817 , n44502 , n44504 );
xor ( n44818 , n44817 , n44812 );
and ( n44819 , n41032 , n40527 );
and ( n44820 , n41047 , n40525 );
nor ( n44821 , n44819 , n44820 );
xnor ( n44822 , n44821 , n40382 );
and ( n44823 , n41615 , n40258 );
and ( n44824 , n41182 , n40256 );
nor ( n44825 , n44823 , n44824 );
xnor ( n44826 , n44825 , n40169 );
and ( n44827 , n44822 , n44826 );
and ( n44828 , n44731 , n44735 );
and ( n44829 , n44735 , n44738 );
and ( n44830 , n44731 , n44738 );
or ( n44831 , n44828 , n44829 , n44830 );
and ( n44832 , n43019 , n39678 );
and ( n44833 , n42811 , n39676 );
nor ( n44834 , n44832 , n44833 );
xnor ( n44835 , n44834 , n39643 );
xor ( n44836 , n44831 , n44835 );
xor ( n44837 , n44530 , n44534 );
xor ( n44838 , n44837 , n44537 );
xor ( n44839 , n44836 , n44838 );
and ( n44840 , n44826 , n44839 );
and ( n44841 , n44822 , n44839 );
or ( n44842 , n44827 , n44840 , n44841 );
xor ( n44843 , n44623 , n44627 );
xor ( n44844 , n44843 , n44632 );
and ( n44845 , n44842 , n44844 );
xor ( n44846 , n44754 , n44797 );
xor ( n44847 , n44846 , n44800 );
and ( n44848 , n44844 , n44847 );
and ( n44849 , n44842 , n44847 );
or ( n44850 , n44845 , n44848 , n44849 );
and ( n44851 , n39948 , n41984 );
and ( n44852 , n39867 , n41982 );
nor ( n44853 , n44851 , n44852 );
xnor ( n44854 , n44853 , n41687 );
and ( n44855 , n44850 , n44854 );
and ( n44856 , n40148 , n41622 );
and ( n44857 , n40009 , n41620 );
nor ( n44858 , n44856 , n44857 );
xnor ( n44859 , n44858 , n41194 );
and ( n44860 , n44854 , n44859 );
and ( n44861 , n44850 , n44859 );
or ( n44862 , n44855 , n44860 , n44861 );
and ( n44863 , n40738 , n40746 );
and ( n44864 , n40492 , n40744 );
nor ( n44865 , n44863 , n44864 );
xnor ( n44866 , n44865 , n40501 );
and ( n44867 , n41047 , n40527 );
and ( n44868 , n40869 , n40525 );
nor ( n44869 , n44867 , n44868 );
xnor ( n44870 , n44869 , n40382 );
and ( n44871 , n44866 , n44870 );
and ( n44872 , n44831 , n44835 );
and ( n44873 , n44835 , n44838 );
and ( n44874 , n44831 , n44838 );
or ( n44875 , n44872 , n44873 , n44874 );
and ( n44876 , n41816 , n39896 );
and ( n44877 , n41807 , n39894 );
nor ( n44878 , n44876 , n44877 );
xnor ( n44879 , n44878 , n39857 );
xor ( n44880 , n44875 , n44879 );
xor ( n44881 , n44540 , n44544 );
xor ( n44882 , n44881 , n44547 );
xor ( n44883 , n44880 , n44882 );
and ( n44884 , n44870 , n44883 );
and ( n44885 , n44866 , n44883 );
or ( n44886 , n44871 , n44884 , n44885 );
and ( n44887 , n40373 , n41055 );
and ( n44888 , n40388 , n41053 );
nor ( n44889 , n44887 , n44888 );
xnor ( n44890 , n44889 , n40728 );
and ( n44891 , n44886 , n44890 );
xor ( n44892 , n44635 , n44639 );
xor ( n44893 , n44892 , n44642 );
and ( n44894 , n44890 , n44893 );
and ( n44895 , n44886 , n44893 );
or ( n44896 , n44891 , n44894 , n44895 );
and ( n44897 , n44862 , n44896 );
xor ( n44898 , n44507 , n44618 );
xor ( n44899 , n44898 , n44809 );
and ( n44900 , n44897 , n44899 );
xor ( n44901 , n44508 , n44510 );
xor ( n44902 , n44901 , n44550 );
and ( n44903 , n44875 , n44879 );
and ( n44904 , n44879 , n44882 );
and ( n44905 , n44875 , n44882 );
or ( n44906 , n44903 , n44904 , n44905 );
and ( n44907 , n44902 , n44906 );
xor ( n44908 , n44803 , n44805 );
and ( n44909 , n44906 , n44908 );
and ( n44910 , n44902 , n44908 );
or ( n44911 , n44907 , n44909 , n44910 );
xor ( n44912 , n44645 , n44647 );
xor ( n44913 , n44912 , n44806 );
and ( n44914 , n44911 , n44913 );
xor ( n44915 , n44862 , n44896 );
and ( n44916 , n44913 , n44915 );
and ( n44917 , n44911 , n44915 );
or ( n44918 , n44914 , n44916 , n44917 );
and ( n44919 , n44899 , n44918 );
and ( n44920 , n44897 , n44918 );
or ( n44921 , n44900 , n44919 , n44920 );
and ( n44922 , n44818 , n44921 );
xor ( n44923 , n44897 , n44899 );
xor ( n44924 , n44923 , n44918 );
and ( n44925 , n41816 , n40053 );
and ( n44926 , n41807 , n40051 );
nor ( n44927 , n44925 , n44926 );
xnor ( n44928 , n44927 , n39999 );
and ( n44929 , n42048 , n39896 );
and ( n44930 , n42061 , n39894 );
nor ( n44931 , n44929 , n44930 );
xnor ( n44932 , n44931 , n39857 );
and ( n44933 , n44928 , n44932 );
xor ( n44934 , n44777 , n44781 );
xor ( n44935 , n44934 , n44784 );
and ( n44936 , n44932 , n44935 );
and ( n44937 , n44928 , n44935 );
or ( n44938 , n44933 , n44936 , n44937 );
and ( n44939 , n40869 , n40746 );
and ( n44940 , n40738 , n40744 );
nor ( n44941 , n44939 , n44940 );
xnor ( n44942 , n44941 , n40501 );
and ( n44943 , n44938 , n44942 );
xor ( n44944 , n44787 , n44791 );
xor ( n44945 , n44944 , n44794 );
and ( n44946 , n44942 , n44945 );
and ( n44947 , n44938 , n44945 );
or ( n44948 , n44943 , n44946 , n44947 );
and ( n44949 , n40388 , n41292 );
and ( n44950 , n40186 , n41290 );
nor ( n44951 , n44949 , n44950 );
xnor ( n44952 , n44951 , n41041 );
and ( n44953 , n44948 , n44952 );
and ( n44954 , n40507 , n41055 );
and ( n44955 , n40373 , n41053 );
nor ( n44956 , n44954 , n44955 );
xnor ( n44957 , n44956 , n40728 );
and ( n44958 , n44952 , n44957 );
and ( n44959 , n44948 , n44957 );
or ( n44960 , n44953 , n44958 , n44959 );
and ( n44961 , n39867 , n42269 );
and ( n44962 , n39795 , n42266 );
nor ( n44963 , n44961 , n44962 );
xnor ( n44964 , n44963 , n41684 );
and ( n44965 , n40197 , n41622 );
and ( n44966 , n40148 , n41620 );
nor ( n44967 , n44965 , n44966 );
xnor ( n44968 , n44967 , n41194 );
and ( n44969 , n44964 , n44968 );
xor ( n44970 , n44842 , n44844 );
xor ( n44971 , n44970 , n44847 );
and ( n44972 , n44968 , n44971 );
and ( n44973 , n44964 , n44971 );
or ( n44974 , n44969 , n44972 , n44973 );
and ( n44975 , n44960 , n44974 );
xor ( n44976 , n44886 , n44890 );
xor ( n44977 , n44976 , n44893 );
and ( n44978 , n44974 , n44977 );
and ( n44979 , n44960 , n44977 );
or ( n44980 , n44975 , n44978 , n44979 );
xor ( n44981 , n44911 , n44913 );
xor ( n44982 , n44981 , n44915 );
and ( n44983 , n44980 , n44982 );
and ( n44984 , n41615 , n40527 );
and ( n44985 , n41182 , n40525 );
nor ( n44986 , n44984 , n44985 );
xnor ( n44987 , n44986 , n40382 );
xor ( n44988 , n39268 , n39270 );
buf ( n572292 , n44988 );
buf ( n572293 , n572292 );
buf ( n44991 , n572293 );
and ( n44992 , n44991 , n39373 );
not ( n44993 , n44992 );
and ( n44994 , n44993 , n39380 );
and ( n44995 , n44991 , n39375 );
xor ( n44996 , n39267 , n39271 );
buf ( n572300 , n44996 );
buf ( n572301 , n572300 );
buf ( n44999 , n572301 );
and ( n45000 , n44999 , n39373 );
nor ( n45001 , n44995 , n45000 );
xnor ( n45002 , n45001 , n39380 );
and ( n45003 , n44994 , n45002 );
and ( n45004 , n44999 , n39375 );
xor ( n45005 , n39262 , n39273 );
buf ( n572309 , n45005 );
buf ( n572310 , n572309 );
buf ( n45008 , n572310 );
and ( n45009 , n45008 , n39373 );
nor ( n45010 , n45004 , n45009 );
xnor ( n45011 , n45010 , n39380 );
and ( n45012 , n45003 , n45011 );
and ( n45013 , n44991 , n39367 );
and ( n45014 , n45011 , n45013 );
and ( n45015 , n45003 , n45013 );
or ( n45016 , n45012 , n45014 , n45015 );
and ( n45017 , n45008 , n39375 );
xor ( n45018 , n39261 , n39274 );
buf ( n572322 , n45018 );
buf ( n572323 , n572322 );
buf ( n45021 , n572323 );
and ( n45022 , n45021 , n39373 );
nor ( n45023 , n45017 , n45022 );
xnor ( n45024 , n45023 , n39380 );
and ( n45025 , n45016 , n45024 );
and ( n45026 , n44999 , n39367 );
and ( n45027 , n45024 , n45026 );
and ( n45028 , n45016 , n45026 );
or ( n45029 , n45025 , n45027 , n45028 );
and ( n45030 , n45021 , n39375 );
xor ( n45031 , n39256 , n39276 );
buf ( n572335 , n45031 );
buf ( n572336 , n572335 );
buf ( n45034 , n572336 );
and ( n45035 , n45034 , n39373 );
nor ( n45036 , n45030 , n45035 );
xnor ( n45037 , n45036 , n39380 );
and ( n45038 , n45029 , n45037 );
and ( n45039 , n45008 , n39367 );
and ( n45040 , n45037 , n45039 );
and ( n45041 , n45029 , n45039 );
or ( n45042 , n45038 , n45040 , n45041 );
and ( n45043 , n45034 , n39375 );
xor ( n45044 , n39243 , n39278 );
buf ( n572348 , n45044 );
buf ( n572349 , n572348 );
buf ( n45047 , n572349 );
and ( n45048 , n45047 , n39373 );
nor ( n45049 , n45043 , n45048 );
xnor ( n45050 , n45049 , n39380 );
and ( n45051 , n45042 , n45050 );
and ( n45052 , n45021 , n39367 );
and ( n45053 , n45050 , n45052 );
and ( n45054 , n45042 , n45052 );
or ( n45055 , n45051 , n45053 , n45054 );
and ( n45056 , n45047 , n39375 );
xor ( n45057 , n39241 , n39279 );
buf ( n572361 , n45057 );
buf ( n572362 , n572361 );
buf ( n45060 , n572362 );
and ( n45061 , n45060 , n39373 );
nor ( n45062 , n45056 , n45061 );
xnor ( n45063 , n45062 , n39380 );
and ( n45064 , n45055 , n45063 );
and ( n45065 , n45034 , n39367 );
and ( n45066 , n45063 , n45065 );
and ( n45067 , n45055 , n45065 );
or ( n45068 , n45064 , n45066 , n45067 );
and ( n45069 , n45060 , n39375 );
xor ( n45070 , n39239 , n39280 );
buf ( n572374 , n45070 );
buf ( n572375 , n572374 );
buf ( n45073 , n572375 );
and ( n45074 , n45073 , n39373 );
nor ( n45075 , n45069 , n45074 );
xnor ( n45076 , n45075 , n39380 );
and ( n45077 , n45068 , n45076 );
and ( n45078 , n45047 , n39367 );
and ( n45079 , n45076 , n45078 );
and ( n45080 , n45068 , n45078 );
or ( n45081 , n45077 , n45079 , n45080 );
and ( n45082 , n45073 , n39375 );
xor ( n45083 , n39180 , n39282 );
buf ( n572387 , n45083 );
buf ( n572388 , n572387 );
buf ( n45086 , n572388 );
and ( n45087 , n45086 , n39373 );
nor ( n45088 , n45082 , n45087 );
xnor ( n45089 , n45088 , n39380 );
and ( n45090 , n45081 , n45089 );
and ( n45091 , n45060 , n39367 );
and ( n45092 , n45089 , n45091 );
and ( n45093 , n45081 , n45091 );
or ( n45094 , n45090 , n45092 , n45093 );
and ( n45095 , n45086 , n39375 );
xor ( n45096 , n39148 , n39284 );
buf ( n572400 , n45096 );
buf ( n572401 , n572400 );
buf ( n45099 , n572401 );
and ( n45100 , n45099 , n39373 );
nor ( n45101 , n45095 , n45100 );
xnor ( n45102 , n45101 , n39380 );
and ( n45103 , n45094 , n45102 );
and ( n45104 , n45073 , n39367 );
and ( n45105 , n45102 , n45104 );
and ( n45106 , n45094 , n45104 );
or ( n45107 , n45103 , n45105 , n45106 );
and ( n45108 , n45099 , n39375 );
xor ( n45109 , n39143 , n39286 );
buf ( n572413 , n45109 );
buf ( n572414 , n572413 );
buf ( n45112 , n572414 );
and ( n45113 , n45112 , n39373 );
nor ( n45114 , n45108 , n45113 );
xnor ( n45115 , n45114 , n39380 );
and ( n45116 , n45107 , n45115 );
and ( n45117 , n45086 , n39367 );
and ( n45118 , n45115 , n45117 );
and ( n45119 , n45107 , n45117 );
or ( n45120 , n45116 , n45118 , n45119 );
and ( n45121 , n45112 , n39375 );
xor ( n45122 , n39141 , n39287 );
buf ( n572426 , n45122 );
buf ( n572427 , n572426 );
buf ( n45125 , n572427 );
and ( n45126 , n45125 , n39373 );
nor ( n45127 , n45121 , n45126 );
xnor ( n45128 , n45127 , n39380 );
and ( n45129 , n45120 , n45128 );
and ( n45130 , n45099 , n39367 );
and ( n45131 , n45128 , n45130 );
and ( n45132 , n45120 , n45130 );
or ( n45133 , n45129 , n45131 , n45132 );
and ( n45134 , n45125 , n39375 );
xor ( n45135 , n39138 , n39289 );
buf ( n572439 , n45135 );
buf ( n572440 , n572439 );
buf ( n45138 , n572440 );
and ( n45139 , n45138 , n39373 );
nor ( n45140 , n45134 , n45139 );
xnor ( n45141 , n45140 , n39380 );
and ( n45142 , n45133 , n45141 );
and ( n45143 , n45112 , n39367 );
and ( n45144 , n45141 , n45143 );
and ( n45145 , n45133 , n45143 );
or ( n45146 , n45142 , n45144 , n45145 );
and ( n45147 , n45138 , n39375 );
xor ( n45148 , n38972 , n39291 );
buf ( n572452 , n45148 );
buf ( n572453 , n572452 );
buf ( n45151 , n572453 );
and ( n45152 , n45151 , n39373 );
nor ( n45153 , n45147 , n45152 );
xnor ( n45154 , n45153 , n39380 );
and ( n45155 , n45146 , n45154 );
and ( n45156 , n45125 , n39367 );
and ( n45157 , n45154 , n45156 );
and ( n45158 , n45146 , n45156 );
or ( n45159 , n45155 , n45157 , n45158 );
and ( n45160 , n45151 , n39375 );
xor ( n45161 , n38971 , n39292 );
buf ( n572465 , n45161 );
buf ( n572466 , n572465 );
buf ( n45164 , n572466 );
and ( n45165 , n45164 , n39373 );
nor ( n45166 , n45160 , n45165 );
xnor ( n45167 , n45166 , n39380 );
and ( n45168 , n45159 , n45167 );
and ( n45169 , n45138 , n39367 );
and ( n45170 , n45167 , n45169 );
and ( n45171 , n45159 , n45169 );
or ( n45172 , n45168 , n45170 , n45171 );
and ( n45173 , n45164 , n39375 );
and ( n45174 , n44665 , n39373 );
nor ( n45175 , n45173 , n45174 );
xnor ( n45176 , n45175 , n39380 );
and ( n45177 , n45172 , n45176 );
and ( n45178 , n45151 , n39367 );
and ( n45179 , n45176 , n45178 );
and ( n45180 , n45172 , n45178 );
or ( n45181 , n45177 , n45179 , n45180 );
and ( n45182 , n44458 , n39480 );
and ( n45183 , n44357 , n39478 );
nor ( n45184 , n45182 , n45183 );
xnor ( n45185 , n45184 , n39462 );
and ( n45186 , n45181 , n45185 );
and ( n45187 , n44565 , n39396 );
and ( n45188 , n44520 , n39394 );
nor ( n45189 , n45187 , n45188 );
xnor ( n45190 , n45189 , n39401 );
and ( n45191 , n44665 , n39375 );
and ( n45192 , n44656 , n39373 );
nor ( n45193 , n45191 , n45192 );
xnor ( n45194 , n45193 , n39380 );
xor ( n45195 , n45190 , n45194 );
and ( n45196 , n45164 , n39367 );
xor ( n45197 , n45195 , n45196 );
and ( n45198 , n45185 , n45197 );
and ( n45199 , n45181 , n45197 );
or ( n45200 , n45186 , n45198 , n45199 );
and ( n45201 , n44264 , n39539 );
and ( n45202 , n43437 , n39537 );
nor ( n45203 , n45201 , n45202 );
xnor ( n45204 , n45203 , n39522 );
and ( n45205 , n45200 , n45204 );
and ( n45206 , n45190 , n45194 );
and ( n45207 , n45194 , n45196 );
and ( n45208 , n45190 , n45196 );
or ( n45209 , n45206 , n45207 , n45208 );
and ( n45210 , n44357 , n39480 );
and ( n45211 , n44347 , n39478 );
nor ( n45212 , n45210 , n45211 );
xnor ( n45213 , n45212 , n39462 );
xor ( n45214 , n45209 , n45213 );
xor ( n45215 , n44652 , n44660 );
xor ( n45216 , n45215 , n44666 );
xor ( n45217 , n45214 , n45216 );
and ( n45218 , n45204 , n45217 );
and ( n45219 , n45200 , n45217 );
or ( n45220 , n45205 , n45218 , n45219 );
and ( n45221 , n43437 , n39539 );
and ( n45222 , n43428 , n39537 );
nor ( n45223 , n45221 , n45222 );
xnor ( n45224 , n45223 , n39522 );
and ( n45225 , n45220 , n45224 );
buf ( n45226 , n557784 );
not ( n45227 , n45226 );
and ( n45228 , n45224 , n45227 );
and ( n45229 , n45220 , n45227 );
or ( n45230 , n45225 , n45228 , n45229 );
and ( n45231 , n43027 , n39760 );
and ( n45232 , n43019 , n39758 );
nor ( n45233 , n45231 , n45232 );
xnor ( n45234 , n45233 , n39742 );
and ( n45235 , n45230 , n45234 );
xor ( n45236 , n44688 , n44692 );
xor ( n45237 , n45236 , n44697 );
and ( n45238 , n45234 , n45237 );
and ( n45239 , n45230 , n45237 );
or ( n45240 , n45235 , n45238 , n45239 );
and ( n45241 , n42456 , n39896 );
and ( n45242 , n42048 , n39894 );
nor ( n45243 , n45241 , n45242 );
xnor ( n45244 , n45243 , n39857 );
xor ( n45245 , n45240 , n45244 );
xor ( n45246 , n44700 , n44704 );
xor ( n45247 , n45246 , n44707 );
xor ( n45248 , n45245 , n45247 );
and ( n45249 , n44987 , n45248 );
and ( n45250 , n45209 , n45213 );
and ( n45251 , n45213 , n45216 );
and ( n45252 , n45209 , n45216 );
or ( n45253 , n45250 , n45251 , n45252 );
and ( n45254 , n43200 , n39678 );
and ( n45255 , n43192 , n39676 );
nor ( n45256 , n45254 , n45255 );
xnor ( n45257 , n45256 , n39643 );
and ( n45258 , n45253 , n45257 );
xor ( n45259 , n44669 , n44673 );
xor ( n45260 , n45259 , n44685 );
and ( n45261 , n45257 , n45260 );
and ( n45262 , n45253 , n45260 );
or ( n45263 , n45258 , n45261 , n45262 );
buf ( n45264 , n557783 );
not ( n45265 , n45264 );
and ( n45266 , n45263 , n45265 );
xor ( n45267 , n44755 , n44759 );
xor ( n45268 , n45267 , n44764 );
and ( n45269 , n45265 , n45268 );
and ( n45270 , n45263 , n45268 );
or ( n45271 , n45266 , n45269 , n45270 );
and ( n45272 , n43019 , n39760 );
and ( n45273 , n42811 , n39758 );
nor ( n45274 , n45272 , n45273 );
xnor ( n45275 , n45274 , n39742 );
xor ( n45276 , n45271 , n45275 );
xor ( n45277 , n44767 , n44771 );
xor ( n45278 , n45277 , n44774 );
xor ( n45279 , n45276 , n45278 );
and ( n45280 , n45248 , n45279 );
and ( n45281 , n44987 , n45279 );
or ( n45282 , n45249 , n45280 , n45281 );
and ( n45283 , n40507 , n41292 );
and ( n45284 , n40373 , n41290 );
nor ( n45285 , n45283 , n45284 );
xnor ( n45286 , n45285 , n41041 );
and ( n45287 , n45282 , n45286 );
and ( n45288 , n45271 , n45275 );
and ( n45289 , n45275 , n45278 );
and ( n45290 , n45271 , n45278 );
or ( n45291 , n45288 , n45289 , n45290 );
and ( n45292 , n41182 , n40527 );
and ( n45293 , n41032 , n40525 );
nor ( n45294 , n45292 , n45293 );
xnor ( n45295 , n45294 , n40382 );
xor ( n45296 , n45291 , n45295 );
and ( n45297 , n41692 , n40258 );
and ( n45298 , n41615 , n40256 );
nor ( n45299 , n45297 , n45298 );
xnor ( n45300 , n45299 , n40169 );
xor ( n45301 , n45296 , n45300 );
and ( n45302 , n45286 , n45301 );
and ( n45303 , n45282 , n45301 );
or ( n45304 , n45287 , n45302 , n45303 );
and ( n45305 , n39948 , n42269 );
and ( n45306 , n39867 , n42266 );
nor ( n45307 , n45305 , n45306 );
xnor ( n45308 , n45307 , n41684 );
and ( n45309 , n45304 , n45308 );
and ( n45310 , n40186 , n41622 );
and ( n45311 , n40197 , n41620 );
nor ( n45312 , n45310 , n45311 );
xnor ( n45313 , n45312 , n41194 );
and ( n45314 , n45308 , n45313 );
and ( n45315 , n45304 , n45313 );
or ( n45316 , n45309 , n45314 , n45315 );
and ( n45317 , n45291 , n45295 );
and ( n45318 , n45295 , n45300 );
and ( n45319 , n45291 , n45300 );
or ( n45320 , n45317 , n45318 , n45319 );
and ( n45321 , n40492 , n41055 );
and ( n45322 , n40507 , n41053 );
nor ( n45323 , n45321 , n45322 );
xnor ( n45324 , n45323 , n40728 );
and ( n45325 , n45320 , n45324 );
xor ( n45326 , n44742 , n44746 );
xor ( n45327 , n45326 , n44751 );
and ( n45328 , n45324 , n45327 );
and ( n45329 , n45320 , n45327 );
or ( n45330 , n45325 , n45328 , n45329 );
and ( n45331 , n40009 , n41984 );
and ( n45332 , n39948 , n41982 );
nor ( n45333 , n45331 , n45332 );
xnor ( n45334 , n45333 , n41687 );
xor ( n45335 , n45330 , n45334 );
xor ( n45336 , n44866 , n44870 );
xor ( n45337 , n45336 , n44883 );
xor ( n45338 , n45335 , n45337 );
and ( n45339 , n45316 , n45338 );
xor ( n45340 , n44964 , n44968 );
xor ( n45341 , n45340 , n44971 );
and ( n45342 , n45338 , n45341 );
and ( n45343 , n45316 , n45341 );
or ( n45344 , n45339 , n45342 , n45343 );
xor ( n45345 , n44850 , n44854 );
xor ( n45346 , n45345 , n44859 );
and ( n45347 , n45344 , n45346 );
xor ( n45348 , n44960 , n44974 );
xor ( n45349 , n45348 , n44977 );
and ( n45350 , n45346 , n45349 );
and ( n45351 , n45344 , n45349 );
or ( n45352 , n45347 , n45350 , n45351 );
and ( n45353 , n44982 , n45352 );
and ( n45354 , n44980 , n45352 );
or ( n45355 , n44983 , n45353 , n45354 );
and ( n45356 , n44924 , n45355 );
and ( n45357 , n40738 , n41055 );
and ( n45358 , n40492 , n41053 );
nor ( n45359 , n45357 , n45358 );
xnor ( n45360 , n45359 , n40728 );
and ( n45361 , n41047 , n40746 );
and ( n45362 , n40869 , n40744 );
nor ( n45363 , n45361 , n45362 );
xnor ( n45364 , n45363 , n40501 );
and ( n45365 , n45360 , n45364 );
xor ( n45366 , n44928 , n44932 );
xor ( n45367 , n45366 , n44935 );
and ( n45368 , n45364 , n45367 );
and ( n45369 , n45360 , n45367 );
or ( n45370 , n45365 , n45368 , n45369 );
xor ( n45371 , n45320 , n45324 );
xor ( n45372 , n45371 , n45327 );
and ( n45373 , n45370 , n45372 );
xor ( n45374 , n44938 , n44942 );
xor ( n45375 , n45374 , n44945 );
and ( n45376 , n45372 , n45375 );
and ( n45377 , n45370 , n45375 );
or ( n45378 , n45373 , n45376 , n45377 );
and ( n45379 , n44520 , n39480 );
and ( n45380 , n44458 , n39478 );
nor ( n45381 , n45379 , n45380 );
xnor ( n45382 , n45381 , n39462 );
and ( n45383 , n44656 , n39396 );
and ( n45384 , n44565 , n39394 );
nor ( n45385 , n45383 , n45384 );
xnor ( n45386 , n45385 , n39401 );
and ( n45387 , n45382 , n45386 );
xor ( n45388 , n45172 , n45176 );
xor ( n45389 , n45388 , n45178 );
and ( n45390 , n45386 , n45389 );
and ( n45391 , n45382 , n45389 );
or ( n45392 , n45387 , n45390 , n45391 );
and ( n45393 , n44347 , n39539 );
and ( n45394 , n44264 , n39537 );
nor ( n45395 , n45393 , n45394 );
xnor ( n45396 , n45395 , n39522 );
and ( n45397 , n45392 , n45396 );
xor ( n45398 , n45181 , n45185 );
xor ( n45399 , n45398 , n45197 );
and ( n45400 , n45396 , n45399 );
and ( n45401 , n45392 , n45399 );
or ( n45402 , n45397 , n45400 , n45401 );
and ( n45403 , n43192 , n39760 );
and ( n45404 , n43073 , n39758 );
nor ( n45405 , n45403 , n45404 );
xnor ( n45406 , n45405 , n39742 );
and ( n45407 , n45402 , n45406 );
and ( n45408 , n43428 , n39678 );
and ( n45409 , n43200 , n39676 );
nor ( n45410 , n45408 , n45409 );
xnor ( n45411 , n45410 , n39643 );
and ( n45412 , n45406 , n45411 );
and ( n45413 , n45402 , n45411 );
or ( n45414 , n45407 , n45412 , n45413 );
and ( n45415 , n43073 , n39760 );
and ( n45416 , n43027 , n39758 );
nor ( n45417 , n45415 , n45416 );
xnor ( n45418 , n45417 , n39742 );
and ( n45419 , n45414 , n45418 );
xor ( n45420 , n45253 , n45257 );
xor ( n45421 , n45420 , n45260 );
and ( n45422 , n45418 , n45421 );
and ( n45423 , n45414 , n45421 );
or ( n45424 , n45419 , n45422 , n45423 );
and ( n45425 , n42811 , n39896 );
and ( n45426 , n42456 , n39894 );
nor ( n45427 , n45425 , n45426 );
xnor ( n45428 , n45427 , n39857 );
and ( n45429 , n45424 , n45428 );
xor ( n45430 , n45263 , n45265 );
xor ( n45431 , n45430 , n45268 );
and ( n45432 , n45428 , n45431 );
and ( n45433 , n45424 , n45431 );
or ( n45434 , n45429 , n45432 , n45433 );
and ( n45435 , n41807 , n40258 );
and ( n45436 , n41692 , n40256 );
nor ( n45437 , n45435 , n45436 );
xnor ( n45438 , n45437 , n40169 );
and ( n45439 , n45434 , n45438 );
and ( n45440 , n42061 , n40053 );
and ( n45441 , n41816 , n40051 );
nor ( n45442 , n45440 , n45441 );
xnor ( n45443 , n45442 , n39999 );
and ( n45444 , n45438 , n45443 );
and ( n45445 , n45434 , n45443 );
or ( n45446 , n45439 , n45444 , n45445 );
and ( n45447 , n45240 , n45244 );
and ( n45448 , n45244 , n45247 );
and ( n45449 , n45240 , n45247 );
or ( n45450 , n45447 , n45448 , n45449 );
and ( n45451 , n45446 , n45450 );
xor ( n45452 , n44710 , n44714 );
xor ( n45453 , n45452 , n44739 );
and ( n45454 , n45450 , n45453 );
and ( n45455 , n45446 , n45453 );
or ( n45456 , n45451 , n45454 , n45455 );
and ( n45457 , n40373 , n41292 );
and ( n45458 , n40388 , n41290 );
nor ( n45459 , n45457 , n45458 );
xnor ( n45460 , n45459 , n41041 );
and ( n45461 , n45456 , n45460 );
xor ( n45462 , n44822 , n44826 );
xor ( n45463 , n45462 , n44839 );
and ( n45464 , n45460 , n45463 );
and ( n45465 , n45456 , n45463 );
or ( n45466 , n45461 , n45464 , n45465 );
and ( n45467 , n45378 , n45466 );
xor ( n45468 , n44948 , n44952 );
xor ( n45469 , n45468 , n44957 );
and ( n45470 , n45466 , n45469 );
and ( n45471 , n45378 , n45469 );
or ( n45472 , n45467 , n45470 , n45471 );
and ( n45473 , n45330 , n45334 );
and ( n45474 , n45334 , n45337 );
and ( n45475 , n45330 , n45337 );
or ( n45476 , n45473 , n45474 , n45475 );
and ( n45477 , n45472 , n45476 );
xor ( n45478 , n44902 , n44906 );
xor ( n45479 , n45478 , n44908 );
xor ( n45480 , n45344 , n45346 );
xor ( n45481 , n45480 , n45349 );
and ( n45482 , n45479 , n45481 );
xor ( n45483 , n45472 , n45476 );
and ( n45484 , n45481 , n45483 );
and ( n45485 , n45479 , n45483 );
or ( n45486 , n45482 , n45484 , n45485 );
and ( n45487 , n45477 , n45486 );
xor ( n45488 , n44980 , n44982 );
xor ( n45489 , n45488 , n45352 );
and ( n45490 , n45486 , n45489 );
and ( n45491 , n45477 , n45489 );
or ( n45492 , n45487 , n45490 , n45491 );
and ( n45493 , n45355 , n45492 );
and ( n45494 , n44924 , n45492 );
or ( n45495 , n45356 , n45493 , n45494 );
and ( n45496 , n44921 , n45495 );
and ( n45497 , n44818 , n45495 );
or ( n45498 , n44922 , n45496 , n45497 );
and ( n45499 , n44815 , n45498 );
and ( n45500 , n44445 , n45498 );
or ( n45501 , n44816 , n45499 , n45500 );
and ( n45502 , n44443 , n45501 );
xor ( n45503 , n44443 , n45501 );
xor ( n45504 , n44445 , n44815 );
xor ( n45505 , n45504 , n45498 );
xor ( n45506 , n44818 , n44921 );
xor ( n45507 , n45506 , n45495 );
xor ( n45508 , n44924 , n45355 );
xor ( n45509 , n45508 , n45492 );
xor ( n45510 , n45477 , n45486 );
xor ( n45511 , n45510 , n45489 );
xor ( n45512 , n44994 , n45002 );
and ( n45513 , n44991 , n39394 );
not ( n45514 , n45513 );
and ( n45515 , n45514 , n39401 );
and ( n45516 , n44991 , n39396 );
and ( n45517 , n44999 , n39394 );
nor ( n45518 , n45516 , n45517 );
xnor ( n45519 , n45518 , n39401 );
and ( n45520 , n45515 , n45519 );
and ( n45521 , n44999 , n39396 );
and ( n45522 , n45008 , n39394 );
nor ( n45523 , n45521 , n45522 );
xnor ( n45524 , n45523 , n39401 );
and ( n45525 , n45520 , n45524 );
and ( n45526 , n45524 , n44992 );
and ( n45527 , n45520 , n44992 );
or ( n45528 , n45525 , n45526 , n45527 );
and ( n45529 , n45512 , n45528 );
and ( n45530 , n45008 , n39396 );
and ( n45531 , n45021 , n39394 );
nor ( n45532 , n45530 , n45531 );
xnor ( n45533 , n45532 , n39401 );
and ( n45534 , n45528 , n45533 );
and ( n45535 , n45512 , n45533 );
or ( n45536 , n45529 , n45534 , n45535 );
and ( n45537 , n45021 , n39396 );
and ( n45538 , n45034 , n39394 );
nor ( n45539 , n45537 , n45538 );
xnor ( n45540 , n45539 , n39401 );
and ( n45541 , n45536 , n45540 );
xor ( n45542 , n45003 , n45011 );
xor ( n45543 , n45542 , n45013 );
and ( n45544 , n45540 , n45543 );
and ( n45545 , n45536 , n45543 );
or ( n45546 , n45541 , n45544 , n45545 );
and ( n45547 , n45034 , n39396 );
and ( n45548 , n45047 , n39394 );
nor ( n45549 , n45547 , n45548 );
xnor ( n45550 , n45549 , n39401 );
and ( n45551 , n45546 , n45550 );
xor ( n45552 , n45016 , n45024 );
xor ( n45553 , n45552 , n45026 );
and ( n45554 , n45550 , n45553 );
and ( n45555 , n45546 , n45553 );
or ( n45556 , n45551 , n45554 , n45555 );
and ( n45557 , n45047 , n39396 );
and ( n45558 , n45060 , n39394 );
nor ( n45559 , n45557 , n45558 );
xnor ( n45560 , n45559 , n39401 );
and ( n45561 , n45556 , n45560 );
xor ( n45562 , n45029 , n45037 );
xor ( n45563 , n45562 , n45039 );
and ( n45564 , n45560 , n45563 );
and ( n45565 , n45556 , n45563 );
or ( n45566 , n45561 , n45564 , n45565 );
and ( n45567 , n45060 , n39396 );
and ( n45568 , n45073 , n39394 );
nor ( n45569 , n45567 , n45568 );
xnor ( n45570 , n45569 , n39401 );
and ( n45571 , n45566 , n45570 );
xor ( n45572 , n45042 , n45050 );
xor ( n45573 , n45572 , n45052 );
and ( n45574 , n45570 , n45573 );
and ( n45575 , n45566 , n45573 );
or ( n45576 , n45571 , n45574 , n45575 );
and ( n45577 , n45073 , n39396 );
and ( n45578 , n45086 , n39394 );
nor ( n45579 , n45577 , n45578 );
xnor ( n45580 , n45579 , n39401 );
and ( n45581 , n45576 , n45580 );
xor ( n45582 , n45055 , n45063 );
xor ( n45583 , n45582 , n45065 );
and ( n45584 , n45580 , n45583 );
and ( n45585 , n45576 , n45583 );
or ( n45586 , n45581 , n45584 , n45585 );
and ( n45587 , n45086 , n39396 );
and ( n45588 , n45099 , n39394 );
nor ( n45589 , n45587 , n45588 );
xnor ( n45590 , n45589 , n39401 );
and ( n45591 , n45586 , n45590 );
xor ( n45592 , n45068 , n45076 );
xor ( n45593 , n45592 , n45078 );
and ( n45594 , n45590 , n45593 );
and ( n45595 , n45586 , n45593 );
or ( n45596 , n45591 , n45594 , n45595 );
and ( n45597 , n45099 , n39396 );
and ( n45598 , n45112 , n39394 );
nor ( n45599 , n45597 , n45598 );
xnor ( n45600 , n45599 , n39401 );
and ( n45601 , n45596 , n45600 );
xor ( n45602 , n45081 , n45089 );
xor ( n45603 , n45602 , n45091 );
and ( n45604 , n45600 , n45603 );
and ( n45605 , n45596 , n45603 );
or ( n45606 , n45601 , n45604 , n45605 );
and ( n45607 , n45112 , n39396 );
and ( n45608 , n45125 , n39394 );
nor ( n45609 , n45607 , n45608 );
xnor ( n45610 , n45609 , n39401 );
and ( n45611 , n45606 , n45610 );
xor ( n45612 , n45094 , n45102 );
xor ( n45613 , n45612 , n45104 );
and ( n45614 , n45610 , n45613 );
and ( n45615 , n45606 , n45613 );
or ( n45616 , n45611 , n45614 , n45615 );
and ( n45617 , n45125 , n39396 );
and ( n45618 , n45138 , n39394 );
nor ( n45619 , n45617 , n45618 );
xnor ( n45620 , n45619 , n39401 );
and ( n45621 , n45616 , n45620 );
xor ( n45622 , n45107 , n45115 );
xor ( n45623 , n45622 , n45117 );
and ( n45624 , n45620 , n45623 );
and ( n45625 , n45616 , n45623 );
or ( n45626 , n45621 , n45624 , n45625 );
and ( n45627 , n45138 , n39396 );
and ( n45628 , n45151 , n39394 );
nor ( n45629 , n45627 , n45628 );
xnor ( n45630 , n45629 , n39401 );
and ( n45631 , n45626 , n45630 );
xor ( n45632 , n45120 , n45128 );
xor ( n45633 , n45632 , n45130 );
and ( n45634 , n45630 , n45633 );
and ( n45635 , n45626 , n45633 );
or ( n45636 , n45631 , n45634 , n45635 );
and ( n45637 , n45151 , n39396 );
and ( n45638 , n45164 , n39394 );
nor ( n45639 , n45637 , n45638 );
xnor ( n45640 , n45639 , n39401 );
and ( n45641 , n45636 , n45640 );
xor ( n45642 , n45133 , n45141 );
xor ( n45643 , n45642 , n45143 );
and ( n45644 , n45640 , n45643 );
and ( n45645 , n45636 , n45643 );
or ( n45646 , n45641 , n45644 , n45645 );
and ( n45647 , n45164 , n39396 );
and ( n45648 , n44665 , n39394 );
nor ( n45649 , n45647 , n45648 );
xnor ( n45650 , n45649 , n39401 );
and ( n45651 , n45646 , n45650 );
xor ( n45652 , n45146 , n45154 );
xor ( n45653 , n45652 , n45156 );
and ( n45654 , n45650 , n45653 );
and ( n45655 , n45646 , n45653 );
or ( n45656 , n45651 , n45654 , n45655 );
and ( n45657 , n44458 , n39539 );
and ( n45658 , n44357 , n39537 );
nor ( n45659 , n45657 , n45658 );
xnor ( n45660 , n45659 , n39522 );
and ( n45661 , n45656 , n45660 );
and ( n45662 , n44565 , n39480 );
and ( n45663 , n44520 , n39478 );
nor ( n45664 , n45662 , n45663 );
xnor ( n45665 , n45664 , n39462 );
and ( n45666 , n44665 , n39396 );
and ( n45667 , n44656 , n39394 );
nor ( n45668 , n45666 , n45667 );
xnor ( n45669 , n45668 , n39401 );
xor ( n45670 , n45665 , n45669 );
xor ( n45671 , n45159 , n45167 );
xor ( n45672 , n45671 , n45169 );
xor ( n45673 , n45670 , n45672 );
and ( n45674 , n45660 , n45673 );
and ( n45675 , n45656 , n45673 );
or ( n45676 , n45661 , n45674 , n45675 );
and ( n45677 , n44264 , n39678 );
and ( n45678 , n43437 , n39676 );
nor ( n45679 , n45677 , n45678 );
xnor ( n45680 , n45679 , n39643 );
and ( n45681 , n45676 , n45680 );
and ( n45682 , n45665 , n45669 );
and ( n45683 , n45669 , n45672 );
and ( n45684 , n45665 , n45672 );
or ( n45685 , n45682 , n45683 , n45684 );
and ( n45686 , n44357 , n39539 );
and ( n45687 , n44347 , n39537 );
nor ( n45688 , n45686 , n45687 );
xnor ( n45689 , n45688 , n39522 );
xor ( n45690 , n45685 , n45689 );
xor ( n45691 , n45382 , n45386 );
xor ( n45692 , n45691 , n45389 );
xor ( n45693 , n45690 , n45692 );
and ( n45694 , n45680 , n45693 );
and ( n45695 , n45676 , n45693 );
or ( n45696 , n45681 , n45694 , n45695 );
buf ( n45697 , n557786 );
not ( n45698 , n45697 );
and ( n45699 , n45696 , n45698 );
xor ( n45700 , n45392 , n45396 );
xor ( n45701 , n45700 , n45399 );
and ( n45702 , n45698 , n45701 );
and ( n45703 , n45696 , n45701 );
or ( n45704 , n45699 , n45702 , n45703 );
and ( n45705 , n43027 , n39896 );
and ( n45706 , n43019 , n39894 );
nor ( n45707 , n45705 , n45706 );
xnor ( n45708 , n45707 , n39857 );
and ( n45709 , n45704 , n45708 );
xor ( n45710 , n45402 , n45406 );
xor ( n45711 , n45710 , n45411 );
and ( n45712 , n45708 , n45711 );
and ( n45713 , n45704 , n45711 );
or ( n45714 , n45709 , n45712 , n45713 );
and ( n45715 , n42456 , n40053 );
and ( n45716 , n42048 , n40051 );
nor ( n45717 , n45715 , n45716 );
xnor ( n45718 , n45717 , n39999 );
and ( n45719 , n45714 , n45718 );
xor ( n45720 , n45414 , n45418 );
xor ( n45721 , n45720 , n45421 );
and ( n45722 , n45718 , n45721 );
and ( n45723 , n45714 , n45721 );
or ( n45724 , n45719 , n45722 , n45723 );
and ( n45725 , n45685 , n45689 );
and ( n45726 , n45689 , n45692 );
and ( n45727 , n45685 , n45692 );
or ( n45728 , n45725 , n45726 , n45727 );
and ( n45729 , n43200 , n39760 );
and ( n45730 , n43192 , n39758 );
nor ( n45731 , n45729 , n45730 );
xnor ( n45732 , n45731 , n39742 );
and ( n45733 , n45728 , n45732 );
and ( n45734 , n43437 , n39678 );
and ( n45735 , n43428 , n39676 );
nor ( n45736 , n45734 , n45735 );
xnor ( n45737 , n45736 , n39643 );
and ( n45738 , n45732 , n45737 );
and ( n45739 , n45728 , n45737 );
or ( n45740 , n45733 , n45738 , n45739 );
buf ( n45741 , n557785 );
not ( n45742 , n45741 );
and ( n45743 , n45740 , n45742 );
xor ( n45744 , n45200 , n45204 );
xor ( n45745 , n45744 , n45217 );
and ( n45746 , n45742 , n45745 );
and ( n45747 , n45740 , n45745 );
or ( n45748 , n45743 , n45746 , n45747 );
and ( n45749 , n43019 , n39896 );
and ( n45750 , n42811 , n39894 );
nor ( n45751 , n45749 , n45750 );
xnor ( n45752 , n45751 , n39857 );
and ( n45753 , n45748 , n45752 );
xor ( n45754 , n45220 , n45224 );
xor ( n45755 , n45754 , n45227 );
and ( n45756 , n45752 , n45755 );
and ( n45757 , n45748 , n45755 );
or ( n45758 , n45753 , n45756 , n45757 );
and ( n45759 , n41816 , n40258 );
and ( n45760 , n41807 , n40256 );
nor ( n45761 , n45759 , n45760 );
xnor ( n45762 , n45761 , n40169 );
xor ( n45763 , n45758 , n45762 );
xor ( n45764 , n45230 , n45234 );
xor ( n45765 , n45764 , n45237 );
xor ( n45766 , n45763 , n45765 );
and ( n45767 , n45724 , n45766 );
xor ( n45768 , n45424 , n45428 );
xor ( n45769 , n45768 , n45431 );
and ( n45770 , n45766 , n45769 );
and ( n45771 , n45724 , n45769 );
or ( n45772 , n45767 , n45770 , n45771 );
and ( n45773 , n41182 , n40746 );
and ( n45774 , n41032 , n40744 );
nor ( n45775 , n45773 , n45774 );
xnor ( n45776 , n45775 , n40501 );
and ( n45777 , n41692 , n40527 );
and ( n45778 , n41615 , n40525 );
nor ( n45779 , n45777 , n45778 );
xnor ( n45780 , n45779 , n40382 );
and ( n45781 , n45776 , n45780 );
and ( n45782 , n42048 , n40053 );
and ( n45783 , n42061 , n40051 );
nor ( n45784 , n45782 , n45783 );
xnor ( n45785 , n45784 , n39999 );
and ( n45786 , n45780 , n45785 );
and ( n45787 , n45776 , n45785 );
or ( n45788 , n45781 , n45786 , n45787 );
and ( n45789 , n45758 , n45762 );
and ( n45790 , n45762 , n45765 );
and ( n45791 , n45758 , n45765 );
or ( n45792 , n45789 , n45790 , n45791 );
xor ( n45793 , n45788 , n45792 );
and ( n45794 , n41032 , n40746 );
and ( n45795 , n41047 , n40744 );
nor ( n45796 , n45794 , n45795 );
xnor ( n45797 , n45796 , n40501 );
xor ( n45798 , n45793 , n45797 );
and ( n45799 , n45772 , n45798 );
xor ( n45800 , n44987 , n45248 );
xor ( n45801 , n45800 , n45279 );
and ( n45802 , n45798 , n45801 );
and ( n45803 , n45772 , n45801 );
or ( n45804 , n45799 , n45802 , n45803 );
and ( n45805 , n40009 , n42269 );
and ( n45806 , n39948 , n42266 );
nor ( n45807 , n45805 , n45806 );
xnor ( n45808 , n45807 , n41684 );
and ( n45809 , n45804 , n45808 );
and ( n45810 , n40197 , n41984 );
and ( n45811 , n40148 , n41982 );
nor ( n45812 , n45810 , n45811 );
xnor ( n45813 , n45812 , n41687 );
and ( n45814 , n45808 , n45813 );
and ( n45815 , n45804 , n45813 );
or ( n45816 , n45809 , n45814 , n45815 );
and ( n45817 , n40492 , n41292 );
and ( n45818 , n40507 , n41290 );
nor ( n45819 , n45817 , n45818 );
xnor ( n45820 , n45819 , n41041 );
and ( n45821 , n40869 , n41055 );
and ( n45822 , n40738 , n41053 );
nor ( n45823 , n45821 , n45822 );
xnor ( n45824 , n45823 , n40728 );
and ( n45825 , n45820 , n45824 );
xor ( n45826 , n45434 , n45438 );
xor ( n45827 , n45826 , n45443 );
and ( n45828 , n45824 , n45827 );
and ( n45829 , n45820 , n45827 );
or ( n45830 , n45825 , n45828 , n45829 );
and ( n45831 , n40388 , n41622 );
and ( n45832 , n40186 , n41620 );
nor ( n45833 , n45831 , n45832 );
xnor ( n45834 , n45833 , n41194 );
and ( n45835 , n45830 , n45834 );
xor ( n45836 , n45282 , n45286 );
xor ( n45837 , n45836 , n45301 );
and ( n45838 , n45834 , n45837 );
and ( n45839 , n45830 , n45837 );
or ( n45840 , n45835 , n45838 , n45839 );
and ( n45841 , n45816 , n45840 );
xor ( n45842 , n45370 , n45372 );
xor ( n45843 , n45842 , n45375 );
and ( n45844 , n45840 , n45843 );
and ( n45845 , n45816 , n45843 );
or ( n45846 , n45841 , n45844 , n45845 );
and ( n45847 , n45788 , n45792 );
and ( n45848 , n45792 , n45797 );
and ( n45849 , n45788 , n45797 );
or ( n45850 , n45847 , n45848 , n45849 );
xor ( n45851 , n45446 , n45450 );
xor ( n45852 , n45851 , n45453 );
and ( n45853 , n45850 , n45852 );
xor ( n45854 , n45360 , n45364 );
xor ( n45855 , n45854 , n45367 );
and ( n45856 , n45852 , n45855 );
and ( n45857 , n45850 , n45855 );
or ( n45858 , n45853 , n45856 , n45857 );
and ( n45859 , n40148 , n41984 );
and ( n45860 , n40009 , n41982 );
nor ( n45861 , n45859 , n45860 );
xnor ( n45862 , n45861 , n41687 );
and ( n45863 , n45858 , n45862 );
xor ( n45864 , n45456 , n45460 );
xor ( n45865 , n45864 , n45463 );
and ( n45866 , n45862 , n45865 );
and ( n45867 , n45858 , n45865 );
or ( n45868 , n45863 , n45866 , n45867 );
and ( n45869 , n45846 , n45868 );
xor ( n45870 , n45378 , n45466 );
xor ( n45871 , n45870 , n45469 );
and ( n45872 , n45868 , n45871 );
and ( n45873 , n45846 , n45871 );
or ( n45874 , n45869 , n45872 , n45873 );
xor ( n45875 , n45479 , n45481 );
xor ( n45876 , n45875 , n45483 );
and ( n45877 , n45874 , n45876 );
and ( n45878 , n44520 , n39539 );
and ( n45879 , n44458 , n39537 );
nor ( n45880 , n45878 , n45879 );
xnor ( n45881 , n45880 , n39522 );
and ( n45882 , n44656 , n39480 );
and ( n45883 , n44565 , n39478 );
nor ( n45884 , n45882 , n45883 );
xnor ( n45885 , n45884 , n39462 );
and ( n45886 , n45881 , n45885 );
xor ( n45887 , n45646 , n45650 );
xor ( n45888 , n45887 , n45653 );
and ( n45889 , n45885 , n45888 );
and ( n45890 , n45881 , n45888 );
or ( n45891 , n45886 , n45889 , n45890 );
and ( n45892 , n44347 , n39678 );
and ( n45893 , n44264 , n39676 );
nor ( n45894 , n45892 , n45893 );
xnor ( n45895 , n45894 , n39643 );
and ( n45896 , n45891 , n45895 );
xor ( n45897 , n45656 , n45660 );
xor ( n45898 , n45897 , n45673 );
and ( n45899 , n45895 , n45898 );
and ( n45900 , n45891 , n45898 );
or ( n45901 , n45896 , n45899 , n45900 );
and ( n45902 , n43428 , n39760 );
and ( n45903 , n43200 , n39758 );
nor ( n45904 , n45902 , n45903 );
xnor ( n45905 , n45904 , n39742 );
and ( n45906 , n45901 , n45905 );
buf ( n45907 , n557787 );
not ( n45908 , n45907 );
and ( n45909 , n45905 , n45908 );
and ( n45910 , n45901 , n45908 );
or ( n45911 , n45906 , n45909 , n45910 );
and ( n45912 , n43073 , n39896 );
and ( n45913 , n43027 , n39894 );
nor ( n45914 , n45912 , n45913 );
xnor ( n45915 , n45914 , n39857 );
and ( n45916 , n45911 , n45915 );
xor ( n45917 , n45728 , n45732 );
xor ( n45918 , n45917 , n45737 );
and ( n45919 , n45915 , n45918 );
and ( n45920 , n45911 , n45918 );
or ( n45921 , n45916 , n45919 , n45920 );
and ( n45922 , n42811 , n40053 );
and ( n45923 , n42456 , n40051 );
nor ( n45924 , n45922 , n45923 );
xnor ( n45925 , n45924 , n39999 );
and ( n45926 , n45921 , n45925 );
xor ( n45927 , n45740 , n45742 );
xor ( n45928 , n45927 , n45745 );
and ( n45929 , n45925 , n45928 );
and ( n45930 , n45921 , n45928 );
or ( n45931 , n45926 , n45929 , n45930 );
and ( n45932 , n42061 , n40258 );
and ( n45933 , n41816 , n40256 );
nor ( n45934 , n45932 , n45933 );
xnor ( n45935 , n45934 , n40169 );
and ( n45936 , n45931 , n45935 );
xor ( n45937 , n45748 , n45752 );
xor ( n45938 , n45937 , n45755 );
and ( n45939 , n45935 , n45938 );
and ( n45940 , n45931 , n45938 );
or ( n45941 , n45936 , n45939 , n45940 );
and ( n45942 , n40738 , n41292 );
and ( n45943 , n40492 , n41290 );
nor ( n45944 , n45942 , n45943 );
xnor ( n45945 , n45944 , n41041 );
and ( n45946 , n45941 , n45945 );
and ( n45947 , n41047 , n41055 );
and ( n45948 , n40869 , n41053 );
nor ( n45949 , n45947 , n45948 );
xnor ( n45950 , n45949 , n40728 );
and ( n45951 , n45945 , n45950 );
and ( n45952 , n45941 , n45950 );
or ( n45953 , n45946 , n45951 , n45952 );
and ( n45954 , n40373 , n41622 );
and ( n45955 , n40388 , n41620 );
nor ( n45956 , n45954 , n45955 );
xnor ( n45957 , n45956 , n41194 );
and ( n45958 , n45953 , n45957 );
xor ( n45959 , n45820 , n45824 );
xor ( n45960 , n45959 , n45827 );
and ( n45961 , n45957 , n45960 );
and ( n45962 , n45953 , n45960 );
or ( n45963 , n45958 , n45961 , n45962 );
xor ( n45964 , n45830 , n45834 );
xor ( n45965 , n45964 , n45837 );
and ( n45966 , n45963 , n45965 );
xor ( n45967 , n45850 , n45852 );
xor ( n45968 , n45967 , n45855 );
and ( n45969 , n45965 , n45968 );
and ( n45970 , n45963 , n45968 );
or ( n45971 , n45966 , n45969 , n45970 );
xor ( n45972 , n45304 , n45308 );
xor ( n45973 , n45972 , n45313 );
and ( n45974 , n45971 , n45973 );
xor ( n45975 , n45858 , n45862 );
xor ( n45976 , n45975 , n45865 );
and ( n45977 , n45973 , n45976 );
and ( n45978 , n45971 , n45976 );
or ( n45979 , n45974 , n45977 , n45978 );
xor ( n45980 , n45846 , n45868 );
xor ( n45981 , n45980 , n45871 );
and ( n45982 , n45979 , n45981 );
xor ( n45983 , n45316 , n45338 );
xor ( n45984 , n45983 , n45341 );
and ( n45985 , n45981 , n45984 );
and ( n45986 , n45979 , n45984 );
or ( n45987 , n45982 , n45985 , n45986 );
and ( n45988 , n45876 , n45987 );
and ( n45989 , n45874 , n45987 );
or ( n45990 , n45877 , n45988 , n45989 );
and ( n45991 , n45511 , n45990 );
xor ( n45992 , n45511 , n45990 );
xor ( n45993 , n45874 , n45876 );
xor ( n45994 , n45993 , n45987 );
and ( n45995 , n41615 , n40746 );
and ( n45996 , n41182 , n40744 );
nor ( n45997 , n45995 , n45996 );
xnor ( n45998 , n45997 , n40501 );
and ( n45999 , n41807 , n40527 );
and ( n46000 , n41692 , n40525 );
nor ( n46001 , n45999 , n46000 );
xnor ( n46002 , n46001 , n40382 );
and ( n46003 , n45998 , n46002 );
xor ( n46004 , n45714 , n45718 );
xor ( n573308 , n46004 , n45721 );
and ( n573309 , n46002 , n573308 );
and ( n573310 , n45998 , n573308 );
or ( n46005 , n46003 , n573309 , n573310 );
xor ( n46006 , n45776 , n45780 );
xor ( n46007 , n46006 , n45785 );
and ( n46008 , n46005 , n46007 );
xor ( n46009 , n45724 , n45766 );
xor ( n46010 , n46009 , n45769 );
and ( n46011 , n46007 , n46010 );
and ( n46012 , n46005 , n46010 );
or ( n46013 , n46008 , n46011 , n46012 );
and ( n46014 , n40148 , n42269 );
and ( n46015 , n40009 , n42266 );
nor ( n46016 , n46014 , n46015 );
xnor ( n46017 , n46016 , n41684 );
and ( n46018 , n46013 , n46017 );
and ( n46019 , n40186 , n41984 );
and ( n46020 , n40197 , n41982 );
nor ( n46021 , n46019 , n46020 );
xnor ( n46022 , n46021 , n41687 );
and ( n46023 , n46017 , n46022 );
and ( n46024 , n46013 , n46022 );
or ( n46025 , n46018 , n46023 , n46024 );
xor ( n46026 , n45515 , n45519 );
and ( n46027 , n44991 , n39478 );
not ( n46028 , n46027 );
and ( n46029 , n46028 , n39462 );
and ( n46030 , n44991 , n39480 );
and ( n46031 , n44999 , n39478 );
nor ( n46032 , n46030 , n46031 );
xnor ( n46033 , n46032 , n39462 );
and ( n46034 , n46029 , n46033 );
and ( n46035 , n44999 , n39480 );
and ( n46036 , n45008 , n39478 );
nor ( n46037 , n46035 , n46036 );
xnor ( n46038 , n46037 , n39462 );
and ( n46039 , n46034 , n46038 );
and ( n46040 , n46038 , n45513 );
and ( n46041 , n46034 , n45513 );
or ( n46042 , n46039 , n46040 , n46041 );
and ( n46043 , n46026 , n46042 );
and ( n46044 , n45008 , n39480 );
and ( n46045 , n45021 , n39478 );
nor ( n46046 , n46044 , n46045 );
xnor ( n46047 , n46046 , n39462 );
and ( n46048 , n46042 , n46047 );
and ( n46049 , n46026 , n46047 );
or ( n46050 , n46043 , n46048 , n46049 );
and ( n46051 , n45021 , n39480 );
and ( n46052 , n45034 , n39478 );
nor ( n46053 , n46051 , n46052 );
xnor ( n46054 , n46053 , n39462 );
and ( n46055 , n46050 , n46054 );
xor ( n46056 , n45520 , n45524 );
xor ( n46057 , n46056 , n44992 );
and ( n46058 , n46054 , n46057 );
and ( n46059 , n46050 , n46057 );
or ( n46060 , n46055 , n46058 , n46059 );
and ( n46061 , n45034 , n39480 );
and ( n46062 , n45047 , n39478 );
nor ( n46063 , n46061 , n46062 );
xnor ( n46064 , n46063 , n39462 );
and ( n46065 , n46060 , n46064 );
xor ( n46066 , n45512 , n45528 );
xor ( n46067 , n46066 , n45533 );
and ( n46068 , n46064 , n46067 );
and ( n46069 , n46060 , n46067 );
or ( n46070 , n46065 , n46068 , n46069 );
and ( n46071 , n45047 , n39480 );
and ( n46072 , n45060 , n39478 );
nor ( n46073 , n46071 , n46072 );
xnor ( n46074 , n46073 , n39462 );
and ( n46075 , n46070 , n46074 );
xor ( n46076 , n45536 , n45540 );
xor ( n46077 , n46076 , n45543 );
and ( n46078 , n46074 , n46077 );
and ( n46079 , n46070 , n46077 );
or ( n46080 , n46075 , n46078 , n46079 );
and ( n46081 , n45060 , n39480 );
and ( n46082 , n45073 , n39478 );
nor ( n46083 , n46081 , n46082 );
xnor ( n46084 , n46083 , n39462 );
and ( n46085 , n46080 , n46084 );
xor ( n46086 , n45546 , n45550 );
xor ( n46087 , n46086 , n45553 );
and ( n46088 , n46084 , n46087 );
and ( n46089 , n46080 , n46087 );
or ( n46090 , n46085 , n46088 , n46089 );
and ( n46091 , n45073 , n39480 );
and ( n46092 , n45086 , n39478 );
nor ( n46093 , n46091 , n46092 );
xnor ( n46094 , n46093 , n39462 );
and ( n46095 , n46090 , n46094 );
xor ( n46096 , n45556 , n45560 );
xor ( n46097 , n46096 , n45563 );
and ( n46098 , n46094 , n46097 );
and ( n46099 , n46090 , n46097 );
or ( n46100 , n46095 , n46098 , n46099 );
and ( n46101 , n45086 , n39480 );
and ( n46102 , n45099 , n39478 );
nor ( n46103 , n46101 , n46102 );
xnor ( n46104 , n46103 , n39462 );
and ( n46105 , n46100 , n46104 );
xor ( n46106 , n45566 , n45570 );
xor ( n46107 , n46106 , n45573 );
and ( n46108 , n46104 , n46107 );
and ( n46109 , n46100 , n46107 );
or ( n46110 , n46105 , n46108 , n46109 );
and ( n46111 , n45099 , n39480 );
and ( n46112 , n45112 , n39478 );
nor ( n46113 , n46111 , n46112 );
xnor ( n46114 , n46113 , n39462 );
and ( n46115 , n46110 , n46114 );
xor ( n46116 , n45576 , n45580 );
xor ( n46117 , n46116 , n45583 );
and ( n46118 , n46114 , n46117 );
and ( n46119 , n46110 , n46117 );
or ( n46120 , n46115 , n46118 , n46119 );
and ( n46121 , n45112 , n39480 );
and ( n46122 , n45125 , n39478 );
nor ( n46123 , n46121 , n46122 );
xnor ( n46124 , n46123 , n39462 );
and ( n46125 , n46120 , n46124 );
xor ( n46126 , n45586 , n45590 );
xor ( n46127 , n46126 , n45593 );
and ( n46128 , n46124 , n46127 );
and ( n46129 , n46120 , n46127 );
or ( n46130 , n46125 , n46128 , n46129 );
and ( n46131 , n45125 , n39480 );
and ( n46132 , n45138 , n39478 );
nor ( n46133 , n46131 , n46132 );
xnor ( n46134 , n46133 , n39462 );
and ( n46135 , n46130 , n46134 );
xor ( n46136 , n45596 , n45600 );
xor ( n46137 , n46136 , n45603 );
and ( n46138 , n46134 , n46137 );
and ( n46139 , n46130 , n46137 );
or ( n46140 , n46135 , n46138 , n46139 );
and ( n46141 , n45138 , n39480 );
and ( n46142 , n45151 , n39478 );
nor ( n46143 , n46141 , n46142 );
xnor ( n46144 , n46143 , n39462 );
and ( n46145 , n46140 , n46144 );
xor ( n46146 , n45606 , n45610 );
xor ( n46147 , n46146 , n45613 );
and ( n46148 , n46144 , n46147 );
and ( n46149 , n46140 , n46147 );
or ( n46150 , n46145 , n46148 , n46149 );
and ( n46151 , n45151 , n39480 );
and ( n46152 , n45164 , n39478 );
nor ( n46153 , n46151 , n46152 );
xnor ( n46154 , n46153 , n39462 );
and ( n46155 , n46150 , n46154 );
xor ( n46156 , n45616 , n45620 );
xor ( n46157 , n46156 , n45623 );
and ( n46158 , n46154 , n46157 );
and ( n46159 , n46150 , n46157 );
or ( n46160 , n46155 , n46158 , n46159 );
and ( n46161 , n45164 , n39480 );
and ( n46162 , n44665 , n39478 );
nor ( n46163 , n46161 , n46162 );
xnor ( n46164 , n46163 , n39462 );
and ( n46165 , n46160 , n46164 );
xor ( n46166 , n45626 , n45630 );
xor ( n46167 , n46166 , n45633 );
and ( n46168 , n46164 , n46167 );
and ( n46169 , n46160 , n46167 );
or ( n46170 , n46165 , n46168 , n46169 );
and ( n46171 , n44458 , n39678 );
and ( n46172 , n44357 , n39676 );
nor ( n46173 , n46171 , n46172 );
xnor ( n46174 , n46173 , n39643 );
and ( n46175 , n46170 , n46174 );
and ( n46176 , n44565 , n39539 );
and ( n46177 , n44520 , n39537 );
nor ( n46178 , n46176 , n46177 );
xnor ( n46179 , n46178 , n39522 );
and ( n46180 , n44665 , n39480 );
and ( n46181 , n44656 , n39478 );
nor ( n46182 , n46180 , n46181 );
xnor ( n46183 , n46182 , n39462 );
xor ( n46184 , n46179 , n46183 );
xor ( n46185 , n45636 , n45640 );
xor ( n46186 , n46185 , n45643 );
xor ( n46187 , n46184 , n46186 );
and ( n46188 , n46174 , n46187 );
and ( n46189 , n46170 , n46187 );
or ( n46190 , n46175 , n46188 , n46189 );
and ( n46191 , n44264 , n39760 );
and ( n46192 , n43437 , n39758 );
nor ( n46193 , n46191 , n46192 );
xnor ( n46194 , n46193 , n39742 );
and ( n46195 , n46190 , n46194 );
buf ( n46196 , n557789 );
not ( n46197 , n46196 );
and ( n46198 , n46194 , n46197 );
and ( n46199 , n46190 , n46197 );
or ( n46200 , n46195 , n46198 , n46199 );
and ( n46201 , n43437 , n39760 );
and ( n46202 , n43428 , n39758 );
nor ( n46203 , n46201 , n46202 );
xnor ( n46204 , n46203 , n39742 );
and ( n46205 , n46200 , n46204 );
xor ( n46206 , n45891 , n45895 );
xor ( n46207 , n46206 , n45898 );
and ( n46208 , n46204 , n46207 );
and ( n46209 , n46200 , n46207 );
or ( n46210 , n46205 , n46208 , n46209 );
and ( n46211 , n43192 , n39896 );
and ( n46212 , n43073 , n39894 );
nor ( n46213 , n46211 , n46212 );
xnor ( n46214 , n46213 , n39857 );
and ( n46215 , n46210 , n46214 );
xor ( n46216 , n45676 , n45680 );
xor ( n46217 , n46216 , n45693 );
and ( n46218 , n46214 , n46217 );
and ( n46219 , n46210 , n46217 );
or ( n46220 , n46215 , n46218 , n46219 );
and ( n46221 , n43019 , n40053 );
and ( n46222 , n42811 , n40051 );
nor ( n46223 , n46221 , n46222 );
xnor ( n46224 , n46223 , n39999 );
and ( n46225 , n46220 , n46224 );
xor ( n46226 , n45696 , n45698 );
xor ( n46227 , n46226 , n45701 );
and ( n46228 , n46224 , n46227 );
and ( n46229 , n46220 , n46227 );
or ( n46230 , n46225 , n46228 , n46229 );
and ( n46231 , n42048 , n40258 );
and ( n46232 , n42061 , n40256 );
nor ( n46233 , n46231 , n46232 );
xnor ( n46234 , n46233 , n40169 );
and ( n46235 , n46230 , n46234 );
xor ( n46236 , n45704 , n45708 );
xor ( n46237 , n46236 , n45711 );
and ( n46238 , n46234 , n46237 );
and ( n46239 , n46230 , n46237 );
or ( n46240 , n46235 , n46238 , n46239 );
and ( n46241 , n41692 , n40746 );
and ( n46242 , n41615 , n40744 );
nor ( n46243 , n46241 , n46242 );
xnor ( n46244 , n46243 , n40501 );
and ( n46245 , n41816 , n40527 );
and ( n46246 , n41807 , n40525 );
nor ( n46247 , n46245 , n46246 );
xnor ( n46248 , n46247 , n40382 );
and ( n46249 , n46244 , n46248 );
xor ( n46250 , n45921 , n45925 );
xor ( n46251 , n46250 , n45928 );
and ( n46252 , n46248 , n46251 );
and ( n46253 , n46244 , n46251 );
or ( n46254 , n46249 , n46252 , n46253 );
and ( n46255 , n46240 , n46254 );
and ( n46256 , n41032 , n41055 );
and ( n46257 , n41047 , n41053 );
nor ( n46258 , n46256 , n46257 );
xnor ( n46259 , n46258 , n40728 );
and ( n46260 , n46254 , n46259 );
and ( n46261 , n46240 , n46259 );
or ( n46262 , n46255 , n46260 , n46261 );
and ( n46263 , n40492 , n41622 );
and ( n46264 , n40507 , n41620 );
nor ( n46265 , n46263 , n46264 );
xnor ( n46266 , n46265 , n41194 );
and ( n46267 , n40869 , n41292 );
and ( n46268 , n40738 , n41290 );
nor ( n46269 , n46267 , n46268 );
xnor ( n46270 , n46269 , n41041 );
and ( n46271 , n46266 , n46270 );
xor ( n46272 , n45931 , n45935 );
xor ( n46273 , n46272 , n45938 );
and ( n46274 , n46270 , n46273 );
and ( n46275 , n46266 , n46273 );
or ( n46276 , n46271 , n46274 , n46275 );
and ( n46277 , n46262 , n46276 );
and ( n46278 , n40507 , n41622 );
and ( n46279 , n40373 , n41620 );
nor ( n46280 , n46278 , n46279 );
xnor ( n46281 , n46280 , n41194 );
and ( n46282 , n46276 , n46281 );
and ( n46283 , n46262 , n46281 );
or ( n46284 , n46277 , n46282 , n46283 );
xor ( n46285 , n45953 , n45957 );
xor ( n46286 , n46285 , n45960 );
and ( n46287 , n46284 , n46286 );
xor ( n46288 , n45772 , n45798 );
xor ( n46289 , n46288 , n45801 );
and ( n46290 , n46286 , n46289 );
and ( n46291 , n46284 , n46289 );
or ( n46292 , n46287 , n46290 , n46291 );
and ( n46293 , n46025 , n46292 );
xor ( n46294 , n45804 , n45808 );
xor ( n46295 , n46294 , n45813 );
and ( n46296 , n46292 , n46295 );
and ( n46297 , n46025 , n46295 );
or ( n46298 , n46293 , n46296 , n46297 );
xor ( n46299 , n45816 , n45840 );
xor ( n46300 , n46299 , n45843 );
and ( n46301 , n46298 , n46300 );
xor ( n46302 , n45971 , n45973 );
xor ( n46303 , n46302 , n45976 );
and ( n46304 , n46300 , n46303 );
and ( n46305 , n46298 , n46303 );
or ( n46306 , n46301 , n46304 , n46305 );
xor ( n46307 , n45979 , n45981 );
xor ( n46308 , n46307 , n45984 );
and ( n46309 , n46306 , n46308 );
xor ( n46310 , n46298 , n46300 );
xor ( n46311 , n46310 , n46303 );
and ( n46312 , n46179 , n46183 );
and ( n46313 , n46183 , n46186 );
and ( n46314 , n46179 , n46186 );
or ( n46315 , n46312 , n46313 , n46314 );
and ( n46316 , n44357 , n39678 );
and ( n46317 , n44347 , n39676 );
nor ( n46318 , n46316 , n46317 );
xnor ( n46319 , n46318 , n39643 );
and ( n46320 , n46315 , n46319 );
xor ( n46321 , n45881 , n45885 );
xor ( n46322 , n46321 , n45888 );
and ( n46323 , n46319 , n46322 );
and ( n46324 , n46315 , n46322 );
or ( n46325 , n46320 , n46323 , n46324 );
and ( n46326 , n43200 , n39896 );
and ( n46327 , n43192 , n39894 );
nor ( n46328 , n46326 , n46327 );
xnor ( n46329 , n46328 , n39857 );
and ( n46330 , n46325 , n46329 );
buf ( n46331 , n557788 );
not ( n46332 , n46331 );
and ( n46333 , n46329 , n46332 );
and ( n46334 , n46325 , n46332 );
or ( n46335 , n46330 , n46333 , n46334 );
and ( n46336 , n43027 , n40053 );
and ( n46337 , n43019 , n40051 );
nor ( n46338 , n46336 , n46337 );
xnor ( n46339 , n46338 , n39999 );
and ( n46340 , n46335 , n46339 );
xor ( n46341 , n45901 , n45905 );
xor ( n46342 , n46341 , n45908 );
and ( n46343 , n46339 , n46342 );
and ( n46344 , n46335 , n46342 );
or ( n46345 , n46340 , n46343 , n46344 );
and ( n46346 , n42456 , n40258 );
and ( n46347 , n42048 , n40256 );
nor ( n46348 , n46346 , n46347 );
xnor ( n46349 , n46348 , n40169 );
and ( n46350 , n46345 , n46349 );
xor ( n46351 , n45911 , n45915 );
xor ( n46352 , n46351 , n45918 );
and ( n46353 , n46349 , n46352 );
and ( n46354 , n46345 , n46352 );
or ( n46355 , n46350 , n46353 , n46354 );
and ( n46356 , n41182 , n41055 );
and ( n46357 , n41032 , n41053 );
nor ( n46358 , n46356 , n46357 );
xnor ( n46359 , n46358 , n40728 );
and ( n46360 , n46355 , n46359 );
xor ( n46361 , n46230 , n46234 );
xor ( n46362 , n46361 , n46237 );
and ( n46363 , n46359 , n46362 );
and ( n46364 , n46355 , n46362 );
or ( n46365 , n46360 , n46363 , n46364 );
and ( n46366 , n41807 , n40746 );
and ( n46367 , n41692 , n40744 );
nor ( n46368 , n46366 , n46367 );
xnor ( n46369 , n46368 , n40501 );
and ( n46370 , n42061 , n40527 );
and ( n46371 , n41816 , n40525 );
nor ( n46372 , n46370 , n46371 );
xnor ( n46373 , n46372 , n40382 );
and ( n46374 , n46369 , n46373 );
xor ( n46375 , n46220 , n46224 );
xor ( n46376 , n46375 , n46227 );
and ( n46377 , n46373 , n46376 );
and ( n46378 , n46369 , n46376 );
or ( n46379 , n46374 , n46377 , n46378 );
and ( n46380 , n40738 , n41622 );
and ( n46381 , n40492 , n41620 );
nor ( n46382 , n46380 , n46381 );
xnor ( n46383 , n46382 , n41194 );
and ( n46384 , n46379 , n46383 );
xor ( n46385 , n46244 , n46248 );
xor ( n46386 , n46385 , n46251 );
and ( n46387 , n46383 , n46386 );
and ( n46388 , n46379 , n46386 );
or ( n46389 , n46384 , n46387 , n46388 );
and ( n46390 , n46365 , n46389 );
xor ( n46391 , n45998 , n46002 );
xor ( n46392 , n46391 , n573308 );
and ( n46393 , n46389 , n46392 );
and ( n46394 , n46365 , n46392 );
or ( n46395 , n46390 , n46393 , n46394 );
and ( n46396 , n40197 , n42269 );
and ( n46397 , n40148 , n42266 );
nor ( n46398 , n46396 , n46397 );
xnor ( n46399 , n46398 , n41684 );
and ( n46400 , n46395 , n46399 );
xor ( n46401 , n46262 , n46276 );
xor ( n46402 , n46401 , n46281 );
and ( n46403 , n46399 , n46402 );
and ( n46404 , n46395 , n46402 );
or ( n46405 , n46400 , n46403 , n46404 );
and ( n46406 , n40388 , n41984 );
and ( n46407 , n40186 , n41982 );
nor ( n46408 , n46406 , n46407 );
xnor ( n46409 , n46408 , n41687 );
xor ( n46410 , n45941 , n45945 );
xor ( n46411 , n46410 , n45950 );
and ( n46412 , n46409 , n46411 );
xor ( n46413 , n46005 , n46007 );
xor ( n46414 , n46413 , n46010 );
and ( n46415 , n46411 , n46414 );
and ( n46416 , n46409 , n46414 );
or ( n46417 , n46412 , n46415 , n46416 );
and ( n46418 , n46405 , n46417 );
xor ( n46419 , n46013 , n46017 );
xor ( n46420 , n46419 , n46022 );
and ( n46421 , n46417 , n46420 );
and ( n46422 , n46405 , n46420 );
or ( n46423 , n46418 , n46421 , n46422 );
xor ( n46424 , n46025 , n46292 );
xor ( n46425 , n46424 , n46295 );
and ( n46426 , n46423 , n46425 );
xor ( n46427 , n45963 , n45965 );
xor ( n46428 , n46427 , n45968 );
and ( n46429 , n46425 , n46428 );
and ( n46430 , n46423 , n46428 );
or ( n46431 , n46426 , n46429 , n46430 );
and ( n46432 , n46311 , n46431 );
xor ( n46433 , n46423 , n46425 );
xor ( n46434 , n46433 , n46428 );
and ( n46435 , n40373 , n41984 );
and ( n46436 , n40388 , n41982 );
nor ( n46437 , n46435 , n46436 );
xnor ( n46438 , n46437 , n41687 );
xor ( n46439 , n46240 , n46254 );
xor ( n46440 , n46439 , n46259 );
and ( n46441 , n46438 , n46440 );
xor ( n46442 , n46266 , n46270 );
xor ( n46443 , n46442 , n46273 );
and ( n46444 , n46440 , n46443 );
and ( n46445 , n46438 , n46443 );
or ( n573752 , n46441 , n46444 , n46445 );
and ( n46446 , n44520 , n39678 );
and ( n46447 , n44458 , n39676 );
nor ( n46448 , n46446 , n46447 );
xnor ( n46449 , n46448 , n39643 );
and ( n46450 , n44656 , n39539 );
and ( n46451 , n44565 , n39537 );
nor ( n46452 , n46450 , n46451 );
xnor ( n46453 , n46452 , n39522 );
and ( n46454 , n46449 , n46453 );
xor ( n46455 , n46160 , n46164 );
xor ( n46456 , n46455 , n46167 );
and ( n46457 , n46453 , n46456 );
and ( n46458 , n46449 , n46456 );
or ( n46459 , n46454 , n46457 , n46458 );
and ( n46460 , n44347 , n39760 );
and ( n46461 , n44264 , n39758 );
nor ( n46462 , n46460 , n46461 );
xnor ( n46463 , n46462 , n39742 );
and ( n46464 , n46459 , n46463 );
buf ( n46465 , n557790 );
not ( n46466 , n46465 );
and ( n46467 , n46463 , n46466 );
and ( n46468 , n46459 , n46466 );
or ( n46469 , n46464 , n46467 , n46468 );
and ( n46470 , n43428 , n39896 );
and ( n46471 , n43200 , n39894 );
nor ( n46472 , n46470 , n46471 );
xnor ( n46473 , n46472 , n39857 );
and ( n46474 , n46469 , n46473 );
xor ( n46475 , n46315 , n46319 );
xor ( n46476 , n46475 , n46322 );
and ( n46477 , n46473 , n46476 );
and ( n46478 , n46469 , n46476 );
or ( n46479 , n46474 , n46477 , n46478 );
and ( n46480 , n43073 , n40053 );
and ( n46481 , n43027 , n40051 );
nor ( n46482 , n46480 , n46481 );
xnor ( n46483 , n46482 , n39999 );
and ( n46484 , n46479 , n46483 );
xor ( n46485 , n46325 , n46329 );
xor ( n46486 , n46485 , n46332 );
and ( n46487 , n46483 , n46486 );
and ( n46488 , n46479 , n46486 );
or ( n46489 , n46484 , n46487 , n46488 );
and ( n46490 , n42811 , n40258 );
and ( n46491 , n42456 , n40256 );
nor ( n46492 , n46490 , n46491 );
xnor ( n46493 , n46492 , n40169 );
and ( n46494 , n46489 , n46493 );
xor ( n46495 , n46210 , n46214 );
xor ( n46496 , n46495 , n46217 );
and ( n46497 , n46493 , n46496 );
and ( n46498 , n46489 , n46496 );
or ( n46499 , n46494 , n46497 , n46498 );
and ( n46500 , n41615 , n41055 );
and ( n46501 , n41182 , n41053 );
nor ( n46502 , n46500 , n46501 );
xnor ( n46503 , n46502 , n40728 );
and ( n46504 , n46499 , n46503 );
xor ( n46505 , n46345 , n46349 );
xor ( n46506 , n46505 , n46352 );
and ( n46507 , n46503 , n46506 );
and ( n46508 , n46499 , n46506 );
or ( n46509 , n46504 , n46507 , n46508 );
and ( n46510 , n40507 , n41984 );
and ( n46511 , n40373 , n41982 );
nor ( n46512 , n46510 , n46511 );
xnor ( n46513 , n46512 , n41687 );
and ( n46514 , n46509 , n46513 );
and ( n46515 , n41047 , n41292 );
and ( n46516 , n40869 , n41290 );
nor ( n46517 , n46515 , n46516 );
xnor ( n46518 , n46517 , n41041 );
and ( n46519 , n46513 , n46518 );
and ( n46520 , n46509 , n46518 );
or ( n46521 , n46514 , n46519 , n46520 );
and ( n46522 , n40186 , n42269 );
and ( n46523 , n40197 , n42266 );
nor ( n46524 , n46522 , n46523 );
xnor ( n46525 , n46524 , n41684 );
and ( n46526 , n46521 , n46525 );
xor ( n46527 , n46365 , n46389 );
xor ( n46528 , n46527 , n46392 );
and ( n46529 , n46525 , n46528 );
and ( n46530 , n46521 , n46528 );
or ( n46531 , n46526 , n46529 , n46530 );
and ( n46532 , n573752 , n46531 );
xor ( n46533 , n46409 , n46411 );
xor ( n46534 , n46533 , n46414 );
and ( n46535 , n46531 , n46534 );
and ( n46536 , n573752 , n46534 );
or ( n46537 , n46532 , n46535 , n46536 );
xor ( n46538 , n46405 , n46417 );
xor ( n46539 , n46538 , n46420 );
and ( n46540 , n46537 , n46539 );
xor ( n46541 , n46284 , n46286 );
xor ( n46542 , n46541 , n46289 );
and ( n46543 , n46539 , n46542 );
and ( n46544 , n46537 , n46542 );
or ( n46545 , n46540 , n46543 , n46544 );
and ( n46546 , n46434 , n46545 );
xor ( n46547 , n46537 , n46539 );
xor ( n46548 , n46547 , n46542 );
and ( n46549 , n43192 , n40053 );
and ( n46550 , n43073 , n40051 );
nor ( n46551 , n46549 , n46550 );
xnor ( n46552 , n46551 , n39999 );
xor ( n46553 , n46190 , n46194 );
xor ( n46554 , n46553 , n46197 );
and ( n46555 , n46552 , n46554 );
xor ( n46556 , n46469 , n46473 );
xor ( n46557 , n46556 , n46476 );
and ( n46558 , n46554 , n46557 );
and ( n46559 , n46552 , n46557 );
or ( n46560 , n46555 , n46558 , n46559 );
and ( n46561 , n43019 , n40258 );
and ( n46562 , n42811 , n40256 );
nor ( n46563 , n46561 , n46562 );
xnor ( n46564 , n46563 , n40169 );
and ( n46565 , n46560 , n46564 );
xor ( n46566 , n46200 , n46204 );
xor ( n46567 , n46566 , n46207 );
and ( n46568 , n46564 , n46567 );
and ( n46569 , n46560 , n46567 );
or ( n46570 , n46565 , n46568 , n46569 );
and ( n46571 , n41816 , n40746 );
and ( n46572 , n41807 , n40744 );
nor ( n46573 , n46571 , n46572 );
xnor ( n46574 , n46573 , n40501 );
and ( n46575 , n46570 , n46574 );
xor ( n46576 , n46335 , n46339 );
xor ( n46577 , n46576 , n46342 );
and ( n46578 , n46574 , n46577 );
and ( n46579 , n46570 , n46577 );
or ( n46580 , n46575 , n46578 , n46579 );
and ( n46581 , n41182 , n41292 );
and ( n46582 , n41032 , n41290 );
nor ( n46583 , n46581 , n46582 );
xnor ( n46584 , n46583 , n41041 );
and ( n46585 , n42048 , n40527 );
and ( n46586 , n42061 , n40525 );
nor ( n46587 , n46585 , n46586 );
xnor ( n46588 , n46587 , n40382 );
and ( n46589 , n46584 , n46588 );
xor ( n46590 , n46489 , n46493 );
xor ( n46591 , n46590 , n46496 );
and ( n46592 , n46588 , n46591 );
and ( n46593 , n46584 , n46591 );
or ( n46594 , n46589 , n46592 , n46593 );
and ( n46595 , n46580 , n46594 );
and ( n46596 , n41032 , n41292 );
and ( n46597 , n41047 , n41290 );
nor ( n46598 , n46596 , n46597 );
xnor ( n46599 , n46598 , n41041 );
and ( n46600 , n46594 , n46599 );
and ( n46601 , n46580 , n46599 );
or ( n46602 , n46595 , n46600 , n46601 );
and ( n46603 , n40492 , n41984 );
and ( n46604 , n40507 , n41982 );
nor ( n46605 , n46603 , n46604 );
xnor ( n46606 , n46605 , n41687 );
and ( n46607 , n40869 , n41622 );
and ( n46608 , n40738 , n41620 );
nor ( n46609 , n46607 , n46608 );
xnor ( n46610 , n46609 , n41194 );
and ( n46611 , n46606 , n46610 );
xor ( n46612 , n46369 , n46373 );
xor ( n46613 , n46612 , n46376 );
and ( n46614 , n46610 , n46613 );
and ( n46615 , n46606 , n46613 );
or ( n46616 , n46611 , n46614 , n46615 );
and ( n46617 , n46602 , n46616 );
xor ( n46618 , n46355 , n46359 );
xor ( n46619 , n46618 , n46362 );
and ( n46620 , n46616 , n46619 );
and ( n46621 , n46602 , n46619 );
or ( n46622 , n46617 , n46620 , n46621 );
and ( n46623 , n40388 , n42269 );
and ( n46624 , n40186 , n42266 );
nor ( n46625 , n46623 , n46624 );
xnor ( n46626 , n46625 , n41684 );
xor ( n46627 , n46509 , n46513 );
xor ( n46628 , n46627 , n46518 );
and ( n46629 , n46626 , n46628 );
xor ( n46630 , n46379 , n46383 );
xor ( n46631 , n46630 , n46386 );
and ( n46632 , n46628 , n46631 );
and ( n46633 , n46626 , n46631 );
or ( n46634 , n46629 , n46632 , n46633 );
and ( n46635 , n46622 , n46634 );
xor ( n46636 , n46438 , n46440 );
xor ( n46637 , n46636 , n46443 );
and ( n46638 , n46634 , n46637 );
and ( n46639 , n46622 , n46637 );
or ( n46640 , n46635 , n46638 , n46639 );
xor ( n46641 , n46395 , n46399 );
xor ( n46642 , n46641 , n46402 );
and ( n46643 , n46640 , n46642 );
xor ( n46644 , n573752 , n46531 );
xor ( n46645 , n46644 , n46534 );
and ( n46646 , n46642 , n46645 );
and ( n46647 , n46640 , n46645 );
or ( n46648 , n46643 , n46646 , n46647 );
and ( n46649 , n46548 , n46648 );
xor ( n46650 , n46029 , n46033 );
and ( n46651 , n44991 , n39537 );
not ( n46652 , n46651 );
and ( n46653 , n46652 , n39522 );
and ( n46654 , n44991 , n39539 );
and ( n46655 , n44999 , n39537 );
nor ( n46656 , n46654 , n46655 );
xnor ( n46657 , n46656 , n39522 );
and ( n46658 , n46653 , n46657 );
and ( n46659 , n44999 , n39539 );
and ( n46660 , n45008 , n39537 );
nor ( n46661 , n46659 , n46660 );
xnor ( n46662 , n46661 , n39522 );
and ( n46663 , n46658 , n46662 );
and ( n46664 , n46662 , n46027 );
and ( n46665 , n46658 , n46027 );
or ( n46666 , n46663 , n46664 , n46665 );
and ( n46667 , n46650 , n46666 );
and ( n46668 , n45008 , n39539 );
and ( n46669 , n45021 , n39537 );
nor ( n46670 , n46668 , n46669 );
xnor ( n46671 , n46670 , n39522 );
and ( n46672 , n46666 , n46671 );
and ( n46673 , n46650 , n46671 );
or ( n46674 , n46667 , n46672 , n46673 );
and ( n46675 , n45021 , n39539 );
and ( n46676 , n45034 , n39537 );
nor ( n46677 , n46675 , n46676 );
xnor ( n46678 , n46677 , n39522 );
and ( n46679 , n46674 , n46678 );
xor ( n46680 , n46034 , n46038 );
xor ( n46681 , n46680 , n45513 );
and ( n46682 , n46678 , n46681 );
and ( n46683 , n46674 , n46681 );
or ( n46684 , n46679 , n46682 , n46683 );
and ( n46685 , n45034 , n39539 );
and ( n46686 , n45047 , n39537 );
nor ( n46687 , n46685 , n46686 );
xnor ( n46688 , n46687 , n39522 );
and ( n46689 , n46684 , n46688 );
xor ( n46690 , n46026 , n46042 );
xor ( n46691 , n46690 , n46047 );
and ( n46692 , n46688 , n46691 );
and ( n46693 , n46684 , n46691 );
or ( n46694 , n46689 , n46692 , n46693 );
and ( n46695 , n45047 , n39539 );
and ( n46696 , n45060 , n39537 );
nor ( n46697 , n46695 , n46696 );
xnor ( n46698 , n46697 , n39522 );
and ( n46699 , n46694 , n46698 );
xor ( n46700 , n46050 , n46054 );
xor ( n46701 , n46700 , n46057 );
and ( n46702 , n46698 , n46701 );
and ( n46703 , n46694 , n46701 );
or ( n46704 , n46699 , n46702 , n46703 );
and ( n46705 , n45060 , n39539 );
and ( n46706 , n45073 , n39537 );
nor ( n46707 , n46705 , n46706 );
xnor ( n46708 , n46707 , n39522 );
and ( n46709 , n46704 , n46708 );
xor ( n46710 , n46060 , n46064 );
xor ( n46711 , n46710 , n46067 );
and ( n46712 , n46708 , n46711 );
and ( n46713 , n46704 , n46711 );
or ( n46714 , n46709 , n46712 , n46713 );
and ( n46715 , n45073 , n39539 );
and ( n46716 , n45086 , n39537 );
nor ( n46717 , n46715 , n46716 );
xnor ( n46718 , n46717 , n39522 );
and ( n46719 , n46714 , n46718 );
xor ( n46720 , n46070 , n46074 );
xor ( n46721 , n46720 , n46077 );
and ( n46722 , n46718 , n46721 );
and ( n46723 , n46714 , n46721 );
or ( n46724 , n46719 , n46722 , n46723 );
and ( n46725 , n45086 , n39539 );
and ( n46726 , n45099 , n39537 );
nor ( n46727 , n46725 , n46726 );
xnor ( n46728 , n46727 , n39522 );
and ( n46729 , n46724 , n46728 );
xor ( n46730 , n46080 , n46084 );
xor ( n46731 , n46730 , n46087 );
and ( n46732 , n46728 , n46731 );
and ( n46733 , n46724 , n46731 );
or ( n46734 , n46729 , n46732 , n46733 );
and ( n46735 , n45099 , n39539 );
and ( n46736 , n45112 , n39537 );
nor ( n46737 , n46735 , n46736 );
xnor ( n46738 , n46737 , n39522 );
and ( n46739 , n46734 , n46738 );
xor ( n46740 , n46090 , n46094 );
xor ( n46741 , n46740 , n46097 );
and ( n46742 , n46738 , n46741 );
and ( n46743 , n46734 , n46741 );
or ( n46744 , n46739 , n46742 , n46743 );
and ( n46745 , n45112 , n39539 );
and ( n46746 , n45125 , n39537 );
nor ( n46747 , n46745 , n46746 );
xnor ( n46748 , n46747 , n39522 );
and ( n46749 , n46744 , n46748 );
xor ( n46750 , n46100 , n46104 );
xor ( n46751 , n46750 , n46107 );
and ( n46752 , n46748 , n46751 );
and ( n46753 , n46744 , n46751 );
or ( n46754 , n46749 , n46752 , n46753 );
and ( n46755 , n45125 , n39539 );
and ( n46756 , n45138 , n39537 );
nor ( n46757 , n46755 , n46756 );
xnor ( n46758 , n46757 , n39522 );
and ( n46759 , n46754 , n46758 );
xor ( n46760 , n46110 , n46114 );
xor ( n46761 , n46760 , n46117 );
and ( n46762 , n46758 , n46761 );
and ( n46763 , n46754 , n46761 );
or ( n46764 , n46759 , n46762 , n46763 );
and ( n46765 , n45138 , n39539 );
and ( n46766 , n45151 , n39537 );
nor ( n46767 , n46765 , n46766 );
xnor ( n46768 , n46767 , n39522 );
and ( n46769 , n46764 , n46768 );
xor ( n46770 , n46120 , n46124 );
xor ( n46771 , n46770 , n46127 );
and ( n46772 , n46768 , n46771 );
and ( n46773 , n46764 , n46771 );
or ( n46774 , n46769 , n46772 , n46773 );
and ( n46775 , n45151 , n39539 );
and ( n46776 , n45164 , n39537 );
nor ( n46777 , n46775 , n46776 );
xnor ( n46778 , n46777 , n39522 );
and ( n46779 , n46774 , n46778 );
xor ( n46780 , n46130 , n46134 );
xor ( n46781 , n46780 , n46137 );
and ( n46782 , n46778 , n46781 );
and ( n46783 , n46774 , n46781 );
or ( n46784 , n46779 , n46782 , n46783 );
and ( n46785 , n45164 , n39539 );
and ( n46786 , n44665 , n39537 );
nor ( n46787 , n46785 , n46786 );
xnor ( n46788 , n46787 , n39522 );
and ( n46789 , n46784 , n46788 );
xor ( n46790 , n46140 , n46144 );
xor ( n46791 , n46790 , n46147 );
and ( n46792 , n46788 , n46791 );
and ( n46793 , n46784 , n46791 );
or ( n46794 , n46789 , n46792 , n46793 );
and ( n46795 , n44458 , n39760 );
and ( n46796 , n44357 , n39758 );
nor ( n46797 , n46795 , n46796 );
xnor ( n46798 , n46797 , n39742 );
and ( n46799 , n46794 , n46798 );
and ( n46800 , n44565 , n39678 );
and ( n46801 , n44520 , n39676 );
nor ( n46802 , n46800 , n46801 );
xnor ( n46803 , n46802 , n39643 );
and ( n46804 , n44665 , n39539 );
and ( n46805 , n44656 , n39537 );
nor ( n46806 , n46804 , n46805 );
xnor ( n46807 , n46806 , n39522 );
xor ( n46808 , n46803 , n46807 );
xor ( n46809 , n46150 , n46154 );
xor ( n46810 , n46809 , n46157 );
xor ( n46811 , n46808 , n46810 );
and ( n46812 , n46798 , n46811 );
and ( n46813 , n46794 , n46811 );
or ( n46814 , n46799 , n46812 , n46813 );
and ( n46815 , n44264 , n39896 );
and ( n46816 , n43437 , n39894 );
nor ( n46817 , n46815 , n46816 );
xnor ( n46818 , n46817 , n39857 );
and ( n46819 , n46814 , n46818 );
xor ( n46820 , n46449 , n46453 );
xor ( n46821 , n46820 , n46456 );
and ( n46822 , n46818 , n46821 );
and ( n46823 , n46814 , n46821 );
or ( n46824 , n46819 , n46822 , n46823 );
and ( n46825 , n43437 , n39896 );
and ( n46826 , n43428 , n39894 );
nor ( n46827 , n46825 , n46826 );
xnor ( n46828 , n46827 , n39857 );
and ( n46829 , n46824 , n46828 );
xor ( n46830 , n46459 , n46463 );
xor ( n46831 , n46830 , n46466 );
and ( n46832 , n46828 , n46831 );
and ( n46833 , n46824 , n46831 );
or ( n46834 , n46829 , n46832 , n46833 );
and ( n46835 , n46803 , n46807 );
and ( n46836 , n46807 , n46810 );
and ( n46837 , n46803 , n46810 );
or ( n46838 , n46835 , n46836 , n46837 );
and ( n46839 , n44357 , n39760 );
and ( n46840 , n44347 , n39758 );
nor ( n46841 , n46839 , n46840 );
xnor ( n46842 , n46841 , n39742 );
and ( n46843 , n46838 , n46842 );
buf ( n46844 , n557791 );
not ( n46845 , n46844 );
and ( n46846 , n46842 , n46845 );
and ( n46847 , n46838 , n46845 );
or ( n46848 , n46843 , n46846 , n46847 );
and ( n46849 , n43200 , n40053 );
and ( n46850 , n43192 , n40051 );
nor ( n46851 , n46849 , n46850 );
xnor ( n46852 , n46851 , n39999 );
and ( n46853 , n46848 , n46852 );
xor ( n46854 , n46170 , n46174 );
xor ( n46855 , n46854 , n46187 );
and ( n46856 , n46852 , n46855 );
and ( n46857 , n46848 , n46855 );
or ( n46858 , n46853 , n46856 , n46857 );
and ( n46859 , n46834 , n46858 );
and ( n46860 , n43027 , n40258 );
and ( n46861 , n43019 , n40256 );
nor ( n46862 , n46860 , n46861 );
xnor ( n46863 , n46862 , n40169 );
and ( n46864 , n46858 , n46863 );
and ( n46865 , n46834 , n46863 );
or ( n46866 , n46859 , n46864 , n46865 );
and ( n46867 , n42456 , n40527 );
and ( n46868 , n42048 , n40525 );
nor ( n46869 , n46867 , n46868 );
xnor ( n46870 , n46869 , n40382 );
and ( n46871 , n46866 , n46870 );
xor ( n46872 , n46479 , n46483 );
xor ( n46873 , n46872 , n46486 );
and ( n46874 , n46870 , n46873 );
and ( n46875 , n46866 , n46873 );
or ( n46876 , n46871 , n46874 , n46875 );
and ( n46877 , n41692 , n41055 );
and ( n46878 , n41615 , n41053 );
nor ( n46879 , n46877 , n46878 );
xnor ( n46880 , n46879 , n40728 );
and ( n46881 , n46876 , n46880 );
xor ( n46882 , n46570 , n46574 );
xor ( n46883 , n46882 , n46577 );
and ( n46884 , n46880 , n46883 );
and ( n46885 , n46876 , n46883 );
or ( n46886 , n46881 , n46884 , n46885 );
and ( n46887 , n41807 , n41055 );
and ( n46888 , n41692 , n41053 );
nor ( n46889 , n46887 , n46888 );
xnor ( n46890 , n46889 , n40728 );
and ( n46891 , n42061 , n40746 );
and ( n46892 , n41816 , n40744 );
nor ( n46893 , n46891 , n46892 );
xnor ( n46894 , n46893 , n40501 );
and ( n46895 , n46890 , n46894 );
xor ( n46896 , n46560 , n46564 );
xor ( n46897 , n46896 , n46567 );
and ( n46898 , n46894 , n46897 );
and ( n46899 , n46890 , n46897 );
or ( n46900 , n46895 , n46898 , n46899 );
and ( n46901 , n41047 , n41622 );
and ( n46902 , n40869 , n41620 );
nor ( n46903 , n46901 , n46902 );
xnor ( n46904 , n46903 , n41194 );
and ( n46905 , n46900 , n46904 );
xor ( n46906 , n46584 , n46588 );
xor ( n46907 , n46906 , n46591 );
and ( n46908 , n46904 , n46907 );
and ( n46909 , n46900 , n46907 );
or ( n46910 , n46905 , n46908 , n46909 );
and ( n46911 , n46886 , n46910 );
xor ( n46912 , n46499 , n46503 );
xor ( n46913 , n46912 , n46506 );
and ( n46914 , n46910 , n46913 );
and ( n46915 , n46886 , n46913 );
or ( n46916 , n46911 , n46914 , n46915 );
and ( n46917 , n40373 , n42269 );
and ( n46918 , n40388 , n42266 );
nor ( n46919 , n46917 , n46918 );
xnor ( n46920 , n46919 , n41684 );
xor ( n46921 , n46580 , n46594 );
xor ( n46922 , n46921 , n46599 );
and ( n46923 , n46920 , n46922 );
xor ( n46924 , n46606 , n46610 );
xor ( n46925 , n46924 , n46613 );
and ( n46926 , n46922 , n46925 );
and ( n46927 , n46920 , n46925 );
or ( n46928 , n46923 , n46926 , n46927 );
and ( n46929 , n46916 , n46928 );
xor ( n46930 , n46602 , n46616 );
xor ( n46931 , n46930 , n46619 );
and ( n46932 , n46928 , n46931 );
and ( n46933 , n46916 , n46931 );
or ( n46934 , n46929 , n46932 , n46933 );
xor ( n46935 , n46622 , n46634 );
xor ( n46936 , n46935 , n46637 );
and ( n46937 , n46934 , n46936 );
xor ( n46938 , n46521 , n46525 );
xor ( n46939 , n46938 , n46528 );
and ( n46940 , n46936 , n46939 );
and ( n46941 , n46934 , n46939 );
or ( n46942 , n46937 , n46940 , n46941 );
xor ( n46943 , n46640 , n46642 );
xor ( n46944 , n46943 , n46645 );
and ( n46945 , n46942 , n46944 );
xor ( n46946 , n46934 , n46936 );
xor ( n46947 , n46946 , n46939 );
and ( n46948 , n44520 , n39760 );
and ( n46949 , n44458 , n39758 );
nor ( n46950 , n46948 , n46949 );
xnor ( n46951 , n46950 , n39742 );
and ( n46952 , n44656 , n39678 );
and ( n46953 , n44565 , n39676 );
nor ( n46954 , n46952 , n46953 );
xnor ( n46955 , n46954 , n39643 );
and ( n46956 , n46951 , n46955 );
xor ( n46957 , n46784 , n46788 );
xor ( n46958 , n46957 , n46791 );
and ( n46959 , n46955 , n46958 );
and ( n46960 , n46951 , n46958 );
or ( n46961 , n46956 , n46959 , n46960 );
and ( n46962 , n44347 , n39896 );
and ( n46963 , n44264 , n39894 );
nor ( n46964 , n46962 , n46963 );
xnor ( n46965 , n46964 , n39857 );
and ( n46966 , n46961 , n46965 );
buf ( n46967 , n557792 );
not ( n46968 , n46967 );
and ( n46969 , n46965 , n46968 );
and ( n46970 , n46961 , n46968 );
or ( n46971 , n46966 , n46969 , n46970 );
and ( n46972 , n43428 , n40053 );
and ( n46973 , n43200 , n40051 );
nor ( n46974 , n46972 , n46973 );
xnor ( n46975 , n46974 , n39999 );
and ( n46976 , n46971 , n46975 );
xor ( n46977 , n46838 , n46842 );
xor ( n46978 , n46977 , n46845 );
and ( n46979 , n46975 , n46978 );
and ( n46980 , n46971 , n46978 );
or ( n46981 , n46976 , n46979 , n46980 );
and ( n46982 , n43073 , n40258 );
and ( n46983 , n43027 , n40256 );
nor ( n46984 , n46982 , n46983 );
xnor ( n46985 , n46984 , n40169 );
and ( n46986 , n46981 , n46985 );
xor ( n46987 , n46848 , n46852 );
xor ( n46988 , n46987 , n46855 );
and ( n46989 , n46985 , n46988 );
and ( n46990 , n46981 , n46988 );
or ( n46991 , n46986 , n46989 , n46990 );
and ( n46992 , n42811 , n40527 );
and ( n46993 , n42456 , n40525 );
nor ( n46994 , n46992 , n46993 );
xnor ( n46995 , n46994 , n40382 );
and ( n46996 , n46991 , n46995 );
xor ( n46997 , n46552 , n46554 );
xor ( n46998 , n46997 , n46557 );
and ( n46999 , n46995 , n46998 );
and ( n47000 , n46991 , n46998 );
or ( n47001 , n46996 , n46999 , n47000 );
and ( n47002 , n41615 , n41292 );
and ( n47003 , n41182 , n41290 );
nor ( n47004 , n47002 , n47003 );
xnor ( n47005 , n47004 , n41041 );
and ( n47006 , n47001 , n47005 );
xor ( n47007 , n46866 , n46870 );
xor ( n47008 , n47007 , n46873 );
and ( n47009 , n47005 , n47008 );
and ( n47010 , n47001 , n47008 );
or ( n47011 , n47006 , n47009 , n47010 );
and ( n47012 , n40507 , n42269 );
and ( n47013 , n40373 , n42266 );
nor ( n47014 , n47012 , n47013 );
xnor ( n47015 , n47014 , n41684 );
and ( n47016 , n47011 , n47015 );
and ( n47017 , n40738 , n41984 );
and ( n47018 , n40492 , n41982 );
nor ( n47019 , n47017 , n47018 );
xnor ( n47020 , n47019 , n41687 );
and ( n47021 , n47015 , n47020 );
and ( n47022 , n47011 , n47020 );
or ( n47023 , n47016 , n47021 , n47022 );
and ( n47024 , n43192 , n40258 );
and ( n47025 , n43073 , n40256 );
nor ( n47026 , n47024 , n47025 );
xnor ( n47027 , n47026 , n40169 );
xor ( n47028 , n46971 , n46975 );
xor ( n47029 , n47028 , n46978 );
and ( n47030 , n47027 , n47029 );
xor ( n47031 , n46814 , n46818 );
xor ( n47032 , n47031 , n46821 );
and ( n47033 , n47029 , n47032 );
and ( n47034 , n47027 , n47032 );
or ( n47035 , n47030 , n47033 , n47034 );
and ( n47036 , n43019 , n40527 );
and ( n47037 , n42811 , n40525 );
nor ( n47038 , n47036 , n47037 );
xnor ( n47039 , n47038 , n40382 );
and ( n47040 , n47035 , n47039 );
xor ( n47041 , n46824 , n46828 );
xor ( n47042 , n47041 , n46831 );
and ( n47043 , n47039 , n47042 );
and ( n47044 , n47035 , n47042 );
or ( n47045 , n47040 , n47043 , n47044 );
and ( n47046 , n41816 , n41055 );
and ( n47047 , n41807 , n41053 );
nor ( n47048 , n47046 , n47047 );
xnor ( n47049 , n47048 , n40728 );
and ( n47050 , n47045 , n47049 );
xor ( n47051 , n46834 , n46858 );
xor ( n47052 , n47051 , n46863 );
and ( n47053 , n47049 , n47052 );
and ( n47054 , n47045 , n47052 );
or ( n47055 , n47050 , n47053 , n47054 );
and ( n47056 , n41182 , n41622 );
and ( n47057 , n41032 , n41620 );
nor ( n47058 , n47056 , n47057 );
xnor ( n47059 , n47058 , n41194 );
and ( n47060 , n42048 , n40746 );
and ( n47061 , n42061 , n40744 );
nor ( n47062 , n47060 , n47061 );
xnor ( n47063 , n47062 , n40501 );
and ( n47064 , n47059 , n47063 );
xor ( n47065 , n46991 , n46995 );
xor ( n47066 , n47065 , n46998 );
and ( n47067 , n47063 , n47066 );
and ( n47068 , n47059 , n47066 );
or ( n47069 , n47064 , n47067 , n47068 );
and ( n47070 , n47055 , n47069 );
and ( n47071 , n41032 , n41622 );
and ( n47072 , n41047 , n41620 );
nor ( n47073 , n47071 , n47072 );
xnor ( n47074 , n47073 , n41194 );
and ( n47075 , n47069 , n47074 );
and ( n47076 , n47055 , n47074 );
or ( n47077 , n47070 , n47075 , n47076 );
and ( n47078 , n40869 , n41984 );
and ( n47079 , n40738 , n41982 );
nor ( n47080 , n47078 , n47079 );
xnor ( n47081 , n47080 , n41687 );
xor ( n47082 , n47001 , n47005 );
xor ( n47083 , n47082 , n47008 );
and ( n47084 , n47081 , n47083 );
xor ( n47085 , n46890 , n46894 );
xor ( n47086 , n47085 , n46897 );
and ( n47087 , n47083 , n47086 );
and ( n47088 , n47081 , n47086 );
or ( n47089 , n47084 , n47087 , n47088 );
and ( n47090 , n47077 , n47089 );
xor ( n47091 , n46876 , n46880 );
xor ( n47092 , n47091 , n46883 );
and ( n47093 , n47089 , n47092 );
and ( n47094 , n47077 , n47092 );
or ( n47095 , n47090 , n47093 , n47094 );
and ( n47096 , n47023 , n47095 );
xor ( n47097 , n46886 , n46910 );
xor ( n47098 , n47097 , n46913 );
and ( n47099 , n47095 , n47098 );
and ( n47100 , n47023 , n47098 );
or ( n47101 , n47096 , n47099 , n47100 );
xor ( n47102 , n46916 , n46928 );
xor ( n47103 , n47102 , n46931 );
and ( n47104 , n47101 , n47103 );
xor ( n47105 , n46626 , n46628 );
xor ( n47106 , n47105 , n46631 );
and ( n47107 , n47103 , n47106 );
and ( n47108 , n47101 , n47106 );
or ( n47109 , n47104 , n47107 , n47108 );
and ( n47110 , n46947 , n47109 );
xor ( n47111 , n47101 , n47103 );
xor ( n47112 , n47111 , n47106 );
xor ( n47113 , n46653 , n46657 );
and ( n47114 , n44991 , n39676 );
not ( n47115 , n47114 );
and ( n47116 , n47115 , n39643 );
and ( n47117 , n44991 , n39678 );
and ( n47118 , n44999 , n39676 );
nor ( n47119 , n47117 , n47118 );
xnor ( n47120 , n47119 , n39643 );
and ( n47121 , n47116 , n47120 );
and ( n47122 , n44999 , n39678 );
and ( n47123 , n45008 , n39676 );
nor ( n47124 , n47122 , n47123 );
xnor ( n47125 , n47124 , n39643 );
and ( n47126 , n47121 , n47125 );
and ( n47127 , n47125 , n46651 );
and ( n47128 , n47121 , n46651 );
or ( n47129 , n47126 , n47127 , n47128 );
and ( n47130 , n47113 , n47129 );
and ( n47131 , n45008 , n39678 );
and ( n47132 , n45021 , n39676 );
nor ( n47133 , n47131 , n47132 );
xnor ( n47134 , n47133 , n39643 );
and ( n47135 , n47129 , n47134 );
and ( n47136 , n47113 , n47134 );
or ( n47137 , n47130 , n47135 , n47136 );
and ( n47138 , n45021 , n39678 );
and ( n47139 , n45034 , n39676 );
nor ( n47140 , n47138 , n47139 );
xnor ( n47141 , n47140 , n39643 );
and ( n47142 , n47137 , n47141 );
xor ( n47143 , n46658 , n46662 );
xor ( n47144 , n47143 , n46027 );
and ( n47145 , n47141 , n47144 );
and ( n47146 , n47137 , n47144 );
or ( n47147 , n47142 , n47145 , n47146 );
and ( n47148 , n45034 , n39678 );
and ( n47149 , n45047 , n39676 );
nor ( n47150 , n47148 , n47149 );
xnor ( n47151 , n47150 , n39643 );
and ( n47152 , n47147 , n47151 );
xor ( n47153 , n46650 , n46666 );
xor ( n47154 , n47153 , n46671 );
and ( n47155 , n47151 , n47154 );
and ( n47156 , n47147 , n47154 );
or ( n47157 , n47152 , n47155 , n47156 );
and ( n47158 , n45047 , n39678 );
and ( n47159 , n45060 , n39676 );
nor ( n47160 , n47158 , n47159 );
xnor ( n47161 , n47160 , n39643 );
and ( n47162 , n47157 , n47161 );
xor ( n47163 , n46674 , n46678 );
xor ( n47164 , n47163 , n46681 );
and ( n47165 , n47161 , n47164 );
and ( n47166 , n47157 , n47164 );
or ( n47167 , n47162 , n47165 , n47166 );
and ( n47168 , n45060 , n39678 );
and ( n47169 , n45073 , n39676 );
nor ( n47170 , n47168 , n47169 );
xnor ( n47171 , n47170 , n39643 );
and ( n47172 , n47167 , n47171 );
xor ( n47173 , n46684 , n46688 );
xor ( n47174 , n47173 , n46691 );
and ( n47175 , n47171 , n47174 );
and ( n47176 , n47167 , n47174 );
or ( n47177 , n47172 , n47175 , n47176 );
and ( n47178 , n45073 , n39678 );
and ( n47179 , n45086 , n39676 );
nor ( n47180 , n47178 , n47179 );
xnor ( n47181 , n47180 , n39643 );
and ( n47182 , n47177 , n47181 );
xor ( n47183 , n46694 , n46698 );
xor ( n47184 , n47183 , n46701 );
and ( n47185 , n47181 , n47184 );
and ( n47186 , n47177 , n47184 );
or ( n47187 , n47182 , n47185 , n47186 );
and ( n47188 , n45086 , n39678 );
and ( n47189 , n45099 , n39676 );
nor ( n47190 , n47188 , n47189 );
xnor ( n47191 , n47190 , n39643 );
and ( n47192 , n47187 , n47191 );
xor ( n47193 , n46704 , n46708 );
xor ( n47194 , n47193 , n46711 );
and ( n47195 , n47191 , n47194 );
and ( n47196 , n47187 , n47194 );
or ( n47197 , n47192 , n47195 , n47196 );
and ( n47198 , n45099 , n39678 );
and ( n47199 , n45112 , n39676 );
nor ( n47200 , n47198 , n47199 );
xnor ( n47201 , n47200 , n39643 );
and ( n47202 , n47197 , n47201 );
xor ( n47203 , n46714 , n46718 );
xor ( n47204 , n47203 , n46721 );
and ( n47205 , n47201 , n47204 );
and ( n47206 , n47197 , n47204 );
or ( n47207 , n47202 , n47205 , n47206 );
and ( n47208 , n45112 , n39678 );
and ( n47209 , n45125 , n39676 );
nor ( n47210 , n47208 , n47209 );
xnor ( n47211 , n47210 , n39643 );
and ( n47212 , n47207 , n47211 );
xor ( n47213 , n46724 , n46728 );
xor ( n47214 , n47213 , n46731 );
and ( n47215 , n47211 , n47214 );
and ( n47216 , n47207 , n47214 );
or ( n47217 , n47212 , n47215 , n47216 );
and ( n47218 , n45125 , n39678 );
and ( n47219 , n45138 , n39676 );
nor ( n47220 , n47218 , n47219 );
xnor ( n47221 , n47220 , n39643 );
and ( n47222 , n47217 , n47221 );
xor ( n47223 , n46734 , n46738 );
xor ( n47224 , n47223 , n46741 );
and ( n47225 , n47221 , n47224 );
and ( n47226 , n47217 , n47224 );
or ( n47227 , n47222 , n47225 , n47226 );
and ( n47228 , n45138 , n39678 );
and ( n47229 , n45151 , n39676 );
nor ( n47230 , n47228 , n47229 );
xnor ( n47231 , n47230 , n39643 );
and ( n47232 , n47227 , n47231 );
xor ( n47233 , n46744 , n46748 );
xor ( n47234 , n47233 , n46751 );
and ( n47235 , n47231 , n47234 );
and ( n47236 , n47227 , n47234 );
or ( n47237 , n47232 , n47235 , n47236 );
and ( n47238 , n45151 , n39678 );
and ( n47239 , n45164 , n39676 );
nor ( n47240 , n47238 , n47239 );
xnor ( n47241 , n47240 , n39643 );
and ( n47242 , n47237 , n47241 );
xor ( n47243 , n46754 , n46758 );
xor ( n47244 , n47243 , n46761 );
and ( n47245 , n47241 , n47244 );
and ( n47246 , n47237 , n47244 );
or ( n47247 , n47242 , n47245 , n47246 );
and ( n47248 , n45164 , n39678 );
and ( n47249 , n44665 , n39676 );
nor ( n47250 , n47248 , n47249 );
xnor ( n47251 , n47250 , n39643 );
and ( n47252 , n47247 , n47251 );
xor ( n47253 , n46764 , n46768 );
xor ( n47254 , n47253 , n46771 );
and ( n47255 , n47251 , n47254 );
and ( n47256 , n47247 , n47254 );
or ( n47257 , n47252 , n47255 , n47256 );
and ( n47258 , n44458 , n39896 );
and ( n47259 , n44357 , n39894 );
nor ( n47260 , n47258 , n47259 );
xnor ( n47261 , n47260 , n39857 );
and ( n47262 , n47257 , n47261 );
buf ( n47263 , n557794 );
not ( n47264 , n47263 );
and ( n47265 , n47261 , n47264 );
and ( n47266 , n47257 , n47264 );
or ( n47267 , n47262 , n47265 , n47266 );
and ( n47268 , n44264 , n40053 );
and ( n47269 , n43437 , n40051 );
nor ( n47270 , n47268 , n47269 );
xnor ( n47271 , n47270 , n39999 );
and ( n47272 , n47267 , n47271 );
xor ( n47273 , n46951 , n46955 );
xor ( n47274 , n47273 , n46958 );
and ( n47275 , n47271 , n47274 );
and ( n47276 , n47267 , n47274 );
or ( n47277 , n47272 , n47275 , n47276 );
and ( n47278 , n43437 , n40053 );
and ( n47279 , n43428 , n40051 );
nor ( n47280 , n47278 , n47279 );
xnor ( n47281 , n47280 , n39999 );
and ( n47282 , n47277 , n47281 );
xor ( n47283 , n46961 , n46965 );
xor ( n47284 , n47283 , n46968 );
and ( n47285 , n47281 , n47284 );
and ( n47286 , n47277 , n47284 );
or ( n47287 , n47282 , n47285 , n47286 );
and ( n47288 , n44565 , n39760 );
and ( n47289 , n44520 , n39758 );
nor ( n47290 , n47288 , n47289 );
xnor ( n47291 , n47290 , n39742 );
and ( n47292 , n44665 , n39678 );
and ( n47293 , n44656 , n39676 );
nor ( n47294 , n47292 , n47293 );
xnor ( n47295 , n47294 , n39643 );
and ( n47296 , n47291 , n47295 );
xor ( n47297 , n46774 , n46778 );
xor ( n47298 , n47297 , n46781 );
and ( n47299 , n47295 , n47298 );
and ( n47300 , n47291 , n47298 );
or ( n47301 , n47296 , n47299 , n47300 );
and ( n47302 , n44357 , n39896 );
and ( n47303 , n44347 , n39894 );
nor ( n47304 , n47302 , n47303 );
xnor ( n47305 , n47304 , n39857 );
and ( n47306 , n47301 , n47305 );
buf ( n47307 , n557793 );
not ( n47308 , n47307 );
and ( n47309 , n47305 , n47308 );
and ( n47310 , n47301 , n47308 );
or ( n47311 , n47306 , n47309 , n47310 );
and ( n47312 , n43200 , n40258 );
and ( n47313 , n43192 , n40256 );
nor ( n47314 , n47312 , n47313 );
xnor ( n47315 , n47314 , n40169 );
and ( n47316 , n47311 , n47315 );
xor ( n47317 , n46794 , n46798 );
xor ( n47318 , n47317 , n46811 );
and ( n47319 , n47315 , n47318 );
and ( n47320 , n47311 , n47318 );
or ( n47321 , n47316 , n47319 , n47320 );
and ( n47322 , n47287 , n47321 );
and ( n47323 , n43027 , n40527 );
and ( n47324 , n43019 , n40525 );
nor ( n47325 , n47323 , n47324 );
xnor ( n47326 , n47325 , n40382 );
and ( n47327 , n47321 , n47326 );
and ( n47328 , n47287 , n47326 );
or ( n47329 , n47322 , n47327 , n47328 );
xor ( n47330 , n47035 , n47039 );
xor ( n47331 , n47330 , n47042 );
and ( n47332 , n47329 , n47331 );
xor ( n47333 , n46981 , n46985 );
xor ( n47334 , n47333 , n46988 );
and ( n47335 , n47331 , n47334 );
and ( n47336 , n47329 , n47334 );
or ( n47337 , n47332 , n47335 , n47336 );
and ( n47338 , n41692 , n41292 );
and ( n47339 , n41615 , n41290 );
nor ( n47340 , n47338 , n47339 );
xnor ( n47341 , n47340 , n41041 );
and ( n47342 , n47337 , n47341 );
xor ( n47343 , n47045 , n47049 );
xor ( n47344 , n47343 , n47052 );
and ( n47345 , n47341 , n47344 );
and ( n47346 , n47337 , n47344 );
or ( n47347 , n47342 , n47345 , n47346 );
and ( n47348 , n41807 , n41292 );
and ( n47349 , n41692 , n41290 );
nor ( n47350 , n47348 , n47349 );
xnor ( n47351 , n47350 , n41041 );
and ( n47352 , n42061 , n41055 );
and ( n47353 , n41816 , n41053 );
nor ( n47354 , n47352 , n47353 );
xnor ( n47355 , n47354 , n40728 );
and ( n47356 , n47351 , n47355 );
and ( n47357 , n42456 , n40746 );
and ( n47358 , n42048 , n40744 );
nor ( n47359 , n47357 , n47358 );
xnor ( n47360 , n47359 , n40501 );
and ( n47361 , n47355 , n47360 );
and ( n47362 , n47351 , n47360 );
or ( n47363 , n47356 , n47361 , n47362 );
and ( n47364 , n40738 , n42269 );
and ( n47365 , n40492 , n42266 );
nor ( n47366 , n47364 , n47365 );
xnor ( n47367 , n47366 , n41684 );
and ( n47368 , n47363 , n47367 );
xor ( n47369 , n47059 , n47063 );
xor ( n47370 , n47369 , n47066 );
and ( n47371 , n47367 , n47370 );
and ( n47372 , n47363 , n47370 );
or ( n47373 , n47368 , n47371 , n47372 );
and ( n47374 , n47347 , n47373 );
and ( n47375 , n40492 , n42269 );
and ( n47376 , n40507 , n42266 );
nor ( n47377 , n47375 , n47376 );
xnor ( n47378 , n47377 , n41684 );
and ( n47379 , n47373 , n47378 );
and ( n47380 , n47347 , n47378 );
or ( n47381 , n47374 , n47379 , n47380 );
xor ( n47382 , n47011 , n47015 );
xor ( n47383 , n47382 , n47020 );
and ( n47384 , n47381 , n47383 );
xor ( n47385 , n46900 , n46904 );
xor ( n47386 , n47385 , n46907 );
and ( n47387 , n47383 , n47386 );
and ( n47388 , n47381 , n47386 );
or ( n47389 , n47384 , n47387 , n47388 );
xor ( n47390 , n47023 , n47095 );
xor ( n47391 , n47390 , n47098 );
and ( n47392 , n47389 , n47391 );
xor ( n47393 , n46920 , n46922 );
xor ( n47394 , n47393 , n46925 );
and ( n47395 , n47391 , n47394 );
and ( n47396 , n47389 , n47394 );
or ( n47397 , n47392 , n47395 , n47396 );
and ( n47398 , n47112 , n47397 );
xor ( n47399 , n47389 , n47391 );
xor ( n47400 , n47399 , n47394 );
and ( n47401 , n44520 , n39896 );
and ( n47402 , n44458 , n39894 );
nor ( n47403 , n47401 , n47402 );
xnor ( n47404 , n47403 , n39857 );
and ( n47405 , n44656 , n39760 );
and ( n47406 , n44565 , n39758 );
nor ( n47407 , n47405 , n47406 );
xnor ( n47408 , n47407 , n39742 );
and ( n47409 , n47404 , n47408 );
buf ( n47410 , n557795 );
not ( n47411 , n47410 );
and ( n47412 , n47408 , n47411 );
and ( n47413 , n47404 , n47411 );
or ( n47414 , n47409 , n47412 , n47413 );
and ( n47415 , n44347 , n40053 );
and ( n47416 , n44264 , n40051 );
nor ( n47417 , n47415 , n47416 );
xnor ( n47418 , n47417 , n39999 );
and ( n47419 , n47414 , n47418 );
xor ( n47420 , n47291 , n47295 );
xor ( n47421 , n47420 , n47298 );
and ( n47422 , n47418 , n47421 );
and ( n47423 , n47414 , n47421 );
or ( n47424 , n47419 , n47422 , n47423 );
and ( n47425 , n43428 , n40258 );
and ( n47426 , n43200 , n40256 );
nor ( n47427 , n47425 , n47426 );
xnor ( n47428 , n47427 , n40169 );
and ( n47429 , n47424 , n47428 );
xor ( n47430 , n47301 , n47305 );
xor ( n47431 , n47430 , n47308 );
and ( n47432 , n47428 , n47431 );
and ( n47433 , n47424 , n47431 );
or ( n47434 , n47429 , n47432 , n47433 );
and ( n47435 , n43073 , n40527 );
and ( n47436 , n43027 , n40525 );
nor ( n47437 , n47435 , n47436 );
xnor ( n47438 , n47437 , n40382 );
and ( n47439 , n47434 , n47438 );
xor ( n47440 , n47311 , n47315 );
xor ( n47441 , n47440 , n47318 );
and ( n47442 , n47438 , n47441 );
and ( n47443 , n47434 , n47441 );
or ( n47444 , n47439 , n47442 , n47443 );
and ( n47445 , n42811 , n40746 );
and ( n47446 , n42456 , n40744 );
nor ( n47447 , n47445 , n47446 );
xnor ( n47448 , n47447 , n40501 );
and ( n47449 , n47444 , n47448 );
xor ( n47450 , n47027 , n47029 );
xor ( n47451 , n47450 , n47032 );
and ( n47452 , n47448 , n47451 );
and ( n47453 , n47444 , n47451 );
or ( n47454 , n47449 , n47452 , n47453 );
and ( n47455 , n41615 , n41622 );
and ( n47456 , n41182 , n41620 );
nor ( n47457 , n47455 , n47456 );
xnor ( n47458 , n47457 , n41194 );
and ( n47459 , n47454 , n47458 );
xor ( n47460 , n47329 , n47331 );
xor ( n47461 , n47460 , n47334 );
and ( n47462 , n47458 , n47461 );
and ( n47463 , n47454 , n47461 );
or ( n47464 , n47459 , n47462 , n47463 );
and ( n47465 , n41047 , n41984 );
and ( n47466 , n40869 , n41982 );
nor ( n47467 , n47465 , n47466 );
xnor ( n47468 , n47467 , n41687 );
and ( n47469 , n47464 , n47468 );
xor ( n47470 , n47337 , n47341 );
xor ( n47471 , n47470 , n47344 );
and ( n47472 , n47468 , n47471 );
and ( n47473 , n47464 , n47471 );
or ( n47474 , n47469 , n47472 , n47473 );
xor ( n47475 , n47055 , n47069 );
xor ( n47476 , n47475 , n47074 );
and ( n47477 , n47474 , n47476 );
xor ( n47478 , n47081 , n47083 );
xor ( n47479 , n47478 , n47086 );
and ( n47480 , n47476 , n47479 );
and ( n47481 , n47474 , n47479 );
or ( n47482 , n47477 , n47480 , n47481 );
xor ( n47483 , n47077 , n47089 );
xor ( n47484 , n47483 , n47092 );
and ( n47485 , n47482 , n47484 );
xor ( n47486 , n47381 , n47383 );
xor ( n47487 , n47486 , n47386 );
and ( n47488 , n47484 , n47487 );
and ( n47489 , n47482 , n47487 );
or ( n47490 , n47485 , n47488 , n47489 );
and ( n47491 , n47400 , n47490 );
xor ( n47492 , n47482 , n47484 );
xor ( n47493 , n47492 , n47487 );
and ( n47494 , n41692 , n41622 );
and ( n47495 , n41615 , n41620 );
nor ( n47496 , n47494 , n47495 );
xnor ( n47497 , n47496 , n41194 );
and ( n47498 , n41816 , n41292 );
and ( n47499 , n41807 , n41290 );
nor ( n47500 , n47498 , n47499 );
xnor ( n47501 , n47500 , n41041 );
and ( n47502 , n47497 , n47501 );
and ( n47503 , n42048 , n41055 );
and ( n47504 , n42061 , n41053 );
nor ( n47505 , n47503 , n47504 );
xnor ( n47506 , n47505 , n40728 );
and ( n47507 , n47501 , n47506 );
and ( n47508 , n47497 , n47506 );
or ( n47509 , n47502 , n47507 , n47508 );
and ( n47510 , n44565 , n39896 );
and ( n47511 , n44520 , n39894 );
nor ( n47512 , n47510 , n47511 );
xnor ( n47513 , n47512 , n39857 );
and ( n47514 , n44665 , n39760 );
and ( n47515 , n44656 , n39758 );
nor ( n47516 , n47514 , n47515 );
xnor ( n47517 , n47516 , n39742 );
and ( n47518 , n47513 , n47517 );
xor ( n47519 , n47237 , n47241 );
xor ( n47520 , n47519 , n47244 );
and ( n47521 , n47517 , n47520 );
and ( n47522 , n47513 , n47520 );
or ( n47523 , n47518 , n47521 , n47522 );
and ( n47524 , n44357 , n40053 );
and ( n47525 , n44347 , n40051 );
nor ( n47526 , n47524 , n47525 );
xnor ( n47527 , n47526 , n39999 );
and ( n47528 , n47523 , n47527 );
xor ( n47529 , n47247 , n47251 );
xor ( n47530 , n47529 , n47254 );
and ( n47531 , n47527 , n47530 );
and ( n47532 , n47523 , n47530 );
or ( n47533 , n47528 , n47531 , n47532 );
xor ( n47534 , n47257 , n47261 );
xor ( n47535 , n47534 , n47264 );
and ( n47536 , n47533 , n47535 );
xor ( n47537 , n47414 , n47418 );
xor ( n47538 , n47537 , n47421 );
and ( n47539 , n47535 , n47538 );
and ( n47540 , n47533 , n47538 );
or ( n47541 , n47536 , n47539 , n47540 );
and ( n47542 , n43192 , n40527 );
and ( n47543 , n43073 , n40525 );
nor ( n47544 , n47542 , n47543 );
xnor ( n47545 , n47544 , n40382 );
and ( n47546 , n47541 , n47545 );
xor ( n47547 , n47267 , n47271 );
xor ( n47548 , n47547 , n47274 );
and ( n47549 , n47545 , n47548 );
and ( n47550 , n47541 , n47548 );
or ( n47551 , n47546 , n47549 , n47550 );
and ( n47552 , n43019 , n40746 );
and ( n47553 , n42811 , n40744 );
nor ( n47554 , n47552 , n47553 );
xnor ( n47555 , n47554 , n40501 );
and ( n47556 , n47551 , n47555 );
xor ( n47557 , n47277 , n47281 );
xor ( n47558 , n47557 , n47284 );
and ( n47559 , n47555 , n47558 );
and ( n47560 , n47551 , n47558 );
or ( n47561 , n47556 , n47559 , n47560 );
xor ( n47562 , n47287 , n47321 );
xor ( n47563 , n47562 , n47326 );
and ( n47564 , n47561 , n47563 );
xor ( n47565 , n47444 , n47448 );
xor ( n47566 , n47565 , n47451 );
and ( n47567 , n47563 , n47566 );
and ( n47568 , n47561 , n47566 );
or ( n47569 , n47564 , n47567 , n47568 );
and ( n47570 , n47509 , n47569 );
and ( n47571 , n41032 , n41984 );
and ( n47572 , n41047 , n41982 );
nor ( n47573 , n47571 , n47572 );
xnor ( n47574 , n47573 , n41687 );
and ( n47575 , n47569 , n47574 );
and ( n574883 , n47509 , n47574 );
or ( n47576 , n47570 , n47575 , n574883 );
and ( n47577 , n40869 , n42269 );
and ( n47578 , n40738 , n42266 );
nor ( n47579 , n47577 , n47578 );
xnor ( n47580 , n47579 , n41684 );
xor ( n47581 , n47351 , n47355 );
xor ( n47582 , n47581 , n47360 );
and ( n47583 , n47580 , n47582 );
xor ( n47584 , n47454 , n47458 );
xor ( n47585 , n47584 , n47461 );
and ( n47586 , n47582 , n47585 );
and ( n47587 , n47580 , n47585 );
or ( n47588 , n47583 , n47586 , n47587 );
and ( n47589 , n47576 , n47588 );
xor ( n47590 , n47363 , n47367 );
xor ( n47591 , n47590 , n47370 );
and ( n47592 , n47588 , n47591 );
and ( n47593 , n47576 , n47591 );
or ( n47594 , n47589 , n47592 , n47593 );
xor ( n47595 , n47347 , n47373 );
xor ( n47596 , n47595 , n47378 );
and ( n47597 , n47594 , n47596 );
xor ( n47598 , n47474 , n47476 );
xor ( n47599 , n47598 , n47479 );
and ( n47600 , n47596 , n47599 );
and ( n47601 , n47594 , n47599 );
or ( n47602 , n47597 , n47600 , n47601 );
and ( n47603 , n47493 , n47602 );
xor ( n47604 , n47594 , n47596 );
xor ( n47605 , n47604 , n47599 );
and ( n47606 , n41807 , n41622 );
and ( n47607 , n41692 , n41620 );
nor ( n47608 , n47606 , n47607 );
xnor ( n47609 , n47608 , n41194 );
and ( n47610 , n42061 , n41292 );
and ( n47611 , n41816 , n41290 );
nor ( n47612 , n47610 , n47611 );
xnor ( n47613 , n47612 , n41041 );
and ( n47614 , n47609 , n47613 );
xor ( n47615 , n47551 , n47555 );
xor ( n47616 , n47615 , n47558 );
and ( n47617 , n47613 , n47616 );
and ( n47618 , n47609 , n47616 );
or ( n47619 , n47614 , n47617 , n47618 );
xor ( n47620 , n47116 , n47120 );
and ( n47621 , n44991 , n39758 );
not ( n47622 , n47621 );
and ( n47623 , n47622 , n39742 );
and ( n47624 , n44991 , n39760 );
and ( n47625 , n44999 , n39758 );
nor ( n47626 , n47624 , n47625 );
xnor ( n47627 , n47626 , n39742 );
and ( n47628 , n47623 , n47627 );
and ( n47629 , n44999 , n39760 );
and ( n47630 , n45008 , n39758 );
nor ( n47631 , n47629 , n47630 );
xnor ( n47632 , n47631 , n39742 );
and ( n47633 , n47628 , n47632 );
and ( n47634 , n47632 , n47114 );
and ( n47635 , n47628 , n47114 );
or ( n47636 , n47633 , n47634 , n47635 );
and ( n47637 , n47620 , n47636 );
and ( n47638 , n45008 , n39760 );
and ( n47639 , n45021 , n39758 );
nor ( n47640 , n47638 , n47639 );
xnor ( n47641 , n47640 , n39742 );
and ( n47642 , n47636 , n47641 );
and ( n47643 , n47620 , n47641 );
or ( n47644 , n47637 , n47642 , n47643 );
and ( n47645 , n45021 , n39760 );
and ( n47646 , n45034 , n39758 );
nor ( n47647 , n47645 , n47646 );
xnor ( n47648 , n47647 , n39742 );
and ( n47649 , n47644 , n47648 );
xor ( n47650 , n47121 , n47125 );
xor ( n47651 , n47650 , n46651 );
and ( n47652 , n47648 , n47651 );
and ( n47653 , n47644 , n47651 );
or ( n47654 , n47649 , n47652 , n47653 );
and ( n47655 , n45034 , n39760 );
and ( n47656 , n45047 , n39758 );
nor ( n47657 , n47655 , n47656 );
xnor ( n47658 , n47657 , n39742 );
and ( n47659 , n47654 , n47658 );
xor ( n47660 , n47113 , n47129 );
xor ( n47661 , n47660 , n47134 );
and ( n47662 , n47658 , n47661 );
and ( n47663 , n47654 , n47661 );
or ( n47664 , n47659 , n47662 , n47663 );
and ( n47665 , n45047 , n39760 );
and ( n47666 , n45060 , n39758 );
nor ( n47667 , n47665 , n47666 );
xnor ( n47668 , n47667 , n39742 );
and ( n47669 , n47664 , n47668 );
xor ( n47670 , n47137 , n47141 );
xor ( n47671 , n47670 , n47144 );
and ( n47672 , n47668 , n47671 );
and ( n47673 , n47664 , n47671 );
or ( n47674 , n47669 , n47672 , n47673 );
and ( n47675 , n45060 , n39760 );
and ( n47676 , n45073 , n39758 );
nor ( n47677 , n47675 , n47676 );
xnor ( n47678 , n47677 , n39742 );
and ( n47679 , n47674 , n47678 );
xor ( n47680 , n47147 , n47151 );
xor ( n47681 , n47680 , n47154 );
and ( n47682 , n47678 , n47681 );
and ( n47683 , n47674 , n47681 );
or ( n47684 , n47679 , n47682 , n47683 );
and ( n47685 , n45073 , n39760 );
and ( n47686 , n45086 , n39758 );
nor ( n47687 , n47685 , n47686 );
xnor ( n47688 , n47687 , n39742 );
and ( n47689 , n47684 , n47688 );
xor ( n47690 , n47157 , n47161 );
xor ( n47691 , n47690 , n47164 );
and ( n47692 , n47688 , n47691 );
and ( n47693 , n47684 , n47691 );
or ( n47694 , n47689 , n47692 , n47693 );
and ( n47695 , n45086 , n39760 );
and ( n47696 , n45099 , n39758 );
nor ( n47697 , n47695 , n47696 );
xnor ( n47698 , n47697 , n39742 );
and ( n47699 , n47694 , n47698 );
xor ( n47700 , n47167 , n47171 );
xor ( n47701 , n47700 , n47174 );
and ( n47702 , n47698 , n47701 );
and ( n47703 , n47694 , n47701 );
or ( n47704 , n47699 , n47702 , n47703 );
and ( n47705 , n45099 , n39760 );
and ( n47706 , n45112 , n39758 );
nor ( n47707 , n47705 , n47706 );
xnor ( n47708 , n47707 , n39742 );
and ( n47709 , n47704 , n47708 );
xor ( n47710 , n47177 , n47181 );
xor ( n47711 , n47710 , n47184 );
and ( n47712 , n47708 , n47711 );
and ( n47713 , n47704 , n47711 );
or ( n47714 , n47709 , n47712 , n47713 );
and ( n47715 , n45112 , n39760 );
and ( n47716 , n45125 , n39758 );
nor ( n47717 , n47715 , n47716 );
xnor ( n47718 , n47717 , n39742 );
and ( n47719 , n47714 , n47718 );
xor ( n47720 , n47187 , n47191 );
xor ( n47721 , n47720 , n47194 );
and ( n47722 , n47718 , n47721 );
and ( n47723 , n47714 , n47721 );
or ( n47724 , n47719 , n47722 , n47723 );
and ( n47725 , n45125 , n39760 );
and ( n47726 , n45138 , n39758 );
nor ( n47727 , n47725 , n47726 );
xnor ( n47728 , n47727 , n39742 );
and ( n47729 , n47724 , n47728 );
xor ( n47730 , n47197 , n47201 );
xor ( n47731 , n47730 , n47204 );
and ( n47732 , n47728 , n47731 );
and ( n47733 , n47724 , n47731 );
or ( n47734 , n47729 , n47732 , n47733 );
and ( n47735 , n45138 , n39760 );
and ( n47736 , n45151 , n39758 );
nor ( n47737 , n47735 , n47736 );
xnor ( n47738 , n47737 , n39742 );
and ( n47739 , n47734 , n47738 );
xor ( n47740 , n47207 , n47211 );
xor ( n47741 , n47740 , n47214 );
and ( n47742 , n47738 , n47741 );
and ( n47743 , n47734 , n47741 );
or ( n47744 , n47739 , n47742 , n47743 );
and ( n47745 , n45151 , n39760 );
and ( n47746 , n45164 , n39758 );
nor ( n47747 , n47745 , n47746 );
xnor ( n47748 , n47747 , n39742 );
and ( n47749 , n47744 , n47748 );
xor ( n47750 , n47217 , n47221 );
xor ( n47751 , n47750 , n47224 );
and ( n47752 , n47748 , n47751 );
and ( n47753 , n47744 , n47751 );
or ( n47754 , n47749 , n47752 , n47753 );
and ( n47755 , n45164 , n39760 );
and ( n47756 , n44665 , n39758 );
nor ( n47757 , n47755 , n47756 );
xnor ( n47758 , n47757 , n39742 );
and ( n47759 , n47754 , n47758 );
xor ( n47760 , n47227 , n47231 );
xor ( n47761 , n47760 , n47234 );
and ( n47762 , n47758 , n47761 );
and ( n47763 , n47754 , n47761 );
or ( n47764 , n47759 , n47762 , n47763 );
and ( n47765 , n44458 , n40053 );
and ( n47766 , n44357 , n40051 );
nor ( n47767 , n47765 , n47766 );
xnor ( n47768 , n47767 , n39999 );
and ( n47769 , n47764 , n47768 );
buf ( n47770 , n557796 );
not ( n47771 , n47770 );
and ( n47772 , n47768 , n47771 );
and ( n47773 , n47764 , n47771 );
or ( n47774 , n47769 , n47772 , n47773 );
and ( n47775 , n44264 , n40258 );
and ( n47776 , n43437 , n40256 );
nor ( n47777 , n47775 , n47776 );
xnor ( n47778 , n47777 , n40169 );
and ( n47779 , n47774 , n47778 );
xor ( n47780 , n47404 , n47408 );
xor ( n47781 , n47780 , n47411 );
and ( n47782 , n47778 , n47781 );
and ( n47783 , n47774 , n47781 );
or ( n47784 , n47779 , n47782 , n47783 );
and ( n47785 , n43200 , n40527 );
and ( n47786 , n43192 , n40525 );
nor ( n47787 , n47785 , n47786 );
xnor ( n47788 , n47787 , n40382 );
and ( n47789 , n47784 , n47788 );
and ( n47790 , n43437 , n40258 );
and ( n47791 , n43428 , n40256 );
nor ( n47792 , n47790 , n47791 );
xnor ( n47793 , n47792 , n40169 );
and ( n47794 , n47788 , n47793 );
and ( n47795 , n47784 , n47793 );
or ( n47796 , n47789 , n47794 , n47795 );
xor ( n47797 , n47424 , n47428 );
xor ( n47798 , n47797 , n47431 );
and ( n47799 , n47796 , n47798 );
xor ( n47800 , n47541 , n47545 );
xor ( n47801 , n47800 , n47548 );
and ( n47802 , n47798 , n47801 );
and ( n47803 , n47796 , n47801 );
or ( n47804 , n47799 , n47802 , n47803 );
and ( n47805 , n42456 , n41055 );
and ( n47806 , n42048 , n41053 );
nor ( n47807 , n47805 , n47806 );
xnor ( n47808 , n47807 , n40728 );
and ( n47809 , n47804 , n47808 );
xor ( n47810 , n47434 , n47438 );
xor ( n47811 , n47810 , n47441 );
and ( n47812 , n47808 , n47811 );
and ( n47813 , n47804 , n47811 );
or ( n47814 , n47809 , n47812 , n47813 );
and ( n47815 , n47619 , n47814 );
and ( n47816 , n41182 , n41984 );
and ( n47817 , n41032 , n41982 );
nor ( n47818 , n47816 , n47817 );
xnor ( n47819 , n47818 , n41687 );
and ( n47820 , n47814 , n47819 );
and ( n47821 , n47619 , n47819 );
or ( n47822 , n47815 , n47820 , n47821 );
and ( n47823 , n41047 , n42269 );
and ( n47824 , n40869 , n42266 );
nor ( n47825 , n47823 , n47824 );
xnor ( n47826 , n47825 , n41684 );
xor ( n47827 , n47497 , n47501 );
xor ( n47828 , n47827 , n47506 );
and ( n47829 , n47826 , n47828 );
xor ( n47830 , n47561 , n47563 );
xor ( n47831 , n47830 , n47566 );
and ( n47832 , n47828 , n47831 );
and ( n47833 , n47826 , n47831 );
or ( n47834 , n47829 , n47832 , n47833 );
and ( n47835 , n47822 , n47834 );
xor ( n47836 , n47509 , n47569 );
xor ( n47837 , n47836 , n47574 );
and ( n47838 , n47834 , n47837 );
and ( n47839 , n47822 , n47837 );
or ( n47840 , n47835 , n47838 , n47839 );
xor ( n47841 , n47464 , n47468 );
xor ( n47842 , n47841 , n47471 );
and ( n47843 , n47840 , n47842 );
xor ( n47844 , n47576 , n47588 );
xor ( n47845 , n47844 , n47591 );
and ( n47846 , n47842 , n47845 );
and ( n47847 , n47840 , n47845 );
or ( n47848 , n47843 , n47846 , n47847 );
and ( n47849 , n47605 , n47848 );
and ( n47850 , n41692 , n41984 );
and ( n47851 , n41615 , n41982 );
nor ( n47852 , n47850 , n47851 );
xnor ( n47853 , n47852 , n41687 );
and ( n47854 , n42048 , n41292 );
and ( n47855 , n42061 , n41290 );
nor ( n47856 , n47854 , n47855 );
xnor ( n47857 , n47856 , n41041 );
and ( n47858 , n47853 , n47857 );
and ( n47859 , n44520 , n40053 );
and ( n47860 , n44458 , n40051 );
nor ( n47861 , n47859 , n47860 );
xnor ( n47862 , n47861 , n39999 );
and ( n47863 , n44656 , n39896 );
and ( n47864 , n44565 , n39894 );
nor ( n47865 , n47863 , n47864 );
xnor ( n47866 , n47865 , n39857 );
and ( n47867 , n47862 , n47866 );
buf ( n47868 , n557797 );
not ( n47869 , n47868 );
and ( n47870 , n47866 , n47869 );
and ( n47871 , n47862 , n47869 );
or ( n47872 , n47867 , n47870 , n47871 );
and ( n47873 , n44347 , n40258 );
and ( n47874 , n44264 , n40256 );
nor ( n47875 , n47873 , n47874 );
xnor ( n47876 , n47875 , n40169 );
and ( n47877 , n47872 , n47876 );
xor ( n47878 , n47513 , n47517 );
xor ( n47879 , n47878 , n47520 );
and ( n47880 , n47876 , n47879 );
and ( n47881 , n47872 , n47879 );
or ( n47882 , n47877 , n47880 , n47881 );
and ( n47883 , n43428 , n40527 );
and ( n47884 , n43200 , n40525 );
nor ( n47885 , n47883 , n47884 );
xnor ( n47886 , n47885 , n40382 );
and ( n47887 , n47882 , n47886 );
xor ( n47888 , n47523 , n47527 );
xor ( n47889 , n47888 , n47530 );
and ( n47890 , n47886 , n47889 );
and ( n47891 , n47882 , n47889 );
or ( n47892 , n47887 , n47890 , n47891 );
xor ( n47893 , n47784 , n47788 );
xor ( n47894 , n47893 , n47793 );
and ( n47895 , n47892 , n47894 );
xor ( n47896 , n47533 , n47535 );
xor ( n47897 , n47896 , n47538 );
and ( n47898 , n47894 , n47897 );
and ( n47899 , n47892 , n47897 );
or ( n47900 , n47895 , n47898 , n47899 );
and ( n47901 , n42811 , n41055 );
and ( n47902 , n42456 , n41053 );
nor ( n47903 , n47901 , n47902 );
xnor ( n47904 , n47903 , n40728 );
xor ( n47905 , n47900 , n47904 );
and ( n47906 , n43027 , n40746 );
and ( n47907 , n43019 , n40744 );
nor ( n47908 , n47906 , n47907 );
xnor ( n47909 , n47908 , n40501 );
xor ( n47910 , n47905 , n47909 );
and ( n47911 , n47857 , n47910 );
and ( n47912 , n47853 , n47910 );
or ( n47913 , n47858 , n47911 , n47912 );
and ( n47914 , n44565 , n40053 );
and ( n47915 , n44520 , n40051 );
nor ( n47916 , n47914 , n47915 );
xnor ( n47917 , n47916 , n39999 );
and ( n47918 , n44665 , n39896 );
and ( n47919 , n44656 , n39894 );
nor ( n47920 , n47918 , n47919 );
xnor ( n47921 , n47920 , n39857 );
and ( n47922 , n47917 , n47921 );
xor ( n47923 , n47744 , n47748 );
xor ( n47924 , n47923 , n47751 );
and ( n47925 , n47921 , n47924 );
and ( n47926 , n47917 , n47924 );
or ( n47927 , n47922 , n47925 , n47926 );
and ( n47928 , n44357 , n40258 );
and ( n47929 , n44347 , n40256 );
nor ( n47930 , n47928 , n47929 );
xnor ( n47931 , n47930 , n40169 );
and ( n47932 , n47927 , n47931 );
xor ( n47933 , n47754 , n47758 );
xor ( n47934 , n47933 , n47761 );
and ( n47935 , n47931 , n47934 );
and ( n47936 , n47927 , n47934 );
or ( n47937 , n47932 , n47935 , n47936 );
xor ( n47938 , n47764 , n47768 );
xor ( n47939 , n47938 , n47771 );
and ( n47940 , n47937 , n47939 );
xor ( n47941 , n47872 , n47876 );
xor ( n47942 , n47941 , n47879 );
and ( n47943 , n47939 , n47942 );
and ( n47944 , n47937 , n47942 );
or ( n47945 , n47940 , n47943 , n47944 );
and ( n47946 , n43192 , n40746 );
and ( n47947 , n43073 , n40744 );
nor ( n47948 , n47946 , n47947 );
xnor ( n47949 , n47948 , n40501 );
and ( n47950 , n47945 , n47949 );
xor ( n47951 , n47774 , n47778 );
xor ( n47952 , n47951 , n47781 );
and ( n47953 , n47949 , n47952 );
and ( n47954 , n47945 , n47952 );
or ( n47955 , n47950 , n47953 , n47954 );
and ( n47956 , n43019 , n41055 );
and ( n47957 , n42811 , n41053 );
nor ( n47958 , n47956 , n47957 );
xnor ( n47959 , n47958 , n40728 );
and ( n47960 , n47955 , n47959 );
and ( n47961 , n43073 , n40746 );
and ( n47962 , n43027 , n40744 );
nor ( n47963 , n47961 , n47962 );
xnor ( n47964 , n47963 , n40501 );
and ( n47965 , n47959 , n47964 );
and ( n47966 , n47955 , n47964 );
or ( n47967 , n47960 , n47965 , n47966 );
and ( n47968 , n41816 , n41622 );
and ( n47969 , n41807 , n41620 );
nor ( n47970 , n47968 , n47969 );
xnor ( n47971 , n47970 , n41194 );
and ( n47972 , n47967 , n47971 );
xor ( n47973 , n47796 , n47798 );
xor ( n47974 , n47973 , n47801 );
and ( n47975 , n47971 , n47974 );
and ( n47976 , n47967 , n47974 );
or ( n47977 , n47972 , n47975 , n47976 );
and ( n47978 , n47913 , n47977 );
and ( n47979 , n41032 , n42269 );
and ( n47980 , n41047 , n42266 );
nor ( n47981 , n47979 , n47980 );
xnor ( n47982 , n47981 , n41684 );
and ( n47983 , n47977 , n47982 );
and ( n47984 , n47913 , n47982 );
or ( n47985 , n47978 , n47983 , n47984 );
and ( n47986 , n47900 , n47904 );
and ( n47987 , n47904 , n47909 );
and ( n47988 , n47900 , n47909 );
or ( n47989 , n47986 , n47987 , n47988 );
and ( n47990 , n41615 , n41984 );
and ( n47991 , n41182 , n41982 );
nor ( n47992 , n47990 , n47991 );
xnor ( n47993 , n47992 , n41687 );
and ( n47994 , n47989 , n47993 );
xor ( n47995 , n47804 , n47808 );
xor ( n47996 , n47995 , n47811 );
and ( n47997 , n47993 , n47996 );
and ( n47998 , n47989 , n47996 );
or ( n47999 , n47994 , n47997 , n47998 );
and ( n48000 , n47985 , n47999 );
xor ( n48001 , n47619 , n47814 );
xor ( n48002 , n48001 , n47819 );
and ( n48003 , n47999 , n48002 );
and ( n48004 , n47985 , n48002 );
or ( n48005 , n48000 , n48003 , n48004 );
xor ( n48006 , n47822 , n47834 );
xor ( n48007 , n48006 , n47837 );
and ( n48008 , n48005 , n48007 );
xor ( n48009 , n47580 , n47582 );
xor ( n48010 , n48009 , n47585 );
and ( n48011 , n48007 , n48010 );
and ( n48012 , n48005 , n48010 );
or ( n48013 , n48008 , n48011 , n48012 );
xor ( n48014 , n47840 , n47842 );
xor ( n48015 , n48014 , n47845 );
and ( n48016 , n48013 , n48015 );
xor ( n48017 , n48005 , n48007 );
xor ( n48018 , n48017 , n48010 );
xor ( n48019 , n47623 , n47627 );
and ( n48020 , n44991 , n39894 );
not ( n48021 , n48020 );
and ( n48022 , n48021 , n39857 );
and ( n48023 , n44991 , n39896 );
and ( n48024 , n44999 , n39894 );
nor ( n48025 , n48023 , n48024 );
xnor ( n48026 , n48025 , n39857 );
and ( n48027 , n48022 , n48026 );
and ( n48028 , n44999 , n39896 );
and ( n48029 , n45008 , n39894 );
nor ( n48030 , n48028 , n48029 );
xnor ( n48031 , n48030 , n39857 );
and ( n48032 , n48027 , n48031 );
and ( n48033 , n48031 , n47621 );
and ( n48034 , n48027 , n47621 );
or ( n48035 , n48032 , n48033 , n48034 );
and ( n48036 , n48019 , n48035 );
and ( n48037 , n45008 , n39896 );
and ( n48038 , n45021 , n39894 );
nor ( n48039 , n48037 , n48038 );
xnor ( n48040 , n48039 , n39857 );
and ( n48041 , n48035 , n48040 );
and ( n48042 , n48019 , n48040 );
or ( n48043 , n48036 , n48041 , n48042 );
and ( n48044 , n45021 , n39896 );
and ( n48045 , n45034 , n39894 );
nor ( n48046 , n48044 , n48045 );
xnor ( n48047 , n48046 , n39857 );
and ( n48048 , n48043 , n48047 );
xor ( n48049 , n47628 , n47632 );
xor ( n48050 , n48049 , n47114 );
and ( n48051 , n48047 , n48050 );
and ( n48052 , n48043 , n48050 );
or ( n48053 , n48048 , n48051 , n48052 );
and ( n48054 , n45034 , n39896 );
and ( n48055 , n45047 , n39894 );
nor ( n48056 , n48054 , n48055 );
xnor ( n48057 , n48056 , n39857 );
and ( n48058 , n48053 , n48057 );
xor ( n48059 , n47620 , n47636 );
xor ( n48060 , n48059 , n47641 );
and ( n48061 , n48057 , n48060 );
and ( n48062 , n48053 , n48060 );
or ( n48063 , n48058 , n48061 , n48062 );
and ( n48064 , n45047 , n39896 );
and ( n48065 , n45060 , n39894 );
nor ( n48066 , n48064 , n48065 );
xnor ( n48067 , n48066 , n39857 );
and ( n48068 , n48063 , n48067 );
xor ( n48069 , n47644 , n47648 );
xor ( n48070 , n48069 , n47651 );
and ( n48071 , n48067 , n48070 );
and ( n48072 , n48063 , n48070 );
or ( n48073 , n48068 , n48071 , n48072 );
and ( n48074 , n45060 , n39896 );
and ( n48075 , n45073 , n39894 );
nor ( n48076 , n48074 , n48075 );
xnor ( n48077 , n48076 , n39857 );
and ( n48078 , n48073 , n48077 );
xor ( n48079 , n47654 , n47658 );
xor ( n48080 , n48079 , n47661 );
and ( n48081 , n48077 , n48080 );
and ( n48082 , n48073 , n48080 );
or ( n48083 , n48078 , n48081 , n48082 );
and ( n48084 , n45073 , n39896 );
and ( n48085 , n45086 , n39894 );
nor ( n48086 , n48084 , n48085 );
xnor ( n48087 , n48086 , n39857 );
and ( n48088 , n48083 , n48087 );
xor ( n48089 , n47664 , n47668 );
xor ( n48090 , n48089 , n47671 );
and ( n48091 , n48087 , n48090 );
and ( n48092 , n48083 , n48090 );
or ( n48093 , n48088 , n48091 , n48092 );
and ( n48094 , n45086 , n39896 );
and ( n48095 , n45099 , n39894 );
nor ( n48096 , n48094 , n48095 );
xnor ( n48097 , n48096 , n39857 );
and ( n48098 , n48093 , n48097 );
xor ( n48099 , n47674 , n47678 );
xor ( n48100 , n48099 , n47681 );
and ( n48101 , n48097 , n48100 );
and ( n48102 , n48093 , n48100 );
or ( n48103 , n48098 , n48101 , n48102 );
and ( n48104 , n45099 , n39896 );
and ( n48105 , n45112 , n39894 );
nor ( n48106 , n48104 , n48105 );
xnor ( n48107 , n48106 , n39857 );
and ( n48108 , n48103 , n48107 );
xor ( n48109 , n47684 , n47688 );
xor ( n48110 , n48109 , n47691 );
and ( n48111 , n48107 , n48110 );
and ( n48112 , n48103 , n48110 );
or ( n48113 , n48108 , n48111 , n48112 );
and ( n48114 , n45112 , n39896 );
and ( n48115 , n45125 , n39894 );
nor ( n48116 , n48114 , n48115 );
xnor ( n48117 , n48116 , n39857 );
and ( n48118 , n48113 , n48117 );
xor ( n48119 , n47694 , n47698 );
xor ( n48120 , n48119 , n47701 );
and ( n48121 , n48117 , n48120 );
and ( n48122 , n48113 , n48120 );
or ( n48123 , n48118 , n48121 , n48122 );
and ( n48124 , n45125 , n39896 );
and ( n48125 , n45138 , n39894 );
nor ( n48126 , n48124 , n48125 );
xnor ( n48127 , n48126 , n39857 );
and ( n48128 , n48123 , n48127 );
xor ( n48129 , n47704 , n47708 );
xor ( n48130 , n48129 , n47711 );
and ( n48131 , n48127 , n48130 );
and ( n48132 , n48123 , n48130 );
or ( n48133 , n48128 , n48131 , n48132 );
and ( n48134 , n45138 , n39896 );
and ( n48135 , n45151 , n39894 );
nor ( n48136 , n48134 , n48135 );
xnor ( n48137 , n48136 , n39857 );
and ( n48138 , n48133 , n48137 );
xor ( n48139 , n47714 , n47718 );
xor ( n48140 , n48139 , n47721 );
and ( n48141 , n48137 , n48140 );
and ( n48142 , n48133 , n48140 );
or ( n48143 , n48138 , n48141 , n48142 );
and ( n48144 , n45151 , n39896 );
and ( n48145 , n45164 , n39894 );
nor ( n48146 , n48144 , n48145 );
xnor ( n48147 , n48146 , n39857 );
and ( n48148 , n48143 , n48147 );
xor ( n48149 , n47724 , n47728 );
xor ( n48150 , n48149 , n47731 );
and ( n48151 , n48147 , n48150 );
and ( n48152 , n48143 , n48150 );
or ( n48153 , n48148 , n48151 , n48152 );
and ( n48154 , n45164 , n39896 );
and ( n48155 , n44665 , n39894 );
nor ( n48156 , n48154 , n48155 );
xnor ( n48157 , n48156 , n39857 );
and ( n48158 , n48153 , n48157 );
xor ( n48159 , n47734 , n47738 );
xor ( n48160 , n48159 , n47741 );
and ( n48161 , n48157 , n48160 );
and ( n48162 , n48153 , n48160 );
or ( n48163 , n48158 , n48161 , n48162 );
and ( n48164 , n44458 , n40258 );
and ( n48165 , n44357 , n40256 );
nor ( n48166 , n48164 , n48165 );
xnor ( n48167 , n48166 , n40169 );
and ( n48168 , n48163 , n48167 );
buf ( n48169 , n557798 );
not ( n48170 , n48169 );
and ( n48171 , n48167 , n48170 );
and ( n48172 , n48163 , n48170 );
or ( n48173 , n48168 , n48171 , n48172 );
and ( n48174 , n44264 , n40527 );
and ( n48175 , n43437 , n40525 );
nor ( n48176 , n48174 , n48175 );
xnor ( n48177 , n48176 , n40382 );
and ( n48178 , n48173 , n48177 );
xor ( n48179 , n47862 , n47866 );
xor ( n48180 , n48179 , n47869 );
and ( n48181 , n48177 , n48180 );
and ( n48182 , n48173 , n48180 );
or ( n48183 , n48178 , n48181 , n48182 );
and ( n48184 , n43200 , n40746 );
and ( n48185 , n43192 , n40744 );
nor ( n48186 , n48184 , n48185 );
xnor ( n48187 , n48186 , n40501 );
and ( n48188 , n48183 , n48187 );
and ( n48189 , n43437 , n40527 );
and ( n48190 , n43428 , n40525 );
nor ( n48191 , n48189 , n48190 );
xnor ( n48192 , n48191 , n40382 );
and ( n48193 , n48187 , n48192 );
and ( n48194 , n48183 , n48192 );
or ( n48195 , n48188 , n48193 , n48194 );
and ( n48196 , n43027 , n41055 );
and ( n48197 , n43019 , n41053 );
nor ( n48198 , n48196 , n48197 );
xnor ( n48199 , n48198 , n40728 );
and ( n48200 , n48195 , n48199 );
xor ( n48201 , n47882 , n47886 );
xor ( n48202 , n48201 , n47889 );
and ( n48203 , n48199 , n48202 );
and ( n48204 , n48195 , n48202 );
or ( n48205 , n48200 , n48203 , n48204 );
and ( n48206 , n42456 , n41292 );
and ( n48207 , n42048 , n41290 );
nor ( n48208 , n48206 , n48207 );
xnor ( n48209 , n48208 , n41041 );
and ( n48210 , n48205 , n48209 );
xor ( n48211 , n47892 , n47894 );
xor ( n48212 , n48211 , n47897 );
and ( n48213 , n48209 , n48212 );
and ( n48214 , n48205 , n48212 );
or ( n48215 , n48210 , n48213 , n48214 );
and ( n48216 , n41182 , n42269 );
and ( n48217 , n41032 , n42266 );
nor ( n48218 , n48216 , n48217 );
xnor ( n48219 , n48218 , n41684 );
and ( n48220 , n48215 , n48219 );
xor ( n48221 , n47967 , n47971 );
xor ( n48222 , n48221 , n47974 );
and ( n48223 , n48219 , n48222 );
and ( n48224 , n48215 , n48222 );
or ( n48225 , n48220 , n48223 , n48224 );
xor ( n48226 , n47609 , n47613 );
xor ( n48227 , n48226 , n47616 );
and ( n48228 , n48225 , n48227 );
xor ( n48229 , n47989 , n47993 );
xor ( n48230 , n48229 , n47996 );
and ( n48231 , n48227 , n48230 );
and ( n48232 , n48225 , n48230 );
or ( n48233 , n48228 , n48231 , n48232 );
xor ( n48234 , n47985 , n47999 );
xor ( n48235 , n48234 , n48002 );
and ( n48236 , n48233 , n48235 );
xor ( n48237 , n47826 , n47828 );
xor ( n48238 , n48237 , n47831 );
and ( n48239 , n48235 , n48238 );
and ( n48240 , n48233 , n48238 );
or ( n48241 , n48236 , n48239 , n48240 );
and ( n48242 , n48018 , n48241 );
and ( n48243 , n44520 , n40258 );
and ( n48244 , n44458 , n40256 );
nor ( n48245 , n48243 , n48244 );
xnor ( n48246 , n48245 , n40169 );
and ( n48247 , n44656 , n40053 );
and ( n48248 , n44565 , n40051 );
nor ( n48249 , n48247 , n48248 );
xnor ( n48250 , n48249 , n39999 );
and ( n48251 , n48246 , n48250 );
buf ( n48252 , n557799 );
not ( n48253 , n48252 );
and ( n48254 , n48250 , n48253 );
and ( n48255 , n48246 , n48253 );
or ( n48256 , n48251 , n48254 , n48255 );
and ( n48257 , n44347 , n40527 );
and ( n48258 , n44264 , n40525 );
nor ( n48259 , n48257 , n48258 );
xnor ( n48260 , n48259 , n40382 );
and ( n48261 , n48256 , n48260 );
xor ( n48262 , n47917 , n47921 );
xor ( n48263 , n48262 , n47924 );
and ( n48264 , n48260 , n48263 );
and ( n48265 , n48256 , n48263 );
or ( n48266 , n48261 , n48264 , n48265 );
xor ( n48267 , n48173 , n48177 );
xor ( n48268 , n48267 , n48180 );
and ( n48269 , n48266 , n48268 );
xor ( n48270 , n47927 , n47931 );
xor ( n48271 , n48270 , n47934 );
and ( n48272 , n48268 , n48271 );
and ( n48273 , n48266 , n48271 );
or ( n48274 , n48269 , n48272 , n48273 );
and ( n48275 , n43073 , n41055 );
and ( n48276 , n43027 , n41053 );
nor ( n48277 , n48275 , n48276 );
xnor ( n48278 , n48277 , n40728 );
and ( n48279 , n48274 , n48278 );
xor ( n48280 , n47937 , n47939 );
xor ( n48281 , n48280 , n47942 );
and ( n48282 , n48278 , n48281 );
and ( n48283 , n48274 , n48281 );
or ( n48284 , n48279 , n48282 , n48283 );
and ( n48285 , n42811 , n41292 );
and ( n48286 , n42456 , n41290 );
nor ( n48287 , n48285 , n48286 );
xnor ( n48288 , n48287 , n41041 );
and ( n48289 , n48284 , n48288 );
xor ( n48290 , n47945 , n47949 );
xor ( n48291 , n48290 , n47952 );
and ( n48292 , n48288 , n48291 );
and ( n48293 , n48284 , n48291 );
or ( n48294 , n48289 , n48292 , n48293 );
and ( n48295 , n42061 , n41622 );
and ( n48296 , n41816 , n41620 );
nor ( n48297 , n48295 , n48296 );
xnor ( n48298 , n48297 , n41194 );
and ( n48299 , n48294 , n48298 );
xor ( n48300 , n47955 , n47959 );
xor ( n48301 , n48300 , n47964 );
and ( n48302 , n48298 , n48301 );
and ( n48303 , n48294 , n48301 );
or ( n48304 , n48299 , n48302 , n48303 );
and ( n48305 , n41615 , n42269 );
and ( n48306 , n41182 , n42266 );
nor ( n48307 , n48305 , n48306 );
xnor ( n48308 , n48307 , n41684 );
and ( n48309 , n41807 , n41984 );
and ( n48310 , n41692 , n41982 );
nor ( n48311 , n48309 , n48310 );
xnor ( n48312 , n48311 , n41687 );
and ( n48313 , n48308 , n48312 );
xor ( n48314 , n48205 , n48209 );
xor ( n48315 , n48314 , n48212 );
and ( n48316 , n48312 , n48315 );
and ( n48317 , n48308 , n48315 );
or ( n48318 , n48313 , n48316 , n48317 );
and ( n48319 , n48304 , n48318 );
xor ( n48320 , n47853 , n47857 );
xor ( n48321 , n48320 , n47910 );
and ( n48322 , n48318 , n48321 );
and ( n48323 , n48304 , n48321 );
or ( n48324 , n48319 , n48322 , n48323 );
xor ( n48325 , n47913 , n47977 );
xor ( n48326 , n48325 , n47982 );
and ( n48327 , n48324 , n48326 );
xor ( n48328 , n48225 , n48227 );
xor ( n48329 , n48328 , n48230 );
and ( n48330 , n48326 , n48329 );
and ( n48331 , n48324 , n48329 );
or ( n48332 , n48327 , n48330 , n48331 );
xor ( n48333 , n48233 , n48235 );
xor ( n48334 , n48333 , n48238 );
and ( n48335 , n48332 , n48334 );
xor ( n48336 , n48324 , n48326 );
xor ( n48337 , n48336 , n48329 );
and ( n48338 , n41692 , n42269 );
and ( n48339 , n41615 , n42266 );
nor ( n48340 , n48338 , n48339 );
xnor ( n48341 , n48340 , n41684 );
and ( n48342 , n42048 , n41622 );
and ( n48343 , n42061 , n41620 );
nor ( n48344 , n48342 , n48343 );
xnor ( n48345 , n48344 , n41194 );
and ( n48346 , n48341 , n48345 );
xor ( n48347 , n48284 , n48288 );
xor ( n48348 , n48347 , n48291 );
and ( n48349 , n48345 , n48348 );
and ( n48350 , n48341 , n48348 );
or ( n48351 , n48346 , n48349 , n48350 );
and ( n48352 , n44565 , n40258 );
and ( n48353 , n44520 , n40256 );
nor ( n48354 , n48352 , n48353 );
xnor ( n48355 , n48354 , n40169 );
and ( n48356 , n44665 , n40053 );
and ( n48357 , n44656 , n40051 );
nor ( n48358 , n48356 , n48357 );
xnor ( n48359 , n48358 , n39999 );
and ( n48360 , n48355 , n48359 );
xor ( n48361 , n48143 , n48147 );
xor ( n48362 , n48361 , n48150 );
and ( n48363 , n48359 , n48362 );
and ( n48364 , n48355 , n48362 );
or ( n48365 , n48360 , n48363 , n48364 );
and ( n48366 , n44357 , n40527 );
and ( n48367 , n44347 , n40525 );
nor ( n48368 , n48366 , n48367 );
xnor ( n48369 , n48368 , n40382 );
and ( n48370 , n48365 , n48369 );
xor ( n48371 , n48153 , n48157 );
xor ( n48372 , n48371 , n48160 );
and ( n48373 , n48369 , n48372 );
and ( n48374 , n48365 , n48372 );
or ( n48375 , n48370 , n48373 , n48374 );
xor ( n48376 , n48163 , n48167 );
xor ( n48377 , n48376 , n48170 );
and ( n48378 , n48375 , n48377 );
xor ( n48379 , n48256 , n48260 );
xor ( n48380 , n48379 , n48263 );
and ( n48381 , n48377 , n48380 );
and ( n48382 , n48375 , n48380 );
or ( n48383 , n48378 , n48381 , n48382 );
and ( n48384 , n43192 , n41055 );
and ( n48385 , n43073 , n41053 );
nor ( n48386 , n48384 , n48385 );
xnor ( n48387 , n48386 , n40728 );
and ( n48388 , n48383 , n48387 );
and ( n48389 , n43428 , n40746 );
and ( n48390 , n43200 , n40744 );
nor ( n48391 , n48389 , n48390 );
xnor ( n48392 , n48391 , n40501 );
and ( n48393 , n48387 , n48392 );
and ( n48394 , n48383 , n48392 );
or ( n48395 , n48388 , n48393 , n48394 );
and ( n48396 , n43019 , n41292 );
and ( n48397 , n42811 , n41290 );
nor ( n48398 , n48396 , n48397 );
xnor ( n48399 , n48398 , n41041 );
and ( n48400 , n48395 , n48399 );
xor ( n48401 , n48183 , n48187 );
xor ( n48402 , n48401 , n48192 );
and ( n48403 , n48399 , n48402 );
and ( n48404 , n48395 , n48402 );
or ( n48405 , n48400 , n48403 , n48404 );
and ( n48406 , n41816 , n41984 );
and ( n48407 , n41807 , n41982 );
nor ( n48408 , n48406 , n48407 );
xnor ( n48409 , n48408 , n41687 );
and ( n48410 , n48405 , n48409 );
xor ( n48411 , n48195 , n48199 );
xor ( n48412 , n48411 , n48202 );
and ( n48413 , n48409 , n48412 );
and ( n48414 , n48405 , n48412 );
or ( n48415 , n48410 , n48413 , n48414 );
and ( n48416 , n48351 , n48415 );
xor ( n48417 , n48294 , n48298 );
xor ( n48418 , n48417 , n48301 );
and ( n48419 , n48415 , n48418 );
and ( n48420 , n48351 , n48418 );
or ( n48421 , n48416 , n48419 , n48420 );
xor ( n48422 , n48304 , n48318 );
xor ( n48423 , n48422 , n48321 );
and ( n48424 , n48421 , n48423 );
xor ( n48425 , n48215 , n48219 );
xor ( n48426 , n48425 , n48222 );
and ( n48427 , n48423 , n48426 );
and ( n48428 , n48421 , n48426 );
or ( n48429 , n48424 , n48427 , n48428 );
and ( n48430 , n48337 , n48429 );
xor ( n48431 , n48421 , n48423 );
xor ( n48432 , n48431 , n48426 );
and ( n48433 , n44665 , n40258 );
and ( n48434 , n44656 , n40256 );
nor ( n48435 , n48433 , n48434 );
xnor ( n48436 , n48435 , n40169 );
buf ( n48437 , n557802 );
not ( n48438 , n48437 );
and ( n48439 , n48436 , n48438 );
xor ( n48440 , n48022 , n48026 );
and ( n48441 , n44991 , n40051 );
not ( n48442 , n48441 );
and ( n48443 , n48442 , n39999 );
and ( n48444 , n44991 , n40053 );
and ( n48445 , n44999 , n40051 );
nor ( n48446 , n48444 , n48445 );
xnor ( n48447 , n48446 , n39999 );
and ( n48448 , n48443 , n48447 );
and ( n48449 , n44999 , n40053 );
and ( n48450 , n45008 , n40051 );
nor ( n48451 , n48449 , n48450 );
xnor ( n48452 , n48451 , n39999 );
and ( n48453 , n48448 , n48452 );
and ( n48454 , n48452 , n48020 );
and ( n48455 , n48448 , n48020 );
or ( n48456 , n48453 , n48454 , n48455 );
and ( n48457 , n48440 , n48456 );
and ( n48458 , n45008 , n40053 );
and ( n48459 , n45021 , n40051 );
nor ( n48460 , n48458 , n48459 );
xnor ( n48461 , n48460 , n39999 );
and ( n48462 , n48456 , n48461 );
and ( n48463 , n48440 , n48461 );
or ( n48464 , n48457 , n48462 , n48463 );
and ( n48465 , n45021 , n40053 );
and ( n48466 , n45034 , n40051 );
nor ( n48467 , n48465 , n48466 );
xnor ( n48468 , n48467 , n39999 );
and ( n48469 , n48464 , n48468 );
xor ( n48470 , n48027 , n48031 );
xor ( n48471 , n48470 , n47621 );
and ( n48472 , n48468 , n48471 );
and ( n48473 , n48464 , n48471 );
or ( n48474 , n48469 , n48472 , n48473 );
and ( n48475 , n45034 , n40053 );
and ( n48476 , n45047 , n40051 );
nor ( n48477 , n48475 , n48476 );
xnor ( n48478 , n48477 , n39999 );
and ( n48479 , n48474 , n48478 );
xor ( n48480 , n48019 , n48035 );
xor ( n48481 , n48480 , n48040 );
and ( n48482 , n48478 , n48481 );
and ( n48483 , n48474 , n48481 );
or ( n48484 , n48479 , n48482 , n48483 );
and ( n48485 , n45047 , n40053 );
and ( n48486 , n45060 , n40051 );
nor ( n48487 , n48485 , n48486 );
xnor ( n48488 , n48487 , n39999 );
and ( n48489 , n48484 , n48488 );
xor ( n48490 , n48043 , n48047 );
xor ( n48491 , n48490 , n48050 );
and ( n48492 , n48488 , n48491 );
and ( n48493 , n48484 , n48491 );
or ( n48494 , n48489 , n48492 , n48493 );
and ( n48495 , n45060 , n40053 );
and ( n48496 , n45073 , n40051 );
nor ( n48497 , n48495 , n48496 );
xnor ( n48498 , n48497 , n39999 );
and ( n48499 , n48494 , n48498 );
xor ( n48500 , n48053 , n48057 );
xor ( n48501 , n48500 , n48060 );
and ( n48502 , n48498 , n48501 );
and ( n48503 , n48494 , n48501 );
or ( n48504 , n48499 , n48502 , n48503 );
and ( n48505 , n45073 , n40053 );
and ( n48506 , n45086 , n40051 );
nor ( n48507 , n48505 , n48506 );
xnor ( n48508 , n48507 , n39999 );
and ( n48509 , n48504 , n48508 );
xor ( n48510 , n48063 , n48067 );
xor ( n48511 , n48510 , n48070 );
and ( n48512 , n48508 , n48511 );
and ( n48513 , n48504 , n48511 );
or ( n48514 , n48509 , n48512 , n48513 );
and ( n48515 , n45086 , n40053 );
and ( n48516 , n45099 , n40051 );
nor ( n48517 , n48515 , n48516 );
xnor ( n48518 , n48517 , n39999 );
and ( n48519 , n48514 , n48518 );
xor ( n48520 , n48073 , n48077 );
xor ( n48521 , n48520 , n48080 );
and ( n48522 , n48518 , n48521 );
and ( n48523 , n48514 , n48521 );
or ( n48524 , n48519 , n48522 , n48523 );
and ( n48525 , n45099 , n40053 );
and ( n48526 , n45112 , n40051 );
nor ( n48527 , n48525 , n48526 );
xnor ( n48528 , n48527 , n39999 );
and ( n48529 , n48524 , n48528 );
xor ( n48530 , n48083 , n48087 );
xor ( n48531 , n48530 , n48090 );
and ( n48532 , n48528 , n48531 );
and ( n48533 , n48524 , n48531 );
or ( n48534 , n48529 , n48532 , n48533 );
and ( n48535 , n45112 , n40053 );
and ( n48536 , n45125 , n40051 );
nor ( n48537 , n48535 , n48536 );
xnor ( n48538 , n48537 , n39999 );
and ( n48539 , n48534 , n48538 );
xor ( n48540 , n48093 , n48097 );
xor ( n48541 , n48540 , n48100 );
and ( n48542 , n48538 , n48541 );
and ( n48543 , n48534 , n48541 );
or ( n48544 , n48539 , n48542 , n48543 );
and ( n48545 , n45125 , n40053 );
and ( n48546 , n45138 , n40051 );
nor ( n48547 , n48545 , n48546 );
xnor ( n48548 , n48547 , n39999 );
and ( n48549 , n48544 , n48548 );
xor ( n48550 , n48103 , n48107 );
xor ( n48551 , n48550 , n48110 );
and ( n48552 , n48548 , n48551 );
and ( n48553 , n48544 , n48551 );
or ( n48554 , n48549 , n48552 , n48553 );
and ( n48555 , n45138 , n40053 );
and ( n48556 , n45151 , n40051 );
nor ( n48557 , n48555 , n48556 );
xnor ( n48558 , n48557 , n39999 );
and ( n48559 , n48554 , n48558 );
xor ( n48560 , n48113 , n48117 );
xor ( n48561 , n48560 , n48120 );
and ( n48562 , n48558 , n48561 );
and ( n48563 , n48554 , n48561 );
or ( n48564 , n48559 , n48562 , n48563 );
and ( n48565 , n45151 , n40053 );
and ( n48566 , n45164 , n40051 );
nor ( n48567 , n48565 , n48566 );
xnor ( n48568 , n48567 , n39999 );
xor ( n48569 , n48564 , n48568 );
xor ( n48570 , n48123 , n48127 );
xor ( n48571 , n48570 , n48130 );
xor ( n48572 , n48569 , n48571 );
and ( n48573 , n48438 , n48572 );
and ( n48574 , n48436 , n48572 );
or ( n48575 , n48439 , n48573 , n48574 );
and ( n48576 , n44357 , n40746 );
and ( n48577 , n44347 , n40744 );
nor ( n48578 , n48576 , n48577 );
xnor ( n48579 , n48578 , n40501 );
and ( n48580 , n48575 , n48579 );
and ( n48581 , n45164 , n40053 );
and ( n48582 , n44665 , n40051 );
nor ( n48583 , n48581 , n48582 );
xnor ( n48584 , n48583 , n39999 );
buf ( n48585 , n557801 );
not ( n48586 , n48585 );
xor ( n48587 , n48584 , n48586 );
xor ( n48588 , n48133 , n48137 );
xor ( n48589 , n48588 , n48140 );
xor ( n48590 , n48587 , n48589 );
and ( n48591 , n48579 , n48590 );
and ( n48592 , n48575 , n48590 );
or ( n48593 , n48580 , n48591 , n48592 );
and ( n48594 , n48584 , n48586 );
and ( n48595 , n48586 , n48589 );
and ( n48596 , n48584 , n48589 );
or ( n48597 , n48594 , n48595 , n48596 );
and ( n48598 , n44458 , n40527 );
and ( n48599 , n44357 , n40525 );
nor ( n48600 , n48598 , n48599 );
xnor ( n48601 , n48600 , n40382 );
xor ( n48602 , n48597 , n48601 );
buf ( n48603 , n557800 );
not ( n48604 , n48603 );
xor ( n48605 , n48602 , n48604 );
and ( n48606 , n48593 , n48605 );
and ( n48607 , n48564 , n48568 );
and ( n48608 , n48568 , n48571 );
and ( n48609 , n48564 , n48571 );
or ( n48610 , n48607 , n48608 , n48609 );
and ( n48611 , n44520 , n40527 );
and ( n48612 , n44458 , n40525 );
nor ( n48613 , n48611 , n48612 );
xnor ( n48614 , n48613 , n40382 );
and ( n48615 , n48610 , n48614 );
and ( n48616 , n44656 , n40258 );
and ( n48617 , n44565 , n40256 );
nor ( n48618 , n48616 , n48617 );
xnor ( n48619 , n48618 , n40169 );
and ( n48620 , n48614 , n48619 );
and ( n48621 , n48610 , n48619 );
or ( n48622 , n48615 , n48620 , n48621 );
and ( n48623 , n44347 , n40746 );
and ( n48624 , n44264 , n40744 );
nor ( n48625 , n48623 , n48624 );
xnor ( n48626 , n48625 , n40501 );
xor ( n48627 , n48622 , n48626 );
xor ( n48628 , n48355 , n48359 );
xor ( n48629 , n48628 , n48362 );
xor ( n48630 , n48627 , n48629 );
and ( n48631 , n48605 , n48630 );
and ( n48632 , n48593 , n48630 );
or ( n48633 , n48606 , n48631 , n48632 );
and ( n48634 , n43192 , n41292 );
and ( n48635 , n43073 , n41290 );
nor ( n48636 , n48634 , n48635 );
xnor ( n48637 , n48636 , n41041 );
and ( n48638 , n48633 , n48637 );
and ( n48639 , n48597 , n48601 );
and ( n48640 , n48601 , n48604 );
and ( n48641 , n48597 , n48604 );
or ( n48642 , n48639 , n48640 , n48641 );
and ( n48643 , n44264 , n40746 );
and ( n48644 , n43437 , n40744 );
nor ( n48645 , n48643 , n48644 );
xnor ( n48646 , n48645 , n40501 );
xor ( n48647 , n48642 , n48646 );
xor ( n48648 , n48246 , n48250 );
xor ( n48649 , n48648 , n48253 );
xor ( n48650 , n48647 , n48649 );
and ( n48651 , n48637 , n48650 );
and ( n48652 , n48633 , n48650 );
or ( n48653 , n48638 , n48651 , n48652 );
and ( n48654 , n48622 , n48626 );
and ( n48655 , n48626 , n48629 );
and ( n48656 , n48622 , n48629 );
or ( n48657 , n48654 , n48655 , n48656 );
and ( n48658 , n43428 , n41055 );
and ( n48659 , n43200 , n41053 );
nor ( n48660 , n48658 , n48659 );
xnor ( n48661 , n48660 , n40728 );
and ( n48662 , n48657 , n48661 );
xor ( n48663 , n48365 , n48369 );
xor ( n48664 , n48663 , n48372 );
and ( n48665 , n48661 , n48664 );
and ( n48666 , n48657 , n48664 );
or ( n48667 , n48662 , n48665 , n48666 );
and ( n48668 , n48653 , n48667 );
xor ( n48669 , n48375 , n48377 );
xor ( n48670 , n48669 , n48380 );
and ( n48671 , n48667 , n48670 );
and ( n48672 , n48653 , n48670 );
or ( n48673 , n48668 , n48671 , n48672 );
and ( n48674 , n42811 , n41622 );
and ( n48675 , n42456 , n41620 );
nor ( n48676 , n48674 , n48675 );
xnor ( n48677 , n48676 , n41194 );
and ( n48678 , n48673 , n48677 );
xor ( n48679 , n48383 , n48387 );
xor ( n48680 , n48679 , n48392 );
and ( n48681 , n48677 , n48680 );
and ( n48682 , n48673 , n48680 );
or ( n48683 , n48678 , n48681 , n48682 );
and ( n48684 , n41807 , n42269 );
and ( n48685 , n41692 , n42266 );
nor ( n48686 , n48684 , n48685 );
xnor ( n48687 , n48686 , n41684 );
and ( n48688 , n48683 , n48687 );
xor ( n48689 , n48395 , n48399 );
xor ( n48690 , n48689 , n48402 );
and ( n48691 , n48687 , n48690 );
and ( n48692 , n48683 , n48690 );
or ( n48693 , n48688 , n48691 , n48692 );
and ( n48694 , n48642 , n48646 );
and ( n48695 , n48646 , n48649 );
and ( n48696 , n48642 , n48649 );
or ( n48697 , n48694 , n48695 , n48696 );
and ( n48698 , n43200 , n41055 );
and ( n48699 , n43192 , n41053 );
nor ( n48700 , n48698 , n48699 );
xnor ( n48701 , n48700 , n40728 );
and ( n48702 , n48697 , n48701 );
and ( n48703 , n43437 , n40746 );
and ( n48704 , n43428 , n40744 );
nor ( n48705 , n48703 , n48704 );
xnor ( n48706 , n48705 , n40501 );
and ( n48707 , n48701 , n48706 );
and ( n48708 , n48697 , n48706 );
or ( n48709 , n48702 , n48707 , n48708 );
and ( n48710 , n43027 , n41292 );
and ( n48711 , n43019 , n41290 );
nor ( n48712 , n48710 , n48711 );
xnor ( n48713 , n48712 , n41041 );
and ( n48714 , n48709 , n48713 );
xor ( n48715 , n48266 , n48268 );
xor ( n48716 , n48715 , n48271 );
and ( n48717 , n48713 , n48716 );
and ( n48718 , n48709 , n48716 );
or ( n48719 , n48714 , n48717 , n48718 );
and ( n48720 , n42456 , n41622 );
and ( n48721 , n42048 , n41620 );
nor ( n48722 , n48720 , n48721 );
xnor ( n48723 , n48722 , n41194 );
and ( n48724 , n48719 , n48723 );
xor ( n48725 , n48274 , n48278 );
xor ( n48726 , n48725 , n48281 );
and ( n48727 , n48723 , n48726 );
and ( n48728 , n48719 , n48726 );
or ( n48729 , n48724 , n48727 , n48728 );
and ( n48730 , n48693 , n48729 );
xor ( n48731 , n48405 , n48409 );
xor ( n48732 , n48731 , n48412 );
and ( n48733 , n48729 , n48732 );
and ( n48734 , n48693 , n48732 );
or ( n48735 , n48730 , n48733 , n48734 );
xor ( n48736 , n48351 , n48415 );
xor ( n48737 , n48736 , n48418 );
and ( n48738 , n48735 , n48737 );
xor ( n48739 , n48308 , n48312 );
xor ( n48740 , n48739 , n48315 );
and ( n48741 , n48737 , n48740 );
and ( n48742 , n48735 , n48740 );
or ( n48743 , n48738 , n48741 , n48742 );
and ( n48744 , n48432 , n48743 );
xor ( n48745 , n48735 , n48737 );
xor ( n48746 , n48745 , n48740 );
and ( n48747 , n43019 , n41622 );
and ( n48748 , n42811 , n41620 );
nor ( n48749 , n48747 , n48748 );
xnor ( n48750 , n48749 , n41194 );
and ( n48751 , n43073 , n41292 );
and ( n48752 , n43027 , n41290 );
nor ( n48753 , n48751 , n48752 );
xnor ( n48754 , n48753 , n41041 );
and ( n48755 , n48750 , n48754 );
xor ( n48756 , n48697 , n48701 );
xor ( n48757 , n48756 , n48706 );
and ( n48758 , n48754 , n48757 );
and ( n48759 , n48750 , n48757 );
or ( n48760 , n48755 , n48758 , n48759 );
xor ( n48761 , n48673 , n48677 );
xor ( n48762 , n48761 , n48680 );
and ( n48763 , n48760 , n48762 );
xor ( n48764 , n48709 , n48713 );
xor ( n48765 , n48764 , n48716 );
and ( n48766 , n48762 , n48765 );
and ( n48767 , n48760 , n48765 );
or ( n48768 , n48763 , n48766 , n48767 );
and ( n48769 , n42061 , n41984 );
and ( n48770 , n41816 , n41982 );
nor ( n48771 , n48769 , n48770 );
xnor ( n48772 , n48771 , n41687 );
and ( n48773 , n48768 , n48772 );
xor ( n48774 , n48719 , n48723 );
xor ( n48775 , n48774 , n48726 );
and ( n48776 , n48772 , n48775 );
and ( n48777 , n48768 , n48775 );
or ( n48778 , n48773 , n48776 , n48777 );
xor ( n48779 , n48341 , n48345 );
xor ( n48780 , n48779 , n48348 );
and ( n48781 , n48778 , n48780 );
xor ( n48782 , n48693 , n48729 );
xor ( n48783 , n48782 , n48732 );
and ( n48784 , n48780 , n48783 );
and ( n48785 , n48778 , n48783 );
or ( n48786 , n48781 , n48784 , n48785 );
and ( n48787 , n48746 , n48786 );
xor ( n48788 , n48778 , n48780 );
xor ( n48789 , n48788 , n48783 );
and ( n48790 , n45164 , n40258 );
and ( n48791 , n44665 , n40256 );
nor ( n48792 , n48790 , n48791 );
xnor ( n48793 , n48792 , n40169 );
buf ( n48794 , n557803 );
not ( n48795 , n48794 );
and ( n48796 , n48793 , n48795 );
xor ( n48797 , n48554 , n48558 );
xor ( n48798 , n48797 , n48561 );
and ( n48799 , n48795 , n48798 );
and ( n48800 , n48793 , n48798 );
or ( n48801 , n48796 , n48799 , n48800 );
and ( n48802 , n44565 , n40527 );
and ( n48803 , n44520 , n40525 );
nor ( n48804 , n48802 , n48803 );
xnor ( n48805 , n48804 , n40382 );
and ( n48806 , n48801 , n48805 );
xor ( n48807 , n48436 , n48438 );
xor ( n48808 , n48807 , n48572 );
and ( n48809 , n48805 , n48808 );
and ( n48810 , n48801 , n48808 );
or ( n48811 , n48806 , n48809 , n48810 );
xor ( n48812 , n48610 , n48614 );
xor ( n48813 , n48812 , n48619 );
and ( n48814 , n48811 , n48813 );
xor ( n48815 , n48575 , n48579 );
xor ( n48816 , n48815 , n48590 );
and ( n48817 , n48813 , n48816 );
and ( n48818 , n48811 , n48816 );
or ( n48819 , n48814 , n48817 , n48818 );
and ( n48820 , n43200 , n41292 );
and ( n48821 , n43192 , n41290 );
nor ( n48822 , n48820 , n48821 );
xnor ( n48823 , n48822 , n41041 );
and ( n48824 , n48819 , n48823 );
and ( n48825 , n43437 , n41055 );
and ( n48826 , n43428 , n41053 );
nor ( n48827 , n48825 , n48826 );
xnor ( n48828 , n48827 , n40728 );
and ( n48829 , n48823 , n48828 );
and ( n48830 , n48819 , n48828 );
or ( n48831 , n48824 , n48829 , n48830 );
and ( n48832 , n43027 , n41622 );
and ( n48833 , n43019 , n41620 );
nor ( n48834 , n48832 , n48833 );
xnor ( n48835 , n48834 , n41194 );
and ( n48836 , n48831 , n48835 );
xor ( n48837 , n48657 , n48661 );
xor ( n48838 , n48837 , n48664 );
and ( n48839 , n48835 , n48838 );
and ( n48840 , n48831 , n48838 );
or ( n48841 , n48836 , n48839 , n48840 );
xor ( n48842 , n48750 , n48754 );
xor ( n48843 , n48842 , n48757 );
and ( n48844 , n48841 , n48843 );
xor ( n48845 , n48653 , n48667 );
xor ( n48846 , n48845 , n48670 );
and ( n48847 , n48843 , n48846 );
and ( n48848 , n48841 , n48846 );
or ( n48849 , n48844 , n48847 , n48848 );
and ( n48850 , n41816 , n42269 );
and ( n48851 , n41807 , n42266 );
nor ( n48852 , n48850 , n48851 );
xnor ( n48853 , n48852 , n41684 );
and ( n48854 , n48849 , n48853 );
and ( n48855 , n42048 , n41984 );
and ( n48856 , n42061 , n41982 );
nor ( n48857 , n48855 , n48856 );
xnor ( n48858 , n48857 , n41687 );
and ( n48859 , n48853 , n48858 );
and ( n48860 , n48849 , n48858 );
or ( n48861 , n48854 , n48859 , n48860 );
xor ( n48862 , n48683 , n48687 );
xor ( n48863 , n48862 , n48690 );
and ( n48864 , n48861 , n48863 );
xor ( n48865 , n48768 , n48772 );
xor ( n48866 , n48865 , n48775 );
and ( n48867 , n48863 , n48866 );
and ( n48868 , n48861 , n48866 );
or ( n48869 , n48864 , n48867 , n48868 );
and ( n48870 , n48789 , n48869 );
and ( n48871 , n45151 , n40258 );
and ( n48872 , n45164 , n40256 );
nor ( n48873 , n48871 , n48872 );
xnor ( n48874 , n48873 , n40169 );
buf ( n48875 , n557804 );
not ( n48876 , n48875 );
and ( n48877 , n48874 , n48876 );
xor ( n48878 , n48544 , n48548 );
xor ( n48879 , n48878 , n48551 );
and ( n48880 , n48876 , n48879 );
and ( n48881 , n48874 , n48879 );
or ( n48882 , n48877 , n48880 , n48881 );
and ( n48883 , n44656 , n40527 );
and ( n48884 , n44565 , n40525 );
nor ( n48885 , n48883 , n48884 );
xnor ( n48886 , n48885 , n40382 );
and ( n48887 , n48882 , n48886 );
xor ( n48888 , n48793 , n48795 );
xor ( n48889 , n48888 , n48798 );
and ( n48890 , n48886 , n48889 );
and ( n48891 , n48882 , n48889 );
or ( n48892 , n48887 , n48890 , n48891 );
and ( n48893 , n44347 , n41055 );
and ( n48894 , n44264 , n41053 );
nor ( n48895 , n48893 , n48894 );
xnor ( n48896 , n48895 , n40728 );
and ( n48897 , n48892 , n48896 );
and ( n48898 , n44458 , n40746 );
and ( n48899 , n44357 , n40744 );
nor ( n48900 , n48898 , n48899 );
xnor ( n48901 , n48900 , n40501 );
and ( n48902 , n48896 , n48901 );
and ( n48903 , n48892 , n48901 );
or ( n48904 , n48897 , n48902 , n48903 );
and ( n48905 , n43428 , n41292 );
and ( n48906 , n43200 , n41290 );
nor ( n48907 , n48905 , n48906 );
xnor ( n48908 , n48907 , n41041 );
and ( n48909 , n48904 , n48908 );
and ( n48910 , n44264 , n41055 );
and ( n48911 , n43437 , n41053 );
nor ( n48912 , n48910 , n48911 );
xnor ( n48913 , n48912 , n40728 );
and ( n48914 , n48908 , n48913 );
and ( n48915 , n48904 , n48913 );
or ( n48916 , n48909 , n48914 , n48915 );
xor ( n48917 , n48819 , n48823 );
xor ( n48918 , n48917 , n48828 );
and ( n48919 , n48916 , n48918 );
xor ( n48920 , n48593 , n48605 );
xor ( n48921 , n48920 , n48630 );
and ( n48922 , n48918 , n48921 );
and ( n48923 , n48916 , n48921 );
or ( n48924 , n48919 , n48922 , n48923 );
and ( n48925 , n42811 , n41984 );
and ( n48926 , n42456 , n41982 );
nor ( n48927 , n48925 , n48926 );
xnor ( n48928 , n48927 , n41687 );
and ( n48929 , n48924 , n48928 );
xor ( n48930 , n48633 , n48637 );
xor ( n48931 , n48930 , n48650 );
and ( n48932 , n48928 , n48931 );
and ( n48933 , n48924 , n48931 );
or ( n48934 , n48929 , n48932 , n48933 );
and ( n48935 , n42061 , n42269 );
and ( n48936 , n41816 , n42266 );
nor ( n48937 , n48935 , n48936 );
xnor ( n48938 , n48937 , n41684 );
and ( n48939 , n48934 , n48938 );
and ( n48940 , n42456 , n41984 );
and ( n48941 , n42048 , n41982 );
nor ( n48942 , n48940 , n48941 );
xnor ( n48943 , n48942 , n41687 );
and ( n48944 , n48938 , n48943 );
and ( n48945 , n48934 , n48943 );
or ( n48946 , n48939 , n48944 , n48945 );
xor ( n48947 , n48849 , n48853 );
xor ( n48948 , n48947 , n48858 );
and ( n48949 , n48946 , n48948 );
xor ( n48950 , n48760 , n48762 );
xor ( n48951 , n48950 , n48765 );
and ( n48952 , n48948 , n48951 );
and ( n48953 , n48946 , n48951 );
or ( n48954 , n48949 , n48952 , n48953 );
xor ( n48955 , n48861 , n48863 );
xor ( n48956 , n48955 , n48866 );
and ( n48957 , n48954 , n48956 );
and ( n48958 , n42048 , n42269 );
and ( n48959 , n42061 , n42266 );
nor ( n48960 , n48958 , n48959 );
xnor ( n48961 , n48960 , n41684 );
and ( n48962 , n42456 , n42269 );
and ( n48963 , n42048 , n42266 );
nor ( n48964 , n48962 , n48963 );
xnor ( n48965 , n48964 , n41684 );
and ( n48966 , n43019 , n41984 );
and ( n48967 , n42811 , n41982 );
nor ( n48968 , n48966 , n48967 );
xnor ( n48969 , n48968 , n41687 );
and ( n48970 , n48965 , n48969 );
and ( n48971 , n43073 , n41622 );
and ( n48972 , n43027 , n41620 );
nor ( n48973 , n48971 , n48972 );
xnor ( n48974 , n48973 , n41194 );
and ( n48975 , n48969 , n48974 );
and ( n48976 , n48965 , n48974 );
or ( n48977 , n48970 , n48975 , n48976 );
and ( n48978 , n48961 , n48977 );
and ( n48979 , n42811 , n42269 );
and ( n48980 , n42456 , n42266 );
nor ( n48981 , n48979 , n48980 );
xnor ( n48982 , n48981 , n41684 );
and ( n48983 , n43027 , n41984 );
and ( n48984 , n43019 , n41982 );
nor ( n48985 , n48983 , n48984 );
xnor ( n48986 , n48985 , n41687 );
and ( n48987 , n48982 , n48986 );
xor ( n48988 , n48965 , n48969 );
xor ( n48989 , n48988 , n48974 );
and ( n48990 , n48987 , n48989 );
and ( n48991 , n43192 , n41622 );
and ( n48992 , n43073 , n41620 );
nor ( n48993 , n48991 , n48992 );
xnor ( n48994 , n48993 , n41194 );
xor ( n48995 , n48982 , n48986 );
and ( n48996 , n48994 , n48995 );
and ( n48997 , n43019 , n42269 );
and ( n48998 , n42811 , n42266 );
nor ( n48999 , n48997 , n48998 );
xnor ( n49000 , n48999 , n41684 );
and ( n49001 , n43073 , n41984 );
and ( n49002 , n43027 , n41982 );
nor ( n49003 , n49001 , n49002 );
xnor ( n49004 , n49003 , n41687 );
and ( n49005 , n49000 , n49004 );
and ( n49006 , n43200 , n41622 );
and ( n49007 , n43192 , n41620 );
nor ( n49008 , n49006 , n49007 );
xnor ( n49009 , n49008 , n41194 );
and ( n49010 , n49004 , n49009 );
and ( n49011 , n49000 , n49009 );
or ( n49012 , n49005 , n49010 , n49011 );
and ( n49013 , n48995 , n49012 );
and ( n49014 , n48994 , n49012 );
or ( n49015 , n48996 , n49013 , n49014 );
and ( n49016 , n48989 , n49015 );
and ( n49017 , n48987 , n49015 );
or ( n49018 , n48990 , n49016 , n49017 );
and ( n49019 , n48977 , n49018 );
and ( n49020 , n48961 , n49018 );
or ( n49021 , n48978 , n49019 , n49020 );
xor ( n49022 , n48841 , n48843 );
xor ( n49023 , n49022 , n48846 );
and ( n49024 , n49021 , n49023 );
xor ( n49025 , n48961 , n48977 );
xor ( n49026 , n49025 , n49018 );
xor ( n49027 , n48831 , n48835 );
xor ( n49028 , n49027 , n48838 );
and ( n49029 , n49026 , n49028 );
xor ( n49030 , n48987 , n48989 );
xor ( n49031 , n49030 , n49015 );
and ( n49032 , n43437 , n41292 );
and ( n49033 , n43428 , n41290 );
nor ( n49034 , n49032 , n49033 );
xnor ( n49035 , n49034 , n41041 );
and ( n49036 , n43027 , n42269 );
and ( n49037 , n43019 , n42266 );
nor ( n49038 , n49036 , n49037 );
xnor ( n49039 , n49038 , n41684 );
and ( n49040 , n43192 , n41984 );
and ( n49041 , n43073 , n41982 );
nor ( n49042 , n49040 , n49041 );
xnor ( n49043 , n49042 , n41687 );
and ( n49044 , n49039 , n49043 );
and ( n49045 , n43428 , n41622 );
and ( n49046 , n43200 , n41620 );
nor ( n49047 , n49045 , n49046 );
xnor ( n49048 , n49047 , n41194 );
and ( n49049 , n49043 , n49048 );
and ( n49050 , n49039 , n49048 );
or ( n49051 , n49044 , n49049 , n49050 );
and ( n49052 , n49035 , n49051 );
and ( n49053 , n44264 , n41292 );
and ( n49054 , n43437 , n41290 );
nor ( n49055 , n49053 , n49054 );
xnor ( n49056 , n49055 , n41041 );
and ( n49057 , n44357 , n41055 );
and ( n49058 , n44347 , n41053 );
nor ( n49059 , n49057 , n49058 );
xnor ( n49060 , n49059 , n40728 );
and ( n49061 , n49056 , n49060 );
and ( n49062 , n44520 , n40746 );
and ( n49063 , n44458 , n40744 );
nor ( n49064 , n49062 , n49063 );
xnor ( n49065 , n49064 , n40501 );
and ( n49066 , n49060 , n49065 );
and ( n49067 , n49056 , n49065 );
or ( n49068 , n49061 , n49066 , n49067 );
and ( n49069 , n49051 , n49068 );
and ( n49070 , n49035 , n49068 );
or ( n49071 , n49052 , n49069 , n49070 );
xor ( n49072 , n48994 , n48995 );
xor ( n49073 , n49072 , n49012 );
and ( n49074 , n49071 , n49073 );
xor ( n49075 , n49000 , n49004 );
xor ( n49076 , n49075 , n49009 );
and ( n49077 , n43073 , n42269 );
and ( n49078 , n43027 , n42266 );
nor ( n49079 , n49077 , n49078 );
xnor ( n49080 , n49079 , n41684 );
and ( n49081 , n43200 , n41984 );
and ( n49082 , n43192 , n41982 );
nor ( n49083 , n49081 , n49082 );
xnor ( n49084 , n49083 , n41687 );
and ( n49085 , n49080 , n49084 );
and ( n49086 , n43437 , n41622 );
and ( n49087 , n43428 , n41620 );
nor ( n49088 , n49086 , n49087 );
xnor ( n49089 , n49088 , n41194 );
and ( n49090 , n49084 , n49089 );
and ( n49091 , n49080 , n49089 );
or ( n49092 , n49085 , n49090 , n49091 );
and ( n49093 , n44347 , n41292 );
and ( n49094 , n44264 , n41290 );
nor ( n49095 , n49093 , n49094 );
xnor ( n49096 , n49095 , n41041 );
and ( n49097 , n44458 , n41055 );
and ( n49098 , n44357 , n41053 );
nor ( n49099 , n49097 , n49098 );
xnor ( n49100 , n49099 , n40728 );
and ( n49101 , n49096 , n49100 );
and ( n49102 , n44565 , n40746 );
and ( n49103 , n44520 , n40744 );
nor ( n49104 , n49102 , n49103 );
xnor ( n49105 , n49104 , n40501 );
and ( n49106 , n49100 , n49105 );
and ( n49107 , n49096 , n49105 );
or ( n49108 , n49101 , n49106 , n49107 );
and ( n49109 , n49092 , n49108 );
xor ( n49110 , n49039 , n49043 );
xor ( n49111 , n49110 , n49048 );
and ( n49112 , n49108 , n49111 );
and ( n49113 , n49092 , n49111 );
or ( n49114 , n49109 , n49112 , n49113 );
and ( n49115 , n49076 , n49114 );
xor ( n49116 , n49035 , n49051 );
xor ( n49117 , n49116 , n49068 );
and ( n49118 , n49114 , n49117 );
and ( n49119 , n49076 , n49117 );
or ( n49120 , n49115 , n49118 , n49119 );
and ( n49121 , n49073 , n49120 );
and ( n49122 , n49071 , n49120 );
or ( n49123 , n49074 , n49121 , n49122 );
and ( n49124 , n49031 , n49123 );
xor ( n49125 , n49071 , n49073 );
xor ( n49126 , n49125 , n49120 );
xor ( n49127 , n49056 , n49060 );
xor ( n49128 , n49127 , n49065 );
and ( n49129 , n44665 , n40527 );
and ( n49130 , n44656 , n40525 );
nor ( n49131 , n49129 , n49130 );
xnor ( n49132 , n49131 , n40382 );
and ( n49133 , n43192 , n42269 );
and ( n49134 , n43073 , n42266 );
nor ( n49135 , n49133 , n49134 );
xnor ( n49136 , n49135 , n41684 );
and ( n49137 , n43428 , n41984 );
and ( n49138 , n43200 , n41982 );
nor ( n49139 , n49137 , n49138 );
xnor ( n49140 , n49139 , n41687 );
and ( n49141 , n49136 , n49140 );
and ( n49142 , n44264 , n41622 );
and ( n49143 , n43437 , n41620 );
nor ( n49144 , n49142 , n49143 );
xnor ( n49145 , n49144 , n41194 );
and ( n49146 , n49140 , n49145 );
and ( n49147 , n49136 , n49145 );
or ( n49148 , n49141 , n49146 , n49147 );
and ( n49149 , n49132 , n49148 );
and ( n49150 , n44357 , n41292 );
and ( n49151 , n44347 , n41290 );
nor ( n49152 , n49150 , n49151 );
xnor ( n49153 , n49152 , n41041 );
and ( n49154 , n44520 , n41055 );
and ( n49155 , n44458 , n41053 );
nor ( n49156 , n49154 , n49155 );
xnor ( n49157 , n49156 , n40728 );
and ( n49158 , n49153 , n49157 );
and ( n49159 , n44656 , n40746 );
and ( n49160 , n44565 , n40744 );
nor ( n49161 , n49159 , n49160 );
xnor ( n49162 , n49161 , n40501 );
and ( n49163 , n49157 , n49162 );
and ( n49164 , n49153 , n49162 );
or ( n49165 , n49158 , n49163 , n49164 );
and ( n49166 , n49148 , n49165 );
and ( n49167 , n49132 , n49165 );
or ( n49168 , n49149 , n49166 , n49167 );
and ( n49169 , n49128 , n49168 );
xor ( n49170 , n49092 , n49108 );
xor ( n49171 , n49170 , n49111 );
and ( n49172 , n49168 , n49171 );
and ( n49173 , n49128 , n49171 );
or ( n49174 , n49169 , n49172 , n49173 );
xor ( n49175 , n49076 , n49114 );
xor ( n49176 , n49175 , n49117 );
and ( n49177 , n49174 , n49176 );
xor ( n49178 , n49080 , n49084 );
xor ( n49179 , n49178 , n49089 );
xor ( n49180 , n49096 , n49100 );
xor ( n49181 , n49180 , n49105 );
and ( n49182 , n49179 , n49181 );
and ( n49183 , n45164 , n40527 );
and ( n49184 , n44665 , n40525 );
nor ( n49185 , n49183 , n49184 );
xnor ( n49186 , n49185 , n40382 );
buf ( n49187 , n557805 );
not ( n49188 , n49187 );
and ( n49189 , n49186 , n49188 );
and ( n49190 , n45151 , n40527 );
and ( n49191 , n45164 , n40525 );
nor ( n49192 , n49190 , n49191 );
xnor ( n49193 , n49192 , n40382 );
buf ( n49194 , n557806 );
not ( n49195 , n49194 );
and ( n49196 , n49193 , n49195 );
and ( n49197 , n49188 , n49196 );
and ( n49198 , n49186 , n49196 );
or ( n49199 , n49189 , n49197 , n49198 );
and ( n49200 , n49181 , n49199 );
and ( n49201 , n49179 , n49199 );
or ( n49202 , n49182 , n49200 , n49201 );
xor ( n49203 , n49128 , n49168 );
xor ( n49204 , n49203 , n49171 );
and ( n49205 , n49202 , n49204 );
and ( n49206 , n43200 , n42269 );
and ( n49207 , n43192 , n42266 );
nor ( n49208 , n49206 , n49207 );
xnor ( n49209 , n49208 , n41684 );
and ( n49210 , n43437 , n41984 );
and ( n49211 , n43428 , n41982 );
nor ( n49212 , n49210 , n49211 );
xnor ( n49213 , n49212 , n41687 );
and ( n49214 , n49209 , n49213 );
and ( n49215 , n44347 , n41622 );
and ( n49216 , n44264 , n41620 );
nor ( n49217 , n49215 , n49216 );
xnor ( n49218 , n49217 , n41194 );
and ( n49219 , n49213 , n49218 );
and ( n49220 , n49209 , n49218 );
or ( n49221 , n49214 , n49219 , n49220 );
and ( n49222 , n44458 , n41292 );
and ( n49223 , n44357 , n41290 );
nor ( n49224 , n49222 , n49223 );
xnor ( n49225 , n49224 , n41041 );
and ( n49226 , n44565 , n41055 );
and ( n49227 , n44520 , n41053 );
nor ( n49228 , n49226 , n49227 );
xnor ( n49229 , n49228 , n40728 );
and ( n49230 , n49225 , n49229 );
and ( n49231 , n44665 , n40746 );
and ( n49232 , n44656 , n40744 );
nor ( n49233 , n49231 , n49232 );
xnor ( n49234 , n49233 , n40501 );
and ( n49235 , n49229 , n49234 );
and ( n49236 , n49225 , n49234 );
or ( n49237 , n49230 , n49235 , n49236 );
and ( n49238 , n49221 , n49237 );
xor ( n49239 , n49136 , n49140 );
xor ( n49240 , n49239 , n49145 );
and ( n49241 , n49237 , n49240 );
and ( n49242 , n49221 , n49240 );
or ( n49243 , n49238 , n49241 , n49242 );
xor ( n49244 , n49132 , n49148 );
xor ( n49245 , n49244 , n49165 );
and ( n49246 , n49243 , n49245 );
xor ( n49247 , n49153 , n49157 );
xor ( n49248 , n49247 , n49162 );
xor ( n49249 , n49193 , n49195 );
and ( n49250 , n43428 , n42269 );
and ( n49251 , n43200 , n42266 );
nor ( n49252 , n49250 , n49251 );
xnor ( n49253 , n49252 , n41684 );
and ( n49254 , n44264 , n41984 );
and ( n49255 , n43437 , n41982 );
nor ( n49256 , n49254 , n49255 );
xnor ( n49257 , n49256 , n41687 );
and ( n49258 , n49253 , n49257 );
and ( n49259 , n44357 , n41622 );
and ( n49260 , n44347 , n41620 );
nor ( n49261 , n49259 , n49260 );
xnor ( n49262 , n49261 , n41194 );
and ( n49263 , n49257 , n49262 );
and ( n49264 , n49253 , n49262 );
or ( n49265 , n49258 , n49263 , n49264 );
and ( n49266 , n49249 , n49265 );
and ( n49267 , n44520 , n41292 );
and ( n49268 , n44458 , n41290 );
nor ( n49269 , n49267 , n49268 );
xnor ( n49270 , n49269 , n41041 );
and ( n49271 , n44656 , n41055 );
and ( n49272 , n44565 , n41053 );
nor ( n49273 , n49271 , n49272 );
xnor ( n49274 , n49273 , n40728 );
and ( n49275 , n49270 , n49274 );
and ( n49276 , n45164 , n40746 );
and ( n49277 , n44665 , n40744 );
nor ( n49278 , n49276 , n49277 );
xnor ( n49279 , n49278 , n40501 );
and ( n49280 , n49274 , n49279 );
and ( n49281 , n49270 , n49279 );
or ( n49282 , n49275 , n49280 , n49281 );
and ( n49283 , n49265 , n49282 );
and ( n49284 , n49249 , n49282 );
or ( n49285 , n49266 , n49283 , n49284 );
and ( n49286 , n49248 , n49285 );
xor ( n49287 , n49186 , n49188 );
xor ( n49288 , n49287 , n49196 );
and ( n49289 , n49285 , n49288 );
and ( n49290 , n49248 , n49288 );
or ( n49291 , n49286 , n49289 , n49290 );
and ( n49292 , n49245 , n49291 );
and ( n49293 , n49243 , n49291 );
or ( n49294 , n49246 , n49292 , n49293 );
and ( n49295 , n49204 , n49294 );
and ( n49296 , n49202 , n49294 );
or ( n49297 , n49205 , n49295 , n49296 );
and ( n49298 , n49176 , n49297 );
and ( n49299 , n49174 , n49297 );
or ( n49300 , n49177 , n49298 , n49299 );
and ( n49301 , n49126 , n49300 );
xor ( n49302 , n48904 , n48908 );
xor ( n49303 , n49302 , n48913 );
and ( n49304 , n49300 , n49303 );
and ( n49305 , n49126 , n49303 );
or ( n49306 , n49301 , n49304 , n49305 );
and ( n49307 , n49123 , n49306 );
and ( n49308 , n49031 , n49306 );
or ( n49309 , n49124 , n49307 , n49308 );
and ( n49310 , n49028 , n49309 );
and ( n49311 , n49026 , n49309 );
or ( n49312 , n49029 , n49310 , n49311 );
and ( n49313 , n49023 , n49312 );
and ( n49314 , n49021 , n49312 );
or ( n49315 , n49024 , n49313 , n49314 );
xor ( n49316 , n48946 , n48948 );
xor ( n49317 , n49316 , n48951 );
and ( n49318 , n49315 , n49317 );
xor ( n49319 , n48934 , n48938 );
xor ( n49320 , n49319 , n48943 );
xor ( n49321 , n48924 , n48928 );
xor ( n49322 , n49321 , n48931 );
xor ( n49323 , n48916 , n48918 );
xor ( n49324 , n49323 , n48921 );
xor ( n49325 , n48811 , n48813 );
xor ( n49326 , n49325 , n48816 );
xor ( n49327 , n49174 , n49176 );
xor ( n49328 , n49327 , n49297 );
xor ( n49329 , n49179 , n49181 );
xor ( n49330 , n49329 , n49199 );
xor ( n49331 , n49221 , n49237 );
xor ( n49332 , n49331 , n49240 );
xor ( n49333 , n49209 , n49213 );
xor ( n49334 , n49333 , n49218 );
xor ( n49335 , n49225 , n49229 );
xor ( n49336 , n49335 , n49234 );
and ( n49337 , n49334 , n49336 );
and ( n49338 , n45138 , n40527 );
and ( n49339 , n45151 , n40525 );
nor ( n49340 , n49338 , n49339 );
xnor ( n49341 , n49340 , n40382 );
buf ( n49342 , n557807 );
not ( n49343 , n49342 );
and ( n49344 , n49341 , n49343 );
and ( n49345 , n45151 , n40746 );
and ( n49346 , n45164 , n40744 );
nor ( n49347 , n49345 , n49346 );
xnor ( n49348 , n49347 , n40501 );
buf ( n49349 , n557808 );
not ( n49350 , n49349 );
and ( n49351 , n49348 , n49350 );
and ( n49352 , n49343 , n49351 );
and ( n49353 , n49341 , n49351 );
or ( n49354 , n49344 , n49352 , n49353 );
and ( n49355 , n49336 , n49354 );
and ( n49356 , n49334 , n49354 );
or ( n49357 , n49337 , n49355 , n49356 );
and ( n49358 , n49332 , n49357 );
xor ( n49359 , n49248 , n49285 );
xor ( n49360 , n49359 , n49288 );
and ( n49361 , n49357 , n49360 );
and ( n49362 , n49332 , n49360 );
or ( n49363 , n49358 , n49361 , n49362 );
and ( n49364 , n49330 , n49363 );
xor ( n49365 , n49243 , n49245 );
xor ( n49366 , n49365 , n49291 );
and ( n49367 , n49363 , n49366 );
and ( n49368 , n49330 , n49366 );
or ( n49369 , n49364 , n49367 , n49368 );
xor ( n49370 , n49202 , n49204 );
xor ( n49371 , n49370 , n49294 );
and ( n49372 , n49369 , n49371 );
xor ( n49373 , n49330 , n49363 );
xor ( n49374 , n49373 , n49366 );
and ( n49375 , n43437 , n42269 );
and ( n49376 , n43428 , n42266 );
nor ( n49377 , n49375 , n49376 );
xnor ( n49378 , n49377 , n41684 );
and ( n49379 , n44347 , n41984 );
and ( n49380 , n44264 , n41982 );
nor ( n49381 , n49379 , n49380 );
xnor ( n49382 , n49381 , n41687 );
and ( n49383 , n49378 , n49382 );
and ( n49384 , n44458 , n41622 );
and ( n49385 , n44357 , n41620 );
nor ( n49386 , n49384 , n49385 );
xnor ( n49387 , n49386 , n41194 );
and ( n49388 , n49382 , n49387 );
and ( n49389 , n49378 , n49387 );
or ( n49390 , n49383 , n49388 , n49389 );
and ( n49391 , n44565 , n41292 );
and ( n49392 , n44520 , n41290 );
nor ( n49393 , n49391 , n49392 );
xnor ( n49394 , n49393 , n41041 );
and ( n49395 , n44665 , n41055 );
and ( n49396 , n44656 , n41053 );
nor ( n49397 , n49395 , n49396 );
xnor ( n49398 , n49397 , n40728 );
and ( n49399 , n49394 , n49398 );
and ( n49400 , n45125 , n40527 );
and ( n49401 , n45138 , n40525 );
nor ( n49402 , n49400 , n49401 );
xnor ( n49403 , n49402 , n40382 );
and ( n49404 , n49398 , n49403 );
and ( n49405 , n49394 , n49403 );
or ( n49406 , n49399 , n49404 , n49405 );
and ( n49407 , n49390 , n49406 );
xor ( n49408 , n49253 , n49257 );
xor ( n49409 , n49408 , n49262 );
and ( n49410 , n49406 , n49409 );
and ( n49411 , n49390 , n49409 );
or ( n49412 , n49407 , n49410 , n49411 );
xor ( n49413 , n49249 , n49265 );
xor ( n49414 , n49413 , n49282 );
and ( n49415 , n49412 , n49414 );
xor ( n49416 , n49270 , n49274 );
xor ( n49417 , n49416 , n49279 );
xor ( n49418 , n49348 , n49350 );
and ( n49419 , n44264 , n42269 );
and ( n49420 , n43437 , n42266 );
nor ( n49421 , n49419 , n49420 );
xnor ( n49422 , n49421 , n41684 );
and ( n49423 , n44357 , n41984 );
and ( n49424 , n44347 , n41982 );
nor ( n49425 , n49423 , n49424 );
xnor ( n49426 , n49425 , n41687 );
and ( n49427 , n49422 , n49426 );
and ( n49428 , n44520 , n41622 );
and ( n49429 , n44458 , n41620 );
nor ( n49430 , n49428 , n49429 );
xnor ( n49431 , n49430 , n41194 );
and ( n49432 , n49426 , n49431 );
and ( n49433 , n49422 , n49431 );
or ( n49434 , n49427 , n49432 , n49433 );
and ( n49435 , n49418 , n49434 );
and ( n49436 , n44656 , n41292 );
and ( n49437 , n44565 , n41290 );
nor ( n49438 , n49436 , n49437 );
xnor ( n49439 , n49438 , n41041 );
and ( n49440 , n45164 , n41055 );
and ( n49441 , n44665 , n41053 );
nor ( n49442 , n49440 , n49441 );
xnor ( n49443 , n49442 , n40728 );
and ( n49444 , n49439 , n49443 );
and ( n49445 , n45138 , n40746 );
and ( n49446 , n45151 , n40744 );
nor ( n49447 , n49445 , n49446 );
xnor ( n49448 , n49447 , n40501 );
and ( n49449 , n49443 , n49448 );
and ( n49450 , n49439 , n49448 );
or ( n49451 , n49444 , n49449 , n49450 );
and ( n49452 , n49434 , n49451 );
and ( n49453 , n49418 , n49451 );
or ( n49454 , n49435 , n49452 , n49453 );
and ( n49455 , n49417 , n49454 );
xor ( n49456 , n49341 , n49343 );
xor ( n49457 , n49456 , n49351 );
and ( n49458 , n49454 , n49457 );
and ( n49459 , n49417 , n49457 );
or ( n49460 , n49455 , n49458 , n49459 );
and ( n49461 , n49414 , n49460 );
and ( n49462 , n49412 , n49460 );
or ( n49463 , n49415 , n49461 , n49462 );
xor ( n49464 , n49332 , n49357 );
xor ( n49465 , n49464 , n49360 );
and ( n49466 , n49463 , n49465 );
xor ( n49467 , n49334 , n49336 );
xor ( n49468 , n49467 , n49354 );
xor ( n49469 , n49390 , n49406 );
xor ( n49470 , n49469 , n49409 );
xor ( n49471 , n49378 , n49382 );
xor ( n49472 , n49471 , n49387 );
xor ( n49473 , n49394 , n49398 );
xor ( n49474 , n49473 , n49403 );
and ( n49475 , n49472 , n49474 );
and ( n49476 , n45112 , n40527 );
and ( n49477 , n45125 , n40525 );
nor ( n49478 , n49476 , n49477 );
xnor ( n49479 , n49478 , n40382 );
buf ( n49480 , n557809 );
not ( n49481 , n49480 );
and ( n49482 , n49479 , n49481 );
and ( n49483 , n44347 , n42269 );
and ( n49484 , n44264 , n42266 );
nor ( n49485 , n49483 , n49484 );
xnor ( n49486 , n49485 , n41684 );
and ( n49487 , n44458 , n41984 );
and ( n49488 , n44357 , n41982 );
nor ( n49489 , n49487 , n49488 );
xnor ( n49490 , n49489 , n41687 );
and ( n49491 , n49486 , n49490 );
and ( n49492 , n44565 , n41622 );
and ( n49493 , n44520 , n41620 );
nor ( n49494 , n49492 , n49493 );
xnor ( n49495 , n49494 , n41194 );
and ( n49496 , n49490 , n49495 );
and ( n49497 , n49486 , n49495 );
or ( n49498 , n49491 , n49496 , n49497 );
and ( n49499 , n49481 , n49498 );
and ( n49500 , n49479 , n49498 );
or ( n49501 , n49482 , n49499 , n49500 );
and ( n49502 , n49474 , n49501 );
and ( n49503 , n49472 , n49501 );
or ( n49504 , n49475 , n49502 , n49503 );
and ( n49505 , n49470 , n49504 );
xor ( n49506 , n49417 , n49454 );
xor ( n49507 , n49506 , n49457 );
and ( n49508 , n49504 , n49507 );
and ( n49509 , n49470 , n49507 );
or ( n49510 , n49505 , n49508 , n49509 );
and ( n49511 , n49468 , n49510 );
xor ( n49512 , n49412 , n49414 );
xor ( n49513 , n49512 , n49460 );
and ( n49514 , n49510 , n49513 );
and ( n49515 , n49468 , n49513 );
or ( n49516 , n49511 , n49514 , n49515 );
and ( n49517 , n49465 , n49516 );
and ( n49518 , n49463 , n49516 );
or ( n49519 , n49466 , n49517 , n49518 );
and ( n49520 , n49374 , n49519 );
and ( n49521 , n45138 , n40258 );
and ( n49522 , n45151 , n40256 );
nor ( n49523 , n49521 , n49522 );
xnor ( n49524 , n49523 , n40169 );
xor ( n49525 , n48534 , n48538 );
xor ( n49526 , n49525 , n48541 );
and ( n49527 , n49524 , n49526 );
and ( n49528 , n49519 , n49527 );
and ( n49529 , n49374 , n49527 );
or ( n49530 , n49520 , n49528 , n49529 );
and ( n49531 , n49371 , n49530 );
and ( n49532 , n49369 , n49530 );
or ( n49533 , n49372 , n49531 , n49532 );
and ( n49534 , n49328 , n49533 );
xor ( n49535 , n48892 , n48896 );
xor ( n49536 , n49535 , n48901 );
and ( n49537 , n49533 , n49536 );
and ( n49538 , n49328 , n49536 );
or ( n49539 , n49534 , n49537 , n49538 );
and ( n49540 , n49326 , n49539 );
xor ( n49541 , n48801 , n48805 );
xor ( n49542 , n49541 , n48808 );
xor ( n49543 , n49463 , n49465 );
xor ( n49544 , n49543 , n49516 );
and ( n49545 , n45125 , n40258 );
and ( n49546 , n45138 , n40256 );
nor ( n49547 , n49545 , n49546 );
xnor ( n49548 , n49547 , n40169 );
xor ( n49549 , n48524 , n48528 );
xor ( n49550 , n49549 , n48531 );
and ( n49551 , n49548 , n49550 );
and ( n49552 , n49544 , n49551 );
xor ( n49553 , n49468 , n49510 );
xor ( n49554 , n49553 , n49513 );
and ( n49555 , n44665 , n41292 );
and ( n49556 , n44656 , n41290 );
nor ( n49557 , n49555 , n49556 );
xnor ( n49558 , n49557 , n41041 );
and ( n49559 , n45151 , n41055 );
and ( n49560 , n45164 , n41053 );
nor ( n49561 , n49559 , n49560 );
xnor ( n49562 , n49561 , n40728 );
and ( n49563 , n49558 , n49562 );
and ( n49564 , n45125 , n40746 );
and ( n49565 , n45138 , n40744 );
nor ( n49566 , n49564 , n49565 );
xnor ( n49567 , n49566 , n40501 );
and ( n49568 , n49562 , n49567 );
and ( n49569 , n49558 , n49567 );
or ( n49570 , n49563 , n49568 , n49569 );
and ( n49571 , n45099 , n40527 );
and ( n49572 , n45112 , n40525 );
nor ( n49573 , n49571 , n49572 );
xnor ( n49574 , n49573 , n40382 );
and ( n49575 , n45073 , n40258 );
and ( n49576 , n45086 , n40256 );
nor ( n49577 , n49575 , n49576 );
xnor ( n49578 , n49577 , n40169 );
and ( n49579 , n49574 , n49578 );
buf ( n49580 , n557810 );
not ( n49581 , n49580 );
and ( n49582 , n49578 , n49581 );
and ( n49583 , n49574 , n49581 );
or ( n49584 , n49579 , n49582 , n49583 );
and ( n49585 , n49570 , n49584 );
xor ( n49586 , n49422 , n49426 );
xor ( n49587 , n49586 , n49431 );
and ( n49588 , n49584 , n49587 );
and ( n49589 , n49570 , n49587 );
or ( n49590 , n49585 , n49588 , n49589 );
xor ( n49591 , n49418 , n49434 );
xor ( n49592 , n49591 , n49451 );
and ( n49593 , n49590 , n49592 );
xor ( n49594 , n49439 , n49443 );
xor ( n49595 , n49594 , n49448 );
and ( n49596 , n45138 , n41055 );
and ( n49597 , n45151 , n41053 );
nor ( n49598 , n49596 , n49597 );
xnor ( n49599 , n49598 , n40728 );
buf ( n49600 , n557811 );
not ( n49601 , n49600 );
and ( n49602 , n49599 , n49601 );
and ( n49603 , n44357 , n42269 );
and ( n49604 , n44347 , n42266 );
nor ( n49605 , n49603 , n49604 );
xnor ( n49606 , n49605 , n41684 );
and ( n49607 , n44520 , n41984 );
and ( n49608 , n44458 , n41982 );
nor ( n49609 , n49607 , n49608 );
xnor ( n49610 , n49609 , n41687 );
and ( n49611 , n49606 , n49610 );
and ( n49612 , n44656 , n41622 );
and ( n49613 , n44565 , n41620 );
nor ( n49614 , n49612 , n49613 );
xnor ( n49615 , n49614 , n41194 );
and ( n49616 , n49610 , n49615 );
and ( n49617 , n49606 , n49615 );
or ( n49618 , n49611 , n49616 , n49617 );
and ( n49619 , n49602 , n49618 );
and ( n49620 , n45164 , n41292 );
and ( n49621 , n44665 , n41290 );
nor ( n49622 , n49620 , n49621 );
xnor ( n49623 , n49622 , n41041 );
and ( n49624 , n45112 , n40746 );
and ( n49625 , n45125 , n40744 );
nor ( n49626 , n49624 , n49625 );
xnor ( n49627 , n49626 , n40501 );
and ( n49628 , n49623 , n49627 );
and ( n49629 , n45086 , n40527 );
and ( n49630 , n45099 , n40525 );
nor ( n49631 , n49629 , n49630 );
xnor ( n49632 , n49631 , n40382 );
and ( n49633 , n49627 , n49632 );
and ( n49634 , n49623 , n49632 );
or ( n49635 , n49628 , n49633 , n49634 );
and ( n49636 , n49618 , n49635 );
and ( n49637 , n49602 , n49635 );
or ( n49638 , n49619 , n49636 , n49637 );
and ( n49639 , n49595 , n49638 );
xor ( n49640 , n49486 , n49490 );
xor ( n49641 , n49640 , n49495 );
xor ( n49642 , n49558 , n49562 );
xor ( n49643 , n49642 , n49567 );
and ( n49644 , n49641 , n49643 );
xor ( n49645 , n49574 , n49578 );
xor ( n49646 , n49645 , n49581 );
and ( n49647 , n49643 , n49646 );
and ( n49648 , n49641 , n49646 );
or ( n49649 , n49644 , n49647 , n49648 );
and ( n49650 , n49638 , n49649 );
and ( n49651 , n49595 , n49649 );
or ( n49652 , n49639 , n49650 , n49651 );
and ( n49653 , n49592 , n49652 );
and ( n49654 , n49590 , n49652 );
or ( n49655 , n49593 , n49653 , n49654 );
xor ( n49656 , n49470 , n49504 );
xor ( n49657 , n49656 , n49507 );
and ( n49658 , n49655 , n49657 );
xor ( n49659 , n49472 , n49474 );
xor ( n49660 , n49659 , n49501 );
xor ( n49661 , n49479 , n49481 );
xor ( n49662 , n49661 , n49498 );
xor ( n49663 , n49570 , n49584 );
xor ( n49664 , n49663 , n49587 );
and ( n49665 , n49662 , n49664 );
and ( n49666 , n45060 , n40258 );
and ( n49667 , n45073 , n40256 );
nor ( n49668 , n49666 , n49667 );
xnor ( n49669 , n49668 , n40169 );
xor ( n49670 , n49599 , n49601 );
and ( n49671 , n49669 , n49670 );
and ( n49672 , n44458 , n42269 );
and ( n49673 , n44357 , n42266 );
nor ( n49674 , n49672 , n49673 );
xnor ( n49675 , n49674 , n41684 );
and ( n49676 , n44565 , n41984 );
and ( n49677 , n44520 , n41982 );
nor ( n49678 , n49676 , n49677 );
xnor ( n49679 , n49678 , n41687 );
and ( n576988 , n49675 , n49679 );
and ( n49680 , n44665 , n41622 );
and ( n49681 , n44656 , n41620 );
nor ( n49682 , n49680 , n49681 );
xnor ( n49683 , n49682 , n41194 );
and ( n49684 , n49679 , n49683 );
and ( n49685 , n49675 , n49683 );
or ( n49686 , n576988 , n49684 , n49685 );
and ( n49687 , n49670 , n49686 );
and ( n49688 , n49669 , n49686 );
or ( n49689 , n49671 , n49687 , n49688 );
and ( n49690 , n45151 , n41292 );
and ( n49691 , n45164 , n41290 );
nor ( n49692 , n49690 , n49691 );
xnor ( n49693 , n49692 , n41041 );
and ( n49694 , n45125 , n41055 );
and ( n49695 , n45138 , n41053 );
nor ( n49696 , n49694 , n49695 );
xnor ( n49697 , n49696 , n40728 );
and ( n49698 , n49693 , n49697 );
and ( n49699 , n45099 , n40746 );
and ( n49700 , n45112 , n40744 );
nor ( n49701 , n49699 , n49700 );
xnor ( n49702 , n49701 , n40501 );
and ( n49703 , n49697 , n49702 );
and ( n49704 , n49693 , n49702 );
or ( n49705 , n49698 , n49703 , n49704 );
and ( n49706 , n45073 , n40527 );
and ( n49707 , n45086 , n40525 );
nor ( n49708 , n49706 , n49707 );
xnor ( n49709 , n49708 , n40382 );
and ( n49710 , n45047 , n40258 );
and ( n49711 , n45060 , n40256 );
nor ( n49712 , n49710 , n49711 );
xnor ( n49713 , n49712 , n40169 );
and ( n49714 , n49709 , n49713 );
buf ( n49715 , n557812 );
not ( n49716 , n49715 );
and ( n49717 , n49713 , n49716 );
and ( n49718 , n49709 , n49716 );
or ( n49719 , n49714 , n49717 , n49718 );
and ( n49720 , n49705 , n49719 );
xor ( n49721 , n49606 , n49610 );
xor ( n49722 , n49721 , n49615 );
and ( n49723 , n49719 , n49722 );
and ( n49724 , n49705 , n49722 );
or ( n49725 , n49720 , n49723 , n49724 );
and ( n49726 , n49689 , n49725 );
xor ( n49727 , n49602 , n49618 );
xor ( n49728 , n49727 , n49635 );
and ( n49729 , n49725 , n49728 );
and ( n49730 , n49689 , n49728 );
or ( n49731 , n49726 , n49729 , n49730 );
and ( n49732 , n49664 , n49731 );
and ( n49733 , n49662 , n49731 );
or ( n49734 , n49665 , n49732 , n49733 );
and ( n49735 , n49660 , n49734 );
xor ( n49736 , n49590 , n49592 );
xor ( n49737 , n49736 , n49652 );
and ( n49738 , n49734 , n49737 );
and ( n49739 , n49660 , n49737 );
or ( n49740 , n49735 , n49738 , n49739 );
and ( n49741 , n49657 , n49740 );
and ( n49742 , n49655 , n49740 );
or ( n49743 , n49658 , n49741 , n49742 );
and ( n49744 , n49554 , n49743 );
and ( n49745 , n45112 , n40258 );
and ( n49746 , n45125 , n40256 );
nor ( n49747 , n49745 , n49746 );
xnor ( n49748 , n49747 , n40169 );
xor ( n49749 , n48514 , n48518 );
xor ( n49750 , n49749 , n48521 );
and ( n49751 , n49748 , n49750 );
and ( n49752 , n49743 , n49751 );
and ( n49753 , n49554 , n49751 );
or ( n49754 , n49744 , n49752 , n49753 );
and ( n49755 , n49551 , n49754 );
and ( n49756 , n49544 , n49754 );
or ( n49757 , n49552 , n49755 , n49756 );
xor ( n49758 , n48874 , n48876 );
xor ( n49759 , n49758 , n48879 );
and ( n49760 , n49757 , n49759 );
xor ( n49761 , n49524 , n49526 );
xor ( n49762 , n49655 , n49657 );
xor ( n49763 , n49762 , n49740 );
and ( n49764 , n45099 , n40258 );
and ( n49765 , n45112 , n40256 );
nor ( n49766 , n49764 , n49765 );
xnor ( n49767 , n49766 , n40169 );
xor ( n49768 , n48504 , n48508 );
xor ( n49769 , n49768 , n48511 );
and ( n49770 , n49767 , n49769 );
and ( n49771 , n49763 , n49770 );
xor ( n49772 , n49595 , n49638 );
xor ( n49773 , n49772 , n49649 );
xor ( n49774 , n49641 , n49643 );
xor ( n49775 , n49774 , n49646 );
xor ( n49776 , n49623 , n49627 );
xor ( n49777 , n49776 , n49632 );
and ( n49778 , n44520 , n42269 );
and ( n49779 , n44458 , n42266 );
nor ( n49780 , n49778 , n49779 );
xnor ( n49781 , n49780 , n41684 );
and ( n49782 , n44656 , n41984 );
and ( n49783 , n44565 , n41982 );
nor ( n49784 , n49782 , n49783 );
xnor ( n49785 , n49784 , n41687 );
and ( n49786 , n49781 , n49785 );
and ( n49787 , n45164 , n41622 );
and ( n49788 , n44665 , n41620 );
nor ( n49789 , n49787 , n49788 );
xnor ( n49790 , n49789 , n41194 );
and ( n49791 , n49785 , n49790 );
and ( n49792 , n49781 , n49790 );
or ( n49793 , n49786 , n49791 , n49792 );
and ( n49794 , n45138 , n41292 );
and ( n49795 , n45151 , n41290 );
nor ( n49796 , n49794 , n49795 );
xnor ( n49797 , n49796 , n41041 );
and ( n49798 , n45112 , n41055 );
and ( n49799 , n45125 , n41053 );
nor ( n49800 , n49798 , n49799 );
xnor ( n49801 , n49800 , n40728 );
and ( n49802 , n49797 , n49801 );
and ( n49803 , n45086 , n40746 );
and ( n49804 , n45099 , n40744 );
nor ( n49805 , n49803 , n49804 );
xnor ( n49806 , n49805 , n40501 );
and ( n49807 , n49801 , n49806 );
and ( n49808 , n49797 , n49806 );
or ( n49809 , n49802 , n49807 , n49808 );
and ( n49810 , n49793 , n49809 );
xor ( n49811 , n49675 , n49679 );
xor ( n49812 , n49811 , n49683 );
and ( n49813 , n49809 , n49812 );
and ( n49814 , n49793 , n49812 );
or ( n49815 , n49810 , n49813 , n49814 );
and ( n49816 , n49777 , n49815 );
xor ( n49817 , n49669 , n49670 );
xor ( n49818 , n49817 , n49686 );
and ( n49819 , n49815 , n49818 );
and ( n49820 , n49777 , n49818 );
or ( n49821 , n49816 , n49819 , n49820 );
and ( n49822 , n49775 , n49821 );
xor ( n49823 , n49689 , n49725 );
xor ( n49824 , n49823 , n49728 );
and ( n49825 , n49821 , n49824 );
and ( n49826 , n49775 , n49824 );
or ( n49827 , n49822 , n49825 , n49826 );
and ( n49828 , n49773 , n49827 );
xor ( n49829 , n49662 , n49664 );
xor ( n49830 , n49829 , n49731 );
and ( n49831 , n49827 , n49830 );
and ( n49832 , n49773 , n49830 );
or ( n49833 , n49828 , n49831 , n49832 );
xor ( n49834 , n49660 , n49734 );
xor ( n49835 , n49834 , n49737 );
and ( n49836 , n49833 , n49835 );
and ( n49837 , n45086 , n40258 );
and ( n49838 , n45099 , n40256 );
nor ( n49839 , n49837 , n49838 );
xnor ( n49840 , n49839 , n40169 );
xor ( n49841 , n48494 , n48498 );
xor ( n49842 , n49841 , n48501 );
and ( n49843 , n49840 , n49842 );
and ( n49844 , n49835 , n49843 );
and ( n49845 , n49833 , n49843 );
or ( n49846 , n49836 , n49844 , n49845 );
and ( n49847 , n49770 , n49846 );
and ( n49848 , n49763 , n49846 );
or ( n49849 , n49771 , n49847 , n49848 );
xor ( n49850 , n49548 , n49550 );
and ( n49851 , n49849 , n49850 );
xor ( n49852 , n49748 , n49750 );
xor ( n49853 , n49767 , n49769 );
xor ( n49854 , n49773 , n49827 );
xor ( n49855 , n49854 , n49830 );
xor ( n49856 , n49705 , n49719 );
xor ( n49857 , n49856 , n49722 );
xor ( n49858 , n49693 , n49697 );
xor ( n49859 , n49858 , n49702 );
xor ( n49860 , n49709 , n49713 );
xor ( n49861 , n49860 , n49716 );
and ( n49862 , n49859 , n49861 );
buf ( n49863 , n557813 );
not ( n49864 , n49863 );
and ( n49865 , n44565 , n42269 );
and ( n49866 , n44520 , n42266 );
nor ( n49867 , n49865 , n49866 );
xnor ( n49868 , n49867 , n41684 );
and ( n49869 , n44665 , n41984 );
and ( n49870 , n44656 , n41982 );
nor ( n49871 , n49869 , n49870 );
xnor ( n49872 , n49871 , n41687 );
and ( n49873 , n49868 , n49872 );
and ( n49874 , n49864 , n49873 );
and ( n49875 , n45151 , n41622 );
and ( n49876 , n45164 , n41620 );
nor ( n49877 , n49875 , n49876 );
xnor ( n49878 , n49877 , n41194 );
and ( n49879 , n45125 , n41292 );
and ( n49880 , n45138 , n41290 );
nor ( n49881 , n49879 , n49880 );
xnor ( n49882 , n49881 , n41041 );
and ( n49883 , n49878 , n49882 );
and ( n49884 , n45099 , n41055 );
and ( n49885 , n45112 , n41053 );
nor ( n49886 , n49884 , n49885 );
xnor ( n49887 , n49886 , n40728 );
and ( n49888 , n49882 , n49887 );
and ( n49889 , n49878 , n49887 );
or ( n49890 , n49883 , n49888 , n49889 );
and ( n49891 , n49873 , n49890 );
and ( n49892 , n49864 , n49890 );
or ( n49893 , n49874 , n49891 , n49892 );
and ( n49894 , n49861 , n49893 );
and ( n49895 , n49859 , n49893 );
or ( n49896 , n49862 , n49894 , n49895 );
and ( n49897 , n49857 , n49896 );
xor ( n49898 , n49777 , n49815 );
xor ( n49899 , n49898 , n49818 );
and ( n49900 , n49896 , n49899 );
and ( n49901 , n49857 , n49899 );
or ( n49902 , n49897 , n49900 , n49901 );
xor ( n49903 , n49775 , n49821 );
xor ( n49904 , n49903 , n49824 );
and ( n49905 , n49902 , n49904 );
xor ( n49906 , n48484 , n48488 );
xor ( n49907 , n49906 , n48491 );
and ( n49908 , n49904 , n49907 );
and ( n49909 , n49902 , n49907 );
or ( n49910 , n49905 , n49908 , n49909 );
and ( n49911 , n49855 , n49910 );
xor ( n49912 , n49840 , n49842 );
and ( n49913 , n49910 , n49912 );
and ( n49914 , n49855 , n49912 );
or ( n49915 , n49911 , n49913 , n49914 );
and ( n49916 , n49853 , n49915 );
xor ( n49917 , n49833 , n49835 );
xor ( n49918 , n49917 , n49843 );
and ( n49919 , n49915 , n49918 );
and ( n49920 , n49853 , n49918 );
or ( n49921 , n49916 , n49919 , n49920 );
and ( n49922 , n49852 , n49921 );
xor ( n49923 , n49763 , n49770 );
xor ( n49924 , n49923 , n49846 );
and ( n49925 , n49921 , n49924 );
and ( n49926 , n49852 , n49924 );
or ( n49927 , n49922 , n49925 , n49926 );
and ( n49928 , n49850 , n49927 );
and ( n49929 , n49849 , n49927 );
or ( n49930 , n49851 , n49928 , n49929 );
and ( n49931 , n49761 , n49930 );
xor ( n49932 , n49544 , n49551 );
xor ( n49933 , n49932 , n49754 );
and ( n49934 , n49930 , n49933 );
and ( n49935 , n49761 , n49933 );
or ( n49936 , n49931 , n49934 , n49935 );
and ( n49937 , n49759 , n49936 );
and ( n49938 , n49757 , n49936 );
or ( n49939 , n49760 , n49937 , n49938 );
xor ( n49940 , n49369 , n49371 );
xor ( n49941 , n49940 , n49530 );
and ( n49942 , n49939 , n49941 );
xor ( n49943 , n48882 , n48886 );
xor ( n49944 , n49943 , n48889 );
and ( n49945 , n49941 , n49944 );
and ( n49946 , n49939 , n49944 );
or ( n49947 , n49942 , n49945 , n49946 );
and ( n49948 , n49542 , n49947 );
xor ( n49949 , n49328 , n49533 );
xor ( n49950 , n49949 , n49536 );
and ( n49951 , n49947 , n49950 );
and ( n49952 , n49542 , n49950 );
or ( n49953 , n49948 , n49951 , n49952 );
and ( n49954 , n49539 , n49953 );
and ( n49955 , n49326 , n49953 );
or ( n49956 , n49540 , n49954 , n49955 );
and ( n49957 , n49324 , n49956 );
xor ( n49958 , n49031 , n49123 );
xor ( n49959 , n49958 , n49306 );
and ( n49960 , n49956 , n49959 );
and ( n49961 , n49324 , n49959 );
or ( n49962 , n49957 , n49960 , n49961 );
and ( n49963 , n49322 , n49962 );
xor ( n49964 , n49026 , n49028 );
xor ( n49965 , n49964 , n49309 );
and ( n49966 , n49962 , n49965 );
and ( n49967 , n49322 , n49965 );
or ( n49968 , n49963 , n49966 , n49967 );
and ( n49969 , n49320 , n49968 );
xor ( n49970 , n49021 , n49023 );
xor ( n49971 , n49970 , n49312 );
and ( n49972 , n49968 , n49971 );
and ( n49973 , n49320 , n49971 );
or ( n49974 , n49969 , n49972 , n49973 );
and ( n49975 , n49317 , n49974 );
and ( n49976 , n49315 , n49974 );
or ( n49977 , n49318 , n49975 , n49976 );
and ( n49978 , n48956 , n49977 );
and ( n49979 , n48954 , n49977 );
or ( n49980 , n48957 , n49978 , n49979 );
and ( n49981 , n48869 , n49980 );
and ( n49982 , n48789 , n49980 );
or ( n49983 , n48870 , n49981 , n49982 );
and ( n49984 , n48786 , n49983 );
and ( n49985 , n48746 , n49983 );
or ( n49986 , n48787 , n49984 , n49985 );
and ( n49987 , n48743 , n49986 );
and ( n49988 , n48432 , n49986 );
or ( n49989 , n48744 , n49987 , n49988 );
and ( n49990 , n48429 , n49989 );
and ( n49991 , n48337 , n49989 );
or ( n49992 , n48430 , n49990 , n49991 );
and ( n49993 , n48334 , n49992 );
and ( n49994 , n48332 , n49992 );
or ( n49995 , n48335 , n49993 , n49994 );
and ( n49996 , n48241 , n49995 );
and ( n49997 , n48018 , n49995 );
or ( n49998 , n48242 , n49996 , n49997 );
and ( n49999 , n48015 , n49998 );
and ( n50000 , n48013 , n49998 );
or ( n50001 , n48016 , n49999 , n50000 );
and ( n50002 , n47848 , n50001 );
and ( n50003 , n47605 , n50001 );
or ( n50004 , n47849 , n50002 , n50003 );
and ( n50005 , n47602 , n50004 );
and ( n50006 , n47493 , n50004 );
or ( n50007 , n47603 , n50005 , n50006 );
and ( n50008 , n47490 , n50007 );
and ( n50009 , n47400 , n50007 );
or ( n50010 , n47491 , n50008 , n50009 );
and ( n50011 , n47397 , n50010 );
and ( n50012 , n47112 , n50010 );
or ( n50013 , n47398 , n50011 , n50012 );
and ( n50014 , n47109 , n50013 );
and ( n50015 , n46947 , n50013 );
or ( n50016 , n47110 , n50014 , n50015 );
and ( n50017 , n46944 , n50016 );
and ( n50018 , n46942 , n50016 );
or ( n50019 , n46945 , n50017 , n50018 );
and ( n50020 , n46648 , n50019 );
and ( n50021 , n46548 , n50019 );
or ( n50022 , n46649 , n50020 , n50021 );
and ( n50023 , n46545 , n50022 );
and ( n50024 , n46434 , n50022 );
or ( n50025 , n46546 , n50023 , n50024 );
and ( n50026 , n46431 , n50025 );
and ( n50027 , n46311 , n50025 );
or ( n50028 , n46432 , n50026 , n50027 );
and ( n50029 , n46308 , n50028 );
and ( n50030 , n46306 , n50028 );
or ( n50031 , n46309 , n50029 , n50030 );
and ( n50032 , n45994 , n50031 );
xor ( n50033 , n45994 , n50031 );
xor ( n50034 , n46306 , n46308 );
xor ( n50035 , n50034 , n50028 );
xor ( n50036 , n46311 , n46431 );
xor ( n50037 , n50036 , n50025 );
xor ( n50038 , n46434 , n46545 );
xor ( n50039 , n50038 , n50022 );
xor ( n50040 , n46548 , n46648 );
xor ( n50041 , n50040 , n50019 );
xor ( n50042 , n46942 , n46944 );
xor ( n50043 , n50042 , n50016 );
xor ( n50044 , n46947 , n47109 );
xor ( n50045 , n50044 , n50013 );
xor ( n50046 , n47112 , n47397 );
xor ( n50047 , n50046 , n50010 );
xor ( n50048 , n47400 , n47490 );
xor ( n577358 , n50048 , n50007 );
xor ( n577359 , n47493 , n47602 );
xor ( n577360 , n577359 , n50004 );
xor ( n50049 , n47605 , n47848 );
xor ( n50050 , n50049 , n50001 );
xor ( n50051 , n48013 , n48015 );
xor ( n50052 , n50051 , n49998 );
xor ( n50053 , n48018 , n48241 );
xor ( n50054 , n50053 , n49995 );
xor ( n50055 , n48332 , n48334 );
xor ( n50056 , n50055 , n49992 );
xor ( n50057 , n48337 , n48429 );
xor ( n50058 , n50057 , n49989 );
xor ( n50059 , n48432 , n48743 );
xor ( n50060 , n50059 , n49986 );
xor ( n50061 , n48746 , n48786 );
xor ( n50062 , n50061 , n49983 );
xor ( n50063 , n48789 , n48869 );
xor ( n50064 , n50063 , n49980 );
xor ( n50065 , n48954 , n48956 );
xor ( n50066 , n50065 , n49977 );
xor ( n50067 , n49315 , n49317 );
xor ( n50068 , n50067 , n49974 );
xor ( n50069 , n49320 , n49968 );
xor ( n50070 , n50069 , n49971 );
xor ( n50071 , n49322 , n49962 );
xor ( n50072 , n50071 , n49965 );
xor ( n50073 , n49324 , n49956 );
xor ( n50074 , n50073 , n49959 );
xor ( n50075 , n49126 , n49300 );
xor ( n50076 , n50075 , n49303 );
xor ( n50077 , n49326 , n49539 );
xor ( n50078 , n50077 , n49953 );
and ( n50079 , n50076 , n50078 );
xor ( n50080 , n50076 , n50078 );
xor ( n50081 , n49542 , n49947 );
xor ( n50082 , n50081 , n49950 );
xor ( n50083 , n49939 , n49941 );
xor ( n50084 , n50083 , n49944 );
xor ( n50085 , n49374 , n49519 );
xor ( n50086 , n50085 , n49527 );
xor ( n50087 , n49757 , n49759 );
xor ( n50088 , n50087 , n49936 );
and ( n50089 , n50086 , n50088 );
xor ( n50090 , n50086 , n50088 );
xor ( n50091 , n49761 , n49930 );
xor ( n50092 , n50091 , n49933 );
xor ( n50093 , n49554 , n49743 );
xor ( n50094 , n50093 , n49751 );
xor ( n50095 , n49849 , n49850 );
xor ( n50096 , n50095 , n49927 );
and ( n50097 , n50094 , n50096 );
xor ( n50098 , n50094 , n50096 );
xor ( n50099 , n49852 , n49921 );
xor ( n50100 , n50099 , n49924 );
xor ( n50101 , n49853 , n49915 );
xor ( n50102 , n50101 , n49918 );
xor ( n50103 , n49793 , n49809 );
xor ( n50104 , n50103 , n49812 );
xor ( n50105 , n49781 , n49785 );
xor ( n50106 , n50105 , n49790 );
xor ( n50107 , n49797 , n49801 );
xor ( n50108 , n50107 , n49806 );
and ( n50109 , n50106 , n50108 );
and ( n50110 , n45073 , n40746 );
and ( n50111 , n45086 , n40744 );
nor ( n50112 , n50110 , n50111 );
xnor ( n50113 , n50112 , n40501 );
buf ( n50114 , n557814 );
not ( n50115 , n50114 );
and ( n50116 , n50113 , n50115 );
xor ( n50117 , n49868 , n49872 );
and ( n50118 , n50115 , n50117 );
and ( n50119 , n50113 , n50117 );
or ( n50120 , n50116 , n50118 , n50119 );
and ( n50121 , n50108 , n50120 );
and ( n50122 , n50106 , n50120 );
or ( n50123 , n50109 , n50121 , n50122 );
and ( n50124 , n50104 , n50123 );
xor ( n50125 , n49859 , n49861 );
xor ( n50126 , n50125 , n49893 );
and ( n50127 , n50123 , n50126 );
and ( n50128 , n50104 , n50126 );
or ( n50129 , n50124 , n50127 , n50128 );
xor ( n50130 , n49857 , n49896 );
xor ( n50131 , n50130 , n49899 );
and ( n50132 , n50129 , n50131 );
xor ( n50133 , n48474 , n48478 );
xor ( n50134 , n50133 , n48481 );
and ( n50135 , n50131 , n50134 );
and ( n50136 , n50129 , n50134 );
or ( n50137 , n50132 , n50135 , n50136 );
xor ( n50138 , n48464 , n48468 );
xor ( n50139 , n50138 , n48471 );
and ( n50140 , n44656 , n42269 );
and ( n50141 , n44565 , n42266 );
nor ( n50142 , n50140 , n50141 );
xnor ( n50143 , n50142 , n41684 );
and ( n50144 , n45164 , n41984 );
and ( n50145 , n44665 , n41982 );
nor ( n50146 , n50144 , n50145 );
xnor ( n50147 , n50146 , n41687 );
and ( n50148 , n50143 , n50147 );
and ( n50149 , n45138 , n41622 );
and ( n50150 , n45151 , n41620 );
nor ( n50151 , n50149 , n50150 );
xnor ( n50152 , n50151 , n41194 );
and ( n50153 , n50147 , n50152 );
and ( n50154 , n50143 , n50152 );
or ( n50155 , n50148 , n50153 , n50154 );
and ( n50156 , n45112 , n41292 );
and ( n50157 , n45125 , n41290 );
nor ( n50158 , n50156 , n50157 );
xnor ( n50159 , n50158 , n41041 );
and ( n50160 , n45086 , n41055 );
and ( n50161 , n45099 , n41053 );
nor ( n50162 , n50160 , n50161 );
xnor ( n50163 , n50162 , n40728 );
and ( n50164 , n50159 , n50163 );
and ( n50165 , n45060 , n40746 );
and ( n50166 , n45073 , n40744 );
nor ( n50167 , n50165 , n50166 );
xnor ( n50168 , n50167 , n40501 );
and ( n50169 , n50163 , n50168 );
and ( n50170 , n50159 , n50168 );
or ( n50171 , n50164 , n50169 , n50170 );
and ( n50172 , n50155 , n50171 );
xor ( n50173 , n49878 , n49882 );
xor ( n50174 , n50173 , n49887 );
and ( n50175 , n50171 , n50174 );
and ( n50176 , n50155 , n50174 );
or ( n50177 , n50172 , n50175 , n50176 );
xor ( n50178 , n49864 , n49873 );
xor ( n50179 , n50178 , n49890 );
and ( n50180 , n50177 , n50179 );
and ( n50181 , n45034 , n40527 );
and ( n50182 , n45047 , n40525 );
nor ( n50183 , n50181 , n50182 );
xnor ( n50184 , n50183 , n40382 );
buf ( n50185 , n557815 );
not ( n50186 , n50185 );
and ( n50187 , n50184 , n50186 );
and ( n50188 , n44665 , n42269 );
and ( n50189 , n44656 , n42266 );
nor ( n50190 , n50188 , n50189 );
xnor ( n50191 , n50190 , n41684 );
and ( n50192 , n45151 , n41984 );
and ( n50193 , n45164 , n41982 );
nor ( n50194 , n50192 , n50193 );
xnor ( n50195 , n50194 , n41687 );
and ( n50196 , n50191 , n50195 );
and ( n50197 , n45125 , n41622 );
and ( n50198 , n45138 , n41620 );
nor ( n50199 , n50197 , n50198 );
xnor ( n50200 , n50199 , n41194 );
and ( n50201 , n50195 , n50200 );
and ( n50202 , n50191 , n50200 );
or ( n50203 , n50196 , n50201 , n50202 );
and ( n50204 , n50186 , n50203 );
and ( n50205 , n50184 , n50203 );
or ( n50206 , n50187 , n50204 , n50205 );
and ( n50207 , n45099 , n41292 );
and ( n50208 , n45112 , n41290 );
nor ( n50209 , n50207 , n50208 );
xnor ( n50210 , n50209 , n41041 );
and ( n50211 , n45073 , n41055 );
and ( n50212 , n45086 , n41053 );
nor ( n50213 , n50211 , n50212 );
xnor ( n50214 , n50213 , n40728 );
and ( n50215 , n50210 , n50214 );
and ( n50216 , n45047 , n40746 );
and ( n50217 , n45060 , n40744 );
nor ( n50218 , n50216 , n50217 );
xnor ( n50219 , n50218 , n40501 );
and ( n50220 , n50214 , n50219 );
and ( n50221 , n50210 , n50219 );
or ( n50222 , n50215 , n50220 , n50221 );
xor ( n50223 , n50143 , n50147 );
xor ( n50224 , n50223 , n50152 );
and ( n50225 , n50222 , n50224 );
xor ( n50226 , n50159 , n50163 );
xor ( n50227 , n50226 , n50168 );
and ( n50228 , n50224 , n50227 );
and ( n50229 , n50222 , n50227 );
or ( n50230 , n50225 , n50228 , n50229 );
and ( n50231 , n50206 , n50230 );
xor ( n50232 , n50113 , n50115 );
xor ( n50233 , n50232 , n50117 );
and ( n50234 , n50230 , n50233 );
and ( n50235 , n50206 , n50233 );
or ( n50236 , n50231 , n50234 , n50235 );
and ( n50237 , n50179 , n50236 );
and ( n50238 , n50177 , n50236 );
or ( n50239 , n50180 , n50237 , n50238 );
and ( n50240 , n50139 , n50239 );
xor ( n50241 , n50104 , n50123 );
xor ( n50242 , n50241 , n50126 );
and ( n50243 , n50239 , n50242 );
and ( n50244 , n50139 , n50242 );
or ( n50245 , n50240 , n50243 , n50244 );
xor ( n50246 , n48443 , n48447 );
and ( n50247 , n44991 , n40256 );
not ( n50248 , n50247 );
and ( n50249 , n50248 , n40169 );
and ( n50250 , n44991 , n40258 );
and ( n50251 , n44999 , n40256 );
nor ( n50252 , n50250 , n50251 );
xnor ( n50253 , n50252 , n40169 );
and ( n50254 , n50249 , n50253 );
and ( n50255 , n44999 , n40258 );
and ( n50256 , n45008 , n40256 );
nor ( n50257 , n50255 , n50256 );
xnor ( n50258 , n50257 , n40169 );
and ( n50259 , n50254 , n50258 );
and ( n50260 , n50258 , n48441 );
and ( n50261 , n50254 , n48441 );
or ( n50262 , n50259 , n50260 , n50261 );
and ( n50263 , n50246 , n50262 );
and ( n50264 , n45008 , n40258 );
and ( n50265 , n45021 , n40256 );
nor ( n50266 , n50264 , n50265 );
xnor ( n50267 , n50266 , n40169 );
and ( n50268 , n50262 , n50267 );
and ( n50269 , n50246 , n50267 );
or ( n50270 , n50263 , n50268 , n50269 );
and ( n50271 , n45021 , n40258 );
and ( n50272 , n45034 , n40256 );
nor ( n50273 , n50271 , n50272 );
xnor ( n50274 , n50273 , n40169 );
and ( n50275 , n50270 , n50274 );
xor ( n50276 , n48448 , n48452 );
xor ( n50277 , n50276 , n48020 );
and ( n50278 , n50274 , n50277 );
and ( n50279 , n50270 , n50277 );
or ( n50280 , n50275 , n50278 , n50279 );
and ( n50281 , n45034 , n40258 );
and ( n50282 , n45047 , n40256 );
nor ( n50283 , n50281 , n50282 );
xnor ( n50284 , n50283 , n40169 );
and ( n50285 , n50280 , n50284 );
xor ( n50286 , n48440 , n48456 );
xor ( n50287 , n50286 , n48461 );
and ( n50288 , n50284 , n50287 );
and ( n50289 , n50280 , n50287 );
or ( n50290 , n50285 , n50288 , n50289 );
xor ( n50291 , n50106 , n50108 );
xor ( n50292 , n50291 , n50120 );
xor ( n50293 , n50155 , n50171 );
xor ( n50294 , n50293 , n50174 );
and ( n50295 , n45021 , n40527 );
and ( n50296 , n45034 , n40525 );
nor ( n50297 , n50295 , n50296 );
xnor ( n50298 , n50297 , n40382 );
buf ( n50299 , n557816 );
not ( n50300 , n50299 );
and ( n50301 , n50298 , n50300 );
xor ( n50302 , n50191 , n50195 );
xor ( n50303 , n50302 , n50200 );
and ( n50304 , n50300 , n50303 );
and ( n50305 , n50298 , n50303 );
or ( n50306 , n50301 , n50304 , n50305 );
xor ( n50307 , n50184 , n50186 );
xor ( n50308 , n50307 , n50203 );
and ( n50309 , n50306 , n50308 );
xor ( n50310 , n50222 , n50224 );
xor ( n50311 , n50310 , n50227 );
and ( n50312 , n50308 , n50311 );
and ( n50313 , n50306 , n50311 );
or ( n50314 , n50309 , n50312 , n50313 );
and ( n50315 , n50294 , n50314 );
xor ( n50316 , n50206 , n50230 );
xor ( n50317 , n50316 , n50233 );
and ( n50318 , n50314 , n50317 );
and ( n50319 , n50294 , n50317 );
or ( n50320 , n50315 , n50318 , n50319 );
and ( n50321 , n50292 , n50320 );
xor ( n50322 , n50177 , n50179 );
xor ( n50323 , n50322 , n50236 );
and ( n50324 , n50320 , n50323 );
and ( n50325 , n50292 , n50323 );
or ( n50326 , n50321 , n50324 , n50325 );
and ( n50327 , n50290 , n50326 );
xor ( n50328 , n50139 , n50239 );
xor ( n50329 , n50328 , n50242 );
and ( n50330 , n50326 , n50329 );
and ( n50331 , n50290 , n50329 );
or ( n50332 , n50327 , n50330 , n50331 );
and ( n50333 , n50245 , n50332 );
xor ( n50334 , n50129 , n50131 );
xor ( n50335 , n50334 , n50134 );
and ( n50336 , n50332 , n50335 );
and ( n50337 , n50245 , n50335 );
or ( n50338 , n50333 , n50336 , n50337 );
and ( n50339 , n50137 , n50338 );
xor ( n50340 , n49902 , n49904 );
xor ( n50341 , n50340 , n49907 );
and ( n50342 , n50338 , n50341 );
and ( n50343 , n50137 , n50341 );
or ( n50344 , n50339 , n50342 , n50343 );
xor ( n50345 , n49855 , n49910 );
xor ( n50346 , n50345 , n49912 );
and ( n50347 , n50344 , n50346 );
xor ( n50348 , n50344 , n50346 );
xor ( n50349 , n50137 , n50338 );
xor ( n50350 , n50349 , n50341 );
xor ( n50351 , n50245 , n50332 );
xor ( n50352 , n50351 , n50335 );
and ( n50353 , n45060 , n40527 );
and ( n50354 , n45073 , n40525 );
nor ( n50355 , n50353 , n50354 );
xnor ( n50356 , n50355 , n40382 );
xor ( n50357 , n50280 , n50284 );
xor ( n50358 , n50357 , n50287 );
and ( n50359 , n50356 , n50358 );
xor ( n50360 , n50290 , n50326 );
xor ( n50361 , n50360 , n50329 );
and ( n50362 , n50359 , n50361 );
and ( n50363 , n45047 , n40527 );
and ( n50364 , n45060 , n40525 );
nor ( n50365 , n50363 , n50364 );
xnor ( n50366 , n50365 , n40382 );
xor ( n50367 , n50270 , n50274 );
xor ( n50368 , n50367 , n50277 );
and ( n50369 , n50366 , n50368 );
xor ( n50370 , n50292 , n50320 );
xor ( n50371 , n50370 , n50323 );
and ( n50372 , n50369 , n50371 );
xor ( n50373 , n50356 , n50358 );
and ( n50374 , n50371 , n50373 );
and ( n50375 , n50369 , n50373 );
or ( n50376 , n50372 , n50374 , n50375 );
and ( n50377 , n50361 , n50376 );
and ( n50378 , n50359 , n50376 );
or ( n50379 , n50362 , n50377 , n50378 );
and ( n50380 , n50352 , n50379 );
xor ( n50381 , n50352 , n50379 );
xor ( n50382 , n50359 , n50361 );
xor ( n50383 , n50382 , n50376 );
xor ( n50384 , n50246 , n50262 );
xor ( n50385 , n50384 , n50267 );
xor ( n50386 , n50210 , n50214 );
xor ( n50387 , n50386 , n50219 );
xor ( n50388 , n50254 , n50258 );
xor ( n50389 , n50388 , n48441 );
and ( n50390 , n50387 , n50389 );
xor ( n50391 , n50298 , n50300 );
xor ( n50392 , n50391 , n50303 );
and ( n50393 , n50389 , n50392 );
and ( n50394 , n50387 , n50392 );
or ( n50395 , n50390 , n50393 , n50394 );
and ( n50396 , n50385 , n50395 );
xor ( n50397 , n50306 , n50308 );
xor ( n50398 , n50397 , n50311 );
and ( n50399 , n50395 , n50398 );
and ( n50400 , n50385 , n50398 );
or ( n50401 , n50396 , n50399 , n50400 );
xor ( n50402 , n50294 , n50314 );
xor ( n50403 , n50402 , n50317 );
and ( n50404 , n50401 , n50403 );
xor ( n50405 , n50366 , n50368 );
and ( n50406 , n50403 , n50405 );
and ( n50407 , n50401 , n50405 );
or ( n50408 , n50404 , n50406 , n50407 );
xor ( n50409 , n50369 , n50371 );
xor ( n50410 , n50409 , n50373 );
and ( n50411 , n50408 , n50410 );
xor ( n50412 , n50401 , n50403 );
xor ( n50413 , n50412 , n50405 );
xor ( n50414 , n50385 , n50395 );
xor ( n50415 , n50414 , n50398 );
xor ( n50416 , n50249 , n50253 );
and ( n50417 , n44991 , n40525 );
not ( n50418 , n50417 );
and ( n50419 , n50418 , n40382 );
and ( n50420 , n44991 , n40527 );
and ( n50421 , n44999 , n40525 );
nor ( n50422 , n50420 , n50421 );
xnor ( n50423 , n50422 , n40382 );
and ( n50424 , n50419 , n50423 );
and ( n50425 , n44999 , n40527 );
and ( n50426 , n45008 , n40525 );
nor ( n50427 , n50425 , n50426 );
xnor ( n50428 , n50427 , n40382 );
and ( n50429 , n50424 , n50428 );
and ( n50430 , n50428 , n50247 );
and ( n50431 , n50424 , n50247 );
or ( n50432 , n50429 , n50430 , n50431 );
and ( n50433 , n50416 , n50432 );
and ( n50434 , n45008 , n40527 );
and ( n50435 , n45021 , n40525 );
nor ( n50436 , n50434 , n50435 );
xnor ( n50437 , n50436 , n40382 );
and ( n50438 , n50432 , n50437 );
and ( n50439 , n50416 , n50437 );
or ( n50440 , n50433 , n50438 , n50439 );
xor ( n50441 , n50387 , n50389 );
xor ( n50442 , n50441 , n50392 );
and ( n50443 , n50440 , n50442 );
xor ( n50444 , n50419 , n50423 );
and ( n50445 , n44991 , n40744 );
not ( n50446 , n50445 );
and ( n50447 , n50446 , n40501 );
and ( n50448 , n44991 , n40746 );
and ( n50449 , n44999 , n40744 );
nor ( n50450 , n50448 , n50449 );
xnor ( n50451 , n50450 , n40501 );
and ( n50452 , n50447 , n50451 );
and ( n50453 , n44999 , n40746 );
and ( n50454 , n45008 , n40744 );
nor ( n50455 , n50453 , n50454 );
xnor ( n50456 , n50455 , n40501 );
and ( n50457 , n50452 , n50456 );
and ( n50458 , n50456 , n50417 );
and ( n50459 , n50452 , n50417 );
or ( n50460 , n50457 , n50458 , n50459 );
and ( n50461 , n50444 , n50460 );
and ( n50462 , n45008 , n40746 );
and ( n50463 , n45021 , n40744 );
nor ( n50464 , n50462 , n50463 );
xnor ( n50465 , n50464 , n40501 );
and ( n50466 , n50460 , n50465 );
and ( n50467 , n50444 , n50465 );
or ( n50468 , n50461 , n50466 , n50467 );
and ( n50469 , n45021 , n40746 );
and ( n50470 , n45034 , n40744 );
nor ( n50471 , n50469 , n50470 );
xnor ( n50472 , n50471 , n40501 );
and ( n50473 , n50468 , n50472 );
xor ( n50474 , n50424 , n50428 );
xor ( n50475 , n50474 , n50247 );
and ( n50476 , n50472 , n50475 );
and ( n50477 , n50468 , n50475 );
or ( n50478 , n50473 , n50476 , n50477 );
and ( n50479 , n45034 , n40746 );
and ( n50480 , n45047 , n40744 );
nor ( n50481 , n50479 , n50480 );
xnor ( n50482 , n50481 , n40501 );
and ( n50483 , n50478 , n50482 );
xor ( n50484 , n50416 , n50432 );
xor ( n50485 , n50484 , n50437 );
and ( n50486 , n50482 , n50485 );
and ( n50487 , n50478 , n50485 );
or ( n50488 , n50483 , n50486 , n50487 );
and ( n50489 , n50442 , n50488 );
and ( n50490 , n50440 , n50488 );
or ( n50491 , n50443 , n50489 , n50490 );
and ( n50492 , n50415 , n50491 );
xor ( n50493 , n50440 , n50442 );
xor ( n50494 , n50493 , n50488 );
xor ( n50495 , n50447 , n50451 );
and ( n50496 , n44991 , n41053 );
not ( n50497 , n50496 );
and ( n50498 , n50497 , n40728 );
and ( n50499 , n44991 , n41055 );
and ( n50500 , n44999 , n41053 );
nor ( n50501 , n50499 , n50500 );
xnor ( n50502 , n50501 , n40728 );
and ( n50503 , n50498 , n50502 );
and ( n50504 , n44999 , n41055 );
and ( n50505 , n45008 , n41053 );
nor ( n50506 , n50504 , n50505 );
xnor ( n50507 , n50506 , n40728 );
and ( n50508 , n50503 , n50507 );
and ( n50509 , n50507 , n50445 );
and ( n50510 , n50503 , n50445 );
or ( n50511 , n50508 , n50509 , n50510 );
and ( n50512 , n50495 , n50511 );
and ( n50513 , n45008 , n41055 );
and ( n50514 , n45021 , n41053 );
nor ( n50515 , n50513 , n50514 );
xnor ( n50516 , n50515 , n40728 );
and ( n50517 , n50511 , n50516 );
and ( n50518 , n50495 , n50516 );
or ( n50519 , n50512 , n50517 , n50518 );
and ( n50520 , n45021 , n41055 );
and ( n50521 , n45034 , n41053 );
nor ( n50522 , n50520 , n50521 );
xnor ( n50523 , n50522 , n40728 );
and ( n50524 , n50519 , n50523 );
xor ( n50525 , n50452 , n50456 );
xor ( n50526 , n50525 , n50417 );
and ( n50527 , n50523 , n50526 );
and ( n577840 , n50519 , n50526 );
or ( n50528 , n50524 , n50527 , n577840 );
and ( n50529 , n45034 , n41055 );
and ( n50530 , n45047 , n41053 );
nor ( n50531 , n50529 , n50530 );
xnor ( n50532 , n50531 , n40728 );
and ( n50533 , n50528 , n50532 );
xor ( n50534 , n50444 , n50460 );
xor ( n50535 , n50534 , n50465 );
and ( n50536 , n50532 , n50535 );
and ( n50537 , n50528 , n50535 );
or ( n50538 , n50533 , n50536 , n50537 );
and ( n50539 , n45047 , n41055 );
and ( n50540 , n45060 , n41053 );
nor ( n50541 , n50539 , n50540 );
xnor ( n50542 , n50541 , n40728 );
and ( n50543 , n50538 , n50542 );
xor ( n50544 , n50468 , n50472 );
xor ( n50545 , n50544 , n50475 );
and ( n50546 , n50542 , n50545 );
and ( n50547 , n50538 , n50545 );
or ( n50548 , n50543 , n50546 , n50547 );
and ( n50549 , n45060 , n41055 );
and ( n50550 , n45073 , n41053 );
nor ( n50551 , n50549 , n50550 );
xnor ( n50552 , n50551 , n40728 );
and ( n50553 , n50548 , n50552 );
xor ( n50554 , n50478 , n50482 );
xor ( n50555 , n50554 , n50485 );
and ( n50556 , n50552 , n50555 );
and ( n50557 , n50548 , n50555 );
or ( n50558 , n50553 , n50556 , n50557 );
and ( n50559 , n50494 , n50558 );
and ( n50560 , n45086 , n41292 );
and ( n50561 , n45099 , n41290 );
nor ( n50562 , n50560 , n50561 );
xnor ( n50563 , n50562 , n41041 );
buf ( n50564 , n557817 );
not ( n50565 , n50564 );
and ( n50566 , n50563 , n50565 );
xor ( n50567 , n50548 , n50552 );
xor ( n50568 , n50567 , n50555 );
and ( n50569 , n50565 , n50568 );
and ( n50570 , n50563 , n50568 );
or ( n50571 , n50566 , n50569 , n50570 );
and ( n50572 , n50558 , n50571 );
and ( n50573 , n50494 , n50571 );
or ( n50574 , n50559 , n50572 , n50573 );
and ( n50575 , n50491 , n50574 );
and ( n50576 , n50415 , n50574 );
or ( n50577 , n50492 , n50575 , n50576 );
and ( n50578 , n50413 , n50577 );
xor ( n50579 , n50415 , n50491 );
xor ( n50580 , n50579 , n50574 );
xor ( n50581 , n50498 , n50502 );
and ( n50582 , n44991 , n41290 );
not ( n50583 , n50582 );
and ( n50584 , n50583 , n41041 );
and ( n50585 , n44991 , n41292 );
and ( n50586 , n44999 , n41290 );
nor ( n50587 , n50585 , n50586 );
xnor ( n50588 , n50587 , n41041 );
and ( n50589 , n50584 , n50588 );
and ( n50590 , n44999 , n41292 );
and ( n50591 , n45008 , n41290 );
nor ( n50592 , n50590 , n50591 );
xnor ( n50593 , n50592 , n41041 );
and ( n50594 , n50589 , n50593 );
and ( n50595 , n50593 , n50496 );
and ( n50596 , n50589 , n50496 );
or ( n50597 , n50594 , n50595 , n50596 );
and ( n50598 , n50581 , n50597 );
and ( n50599 , n45008 , n41292 );
and ( n50600 , n45021 , n41290 );
nor ( n50601 , n50599 , n50600 );
xnor ( n50602 , n50601 , n41041 );
and ( n50603 , n50597 , n50602 );
and ( n50604 , n50581 , n50602 );
or ( n50605 , n50598 , n50603 , n50604 );
and ( n50606 , n45021 , n41292 );
and ( n50607 , n45034 , n41290 );
nor ( n50608 , n50606 , n50607 );
xnor ( n50609 , n50608 , n41041 );
and ( n50610 , n50605 , n50609 );
xor ( n50611 , n50503 , n50507 );
xor ( n50612 , n50611 , n50445 );
and ( n50613 , n50609 , n50612 );
and ( n50614 , n50605 , n50612 );
or ( n50615 , n50610 , n50613 , n50614 );
and ( n50616 , n45034 , n41292 );
and ( n50617 , n45047 , n41290 );
nor ( n50618 , n50616 , n50617 );
xnor ( n50619 , n50618 , n41041 );
and ( n50620 , n50615 , n50619 );
xor ( n50621 , n50495 , n50511 );
xor ( n50622 , n50621 , n50516 );
and ( n50623 , n50619 , n50622 );
and ( n50624 , n50615 , n50622 );
or ( n50625 , n50620 , n50623 , n50624 );
and ( n50626 , n45047 , n41292 );
and ( n50627 , n45060 , n41290 );
nor ( n50628 , n50626 , n50627 );
xnor ( n50629 , n50628 , n41041 );
and ( n50630 , n50625 , n50629 );
xor ( n50631 , n50519 , n50523 );
xor ( n50632 , n50631 , n50526 );
and ( n50633 , n50629 , n50632 );
and ( n50634 , n50625 , n50632 );
or ( n50635 , n50630 , n50633 , n50634 );
and ( n50636 , n45060 , n41292 );
and ( n50637 , n45073 , n41290 );
nor ( n50638 , n50636 , n50637 );
xnor ( n50639 , n50638 , n41041 );
and ( n50640 , n50635 , n50639 );
xor ( n50641 , n50528 , n50532 );
xor ( n50642 , n50641 , n50535 );
and ( n50643 , n50639 , n50642 );
and ( n50644 , n50635 , n50642 );
or ( n50645 , n50640 , n50643 , n50644 );
and ( n50646 , n45073 , n41292 );
and ( n50647 , n45086 , n41290 );
nor ( n50648 , n50646 , n50647 );
xnor ( n50649 , n50648 , n41041 );
and ( n50650 , n50645 , n50649 );
xor ( n50651 , n50538 , n50542 );
xor ( n50652 , n50651 , n50545 );
and ( n50653 , n50649 , n50652 );
and ( n50654 , n50645 , n50652 );
or ( n50655 , n50650 , n50653 , n50654 );
and ( n50656 , n45112 , n41622 );
and ( n50657 , n45125 , n41620 );
nor ( n50658 , n50656 , n50657 );
xnor ( n50659 , n50658 , n41194 );
and ( n50660 , n50655 , n50659 );
xor ( n50661 , n50563 , n50565 );
xor ( n50662 , n50661 , n50568 );
and ( n50663 , n50659 , n50662 );
and ( n50664 , n50655 , n50662 );
or ( n50665 , n50660 , n50663 , n50664 );
xor ( n50666 , n50494 , n50558 );
xor ( n50667 , n50666 , n50571 );
and ( n50668 , n50665 , n50667 );
and ( n50669 , n45099 , n41622 );
and ( n50670 , n45112 , n41620 );
nor ( n50671 , n50669 , n50670 );
xnor ( n50672 , n50671 , n41194 );
buf ( n50673 , n557818 );
not ( n50674 , n50673 );
and ( n50675 , n50672 , n50674 );
xor ( n50676 , n50645 , n50649 );
xor ( n50677 , n50676 , n50652 );
and ( n50678 , n50674 , n50677 );
and ( n50679 , n50672 , n50677 );
or ( n50680 , n50675 , n50678 , n50679 );
and ( n50681 , n45138 , n41984 );
and ( n50682 , n45151 , n41982 );
nor ( n50683 , n50681 , n50682 );
xnor ( n50684 , n50683 , n41687 );
and ( n50685 , n50680 , n50684 );
xor ( n50686 , n50655 , n50659 );
xor ( n50687 , n50686 , n50662 );
and ( n50688 , n50684 , n50687 );
and ( n50689 , n50680 , n50687 );
or ( n50690 , n50685 , n50688 , n50689 );
and ( n50691 , n50667 , n50690 );
and ( n50692 , n50665 , n50690 );
or ( n50693 , n50668 , n50691 , n50692 );
and ( n50694 , n50580 , n50693 );
xor ( n50695 , n50665 , n50667 );
xor ( n50696 , n50695 , n50690 );
and ( n50697 , n45086 , n41622 );
and ( n50698 , n45099 , n41620 );
nor ( n50699 , n50697 , n50698 );
xnor ( n50700 , n50699 , n41194 );
buf ( n50701 , n557819 );
not ( n50702 , n50701 );
and ( n50703 , n50700 , n50702 );
xor ( n50704 , n50635 , n50639 );
xor ( n50705 , n50704 , n50642 );
and ( n50706 , n50702 , n50705 );
and ( n50707 , n50700 , n50705 );
or ( n50708 , n50703 , n50706 , n50707 );
and ( n50709 , n45060 , n41622 );
and ( n50710 , n45073 , n41620 );
nor ( n50711 , n50709 , n50710 );
xnor ( n50712 , n50711 , n41194 );
buf ( n50713 , n557821 );
not ( n50714 , n50713 );
and ( n50715 , n50712 , n50714 );
xor ( n50716 , n50615 , n50619 );
xor ( n50717 , n50716 , n50622 );
and ( n50718 , n50714 , n50717 );
and ( n50719 , n50712 , n50717 );
or ( n50720 , n50715 , n50718 , n50719 );
buf ( n50721 , n557820 );
not ( n50722 , n50721 );
and ( n50723 , n50720 , n50722 );
xor ( n50724 , n50625 , n50629 );
xor ( n50725 , n50724 , n50632 );
and ( n50726 , n50722 , n50725 );
and ( n50727 , n50720 , n50725 );
or ( n50728 , n50723 , n50726 , n50727 );
and ( n50729 , n45112 , n41984 );
and ( n50730 , n45125 , n41982 );
nor ( n50731 , n50729 , n50730 );
xnor ( n50732 , n50731 , n41687 );
and ( n50733 , n50728 , n50732 );
xor ( n50734 , n50700 , n50702 );
xor ( n50735 , n50734 , n50705 );
and ( n50736 , n50732 , n50735 );
and ( n50737 , n50728 , n50735 );
or ( n50738 , n50733 , n50736 , n50737 );
and ( n50739 , n50708 , n50738 );
xor ( n50740 , n50672 , n50674 );
xor ( n50741 , n50740 , n50677 );
and ( n50742 , n50738 , n50741 );
and ( n50743 , n50708 , n50741 );
or ( n50744 , n50739 , n50742 , n50743 );
and ( n50745 , n45047 , n41622 );
and ( n50746 , n45060 , n41620 );
nor ( n50747 , n50745 , n50746 );
xnor ( n50748 , n50747 , n41194 );
buf ( n50749 , n557822 );
not ( n50750 , n50749 );
and ( n50751 , n50748 , n50750 );
xor ( n50752 , n50605 , n50609 );
xor ( n50753 , n50752 , n50612 );
and ( n50754 , n50750 , n50753 );
and ( n50755 , n50748 , n50753 );
or ( n50756 , n50751 , n50754 , n50755 );
xor ( n50757 , n50584 , n50588 );
and ( n50758 , n44991 , n41620 );
not ( n50759 , n50758 );
and ( n50760 , n50759 , n41194 );
and ( n50761 , n44991 , n41622 );
and ( n50762 , n44999 , n41620 );
nor ( n50763 , n50761 , n50762 );
xnor ( n50764 , n50763 , n41194 );
and ( n50765 , n50760 , n50764 );
and ( n50766 , n44999 , n41622 );
and ( n50767 , n45008 , n41620 );
nor ( n50768 , n50766 , n50767 );
xnor ( n50769 , n50768 , n41194 );
and ( n50770 , n50765 , n50769 );
and ( n50771 , n50769 , n50582 );
and ( n50772 , n50765 , n50582 );
or ( n50773 , n50770 , n50771 , n50772 );
and ( n50774 , n50757 , n50773 );
and ( n50775 , n45008 , n41622 );
and ( n50776 , n45021 , n41620 );
nor ( n50777 , n50775 , n50776 );
xnor ( n50778 , n50777 , n41194 );
and ( n50779 , n50773 , n50778 );
and ( n50780 , n50757 , n50778 );
or ( n50781 , n50774 , n50779 , n50780 );
and ( n50782 , n45021 , n41622 );
and ( n50783 , n45034 , n41620 );
nor ( n50784 , n50782 , n50783 );
xnor ( n50785 , n50784 , n41194 );
and ( n50786 , n50781 , n50785 );
xor ( n50787 , n50589 , n50593 );
xor ( n50788 , n50787 , n50496 );
and ( n50789 , n50785 , n50788 );
and ( n50790 , n50781 , n50788 );
or ( n50791 , n50786 , n50789 , n50790 );
and ( n50792 , n45034 , n41622 );
and ( n50793 , n45047 , n41620 );
nor ( n50794 , n50792 , n50793 );
xnor ( n50795 , n50794 , n41194 );
and ( n50796 , n50791 , n50795 );
xor ( n50797 , n50581 , n50597 );
xor ( n50798 , n50797 , n50602 );
and ( n50799 , n50795 , n50798 );
and ( n50800 , n50791 , n50798 );
or ( n50801 , n50796 , n50799 , n50800 );
xor ( n50802 , n50760 , n50764 );
and ( n50803 , n44991 , n41982 );
not ( n50804 , n50803 );
and ( n50805 , n50804 , n41687 );
and ( n50806 , n44991 , n41984 );
and ( n50807 , n44999 , n41982 );
nor ( n50808 , n50806 , n50807 );
xnor ( n50809 , n50808 , n41687 );
and ( n50810 , n50805 , n50809 );
and ( n50811 , n50810 , n50758 );
buf ( n50812 , n557828 );
not ( n50813 , n50812 );
and ( n50814 , n50758 , n50813 );
and ( n50815 , n50810 , n50813 );
or ( n50816 , n50811 , n50814 , n50815 );
and ( n50817 , n50802 , n50816 );
buf ( n50818 , n557827 );
not ( n50819 , n50818 );
and ( n50820 , n50816 , n50819 );
and ( n50821 , n50802 , n50819 );
or ( n50822 , n50817 , n50820 , n50821 );
buf ( n50823 , n557826 );
not ( n50824 , n50823 );
and ( n50825 , n50822 , n50824 );
xor ( n50826 , n50765 , n50769 );
xor ( n50827 , n50826 , n50582 );
and ( n50828 , n50824 , n50827 );
and ( n50829 , n50822 , n50827 );
or ( n50830 , n50825 , n50828 , n50829 );
buf ( n50831 , n557825 );
not ( n50832 , n50831 );
and ( n50833 , n50830 , n50832 );
xor ( n50834 , n50757 , n50773 );
xor ( n50835 , n50834 , n50778 );
and ( n50836 , n50832 , n50835 );
and ( n50837 , n50830 , n50835 );
or ( n50838 , n50833 , n50836 , n50837 );
buf ( n50839 , n557824 );
not ( n50840 , n50839 );
and ( n50841 , n50838 , n50840 );
xor ( n50842 , n50781 , n50785 );
xor ( n50843 , n50842 , n50788 );
and ( n50844 , n50840 , n50843 );
and ( n50845 , n50838 , n50843 );
or ( n50846 , n50841 , n50844 , n50845 );
buf ( n50847 , n557823 );
not ( n50848 , n50847 );
and ( n50849 , n50846 , n50848 );
xor ( n50850 , n50791 , n50795 );
xor ( n50851 , n50850 , n50798 );
and ( n50852 , n50848 , n50851 );
and ( n50853 , n50846 , n50851 );
or ( n50854 , n50849 , n50852 , n50853 );
and ( n50855 , n50801 , n50854 );
xor ( n50856 , n50748 , n50750 );
xor ( n50857 , n50856 , n50753 );
and ( n50858 , n50854 , n50857 );
and ( n50859 , n50801 , n50857 );
or ( n50860 , n50855 , n50858 , n50859 );
and ( n50861 , n50756 , n50860 );
xor ( n50862 , n50712 , n50714 );
xor ( n50863 , n50862 , n50717 );
and ( n50864 , n50860 , n50863 );
and ( n50865 , n50756 , n50863 );
or ( n50866 , n50861 , n50864 , n50865 );
and ( n50867 , n45073 , n41622 );
and ( n50868 , n45086 , n41620 );
nor ( n50869 , n50867 , n50868 );
xnor ( n50870 , n50869 , n41194 );
and ( n50871 , n50866 , n50870 );
xor ( n50872 , n50720 , n50722 );
xor ( n50873 , n50872 , n50725 );
and ( n50874 , n50870 , n50873 );
and ( n50875 , n50866 , n50873 );
or ( n50876 , n50871 , n50874 , n50875 );
xor ( n50877 , n50805 , n50809 );
and ( n50878 , n44991 , n42266 );
not ( n50879 , n50878 );
and ( n50880 , n50879 , n41684 );
buf ( n50881 , n557831 );
not ( n50882 , n50881 );
and ( n50883 , n50880 , n50882 );
and ( n50884 , n50883 , n50803 );
buf ( n50885 , n557830 );
not ( n50886 , n50885 );
and ( n50887 , n50803 , n50886 );
and ( n50888 , n50883 , n50886 );
or ( n50889 , n50884 , n50887 , n50888 );
and ( n50890 , n50877 , n50889 );
buf ( n50891 , n557829 );
not ( n50892 , n50891 );
and ( n50893 , n50889 , n50892 );
and ( n50894 , n50877 , n50892 );
or ( n50895 , n50890 , n50893 , n50894 );
and ( n50896 , n44999 , n41984 );
and ( n50897 , n45008 , n41982 );
nor ( n50898 , n50896 , n50897 );
xnor ( n50899 , n50898 , n41687 );
and ( n50900 , n50895 , n50899 );
xor ( n50901 , n50810 , n50758 );
xor ( n50902 , n50901 , n50813 );
and ( n50903 , n50899 , n50902 );
and ( n50904 , n50895 , n50902 );
or ( n50905 , n50900 , n50903 , n50904 );
and ( n50906 , n45008 , n41984 );
and ( n50907 , n45021 , n41982 );
nor ( n50908 , n50906 , n50907 );
xnor ( n50909 , n50908 , n41687 );
and ( n50910 , n50905 , n50909 );
xor ( n50911 , n50802 , n50816 );
xor ( n50912 , n50911 , n50819 );
and ( n50913 , n50909 , n50912 );
and ( n50914 , n50905 , n50912 );
or ( n50915 , n50910 , n50913 , n50914 );
and ( n50916 , n45021 , n41984 );
and ( n50917 , n45034 , n41982 );
nor ( n50918 , n50916 , n50917 );
xnor ( n50919 , n50918 , n41687 );
and ( n50920 , n50915 , n50919 );
xor ( n50921 , n50822 , n50824 );
xor ( n50922 , n50921 , n50827 );
and ( n50923 , n50919 , n50922 );
and ( n50924 , n50915 , n50922 );
or ( n50925 , n50920 , n50923 , n50924 );
and ( n50926 , n45034 , n41984 );
and ( n50927 , n45047 , n41982 );
nor ( n50928 , n50926 , n50927 );
xnor ( n50929 , n50928 , n41687 );
and ( n50930 , n50925 , n50929 );
xor ( n50931 , n50830 , n50832 );
xor ( n50932 , n50931 , n50835 );
and ( n50933 , n50929 , n50932 );
and ( n50934 , n50925 , n50932 );
or ( n50935 , n50930 , n50933 , n50934 );
and ( n50936 , n45047 , n41984 );
and ( n50937 , n45060 , n41982 );
nor ( n50938 , n50936 , n50937 );
xnor ( n50939 , n50938 , n41687 );
and ( n50940 , n50935 , n50939 );
xor ( n50941 , n50838 , n50840 );
xor ( n50942 , n50941 , n50843 );
and ( n50943 , n50939 , n50942 );
and ( n50944 , n50935 , n50942 );
or ( n50945 , n50940 , n50943 , n50944 );
and ( n50946 , n45060 , n41984 );
and ( n50947 , n45073 , n41982 );
nor ( n50948 , n50946 , n50947 );
xnor ( n50949 , n50948 , n41687 );
and ( n50950 , n50945 , n50949 );
xor ( n50951 , n50846 , n50848 );
xor ( n50952 , n50951 , n50851 );
and ( n50953 , n50949 , n50952 );
and ( n50954 , n50945 , n50952 );
or ( n50955 , n50950 , n50953 , n50954 );
and ( n50956 , n45073 , n41984 );
and ( n50957 , n45086 , n41982 );
nor ( n50958 , n50956 , n50957 );
xnor ( n50959 , n50958 , n41687 );
and ( n50960 , n50955 , n50959 );
xor ( n50961 , n50801 , n50854 );
xor ( n50962 , n50961 , n50857 );
and ( n50963 , n50959 , n50962 );
and ( n50964 , n50955 , n50962 );
or ( n50965 , n50960 , n50963 , n50964 );
and ( n50966 , n45086 , n41984 );
and ( n50967 , n45099 , n41982 );
nor ( n50968 , n50966 , n50967 );
xnor ( n50969 , n50968 , n41687 );
and ( n50970 , n50965 , n50969 );
xor ( n50971 , n50756 , n50860 );
xor ( n50972 , n50971 , n50863 );
and ( n50973 , n50969 , n50972 );
and ( n50974 , n50965 , n50972 );
or ( n50975 , n50970 , n50973 , n50974 );
and ( n50976 , n45099 , n41984 );
and ( n50977 , n45112 , n41982 );
nor ( n50978 , n50976 , n50977 );
xnor ( n50979 , n50978 , n41687 );
and ( n50980 , n50975 , n50979 );
xor ( n50981 , n50866 , n50870 );
xor ( n50982 , n50981 , n50873 );
and ( n50983 , n50979 , n50982 );
and ( n50984 , n50975 , n50982 );
or ( n50985 , n50980 , n50983 , n50984 );
and ( n50986 , n50876 , n50985 );
xor ( n50987 , n50728 , n50732 );
xor ( n50988 , n50987 , n50735 );
and ( n50989 , n50985 , n50988 );
and ( n50990 , n50876 , n50988 );
or ( n50991 , n50986 , n50989 , n50990 );
and ( n50992 , n45125 , n41984 );
and ( n50993 , n45138 , n41982 );
nor ( n50994 , n50992 , n50993 );
xnor ( n50995 , n50994 , n41687 );
and ( n50996 , n50991 , n50995 );
xor ( n50997 , n50708 , n50738 );
xor ( n50998 , n50997 , n50741 );
and ( n50999 , n50995 , n50998 );
and ( n51000 , n50991 , n50998 );
or ( n51001 , n50996 , n50999 , n51000 );
and ( n51002 , n50744 , n51001 );
xor ( n51003 , n50680 , n50684 );
xor ( n51004 , n51003 , n50687 );
and ( n51005 , n51001 , n51004 );
and ( n51006 , n50744 , n51004 );
or ( n51007 , n51002 , n51005 , n51006 );
and ( n51008 , n50696 , n51007 );
and ( n51009 , n45164 , n42269 );
and ( n51010 , n44665 , n42266 );
nor ( n51011 , n51009 , n51010 );
xnor ( n51012 , n51011 , n41684 );
xor ( n51013 , n50744 , n51001 );
xor ( n51014 , n51013 , n51004 );
and ( n51015 , n51012 , n51014 );
and ( n51016 , n45151 , n42269 );
and ( n51017 , n45164 , n42266 );
nor ( n51018 , n51016 , n51017 );
xnor ( n51019 , n51018 , n41684 );
xor ( n51020 , n50991 , n50995 );
xor ( n51021 , n51020 , n50998 );
and ( n51022 , n51019 , n51021 );
and ( n51023 , n45138 , n42269 );
and ( n51024 , n45151 , n42266 );
nor ( n51025 , n51023 , n51024 );
xnor ( n51026 , n51025 , n41684 );
xor ( n51027 , n50876 , n50985 );
xor ( n51028 , n51027 , n50988 );
and ( n51029 , n51026 , n51028 );
and ( n51030 , n45125 , n42269 );
and ( n51031 , n45138 , n42266 );
nor ( n51032 , n51030 , n51031 );
xnor ( n51033 , n51032 , n41684 );
xor ( n51034 , n50975 , n50979 );
xor ( n51035 , n51034 , n50982 );
and ( n51036 , n51033 , n51035 );
and ( n51037 , n45112 , n42269 );
and ( n51038 , n45125 , n42266 );
nor ( n51039 , n51037 , n51038 );
xnor ( n51040 , n51039 , n41684 );
xor ( n51041 , n50965 , n50969 );
xor ( n51042 , n51041 , n50972 );
and ( n51043 , n51040 , n51042 );
and ( n51044 , n45099 , n42269 );
and ( n51045 , n45112 , n42266 );
nor ( n51046 , n51044 , n51045 );
xnor ( n51047 , n51046 , n41684 );
xor ( n51048 , n50955 , n50959 );
xor ( n51049 , n51048 , n50962 );
and ( n51050 , n51047 , n51049 );
and ( n51051 , n45086 , n42269 );
and ( n51052 , n45099 , n42266 );
nor ( n51053 , n51051 , n51052 );
xnor ( n51054 , n51053 , n41684 );
xor ( n51055 , n50945 , n50949 );
xor ( n51056 , n51055 , n50952 );
and ( n51057 , n51054 , n51056 );
and ( n51058 , n45073 , n42269 );
and ( n51059 , n45086 , n42266 );
nor ( n51060 , n51058 , n51059 );
xnor ( n51061 , n51060 , n41684 );
xor ( n51062 , n50935 , n50939 );
xor ( n51063 , n51062 , n50942 );
and ( n51064 , n51061 , n51063 );
and ( n51065 , n45060 , n42269 );
and ( n51066 , n45073 , n42266 );
nor ( n51067 , n51065 , n51066 );
xnor ( n51068 , n51067 , n41684 );
xor ( n51069 , n50925 , n50929 );
xor ( n51070 , n51069 , n50932 );
and ( n51071 , n51068 , n51070 );
and ( n51072 , n45047 , n42269 );
and ( n51073 , n45060 , n42266 );
nor ( n51074 , n51072 , n51073 );
xnor ( n51075 , n51074 , n41684 );
xor ( n51076 , n50915 , n50919 );
xor ( n51077 , n51076 , n50922 );
and ( n51078 , n51075 , n51077 );
and ( n51079 , n45034 , n42269 );
and ( n51080 , n45047 , n42266 );
nor ( n51081 , n51079 , n51080 );
xnor ( n51082 , n51081 , n41684 );
xor ( n51083 , n50905 , n50909 );
xor ( n51084 , n51083 , n50912 );
and ( n51085 , n51082 , n51084 );
and ( n51086 , n45021 , n42269 );
and ( n51087 , n45034 , n42266 );
nor ( n51088 , n51086 , n51087 );
xnor ( n51089 , n51088 , n41684 );
xor ( n51090 , n50895 , n50899 );
xor ( n51091 , n51090 , n50902 );
and ( n51092 , n51089 , n51091 );
and ( n51093 , n45008 , n42269 );
and ( n51094 , n45021 , n42266 );
nor ( n51095 , n51093 , n51094 );
xnor ( n51096 , n51095 , n41684 );
xor ( n51097 , n50877 , n50889 );
xor ( n51098 , n51097 , n50892 );
and ( n51099 , n51096 , n51098 );
and ( n51100 , n44999 , n42269 );
and ( n51101 , n45008 , n42266 );
nor ( n51102 , n51100 , n51101 );
xnor ( n51103 , n51102 , n41684 );
xor ( n51104 , n50883 , n50803 );
xor ( n51105 , n51104 , n50886 );
and ( n51106 , n51103 , n51105 );
and ( n51107 , n44991 , n42269 );
and ( n51108 , n44999 , n42266 );
nor ( n51109 , n51107 , n51108 );
xnor ( n51110 , n51109 , n41684 );
xor ( n51111 , n50880 , n50882 );
and ( n51112 , n51110 , n51111 );
buf ( n51113 , n557832 );
not ( n51114 , n51113 );
or ( n51115 , n50878 , n51114 );
and ( n51116 , n51111 , n51115 );
and ( n51117 , n51110 , n51115 );
or ( n51118 , n51112 , n51116 , n51117 );
and ( n51119 , n51105 , n51118 );
and ( n51120 , n51103 , n51118 );
or ( n51121 , n51106 , n51119 , n51120 );
and ( n51122 , n51098 , n51121 );
and ( n51123 , n51096 , n51121 );
or ( n51124 , n51099 , n51122 , n51123 );
and ( n51125 , n51091 , n51124 );
and ( n51126 , n51089 , n51124 );
or ( n51127 , n51092 , n51125 , n51126 );
and ( n51128 , n51084 , n51127 );
and ( n51129 , n51082 , n51127 );
or ( n51130 , n51085 , n51128 , n51129 );
and ( n51131 , n51077 , n51130 );
and ( n51132 , n51075 , n51130 );
or ( n51133 , n51078 , n51131 , n51132 );
and ( n51134 , n51070 , n51133 );
and ( n51135 , n51068 , n51133 );
or ( n51136 , n51071 , n51134 , n51135 );
and ( n51137 , n51063 , n51136 );
and ( n51138 , n51061 , n51136 );
or ( n51139 , n51064 , n51137 , n51138 );
and ( n51140 , n51056 , n51139 );
and ( n51141 , n51054 , n51139 );
or ( n51142 , n51057 , n51140 , n51141 );
and ( n51143 , n51049 , n51142 );
and ( n51144 , n51047 , n51142 );
or ( n51145 , n51050 , n51143 , n51144 );
and ( n51146 , n51042 , n51145 );
and ( n51147 , n51040 , n51145 );
or ( n51148 , n51043 , n51146 , n51147 );
and ( n51149 , n51035 , n51148 );
and ( n51150 , n51033 , n51148 );
or ( n51151 , n51036 , n51149 , n51150 );
and ( n51152 , n51028 , n51151 );
and ( n51153 , n51026 , n51151 );
or ( n51154 , n51029 , n51152 , n51153 );
and ( n51155 , n51021 , n51154 );
and ( n51156 , n51019 , n51154 );
or ( n51157 , n51022 , n51155 , n51156 );
and ( n51158 , n51014 , n51157 );
and ( n51159 , n51012 , n51157 );
or ( n51160 , n51015 , n51158 , n51159 );
and ( n51161 , n51007 , n51160 );
and ( n51162 , n50696 , n51160 );
or ( n51163 , n51008 , n51161 , n51162 );
and ( n51164 , n50693 , n51163 );
and ( n51165 , n50580 , n51163 );
or ( n51166 , n50694 , n51164 , n51165 );
and ( n51167 , n50577 , n51166 );
and ( n51168 , n50413 , n51166 );
or ( n51169 , n50578 , n51167 , n51168 );
and ( n51170 , n50410 , n51169 );
and ( n51171 , n50408 , n51169 );
or ( n51172 , n50411 , n51170 , n51171 );
and ( n51173 , n50383 , n51172 );
and ( n51174 , n50381 , n51173 );
or ( n51175 , n50380 , n51174 );
and ( n51176 , n50350 , n51175 );
and ( n51177 , n50348 , n51176 );
or ( n51178 , n50347 , n51177 );
and ( n51179 , n50102 , n51178 );
and ( n51180 , n50100 , n51179 );
and ( n51181 , n50098 , n51180 );
or ( n51182 , n50097 , n51181 );
and ( n51183 , n50092 , n51182 );
and ( n51184 , n50090 , n51183 );
or ( n51185 , n50089 , n51184 );
and ( n51186 , n50084 , n51185 );
and ( n51187 , n50082 , n51186 );
and ( n51188 , n50080 , n51187 );
or ( n51189 , n50079 , n51188 );
and ( n51190 , n50074 , n51189 );
and ( n51191 , n50072 , n51190 );
and ( n51192 , n50070 , n51191 );
and ( n51193 , n50068 , n51192 );
and ( n51194 , n50066 , n51193 );
and ( n51195 , n50064 , n51194 );
and ( n51196 , n50062 , n51195 );
and ( n51197 , n50060 , n51196 );
and ( n51198 , n50058 , n51197 );
and ( n51199 , n50056 , n51198 );
and ( n51200 , n50054 , n51199 );
and ( n51201 , n50052 , n51200 );
and ( n51202 , n50050 , n51201 );
and ( n51203 , n577360 , n51202 );
and ( n51204 , n577358 , n51203 );
and ( n51205 , n50047 , n51204 );
and ( n51206 , n50045 , n51205 );
and ( n51207 , n50043 , n51206 );
and ( n51208 , n50041 , n51207 );
and ( n51209 , n50039 , n51208 );
and ( n51210 , n50037 , n51209 );
and ( n51211 , n50035 , n51210 );
and ( n51212 , n50033 , n51211 );
or ( n51213 , n50032 , n51212 );
and ( n51214 , n45992 , n51213 );
or ( n51215 , n45991 , n51214 );
and ( n51216 , n45509 , n51215 );
and ( n51217 , n45507 , n51216 );
and ( n51218 , n45505 , n51217 );
and ( n51219 , n45503 , n51218 );
or ( n51220 , n45502 , n51219 );
and ( n51221 , n44441 , n51220 );
and ( n51222 , n44439 , n51221 );
or ( n51223 , n44438 , n51222 );
and ( n51224 , n44433 , n51223 );
and ( n51225 , n44431 , n51224 );
and ( n51226 , n44429 , n51225 );
or ( n51227 , n44428 , n51226 );
and ( n51228 , n44053 , n51227 );
and ( n51229 , n44051 , n51228 );
and ( n51230 , n44049 , n51229 );
and ( n51231 , n44048 , n51230 );
or ( n51232 , n44047 , n51231 );
and ( n51233 , n44045 , n51232 );
and ( n51234 , n44044 , n51233 );
and ( n51235 , n44043 , n51234 );
or ( n51236 , n44042 , n51235 );
and ( n51237 , n43134 , n51236 );
or ( n51238 , n43133 , n51237 );
and ( n51239 , n42231 , n51238 );
and ( n51240 , n42229 , n51239 );
and ( n51241 , n42227 , n51240 );
and ( n51242 , n42226 , n51241 );
or ( n51243 , n42225 , n51242 );
and ( n51244 , n42223 , n51243 );
and ( n51245 , n42222 , n51244 );
and ( n51246 , n42221 , n51245 );
and ( n51247 , n42220 , n51246 );
and ( n51248 , n42219 , n51247 );
and ( n51249 , n42218 , n51248 );
and ( n51250 , n42217 , n51249 );
and ( n51251 , n42216 , n51250 );
and ( n51252 , n42215 , n51251 );
and ( n51253 , n42214 , n51252 );
and ( n51254 , n42213 , n51253 );
and ( n51255 , n42212 , n51254 );
and ( n51256 , n42211 , n51255 );
and ( n51257 , n42210 , n51256 );
and ( n51258 , n42209 , n51257 );
and ( n51259 , n42208 , n51258 );
and ( n51260 , n42207 , n51259 );
and ( n51261 , n42206 , n51260 );
and ( n51262 , n42205 , n51261 );
and ( n51263 , n42204 , n51262 );
and ( n51264 , n42203 , n51263 );
and ( n51265 , n42201 , n51264 );
or ( n51266 , n42200 , n51265 );
not ( n51267 , n51266 );
buf ( n51268 , n51267 );
buf ( n578582 , n51268 );
buf ( n51270 , n51267 );
buf ( n578584 , n51270 );
buf ( n51272 , n51267 );
buf ( n578586 , n51272 );
buf ( n51274 , n51267 );
buf ( n578588 , n51274 );
buf ( n51276 , n51267 );
buf ( n578590 , n51276 );
buf ( n51278 , n51267 );
buf ( n578592 , n51278 );
buf ( n51280 , n51267 );
buf ( n578594 , n51280 );
buf ( n51282 , n51267 );
buf ( n578596 , n51282 );
buf ( n51284 , n51267 );
buf ( n578598 , n51284 );
buf ( n51286 , n51267 );
buf ( n578600 , n51286 );
buf ( n51288 , n51267 );
buf ( n578602 , n51288 );
buf ( n51290 , n51267 );
buf ( n578604 , n51290 );
buf ( n51292 , n51267 );
buf ( n578606 , n51292 );
buf ( n51294 , n51267 );
buf ( n578608 , n51294 );
buf ( n51296 , n51267 );
buf ( n578610 , n51296 );
buf ( n51298 , n51267 );
buf ( n578612 , n51298 );
buf ( n51300 , n51267 );
buf ( n578614 , n51300 );
buf ( n51302 , n51267 );
buf ( n578616 , n51302 );
buf ( n51304 , n51267 );
buf ( n578618 , n51304 );
buf ( n51306 , n51267 );
buf ( n578620 , n51306 );
buf ( n51308 , n51267 );
buf ( n578622 , n51308 );
buf ( n51310 , n51267 );
buf ( n578624 , n51310 );
buf ( n51312 , n51267 );
buf ( n578626 , n51312 );
buf ( n51314 , n51267 );
buf ( n578628 , n51314 );
buf ( n51316 , n51267 );
buf ( n578630 , n51316 );
buf ( n51318 , n51267 );
buf ( n578632 , n51318 );
buf ( n51320 , n51267 );
buf ( n578634 , n51320 );
buf ( n51322 , n51267 );
buf ( n578636 , n51322 );
buf ( n51324 , n51267 );
buf ( n578638 , n51324 );
buf ( n578639 , n51267 );
xor ( n51327 , n42201 , n51264 );
buf ( n578641 , n51327 );
xor ( n51329 , n42203 , n51263 );
buf ( n578643 , n51329 );
xor ( n51331 , n42204 , n51262 );
buf ( n578645 , n51331 );
xor ( n51333 , n42205 , n51261 );
buf ( n578647 , n51333 );
xor ( n51335 , n42206 , n51260 );
buf ( n578649 , n51335 );
xor ( n51337 , n42207 , n51259 );
buf ( n578651 , n51337 );
xor ( n51339 , n42208 , n51258 );
buf ( n578653 , n51339 );
xor ( n51341 , n42209 , n51257 );
buf ( n578655 , n51341 );
xor ( n51343 , n42210 , n51256 );
buf ( n578657 , n51343 );
xor ( n51345 , n42211 , n51255 );
buf ( n578659 , n51345 );
xor ( n51347 , n42212 , n51254 );
buf ( n578661 , n51347 );
xor ( n51349 , n42213 , n51253 );
buf ( n578663 , n51349 );
xor ( n51351 , n42214 , n51252 );
buf ( n578665 , n51351 );
xor ( n51353 , n42215 , n51251 );
buf ( n578667 , n51353 );
xor ( n51355 , n42216 , n51250 );
buf ( n578669 , n51355 );
xor ( n51357 , n42217 , n51249 );
buf ( n578671 , n51357 );
xor ( n51359 , n42218 , n51248 );
buf ( n578673 , n51359 );
xor ( n51361 , n42219 , n51247 );
buf ( n578675 , n51361 );
xor ( n51363 , n42220 , n51246 );
buf ( n578677 , n51363 );
xor ( n51365 , n42221 , n51245 );
buf ( n578679 , n51365 );
xor ( n578680 , n42222 , n51244 );
buf ( n578681 , n578680 );
xor ( n578682 , n42223 , n51243 );
buf ( n578683 , n578682 );
xor ( n51368 , n42226 , n51241 );
buf ( n578685 , n51368 );
xor ( n51370 , n42227 , n51240 );
buf ( n578687 , n51370 );
xor ( n51372 , n42229 , n51239 );
buf ( n578689 , n51372 );
xor ( n51374 , n42231 , n51238 );
buf ( n578691 , n51374 );
xor ( n51376 , n43134 , n51236 );
buf ( n578693 , n51376 );
xor ( n51378 , n44043 , n51234 );
buf ( n578695 , n51378 );
xor ( n51380 , n44044 , n51233 );
buf ( n578697 , n51380 );
xor ( n51382 , n44045 , n51232 );
buf ( n578699 , n51382 );
xor ( n51384 , n44048 , n51230 );
buf ( n578701 , n51384 );
xor ( n51386 , n44049 , n51229 );
buf ( n578703 , n51386 );
xor ( n51388 , n44051 , n51228 );
buf ( n578705 , n51388 );
xor ( n51390 , n44053 , n51227 );
buf ( n578707 , n51390 );
xor ( n51392 , n44429 , n51225 );
buf ( n578709 , n51392 );
xor ( n51394 , n44431 , n51224 );
buf ( n578711 , n51394 );
xor ( n51396 , n44433 , n51223 );
buf ( n578713 , n51396 );
xor ( n51398 , n44439 , n51221 );
buf ( n578715 , n51398 );
xor ( n51400 , n44441 , n51220 );
buf ( n578717 , n51400 );
xor ( n51402 , n45503 , n51218 );
buf ( n578719 , n51402 );
xor ( n51404 , n45505 , n51217 );
buf ( n578721 , n51404 );
xor ( n51406 , n45507 , n51216 );
buf ( n578723 , n51406 );
xor ( n51408 , n45509 , n51215 );
buf ( n578725 , n51408 );
xor ( n51410 , n45992 , n51213 );
buf ( n578727 , n51410 );
xor ( n51412 , n50033 , n51211 );
buf ( n578729 , n51412 );
xor ( n51414 , n50035 , n51210 );
buf ( n578731 , n51414 );
xor ( n51416 , n50037 , n51209 );
buf ( n578733 , n51416 );
xor ( n51418 , n50039 , n51208 );
buf ( n578735 , n51418 );
xor ( n51420 , n50041 , n51207 );
buf ( n578737 , n51420 );
xor ( n51422 , n50043 , n51206 );
buf ( n578739 , n51422 );
xor ( n51424 , n50045 , n51205 );
buf ( n578741 , n51424 );
xor ( n51426 , n50047 , n51204 );
buf ( n578743 , n51426 );
xor ( n51428 , n577358 , n51203 );
buf ( n578745 , n51428 );
xor ( n51430 , n577360 , n51202 );
buf ( n578747 , n51430 );
xor ( n51432 , n50050 , n51201 );
buf ( n578749 , n51432 );
xor ( n51434 , n50052 , n51200 );
buf ( n578751 , n51434 );
xor ( n51436 , n50054 , n51199 );
buf ( n578753 , n51436 );
xor ( n51438 , n50056 , n51198 );
buf ( n578755 , n51438 );
xor ( n51440 , n50058 , n51197 );
buf ( n578757 , n51440 );
xor ( n51442 , n50060 , n51196 );
buf ( n578759 , n51442 );
xor ( n51444 , n50062 , n51195 );
buf ( n578761 , n51444 );
xor ( n51446 , n50064 , n51194 );
buf ( n578763 , n51446 );
xor ( n51448 , n50066 , n51193 );
buf ( n578765 , n51448 );
xor ( n51450 , n50068 , n51192 );
buf ( n578767 , n51450 );
xor ( n51452 , n50070 , n51191 );
buf ( n578769 , n51452 );
xor ( n51454 , n50072 , n51190 );
buf ( n578771 , n51454 );
xor ( n51456 , n50074 , n51189 );
buf ( n578773 , n51456 );
xor ( n51458 , n50080 , n51187 );
buf ( n578775 , n51458 );
xor ( n51460 , n50082 , n51186 );
buf ( n578777 , n51460 );
xor ( n51462 , n50084 , n51185 );
buf ( n578779 , n51462 );
xor ( n51464 , n50090 , n51183 );
buf ( n578781 , n51464 );
xor ( n51466 , n50092 , n51182 );
buf ( n578783 , n51466 );
xor ( n51468 , n50098 , n51180 );
buf ( n578785 , n51468 );
xor ( n51470 , n50100 , n51179 );
buf ( n578787 , n51470 );
xor ( n51472 , n50102 , n51178 );
buf ( n578789 , n51472 );
xor ( n51474 , n50348 , n51176 );
buf ( n578791 , n51474 );
xor ( n51476 , n50350 , n51175 );
buf ( n578793 , n51476 );
xor ( n51478 , n50381 , n51173 );
buf ( n578795 , n51478 );
xor ( n51480 , n50383 , n51172 );
buf ( n578797 , n51480 );
xor ( n51482 , n50408 , n50410 );
xor ( n51483 , n51482 , n51169 );
buf ( n578800 , n51483 );
xor ( n51485 , n50413 , n50577 );
xor ( n51486 , n51485 , n51166 );
buf ( n578803 , n51486 );
xor ( n51488 , n50580 , n50693 );
xor ( n51489 , n51488 , n51163 );
buf ( n578806 , n51489 );
xor ( n51491 , n50696 , n51007 );
xor ( n51492 , n51491 , n51160 );
buf ( n578809 , n51492 );
xor ( n51494 , n51012 , n51014 );
xor ( n51495 , n51494 , n51157 );
buf ( n578812 , n51495 );
xor ( n51497 , n51019 , n51021 );
xor ( n51498 , n51497 , n51154 );
buf ( n578815 , n51498 );
xor ( n51500 , n51026 , n51028 );
xor ( n51501 , n51500 , n51151 );
buf ( n578818 , n51501 );
xor ( n51503 , n51033 , n51035 );
xor ( n51504 , n51503 , n51148 );
buf ( n578821 , n51504 );
xor ( n51506 , n51040 , n51042 );
xor ( n51507 , n51506 , n51145 );
buf ( n578824 , n51507 );
xor ( n51509 , n51047 , n51049 );
xor ( n51510 , n51509 , n51142 );
buf ( n578827 , n51510 );
xor ( n51512 , n51054 , n51056 );
xor ( n51513 , n51512 , n51139 );
buf ( n578830 , n51513 );
xor ( n51515 , n51061 , n51063 );
xor ( n51516 , n51515 , n51136 );
buf ( n578833 , n51516 );
xor ( n51518 , n51068 , n51070 );
xor ( n51519 , n51518 , n51133 );
buf ( n578836 , n51519 );
xor ( n51521 , n51075 , n51077 );
xor ( n51522 , n51521 , n51130 );
buf ( n578839 , n51522 );
xor ( n51524 , n51082 , n51084 );
xor ( n51525 , n51524 , n51127 );
buf ( n578842 , n51525 );
xor ( n51527 , n51089 , n51091 );
xor ( n51528 , n51527 , n51124 );
buf ( n578845 , n51528 );
xor ( n51530 , n51096 , n51098 );
xor ( n51531 , n51530 , n51121 );
buf ( n578848 , n51531 );
xor ( n51533 , n51103 , n51105 );
xor ( n51534 , n51533 , n51118 );
buf ( n578851 , n51534 );
xor ( n51536 , n51110 , n51111 );
xor ( n51537 , n51536 , n51115 );
buf ( n578854 , n51537 );
xnor ( n51539 , n50878 , n51114 );
buf ( n578856 , n51539 );
buf ( n578857 , n557576 );
buf ( n578858 , n557579 );
buf ( n578859 , n557582 );
buf ( n578860 , n557585 );
buf ( n578861 , n557588 );
buf ( n578862 , n557591 );
buf ( n578863 , n557594 );
buf ( n578864 , n557597 );
buf ( n578865 , n557600 );
buf ( n578866 , n557603 );
buf ( n578867 , n557606 );
buf ( n578868 , n557609 );
buf ( n578869 , n557612 );
buf ( n578870 , n557615 );
buf ( n578871 , n557618 );
buf ( n578872 , n557621 );
buf ( n578873 , n557624 );
buf ( n578874 , n557627 );
buf ( n578875 , n557630 );
buf ( n578876 , n557633 );
buf ( n578877 , n557636 );
buf ( n578878 , n557639 );
buf ( n578879 , n557642 );
buf ( n578880 , n557645 );
buf ( n578881 , n557648 );
buf ( n578882 , n557651 );
buf ( n578883 , n557654 );
buf ( n578884 , n557657 );
buf ( n578885 , n557660 );
buf ( n578886 , n557663 );
buf ( n578887 , n557666 );
buf ( n578888 , n557669 );
buf ( n578889 , n557672 );
buf ( n578890 , n557675 );
buf ( n578891 , n557678 );
buf ( n578892 , n557681 );
buf ( n578893 , n557684 );
buf ( n578894 , n557687 );
buf ( n578895 , n557690 );
buf ( n578896 , n557693 );
buf ( n578897 , n557696 );
buf ( n578898 , n557699 );
buf ( n578899 , n557702 );
buf ( n578900 , n557705 );
buf ( n578901 , n557708 );
buf ( n578902 , n557711 );
buf ( n578903 , n557714 );
buf ( n578904 , n557717 );
buf ( n578905 , n557720 );
buf ( n578906 , n557723 );
buf ( n578907 , n557726 );
buf ( n578908 , n557729 );
buf ( n578909 , n557732 );
buf ( n578910 , n557735 );
buf ( n578911 , n557738 );
buf ( n578912 , n557741 );
buf ( n578913 , n557744 );
buf ( n578914 , n557747 );
buf ( n578915 , n557750 );
buf ( n578916 , n557753 );
buf ( n578917 , n557756 );
buf ( n578918 , n557759 );
buf ( n578919 , n557762 );
buf ( n578920 , n557765 );
buf ( n578921 , n557767 );
buf ( n578922 , n1218 );
buf ( n578923 , n1186 );
and ( n51608 , n578922 , n578923 );
buf ( n578925 , n1219 );
buf ( n578926 , n1187 );
and ( n51611 , n578925 , n578926 );
buf ( n578928 , n1220 );
buf ( n578929 , n1188 );
and ( n51614 , n578928 , n578929 );
buf ( n578931 , n1221 );
buf ( n578932 , n1189 );
and ( n51617 , n578931 , n578932 );
buf ( n578934 , n1222 );
buf ( n578935 , n1190 );
and ( n51620 , n578934 , n578935 );
buf ( n578937 , n1223 );
buf ( n578938 , n1191 );
and ( n51623 , n578937 , n578938 );
buf ( n578940 , n1224 );
buf ( n578941 , n1192 );
and ( n51626 , n578940 , n578941 );
buf ( n578943 , n1225 );
buf ( n578944 , n1193 );
and ( n51629 , n578943 , n578944 );
buf ( n578946 , n1226 );
buf ( n578947 , n1194 );
and ( n51632 , n578946 , n578947 );
buf ( n578949 , n1227 );
buf ( n578950 , n1195 );
and ( n51635 , n578949 , n578950 );
buf ( n578952 , n1228 );
buf ( n578953 , n1196 );
and ( n51638 , n578952 , n578953 );
buf ( n578955 , n1229 );
buf ( n578956 , n1197 );
and ( n51641 , n578955 , n578956 );
buf ( n578958 , n1230 );
buf ( n578959 , n1198 );
and ( n51644 , n578958 , n578959 );
buf ( n578961 , n1231 );
buf ( n578962 , n1199 );
and ( n51647 , n578961 , n578962 );
buf ( n578964 , n1232 );
buf ( n578965 , n1200 );
and ( n51650 , n578964 , n578965 );
buf ( n578967 , n1233 );
buf ( n578968 , n1201 );
and ( n51653 , n578967 , n578968 );
buf ( n578970 , n1234 );
buf ( n578971 , n1202 );
and ( n51656 , n578970 , n578971 );
buf ( n578973 , n1235 );
buf ( n578974 , n1203 );
and ( n51659 , n578973 , n578974 );
buf ( n578976 , n1236 );
buf ( n578977 , n1204 );
and ( n51662 , n578976 , n578977 );
buf ( n578979 , n1237 );
buf ( n578980 , n1205 );
and ( n51665 , n578979 , n578980 );
buf ( n578982 , n1238 );
buf ( n578983 , n1206 );
and ( n51668 , n578982 , n578983 );
buf ( n578985 , n1239 );
buf ( n578986 , n1207 );
and ( n51671 , n578985 , n578986 );
buf ( n578988 , n1240 );
buf ( n578989 , n1208 );
and ( n51674 , n578988 , n578989 );
buf ( n578991 , n1241 );
buf ( n578992 , n1209 );
and ( n51677 , n578991 , n578992 );
buf ( n578994 , n1242 );
buf ( n578995 , n1210 );
and ( n51680 , n578994 , n578995 );
buf ( n578997 , n1243 );
buf ( n578998 , n1211 );
and ( n51683 , n578997 , n578998 );
buf ( n579000 , n1244 );
buf ( n579001 , n1212 );
and ( n51686 , n579000 , n579001 );
buf ( n579003 , n1245 );
buf ( n579004 , n1213 );
and ( n51689 , n579003 , n579004 );
buf ( n579006 , n1246 );
buf ( n579007 , n1214 );
and ( n51692 , n579006 , n579007 );
buf ( n579009 , n1247 );
buf ( n579010 , n1215 );
and ( n51695 , n579009 , n579010 );
buf ( n579012 , n1248 );
buf ( n579013 , n1216 );
and ( n51698 , n579012 , n579013 );
buf ( n579015 , n1249 );
buf ( n579016 , n1217 );
and ( n51701 , n579015 , n579016 );
and ( n51702 , n579013 , n51701 );
and ( n51703 , n579012 , n51701 );
or ( n51704 , n51698 , n51702 , n51703 );
and ( n51705 , n579010 , n51704 );
and ( n51706 , n579009 , n51704 );
or ( n51707 , n51695 , n51705 , n51706 );
and ( n51708 , n579007 , n51707 );
and ( n51709 , n579006 , n51707 );
or ( n51710 , n51692 , n51708 , n51709 );
and ( n51711 , n579004 , n51710 );
and ( n51712 , n579003 , n51710 );
or ( n51713 , n51689 , n51711 , n51712 );
and ( n51714 , n579001 , n51713 );
and ( n51715 , n579000 , n51713 );
or ( n51716 , n51686 , n51714 , n51715 );
and ( n51717 , n578998 , n51716 );
and ( n51718 , n578997 , n51716 );
or ( n51719 , n51683 , n51717 , n51718 );
and ( n51720 , n578995 , n51719 );
and ( n51721 , n578994 , n51719 );
or ( n51722 , n51680 , n51720 , n51721 );
and ( n51723 , n578992 , n51722 );
and ( n51724 , n578991 , n51722 );
or ( n51725 , n51677 , n51723 , n51724 );
and ( n51726 , n578989 , n51725 );
and ( n51727 , n578988 , n51725 );
or ( n51728 , n51674 , n51726 , n51727 );
and ( n51729 , n578986 , n51728 );
and ( n51730 , n578985 , n51728 );
or ( n51731 , n51671 , n51729 , n51730 );
and ( n51732 , n578983 , n51731 );
and ( n51733 , n578982 , n51731 );
or ( n51734 , n51668 , n51732 , n51733 );
and ( n51735 , n578980 , n51734 );
and ( n51736 , n578979 , n51734 );
or ( n51737 , n51665 , n51735 , n51736 );
and ( n51738 , n578977 , n51737 );
and ( n51739 , n578976 , n51737 );
or ( n51740 , n51662 , n51738 , n51739 );
and ( n51741 , n578974 , n51740 );
and ( n51742 , n578973 , n51740 );
or ( n51743 , n51659 , n51741 , n51742 );
and ( n51744 , n578971 , n51743 );
and ( n51745 , n578970 , n51743 );
or ( n51746 , n51656 , n51744 , n51745 );
and ( n51747 , n578968 , n51746 );
and ( n51748 , n578967 , n51746 );
or ( n51749 , n51653 , n51747 , n51748 );
and ( n51750 , n578965 , n51749 );
and ( n51751 , n578964 , n51749 );
or ( n51752 , n51650 , n51750 , n51751 );
and ( n51753 , n578962 , n51752 );
and ( n51754 , n578961 , n51752 );
or ( n51755 , n51647 , n51753 , n51754 );
and ( n51756 , n578959 , n51755 );
and ( n51757 , n578958 , n51755 );
or ( n51758 , n51644 , n51756 , n51757 );
and ( n51759 , n578956 , n51758 );
and ( n51760 , n578955 , n51758 );
or ( n51761 , n51641 , n51759 , n51760 );
and ( n51762 , n578953 , n51761 );
and ( n51763 , n578952 , n51761 );
or ( n51764 , n51638 , n51762 , n51763 );
and ( n51765 , n578950 , n51764 );
and ( n51766 , n578949 , n51764 );
or ( n51767 , n51635 , n51765 , n51766 );
and ( n51768 , n578947 , n51767 );
and ( n51769 , n578946 , n51767 );
or ( n51770 , n51632 , n51768 , n51769 );
and ( n51771 , n578944 , n51770 );
and ( n51772 , n578943 , n51770 );
or ( n51773 , n51629 , n51771 , n51772 );
and ( n51774 , n578941 , n51773 );
and ( n51775 , n578940 , n51773 );
or ( n51776 , n51626 , n51774 , n51775 );
and ( n51777 , n578938 , n51776 );
and ( n51778 , n578937 , n51776 );
or ( n51779 , n51623 , n51777 , n51778 );
and ( n51780 , n578935 , n51779 );
and ( n51781 , n578934 , n51779 );
or ( n51782 , n51620 , n51780 , n51781 );
and ( n51783 , n578932 , n51782 );
and ( n51784 , n578931 , n51782 );
or ( n51785 , n51617 , n51783 , n51784 );
and ( n51786 , n578929 , n51785 );
and ( n51787 , n578928 , n51785 );
or ( n51788 , n51614 , n51786 , n51787 );
and ( n51789 , n578926 , n51788 );
and ( n51790 , n578925 , n51788 );
or ( n51791 , n51611 , n51789 , n51790 );
and ( n51792 , n578923 , n51791 );
and ( n51793 , n578922 , n51791 );
or ( n51794 , n51608 , n51792 , n51793 );
buf ( n579111 , n51794 );
buf ( n579112 , n579111 );
xor ( n51797 , n578922 , n578923 );
xor ( n51798 , n51797 , n51791 );
buf ( n579115 , n51798 );
buf ( n579116 , n579115 );
xor ( n51801 , n578925 , n578926 );
xor ( n51802 , n51801 , n51788 );
buf ( n579119 , n51802 );
buf ( n579120 , n579119 );
xor ( n51805 , n578928 , n578929 );
xor ( n51806 , n51805 , n51785 );
buf ( n579123 , n51806 );
buf ( n579124 , n579123 );
xor ( n51809 , n578931 , n578932 );
xor ( n51810 , n51809 , n51782 );
buf ( n579127 , n51810 );
buf ( n579128 , n579127 );
xor ( n51813 , n578934 , n578935 );
xor ( n51814 , n51813 , n51779 );
buf ( n579131 , n51814 );
buf ( n579132 , n579131 );
xor ( n51817 , n578937 , n578938 );
xor ( n51818 , n51817 , n51776 );
buf ( n579135 , n51818 );
buf ( n579136 , n579135 );
xor ( n51821 , n578940 , n578941 );
xor ( n51822 , n51821 , n51773 );
buf ( n579139 , n51822 );
buf ( n579140 , n579139 );
xor ( n51825 , n578943 , n578944 );
xor ( n51826 , n51825 , n51770 );
buf ( n579143 , n51826 );
buf ( n579144 , n579143 );
xor ( n51829 , n578946 , n578947 );
xor ( n51830 , n51829 , n51767 );
buf ( n579147 , n51830 );
buf ( n579148 , n579147 );
xor ( n51833 , n578949 , n578950 );
xor ( n51834 , n51833 , n51764 );
buf ( n579151 , n51834 );
buf ( n579152 , n579151 );
xor ( n51837 , n578952 , n578953 );
xor ( n51838 , n51837 , n51761 );
buf ( n579155 , n51838 );
buf ( n579156 , n579155 );
xor ( n51841 , n578955 , n578956 );
xor ( n51842 , n51841 , n51758 );
buf ( n579159 , n51842 );
buf ( n579160 , n579159 );
xor ( n51845 , n578958 , n578959 );
xor ( n51846 , n51845 , n51755 );
buf ( n579163 , n51846 );
buf ( n579164 , n579163 );
xor ( n51849 , n578961 , n578962 );
xor ( n51850 , n51849 , n51752 );
buf ( n579167 , n51850 );
buf ( n579168 , n579167 );
xor ( n51853 , n578964 , n578965 );
xor ( n51854 , n51853 , n51749 );
buf ( n579171 , n51854 );
buf ( n579172 , n579171 );
xor ( n51857 , n578967 , n578968 );
xor ( n51858 , n51857 , n51746 );
buf ( n579175 , n51858 );
buf ( n579176 , n579175 );
xor ( n51861 , n578970 , n578971 );
xor ( n51862 , n51861 , n51743 );
buf ( n579179 , n51862 );
buf ( n579180 , n579179 );
xor ( n51865 , n578973 , n578974 );
xor ( n51866 , n51865 , n51740 );
buf ( n579183 , n51866 );
buf ( n579184 , n579183 );
xor ( n51869 , n578976 , n578977 );
xor ( n51870 , n51869 , n51737 );
buf ( n579187 , n51870 );
buf ( n579188 , n579187 );
xor ( n51873 , n578979 , n578980 );
xor ( n51874 , n51873 , n51734 );
buf ( n579191 , n51874 );
buf ( n579192 , n579191 );
xor ( n51877 , n578982 , n578983 );
xor ( n51878 , n51877 , n51731 );
buf ( n579195 , n51878 );
buf ( n579196 , n579195 );
xor ( n51881 , n578985 , n578986 );
xor ( n51882 , n51881 , n51728 );
buf ( n579199 , n51882 );
buf ( n579200 , n579199 );
xor ( n51885 , n578988 , n578989 );
xor ( n51886 , n51885 , n51725 );
buf ( n579203 , n51886 );
buf ( n579204 , n579203 );
xor ( n51889 , n578991 , n578992 );
xor ( n51890 , n51889 , n51722 );
buf ( n579207 , n51890 );
buf ( n579208 , n579207 );
xor ( n51893 , n578994 , n578995 );
xor ( n51894 , n51893 , n51719 );
buf ( n579211 , n51894 );
buf ( n579212 , n579211 );
xor ( n51897 , n578997 , n578998 );
xor ( n51898 , n51897 , n51716 );
buf ( n579215 , n51898 );
buf ( n579216 , n579215 );
xor ( n51901 , n579000 , n579001 );
xor ( n51902 , n51901 , n51713 );
buf ( n579219 , n51902 );
buf ( n579220 , n579219 );
xor ( n51905 , n579003 , n579004 );
xor ( n51906 , n51905 , n51710 );
buf ( n579223 , n51906 );
buf ( n579224 , n579223 );
xor ( n51909 , n579006 , n579007 );
xor ( n51910 , n51909 , n51707 );
buf ( n579227 , n51910 );
buf ( n579228 , n579227 );
xor ( n51913 , n579009 , n579010 );
xor ( n51914 , n51913 , n51704 );
buf ( n579231 , n51914 );
buf ( n579232 , n579231 );
xor ( n51917 , n579012 , n579013 );
xor ( n51918 , n51917 , n51701 );
buf ( n579235 , n51918 );
buf ( n579236 , n579235 );
xor ( n51921 , n579015 , n579016 );
buf ( n579238 , n51921 );
buf ( n579239 , n579238 );
buf ( n51924 , n578857 );
buf ( n51925 , n579112 );
buf ( n51926 , n579116 );
xor ( n51927 , n51925 , n51926 );
not ( n51928 , n51927 );
and ( n51929 , n51925 , n51928 );
and ( n51930 , n51924 , n51929 );
buf ( n51931 , n579120 );
xor ( n51932 , n51926 , n51931 );
buf ( n51933 , n579124 );
xor ( n51934 , n51931 , n51933 );
not ( n51935 , n51934 );
and ( n51936 , n51932 , n51935 );
and ( n51937 , n51924 , n51936 );
not ( n51938 , n51937 );
and ( n51939 , n51931 , n51933 );
not ( n51940 , n51939 );
and ( n51941 , n51926 , n51940 );
xnor ( n51942 , n51938 , n51941 );
buf ( n51943 , n51942 );
not ( n51944 , n51941 );
and ( n51945 , n51943 , n51944 );
buf ( n51946 , n578858 );
and ( n51947 , n51946 , n51929 );
and ( n51948 , n51924 , n51927 );
nor ( n51949 , n51947 , n51948 );
not ( n51950 , n51949 );
and ( n51951 , n51944 , n51950 );
and ( n51952 , n51943 , n51950 );
or ( n51953 , n51945 , n51951 , n51952 );
xor ( n51954 , n51930 , n51953 );
buf ( n51955 , n579128 );
buf ( n51956 , n579132 );
and ( n51957 , n51955 , n51956 );
not ( n51958 , n51957 );
and ( n51959 , n51933 , n51958 );
not ( n51960 , n51959 );
and ( n51961 , n51946 , n51936 );
and ( n51962 , n51924 , n51934 );
nor ( n51963 , n51961 , n51962 );
xnor ( n51964 , n51963 , n51941 );
and ( n579281 , n51960 , n51964 );
buf ( n51965 , n578860 );
and ( n51966 , n51965 , n51929 );
buf ( n51967 , n578859 );
and ( n51968 , n51967 , n51927 );
nor ( n51969 , n51966 , n51968 );
not ( n51970 , n51969 );
and ( n51971 , n51964 , n51970 );
and ( n51972 , n51960 , n51970 );
or ( n51973 , n579281 , n51971 , n51972 );
not ( n51974 , n51942 );
and ( n51975 , n51973 , n51974 );
and ( n51976 , n51967 , n51929 );
and ( n51977 , n51946 , n51927 );
nor ( n51978 , n51976 , n51977 );
not ( n51979 , n51978 );
and ( n51980 , n51974 , n51979 );
and ( n51981 , n51973 , n51979 );
or ( n51982 , n51975 , n51980 , n51981 );
xor ( n51983 , n51943 , n51944 );
xor ( n51984 , n51983 , n51950 );
and ( n51985 , n51982 , n51984 );
xor ( n51986 , n51973 , n51974 );
xor ( n51987 , n51986 , n51979 );
xor ( n51988 , n51933 , n51955 );
xor ( n51989 , n51955 , n51956 );
not ( n51990 , n51989 );
and ( n51991 , n51988 , n51990 );
and ( n51992 , n51924 , n51991 );
not ( n51993 , n51992 );
xnor ( n51994 , n51993 , n51959 );
and ( n51995 , n51967 , n51936 );
and ( n51996 , n51946 , n51934 );
nor ( n51997 , n51995 , n51996 );
xnor ( n51998 , n51997 , n51941 );
and ( n51999 , n51994 , n51998 );
buf ( n52000 , n578861 );
and ( n52001 , n52000 , n51929 );
and ( n52002 , n51965 , n51927 );
nor ( n52003 , n52001 , n52002 );
and ( n52004 , n51998 , n52003 );
and ( n52005 , n51994 , n52003 );
or ( n52006 , n51999 , n52004 , n52005 );
not ( n52007 , n52003 );
buf ( n52008 , n52007 );
and ( n52009 , n52006 , n52008 );
xor ( n52010 , n51960 , n51964 );
xor ( n52011 , n52010 , n51970 );
and ( n52012 , n52008 , n52011 );
and ( n52013 , n52006 , n52011 );
or ( n52014 , n52009 , n52012 , n52013 );
and ( n52015 , n51987 , n52014 );
xor ( n52016 , n52006 , n52008 );
xor ( n52017 , n52016 , n52011 );
buf ( n52018 , n579136 );
buf ( n52019 , n579140 );
and ( n52020 , n52018 , n52019 );
not ( n52021 , n52020 );
and ( n52022 , n51956 , n52021 );
not ( n52023 , n52022 );
and ( n52024 , n51965 , n51936 );
and ( n52025 , n51967 , n51934 );
nor ( n52026 , n52024 , n52025 );
xnor ( n52027 , n52026 , n51941 );
and ( n52028 , n52023 , n52027 );
buf ( n52029 , n578862 );
and ( n52030 , n52029 , n51929 );
and ( n52031 , n52000 , n51927 );
nor ( n52032 , n52030 , n52031 );
not ( n52033 , n52032 );
and ( n52034 , n52027 , n52033 );
and ( n52035 , n52023 , n52033 );
or ( n52036 , n52028 , n52034 , n52035 );
buf ( n52037 , n578863 );
and ( n52038 , n52037 , n51929 );
and ( n52039 , n52029 , n51927 );
nor ( n52040 , n52038 , n52039 );
not ( n52041 , n52040 );
buf ( n52042 , n52041 );
and ( n52043 , n51946 , n51991 );
and ( n52044 , n51924 , n51989 );
nor ( n52045 , n52043 , n52044 );
xnor ( n52046 , n52045 , n51959 );
and ( n52047 , n52042 , n52046 );
xor ( n52048 , n52023 , n52027 );
xor ( n52049 , n52048 , n52033 );
and ( n52050 , n52046 , n52049 );
and ( n52051 , n52042 , n52049 );
or ( n52052 , n52047 , n52050 , n52051 );
and ( n52053 , n52036 , n52052 );
xor ( n52054 , n51994 , n51998 );
xor ( n52055 , n52054 , n52003 );
and ( n52056 , n52052 , n52055 );
and ( n52057 , n52036 , n52055 );
or ( n52058 , n52053 , n52056 , n52057 );
and ( n52059 , n52017 , n52058 );
xor ( n52060 , n52036 , n52052 );
xor ( n52061 , n52060 , n52055 );
xor ( n52062 , n51956 , n52018 );
xor ( n52063 , n52018 , n52019 );
not ( n52064 , n52063 );
and ( n52065 , n52062 , n52064 );
and ( n52066 , n51924 , n52065 );
not ( n52067 , n52066 );
xnor ( n52068 , n52067 , n52022 );
and ( n52069 , n51967 , n51991 );
and ( n52070 , n51946 , n51989 );
nor ( n52071 , n52069 , n52070 );
xnor ( n52072 , n52071 , n51959 );
and ( n52073 , n52068 , n52072 );
and ( n52074 , n52000 , n51936 );
and ( n52075 , n51965 , n51934 );
nor ( n52076 , n52074 , n52075 );
xnor ( n52077 , n52076 , n51941 );
and ( n52078 , n52072 , n52077 );
and ( n52079 , n52068 , n52077 );
or ( n52080 , n52073 , n52078 , n52079 );
buf ( n52081 , n579144 );
buf ( n52082 , n579148 );
and ( n52083 , n52081 , n52082 );
not ( n52084 , n52083 );
and ( n52085 , n52019 , n52084 );
not ( n52086 , n52085 );
and ( n52087 , n52029 , n51936 );
and ( n52088 , n52000 , n51934 );
nor ( n52089 , n52087 , n52088 );
xnor ( n52090 , n52089 , n51941 );
and ( n52091 , n52086 , n52090 );
buf ( n52092 , n578864 );
and ( n52093 , n52092 , n51929 );
and ( n52094 , n52037 , n51927 );
nor ( n52095 , n52093 , n52094 );
not ( n52096 , n52095 );
and ( n52097 , n52090 , n52096 );
and ( n52098 , n52086 , n52096 );
or ( n52099 , n52091 , n52097 , n52098 );
and ( n52100 , n52099 , n52040 );
xor ( n52101 , n52068 , n52072 );
xor ( n52102 , n52101 , n52077 );
and ( n52103 , n52040 , n52102 );
and ( n52104 , n52099 , n52102 );
or ( n52105 , n52100 , n52103 , n52104 );
and ( n52106 , n52080 , n52105 );
xor ( n52107 , n52042 , n52046 );
xor ( n52108 , n52107 , n52049 );
and ( n52109 , n52105 , n52108 );
and ( n52110 , n52080 , n52108 );
or ( n52111 , n52106 , n52109 , n52110 );
and ( n52112 , n52061 , n52111 );
xor ( n52113 , n52080 , n52105 );
xor ( n52114 , n52113 , n52108 );
buf ( n52115 , n578865 );
and ( n52116 , n52115 , n51929 );
and ( n52117 , n52092 , n51927 );
nor ( n52118 , n52116 , n52117 );
not ( n52119 , n52118 );
buf ( n52120 , n52119 );
and ( n52121 , n51946 , n52065 );
and ( n52122 , n51924 , n52063 );
nor ( n52123 , n52121 , n52122 );
xnor ( n52124 , n52123 , n52022 );
and ( n52125 , n52120 , n52124 );
and ( n52126 , n51965 , n51991 );
and ( n52127 , n51967 , n51989 );
nor ( n52128 , n52126 , n52127 );
xnor ( n52129 , n52128 , n51959 );
and ( n52130 , n52124 , n52129 );
and ( n52131 , n52120 , n52129 );
or ( n52132 , n52125 , n52130 , n52131 );
buf ( n52133 , n579152 );
buf ( n52134 , n579156 );
and ( n52135 , n52133 , n52134 );
not ( n52136 , n52135 );
and ( n52137 , n52082 , n52136 );
not ( n52138 , n52137 );
and ( n52139 , n52092 , n51936 );
and ( n52140 , n52037 , n51934 );
nor ( n52141 , n52139 , n52140 );
xnor ( n52142 , n52141 , n51941 );
and ( n52143 , n52138 , n52142 );
buf ( n52144 , n578866 );
and ( n52145 , n52144 , n51929 );
and ( n52146 , n52115 , n51927 );
nor ( n52147 , n52145 , n52146 );
not ( n52148 , n52147 );
and ( n52149 , n52142 , n52148 );
and ( n52150 , n52138 , n52148 );
or ( n52151 , n52143 , n52149 , n52150 );
xor ( n52152 , n52019 , n52081 );
xor ( n52153 , n52081 , n52082 );
not ( n52154 , n52153 );
and ( n52155 , n52152 , n52154 );
and ( n52156 , n51924 , n52155 );
not ( n52157 , n52156 );
xnor ( n52158 , n52157 , n52085 );
and ( n52159 , n52151 , n52158 );
and ( n52160 , n51967 , n52065 );
and ( n52161 , n51946 , n52063 );
nor ( n52162 , n52160 , n52161 );
xnor ( n52163 , n52162 , n52022 );
and ( n52164 , n52158 , n52163 );
and ( n52165 , n52151 , n52163 );
or ( n52166 , n52159 , n52164 , n52165 );
and ( n52167 , n52000 , n51991 );
and ( n52168 , n51965 , n51989 );
nor ( n52169 , n52167 , n52168 );
xnor ( n52170 , n52169 , n51959 );
and ( n52171 , n52037 , n51936 );
and ( n52172 , n52029 , n51934 );
nor ( n52173 , n52171 , n52172 );
xnor ( n52174 , n52173 , n51941 );
and ( n52175 , n52170 , n52174 );
and ( n52176 , n52174 , n52118 );
and ( n52177 , n52170 , n52118 );
or ( n52178 , n52175 , n52176 , n52177 );
and ( n52179 , n52166 , n52178 );
xor ( n52180 , n52086 , n52090 );
xor ( n52181 , n52180 , n52096 );
and ( n52182 , n52178 , n52181 );
and ( n52183 , n52166 , n52181 );
or ( n52184 , n52179 , n52182 , n52183 );
and ( n52185 , n52132 , n52184 );
xor ( n52186 , n52099 , n52040 );
xor ( n52187 , n52186 , n52102 );
and ( n52188 , n52184 , n52187 );
and ( n52189 , n52132 , n52187 );
or ( n52190 , n52185 , n52188 , n52189 );
and ( n52191 , n52114 , n52190 );
xor ( n52192 , n52132 , n52184 );
xor ( n52193 , n52192 , n52187 );
buf ( n52194 , n578867 );
and ( n52195 , n52194 , n51929 );
and ( n52196 , n52144 , n51927 );
nor ( n52197 , n52195 , n52196 );
not ( n52198 , n52197 );
buf ( n52199 , n52198 );
and ( n52200 , n51965 , n52065 );
and ( n52201 , n51967 , n52063 );
nor ( n52202 , n52200 , n52201 );
xnor ( n52203 , n52202 , n52022 );
and ( n52204 , n52199 , n52203 );
and ( n52205 , n52029 , n51991 );
and ( n52206 , n52000 , n51989 );
nor ( n52207 , n52205 , n52206 );
xnor ( n52208 , n52207 , n51959 );
and ( n52209 , n52203 , n52208 );
and ( n52210 , n52199 , n52208 );
or ( n52211 , n52204 , n52209 , n52210 );
and ( n52212 , n52037 , n51991 );
and ( n52213 , n52029 , n51989 );
nor ( n52214 , n52212 , n52213 );
xnor ( n52215 , n52214 , n51959 );
and ( n52216 , n52115 , n51936 );
and ( n52217 , n52092 , n51934 );
nor ( n52218 , n52216 , n52217 );
xnor ( n52219 , n52218 , n51941 );
and ( n52220 , n52215 , n52219 );
and ( n52221 , n52219 , n52197 );
and ( n52222 , n52215 , n52197 );
or ( n52223 , n52220 , n52221 , n52222 );
and ( n52224 , n51946 , n52155 );
and ( n52225 , n51924 , n52153 );
nor ( n52226 , n52224 , n52225 );
xnor ( n52227 , n52226 , n52085 );
and ( n52228 , n52223 , n52227 );
xor ( n52229 , n52138 , n52142 );
xor ( n52230 , n52229 , n52148 );
and ( n52231 , n52227 , n52230 );
and ( n52232 , n52223 , n52230 );
or ( n52233 , n52228 , n52231 , n52232 );
and ( n52234 , n52211 , n52233 );
xor ( n52235 , n52170 , n52174 );
xor ( n52236 , n52235 , n52118 );
and ( n52237 , n52233 , n52236 );
and ( n52238 , n52211 , n52236 );
or ( n52239 , n52234 , n52237 , n52238 );
xor ( n52240 , n52120 , n52124 );
xor ( n52241 , n52240 , n52129 );
and ( n52242 , n52239 , n52241 );
xor ( n52243 , n52166 , n52178 );
xor ( n52244 , n52243 , n52181 );
and ( n52245 , n52241 , n52244 );
and ( n52246 , n52239 , n52244 );
or ( n52247 , n52242 , n52245 , n52246 );
and ( n52248 , n52193 , n52247 );
xor ( n52249 , n52239 , n52241 );
xor ( n52250 , n52249 , n52244 );
buf ( n52251 , n579160 );
buf ( n52252 , n579164 );
and ( n52253 , n52251 , n52252 );
not ( n52254 , n52253 );
and ( n52255 , n52134 , n52254 );
not ( n52256 , n52255 );
and ( n52257 , n52092 , n51991 );
and ( n52258 , n52037 , n51989 );
nor ( n52259 , n52257 , n52258 );
xnor ( n52260 , n52259 , n51959 );
and ( n52261 , n52256 , n52260 );
buf ( n52262 , n578868 );
and ( n52263 , n52262 , n51929 );
and ( n52264 , n52194 , n51927 );
nor ( n52265 , n52263 , n52264 );
not ( n52266 , n52265 );
and ( n52267 , n52260 , n52266 );
and ( n52268 , n52256 , n52266 );
or ( n52269 , n52261 , n52267 , n52268 );
xor ( n52270 , n52082 , n52133 );
xor ( n52271 , n52133 , n52134 );
not ( n52272 , n52271 );
and ( n52273 , n52270 , n52272 );
and ( n52274 , n51924 , n52273 );
not ( n52275 , n52274 );
xnor ( n52276 , n52275 , n52137 );
and ( n52277 , n52269 , n52276 );
and ( n52278 , n52000 , n52065 );
and ( n52279 , n51965 , n52063 );
nor ( n52280 , n52278 , n52279 );
xnor ( n52281 , n52280 , n52022 );
and ( n52282 , n52276 , n52281 );
and ( n52283 , n52269 , n52281 );
or ( n52284 , n52277 , n52282 , n52283 );
xor ( n52285 , n52199 , n52203 );
xor ( n52286 , n52285 , n52208 );
and ( n52287 , n52284 , n52286 );
xor ( n52288 , n52223 , n52227 );
xor ( n52289 , n52288 , n52230 );
and ( n52290 , n52286 , n52289 );
and ( n52291 , n52284 , n52289 );
or ( n52292 , n52287 , n52290 , n52291 );
xor ( n52293 , n52151 , n52158 );
xor ( n52294 , n52293 , n52163 );
and ( n52295 , n52292 , n52294 );
xor ( n52296 , n52211 , n52233 );
xor ( n52297 , n52296 , n52236 );
and ( n52298 , n52294 , n52297 );
and ( n52299 , n52292 , n52297 );
or ( n52300 , n52295 , n52298 , n52299 );
and ( n52301 , n52250 , n52300 );
xor ( n52302 , n52292 , n52294 );
xor ( n52303 , n52302 , n52297 );
buf ( n52304 , n578869 );
and ( n52305 , n52304 , n51929 );
and ( n52306 , n52262 , n51927 );
nor ( n52307 , n52305 , n52306 );
not ( n52308 , n52307 );
buf ( n52309 , n52308 );
and ( n52310 , n52029 , n52065 );
and ( n52311 , n52000 , n52063 );
nor ( n52312 , n52310 , n52311 );
xnor ( n52313 , n52312 , n52022 );
and ( n52314 , n52309 , n52313 );
and ( n52315 , n52144 , n51936 );
and ( n52316 , n52115 , n51934 );
nor ( n52317 , n52315 , n52316 );
xnor ( n52318 , n52317 , n51941 );
and ( n52319 , n52313 , n52318 );
and ( n52320 , n52309 , n52318 );
or ( n52321 , n52314 , n52319 , n52320 );
and ( n52322 , n51967 , n52155 );
and ( n52323 , n51946 , n52153 );
nor ( n52324 , n52322 , n52323 );
xnor ( n52325 , n52324 , n52085 );
and ( n52326 , n52321 , n52325 );
xor ( n52327 , n52215 , n52219 );
xor ( n52328 , n52327 , n52197 );
and ( n52329 , n52325 , n52328 );
and ( n52330 , n52321 , n52328 );
or ( n52331 , n52326 , n52329 , n52330 );
and ( n52332 , n51946 , n52273 );
and ( n52333 , n51924 , n52271 );
nor ( n52334 , n52332 , n52333 );
xnor ( n52335 , n52334 , n52137 );
and ( n52336 , n51965 , n52155 );
and ( n52337 , n51967 , n52153 );
nor ( n52338 , n52336 , n52337 );
xnor ( n52339 , n52338 , n52085 );
and ( n52340 , n52335 , n52339 );
xor ( n52341 , n52256 , n52260 );
xor ( n52342 , n52341 , n52266 );
and ( n52343 , n52339 , n52342 );
and ( n52344 , n52335 , n52342 );
or ( n52345 , n52340 , n52343 , n52344 );
xor ( n52346 , n52269 , n52276 );
xor ( n52347 , n52346 , n52281 );
and ( n52348 , n52345 , n52347 );
xor ( n52349 , n52321 , n52325 );
xor ( n52350 , n52349 , n52328 );
and ( n52351 , n52347 , n52350 );
and ( n52352 , n52345 , n52350 );
or ( n52353 , n52348 , n52351 , n52352 );
and ( n52354 , n52331 , n52353 );
xor ( n52355 , n52284 , n52286 );
xor ( n52356 , n52355 , n52289 );
and ( n52357 , n52353 , n52356 );
and ( n52358 , n52331 , n52356 );
or ( n52359 , n52354 , n52357 , n52358 );
and ( n52360 , n52303 , n52359 );
xor ( n52361 , n52331 , n52353 );
xor ( n52362 , n52361 , n52356 );
and ( n52363 , n52037 , n52065 );
and ( n52364 , n52029 , n52063 );
nor ( n52365 , n52363 , n52364 );
xnor ( n52366 , n52365 , n52022 );
and ( n52367 , n52115 , n51991 );
and ( n52368 , n52092 , n51989 );
nor ( n52369 , n52367 , n52368 );
xnor ( n52370 , n52369 , n51959 );
and ( n52371 , n52366 , n52370 );
and ( n52372 , n52194 , n51936 );
and ( n52373 , n52144 , n51934 );
nor ( n52374 , n52372 , n52373 );
xnor ( n52375 , n52374 , n51941 );
and ( n52376 , n52370 , n52375 );
and ( n52377 , n52366 , n52375 );
or ( n52378 , n52371 , n52376 , n52377 );
buf ( n52379 , n579168 );
buf ( n52380 , n579172 );
and ( n52381 , n52379 , n52380 );
not ( n52382 , n52381 );
and ( n52383 , n52252 , n52382 );
not ( n52384 , n52383 );
and ( n52385 , n52262 , n51936 );
and ( n52386 , n52194 , n51934 );
nor ( n52387 , n52385 , n52386 );
xnor ( n52388 , n52387 , n51941 );
and ( n52389 , n52384 , n52388 );
buf ( n52390 , n578870 );
and ( n52391 , n52390 , n51929 );
and ( n52392 , n52304 , n51927 );
nor ( n52393 , n52391 , n52392 );
not ( n52394 , n52393 );
and ( n52395 , n52388 , n52394 );
and ( n52396 , n52384 , n52394 );
or ( n52397 , n52389 , n52395 , n52396 );
and ( n52398 , n52000 , n52155 );
and ( n52399 , n51965 , n52153 );
nor ( n52400 , n52398 , n52399 );
xnor ( n52401 , n52400 , n52085 );
and ( n52402 , n52397 , n52401 );
and ( n52403 , n52401 , n52307 );
and ( n52404 , n52397 , n52307 );
or ( n52405 , n52402 , n52403 , n52404 );
and ( n52406 , n52378 , n52405 );
xor ( n52407 , n52309 , n52313 );
xor ( n52408 , n52407 , n52318 );
and ( n52409 , n52405 , n52408 );
and ( n52410 , n52378 , n52408 );
or ( n52411 , n52406 , n52409 , n52410 );
and ( n52412 , n52194 , n51991 );
and ( n52413 , n52144 , n51989 );
nor ( n52414 , n52412 , n52413 );
xnor ( n52415 , n52414 , n51959 );
buf ( n52416 , n52415 );
and ( n52417 , n52092 , n52065 );
and ( n52418 , n52037 , n52063 );
nor ( n52419 , n52417 , n52418 );
xnor ( n52420 , n52419 , n52022 );
and ( n52421 , n52416 , n52420 );
and ( n52422 , n52144 , n51991 );
and ( n52423 , n52115 , n51989 );
nor ( n52424 , n52422 , n52423 );
xnor ( n52425 , n52424 , n51959 );
and ( n52426 , n52420 , n52425 );
and ( n52427 , n52416 , n52425 );
or ( n52428 , n52421 , n52426 , n52427 );
xor ( n52429 , n52134 , n52251 );
xor ( n52430 , n52251 , n52252 );
not ( n52431 , n52430 );
and ( n52432 , n52429 , n52431 );
and ( n52433 , n51924 , n52432 );
not ( n52434 , n52433 );
xnor ( n52435 , n52434 , n52255 );
and ( n52436 , n52428 , n52435 );
and ( n52437 , n51967 , n52273 );
and ( n52438 , n51946 , n52271 );
nor ( n52439 , n52437 , n52438 );
xnor ( n52440 , n52439 , n52137 );
and ( n52441 , n52435 , n52440 );
and ( n52442 , n52428 , n52440 );
or ( n52443 , n52436 , n52441 , n52442 );
and ( n52444 , n51965 , n52273 );
and ( n52445 , n51967 , n52271 );
nor ( n52446 , n52444 , n52445 );
xnor ( n52447 , n52446 , n52137 );
and ( n52448 , n52029 , n52155 );
and ( n52449 , n52000 , n52153 );
nor ( n52450 , n52448 , n52449 );
xnor ( n52451 , n52450 , n52085 );
and ( n52452 , n52447 , n52451 );
xor ( n52453 , n52384 , n52388 );
xor ( n52454 , n52453 , n52394 );
and ( n52455 , n52451 , n52454 );
and ( n52456 , n52447 , n52454 );
or ( n52457 , n52452 , n52455 , n52456 );
xor ( n52458 , n52366 , n52370 );
xor ( n52459 , n52458 , n52375 );
and ( n52460 , n52457 , n52459 );
xor ( n52461 , n52397 , n52401 );
xor ( n52462 , n52461 , n52307 );
and ( n52463 , n52459 , n52462 );
and ( n52464 , n52457 , n52462 );
or ( n52465 , n52460 , n52463 , n52464 );
and ( n52466 , n52443 , n52465 );
xor ( n52467 , n52335 , n52339 );
xor ( n52468 , n52467 , n52342 );
and ( n52469 , n52465 , n52468 );
and ( n52470 , n52443 , n52468 );
or ( n52471 , n52466 , n52469 , n52470 );
and ( n52472 , n52411 , n52471 );
xor ( n52473 , n52345 , n52347 );
xor ( n52474 , n52473 , n52350 );
and ( n52475 , n52471 , n52474 );
and ( n52476 , n52411 , n52474 );
or ( n52477 , n52472 , n52475 , n52476 );
and ( n52478 , n52362 , n52477 );
and ( n52479 , n52115 , n52065 );
and ( n52480 , n52092 , n52063 );
nor ( n52481 , n52479 , n52480 );
xnor ( n52482 , n52481 , n52022 );
and ( n52483 , n52304 , n51936 );
and ( n52484 , n52262 , n51934 );
nor ( n52485 , n52483 , n52484 );
xnor ( n52486 , n52485 , n51941 );
and ( n52487 , n52482 , n52486 );
buf ( n52488 , n578871 );
and ( n52489 , n52488 , n51929 );
and ( n52490 , n52390 , n51927 );
nor ( n52491 , n52489 , n52490 );
not ( n52492 , n52491 );
and ( n52493 , n52486 , n52492 );
and ( n52494 , n52482 , n52492 );
or ( n52495 , n52487 , n52493 , n52494 );
and ( n52496 , n51946 , n52432 );
and ( n52497 , n51924 , n52430 );
nor ( n52498 , n52496 , n52497 );
xnor ( n52499 , n52498 , n52255 );
and ( n52500 , n52495 , n52499 );
xor ( n52501 , n52416 , n52420 );
xor ( n52502 , n52501 , n52425 );
and ( n52503 , n52499 , n52502 );
and ( n52504 , n52495 , n52502 );
or ( n52505 , n52500 , n52503 , n52504 );
xor ( n52506 , n52252 , n52379 );
xor ( n52507 , n52379 , n52380 );
not ( n52508 , n52507 );
and ( n52509 , n52506 , n52508 );
and ( n52510 , n51924 , n52509 );
not ( n52511 , n52510 );
xnor ( n52512 , n52511 , n52383 );
and ( n52513 , n52037 , n52155 );
and ( n52514 , n52029 , n52153 );
nor ( n52515 , n52513 , n52514 );
xnor ( n52516 , n52515 , n52085 );
and ( n52517 , n52512 , n52516 );
not ( n52518 , n52415 );
and ( n52519 , n52516 , n52518 );
and ( n52520 , n52512 , n52518 );
or ( n52521 , n52517 , n52519 , n52520 );
buf ( n52522 , n579176 );
buf ( n52523 , n579180 );
and ( n52524 , n52522 , n52523 );
not ( n52525 , n52524 );
and ( n52526 , n52380 , n52525 );
not ( n52527 , n52526 );
and ( n52528 , n52390 , n51936 );
and ( n52529 , n52304 , n51934 );
nor ( n52530 , n52528 , n52529 );
xnor ( n52531 , n52530 , n51941 );
and ( n52532 , n52527 , n52531 );
buf ( n52533 , n578872 );
and ( n52534 , n52533 , n51929 );
and ( n52535 , n52488 , n51927 );
nor ( n52536 , n52534 , n52535 );
not ( n52537 , n52536 );
and ( n52538 , n52531 , n52537 );
and ( n52539 , n52527 , n52537 );
or ( n52540 , n52532 , n52538 , n52539 );
and ( n52541 , n52000 , n52273 );
and ( n52542 , n51965 , n52271 );
nor ( n52543 , n52541 , n52542 );
xnor ( n52544 , n52543 , n52137 );
and ( n52545 , n52540 , n52544 );
xor ( n52546 , n52482 , n52486 );
xor ( n52547 , n52546 , n52492 );
and ( n52548 , n52544 , n52547 );
and ( n52549 , n52540 , n52547 );
or ( n52550 , n52545 , n52548 , n52549 );
and ( n52551 , n52521 , n52550 );
xor ( n52552 , n52447 , n52451 );
xor ( n52553 , n52552 , n52454 );
and ( n52554 , n52550 , n52553 );
and ( n52555 , n52521 , n52553 );
or ( n52556 , n52551 , n52554 , n52555 );
and ( n52557 , n52505 , n52556 );
xor ( n52558 , n52428 , n52435 );
xor ( n52559 , n52558 , n52440 );
and ( n52560 , n52556 , n52559 );
and ( n52561 , n52505 , n52559 );
or ( n52562 , n52557 , n52560 , n52561 );
xor ( n52563 , n52378 , n52405 );
xor ( n52564 , n52563 , n52408 );
and ( n52565 , n52562 , n52564 );
xor ( n52566 , n52443 , n52465 );
xor ( n52567 , n52566 , n52468 );
and ( n52568 , n52564 , n52567 );
and ( n52569 , n52562 , n52567 );
or ( n52570 , n52565 , n52568 , n52569 );
xor ( n52571 , n52411 , n52471 );
xor ( n52572 , n52571 , n52474 );
and ( n52573 , n52570 , n52572 );
xor ( n52574 , n52562 , n52564 );
xor ( n52575 , n52574 , n52567 );
and ( n52576 , n52092 , n52155 );
and ( n52577 , n52037 , n52153 );
nor ( n52578 , n52576 , n52577 );
xnor ( n52579 , n52578 , n52085 );
and ( n52580 , n52144 , n52065 );
and ( n52581 , n52115 , n52063 );
nor ( n52582 , n52580 , n52581 );
xnor ( n52583 , n52582 , n52022 );
and ( n52584 , n52579 , n52583 );
and ( n52585 , n52262 , n51991 );
and ( n52586 , n52194 , n51989 );
nor ( n52587 , n52585 , n52586 );
xnor ( n52588 , n52587 , n51959 );
and ( n52589 , n52583 , n52588 );
and ( n52590 , n52579 , n52588 );
or ( n52591 , n52584 , n52589 , n52590 );
and ( n52592 , n52194 , n52065 );
and ( n52593 , n52144 , n52063 );
nor ( n52594 , n52592 , n52593 );
xnor ( n52595 , n52594 , n52022 );
buf ( n52596 , n52595 );
and ( n52597 , n51965 , n52432 );
and ( n52598 , n51967 , n52430 );
nor ( n52599 , n52597 , n52598 );
xnor ( n52600 , n52599 , n52255 );
and ( n52601 , n52596 , n52600 );
and ( n52602 , n52029 , n52273 );
and ( n52603 , n52000 , n52271 );
nor ( n52604 , n52602 , n52603 );
xnor ( n52605 , n52604 , n52137 );
and ( n52606 , n52600 , n52605 );
and ( n52607 , n52596 , n52605 );
or ( n52608 , n52601 , n52606 , n52607 );
and ( n52609 , n52591 , n52608 );
and ( n52610 , n51967 , n52432 );
and ( n52611 , n51946 , n52430 );
nor ( n52612 , n52610 , n52611 );
xnor ( n52613 , n52612 , n52255 );
and ( n52614 , n52608 , n52613 );
and ( n52615 , n52591 , n52613 );
or ( n52616 , n52609 , n52614 , n52615 );
and ( n52617 , n52304 , n51991 );
and ( n52618 , n52262 , n51989 );
nor ( n52619 , n52617 , n52618 );
xnor ( n52620 , n52619 , n51959 );
and ( n52621 , n52488 , n51936 );
and ( n52622 , n52390 , n51934 );
nor ( n52623 , n52621 , n52622 );
xnor ( n52624 , n52623 , n51941 );
and ( n52625 , n52620 , n52624 );
buf ( n52626 , n578873 );
and ( n52627 , n52626 , n51929 );
and ( n52628 , n52533 , n51927 );
nor ( n52629 , n52627 , n52628 );
not ( n52630 , n52629 );
and ( n52631 , n52624 , n52630 );
and ( n52632 , n52620 , n52630 );
or ( n52633 , n52625 , n52631 , n52632 );
and ( n52634 , n51946 , n52509 );
and ( n52635 , n51924 , n52507 );
nor ( n52636 , n52634 , n52635 );
xnor ( n52637 , n52636 , n52383 );
and ( n52638 , n52633 , n52637 );
xor ( n52639 , n52527 , n52531 );
xor ( n52640 , n52639 , n52537 );
and ( n52641 , n52637 , n52640 );
and ( n52642 , n52633 , n52640 );
or ( n52643 , n52638 , n52641 , n52642 );
xor ( n52644 , n52512 , n52516 );
xor ( n52645 , n52644 , n52518 );
and ( n52646 , n52643 , n52645 );
xor ( n52647 , n52540 , n52544 );
xor ( n52648 , n52647 , n52547 );
and ( n52649 , n52645 , n52648 );
and ( n52650 , n52643 , n52648 );
or ( n52651 , n52646 , n52649 , n52650 );
and ( n52652 , n52616 , n52651 );
xor ( n52653 , n52495 , n52499 );
xor ( n52654 , n52653 , n52502 );
and ( n52655 , n52651 , n52654 );
and ( n52656 , n52616 , n52654 );
or ( n52657 , n52652 , n52655 , n52656 );
xor ( n52658 , n52457 , n52459 );
xor ( n52659 , n52658 , n52462 );
and ( n52660 , n52657 , n52659 );
xor ( n52661 , n52505 , n52556 );
xor ( n52662 , n52661 , n52559 );
and ( n52663 , n52659 , n52662 );
and ( n52664 , n52657 , n52662 );
or ( n52665 , n52660 , n52663 , n52664 );
and ( n52666 , n52575 , n52665 );
xor ( n52667 , n52657 , n52659 );
xor ( n52668 , n52667 , n52662 );
buf ( n52669 , n578875 );
and ( n52670 , n52669 , n51929 );
buf ( n52671 , n578874 );
and ( n52672 , n52671 , n51927 );
nor ( n52673 , n52670 , n52672 );
not ( n52674 , n52673 );
buf ( n52675 , n52674 );
buf ( n52676 , n579184 );
buf ( n52677 , n579188 );
and ( n52678 , n52676 , n52677 );
not ( n52679 , n52678 );
and ( n52680 , n52523 , n52679 );
not ( n52681 , n52680 );
and ( n52682 , n52675 , n52681 );
and ( n52683 , n52671 , n51929 );
and ( n52684 , n52626 , n51927 );
nor ( n52685 , n52683 , n52684 );
not ( n52686 , n52685 );
and ( n52687 , n52681 , n52686 );
and ( n52688 , n52675 , n52686 );
or ( n52689 , n52682 , n52687 , n52688 );
and ( n52690 , n52115 , n52155 );
and ( n52691 , n52092 , n52153 );
nor ( n52692 , n52690 , n52691 );
xnor ( n52693 , n52692 , n52085 );
and ( n52694 , n52689 , n52693 );
not ( n52695 , n52595 );
and ( n52696 , n52693 , n52695 );
and ( n580014 , n52689 , n52695 );
or ( n580015 , n52694 , n52696 , n580014 );
xor ( n580016 , n52579 , n52583 );
xor ( n52697 , n580016 , n52588 );
and ( n52698 , n580015 , n52697 );
xor ( n52699 , n52596 , n52600 );
xor ( n52700 , n52699 , n52605 );
and ( n52701 , n52697 , n52700 );
and ( n52702 , n580015 , n52700 );
or ( n52703 , n52698 , n52701 , n52702 );
xor ( n52704 , n52380 , n52522 );
xor ( n52705 , n52522 , n52523 );
not ( n52706 , n52705 );
and ( n52707 , n52704 , n52706 );
and ( n52708 , n51924 , n52707 );
not ( n52709 , n52708 );
xnor ( n52710 , n52709 , n52526 );
and ( n52711 , n52000 , n52432 );
and ( n52712 , n51965 , n52430 );
nor ( n52713 , n52711 , n52712 );
xnor ( n52714 , n52713 , n52255 );
and ( n52715 , n52710 , n52714 );
and ( n52716 , n52037 , n52273 );
and ( n52717 , n52029 , n52271 );
nor ( n52718 , n52716 , n52717 );
xnor ( n52719 , n52718 , n52137 );
and ( n52720 , n52714 , n52719 );
and ( n52721 , n52710 , n52719 );
or ( n52722 , n52715 , n52720 , n52721 );
and ( n52723 , n52262 , n52065 );
and ( n52724 , n52194 , n52063 );
nor ( n52725 , n52723 , n52724 );
xnor ( n52726 , n52725 , n52022 );
and ( n52727 , n52390 , n51991 );
and ( n52728 , n52304 , n51989 );
nor ( n52729 , n52727 , n52728 );
xnor ( n52730 , n52729 , n51959 );
and ( n52731 , n52726 , n52730 );
and ( n52732 , n52533 , n51936 );
and ( n52733 , n52488 , n51934 );
nor ( n52734 , n52732 , n52733 );
xnor ( n52735 , n52734 , n51941 );
and ( n52736 , n52730 , n52735 );
and ( n52737 , n52726 , n52735 );
or ( n52738 , n52731 , n52736 , n52737 );
and ( n52739 , n51967 , n52509 );
and ( n52740 , n51946 , n52507 );
nor ( n52741 , n52739 , n52740 );
xnor ( n52742 , n52741 , n52383 );
and ( n52743 , n52738 , n52742 );
xor ( n52744 , n52620 , n52624 );
xor ( n52745 , n52744 , n52630 );
and ( n52746 , n52742 , n52745 );
and ( n52747 , n52738 , n52745 );
or ( n52748 , n52743 , n52746 , n52747 );
and ( n52749 , n52722 , n52748 );
xor ( n52750 , n52633 , n52637 );
xor ( n52751 , n52750 , n52640 );
and ( n52752 , n52748 , n52751 );
and ( n52753 , n52722 , n52751 );
or ( n52754 , n52749 , n52752 , n52753 );
and ( n52755 , n52703 , n52754 );
xor ( n52756 , n52591 , n52608 );
xor ( n52757 , n52756 , n52613 );
and ( n52758 , n52754 , n52757 );
and ( n52759 , n52703 , n52757 );
or ( n52760 , n52755 , n52758 , n52759 );
xor ( n52761 , n52521 , n52550 );
xor ( n52762 , n52761 , n52553 );
and ( n52763 , n52760 , n52762 );
xor ( n52764 , n52616 , n52651 );
xor ( n52765 , n52764 , n52654 );
and ( n52766 , n52762 , n52765 );
and ( n52767 , n52760 , n52765 );
or ( n52768 , n52763 , n52766 , n52767 );
and ( n52769 , n52668 , n52768 );
xor ( n52770 , n52760 , n52762 );
xor ( n52771 , n52770 , n52765 );
and ( n52772 , n52488 , n51991 );
and ( n52773 , n52390 , n51989 );
nor ( n52774 , n52772 , n52773 );
xnor ( n52775 , n52774 , n51959 );
and ( n52776 , n52626 , n51936 );
and ( n52777 , n52533 , n51934 );
nor ( n52778 , n52776 , n52777 );
xnor ( n52779 , n52778 , n51941 );
and ( n52780 , n52775 , n52779 );
and ( n52781 , n52779 , n52673 );
and ( n52782 , n52775 , n52673 );
or ( n52783 , n52780 , n52781 , n52782 );
and ( n52784 , n51965 , n52509 );
and ( n52785 , n51967 , n52507 );
nor ( n52786 , n52784 , n52785 );
xnor ( n52787 , n52786 , n52383 );
and ( n52788 , n52783 , n52787 );
and ( n52789 , n52029 , n52432 );
and ( n52790 , n52000 , n52430 );
nor ( n52791 , n52789 , n52790 );
xnor ( n52792 , n52791 , n52255 );
and ( n52793 , n52787 , n52792 );
and ( n52794 , n52783 , n52792 );
or ( n52795 , n52788 , n52793 , n52794 );
and ( n52796 , n52092 , n52273 );
and ( n52797 , n52037 , n52271 );
nor ( n52798 , n52796 , n52797 );
xnor ( n52799 , n52798 , n52137 );
and ( n52800 , n52144 , n52155 );
and ( n52801 , n52115 , n52153 );
nor ( n52802 , n52800 , n52801 );
xnor ( n52803 , n52802 , n52085 );
and ( n52804 , n52799 , n52803 );
xor ( n52805 , n52675 , n52681 );
xor ( n52806 , n52805 , n52686 );
and ( n52807 , n52803 , n52806 );
and ( n52808 , n52799 , n52806 );
or ( n52809 , n52804 , n52807 , n52808 );
and ( n52810 , n52795 , n52809 );
xor ( n52811 , n52689 , n52693 );
xor ( n52812 , n52811 , n52695 );
and ( n52813 , n52809 , n52812 );
and ( n52814 , n52795 , n52812 );
or ( n52815 , n52810 , n52813 , n52814 );
buf ( n52816 , n578877 );
and ( n52817 , n52816 , n51929 );
buf ( n52818 , n578876 );
and ( n52819 , n52818 , n51927 );
nor ( n52820 , n52817 , n52819 );
not ( n52821 , n52820 );
buf ( n52822 , n52821 );
buf ( n52823 , n579192 );
buf ( n52824 , n579196 );
and ( n52825 , n52823 , n52824 );
not ( n52826 , n52825 );
and ( n52827 , n52677 , n52826 );
not ( n52828 , n52827 );
and ( n52829 , n52822 , n52828 );
and ( n52830 , n52818 , n51929 );
and ( n52831 , n52669 , n51927 );
nor ( n52832 , n52830 , n52831 );
not ( n52833 , n52832 );
and ( n52834 , n52828 , n52833 );
and ( n52835 , n52822 , n52833 );
or ( n52836 , n52829 , n52834 , n52835 );
and ( n52837 , n52194 , n52155 );
and ( n52838 , n52144 , n52153 );
nor ( n52839 , n52837 , n52838 );
xnor ( n52840 , n52839 , n52085 );
and ( n52841 , n52836 , n52840 );
and ( n52842 , n52304 , n52065 );
and ( n52843 , n52262 , n52063 );
nor ( n52844 , n52842 , n52843 );
xnor ( n52845 , n52844 , n52022 );
and ( n52846 , n52840 , n52845 );
and ( n52847 , n52836 , n52845 );
or ( n52848 , n52841 , n52846 , n52847 );
and ( n52849 , n51946 , n52707 );
and ( n52850 , n51924 , n52705 );
nor ( n52851 , n52849 , n52850 );
xnor ( n52852 , n52851 , n52526 );
and ( n52853 , n52848 , n52852 );
xor ( n52854 , n52726 , n52730 );
xor ( n52855 , n52854 , n52735 );
and ( n52856 , n52852 , n52855 );
and ( n52857 , n52848 , n52855 );
or ( n52858 , n52853 , n52856 , n52857 );
xor ( n52859 , n52710 , n52714 );
xor ( n52860 , n52859 , n52719 );
and ( n52861 , n52858 , n52860 );
xor ( n52862 , n52738 , n52742 );
xor ( n52863 , n52862 , n52745 );
and ( n52864 , n52860 , n52863 );
and ( n52865 , n52858 , n52863 );
or ( n52866 , n52861 , n52864 , n52865 );
and ( n52867 , n52815 , n52866 );
xor ( n52868 , n580015 , n52697 );
xor ( n52869 , n52868 , n52700 );
and ( n52870 , n52866 , n52869 );
and ( n52871 , n52815 , n52869 );
or ( n52872 , n52867 , n52870 , n52871 );
xor ( n52873 , n52703 , n52754 );
xor ( n52874 , n52873 , n52757 );
and ( n52875 , n52872 , n52874 );
xor ( n52876 , n52643 , n52645 );
xor ( n52877 , n52876 , n52648 );
and ( n52878 , n52874 , n52877 );
and ( n52879 , n52872 , n52877 );
or ( n52880 , n52875 , n52878 , n52879 );
and ( n52881 , n52771 , n52880 );
xor ( n52882 , n52872 , n52874 );
xor ( n52883 , n52882 , n52877 );
and ( n52884 , n52000 , n52509 );
and ( n52885 , n51965 , n52507 );
nor ( n52886 , n52884 , n52885 );
xnor ( n52887 , n52886 , n52383 );
and ( n52888 , n52037 , n52432 );
and ( n52889 , n52029 , n52430 );
nor ( n52890 , n52888 , n52889 );
xnor ( n52891 , n52890 , n52255 );
and ( n52892 , n52887 , n52891 );
and ( n52893 , n52115 , n52273 );
and ( n52894 , n52092 , n52271 );
nor ( n52895 , n52893 , n52894 );
xnor ( n52896 , n52895 , n52137 );
and ( n52897 , n52891 , n52896 );
and ( n52898 , n52887 , n52896 );
or ( n52899 , n52892 , n52897 , n52898 );
and ( n52900 , n51967 , n52707 );
and ( n52901 , n51946 , n52705 );
nor ( n52902 , n52900 , n52901 );
xnor ( n52903 , n52902 , n52526 );
xor ( n52904 , n52836 , n52840 );
xor ( n52905 , n52904 , n52845 );
and ( n52906 , n52903 , n52905 );
xor ( n52907 , n52775 , n52779 );
xor ( n52908 , n52907 , n52673 );
and ( n52909 , n52905 , n52908 );
and ( n52910 , n52903 , n52908 );
or ( n52911 , n52906 , n52909 , n52910 );
and ( n52912 , n52899 , n52911 );
xor ( n52913 , n52799 , n52803 );
xor ( n52914 , n52913 , n52806 );
and ( n52915 , n52911 , n52914 );
and ( n52916 , n52899 , n52914 );
or ( n52917 , n52912 , n52915 , n52916 );
and ( n52918 , n52390 , n52065 );
and ( n52919 , n52304 , n52063 );
nor ( n52920 , n52918 , n52919 );
xnor ( n52921 , n52920 , n52022 );
and ( n52922 , n52533 , n51991 );
and ( n52923 , n52488 , n51989 );
nor ( n52924 , n52922 , n52923 );
xnor ( n52925 , n52924 , n51959 );
and ( n52926 , n52921 , n52925 );
and ( n52927 , n52671 , n51936 );
and ( n52928 , n52626 , n51934 );
nor ( n52929 , n52927 , n52928 );
xnor ( n52930 , n52929 , n51941 );
and ( n52931 , n52925 , n52930 );
and ( n52932 , n52921 , n52930 );
or ( n52933 , n52926 , n52931 , n52932 );
buf ( n52934 , n578879 );
and ( n52935 , n52934 , n51929 );
buf ( n52936 , n578878 );
and ( n52937 , n52936 , n51927 );
nor ( n52938 , n52935 , n52937 );
not ( n52939 , n52938 );
buf ( n52940 , n52939 );
buf ( n52941 , n579200 );
buf ( n52942 , n579204 );
and ( n52943 , n52941 , n52942 );
not ( n52944 , n52943 );
and ( n52945 , n52824 , n52944 );
not ( n52946 , n52945 );
and ( n52947 , n52940 , n52946 );
and ( n52948 , n52936 , n51929 );
and ( n52949 , n52816 , n51927 );
nor ( n52950 , n52948 , n52949 );
not ( n52951 , n52950 );
and ( n52952 , n52946 , n52951 );
and ( n52953 , n52940 , n52951 );
or ( n52954 , n52947 , n52952 , n52953 );
and ( n580275 , n52669 , n51936 );
and ( n52955 , n52671 , n51934 );
nor ( n52956 , n580275 , n52955 );
xnor ( n52957 , n52956 , n51941 );
and ( n52958 , n52954 , n52957 );
and ( n52959 , n52957 , n52820 );
and ( n52960 , n52954 , n52820 );
or ( n52961 , n52958 , n52959 , n52960 );
and ( n52962 , n52144 , n52273 );
and ( n52963 , n52115 , n52271 );
nor ( n52964 , n52962 , n52963 );
xnor ( n52965 , n52964 , n52137 );
and ( n52966 , n52961 , n52965 );
and ( n52967 , n52262 , n52155 );
and ( n52968 , n52194 , n52153 );
nor ( n52969 , n52967 , n52968 );
xnor ( n52970 , n52969 , n52085 );
and ( n52971 , n52965 , n52970 );
and ( n52972 , n52961 , n52970 );
or ( n52973 , n52966 , n52971 , n52972 );
and ( n52974 , n52933 , n52973 );
xor ( n52975 , n52523 , n52676 );
xor ( n52976 , n52676 , n52677 );
not ( n52977 , n52976 );
and ( n52978 , n52975 , n52977 );
and ( n52979 , n51924 , n52978 );
not ( n52980 , n52979 );
xnor ( n52981 , n52980 , n52680 );
and ( n52982 , n52973 , n52981 );
and ( n52983 , n52933 , n52981 );
or ( n52984 , n52974 , n52982 , n52983 );
xor ( n52985 , n52783 , n52787 );
xor ( n52986 , n52985 , n52792 );
and ( n52987 , n52984 , n52986 );
xor ( n52988 , n52848 , n52852 );
xor ( n52989 , n52988 , n52855 );
and ( n52990 , n52986 , n52989 );
and ( n52991 , n52984 , n52989 );
or ( n52992 , n52987 , n52990 , n52991 );
and ( n52993 , n52917 , n52992 );
xor ( n52994 , n52795 , n52809 );
xor ( n52995 , n52994 , n52812 );
and ( n52996 , n52992 , n52995 );
and ( n52997 , n52917 , n52995 );
or ( n52998 , n52993 , n52996 , n52997 );
xor ( n52999 , n52722 , n52748 );
xor ( n53000 , n52999 , n52751 );
and ( n53001 , n52998 , n53000 );
xor ( n53002 , n52815 , n52866 );
xor ( n53003 , n53002 , n52869 );
and ( n53004 , n53000 , n53003 );
and ( n53005 , n52998 , n53003 );
or ( n53006 , n53001 , n53004 , n53005 );
and ( n53007 , n52883 , n53006 );
xor ( n53008 , n52998 , n53000 );
xor ( n53009 , n53008 , n53003 );
and ( n53010 , n52194 , n52273 );
and ( n53011 , n52144 , n52271 );
nor ( n53012 , n53010 , n53011 );
xnor ( n53013 , n53012 , n52137 );
and ( n53014 , n52488 , n52065 );
and ( n53015 , n52390 , n52063 );
nor ( n53016 , n53014 , n53015 );
xnor ( n53017 , n53016 , n52022 );
and ( n53018 , n53013 , n53017 );
and ( n53019 , n52626 , n51991 );
and ( n53020 , n52533 , n51989 );
nor ( n53021 , n53019 , n53020 );
xnor ( n53022 , n53021 , n51959 );
and ( n53023 , n53017 , n53022 );
and ( n53024 , n53013 , n53022 );
or ( n53025 , n53018 , n53023 , n53024 );
and ( n53026 , n51965 , n52707 );
and ( n53027 , n51967 , n52705 );
nor ( n53028 , n53026 , n53027 );
xnor ( n53029 , n53028 , n52526 );
and ( n53030 , n53025 , n53029 );
xor ( n53031 , n52921 , n52925 );
xor ( n53032 , n53031 , n52930 );
and ( n53033 , n53029 , n53032 );
and ( n53034 , n53025 , n53032 );
or ( n53035 , n53030 , n53033 , n53034 );
and ( n53036 , n52029 , n52509 );
and ( n53037 , n52000 , n52507 );
nor ( n53038 , n53036 , n53037 );
xnor ( n53039 , n53038 , n52383 );
and ( n53040 , n52092 , n52432 );
and ( n53041 , n52037 , n52430 );
nor ( n53042 , n53040 , n53041 );
xnor ( n53043 , n53042 , n52255 );
and ( n53044 , n53039 , n53043 );
xor ( n53045 , n52822 , n52828 );
xor ( n53046 , n53045 , n52833 );
and ( n53047 , n53043 , n53046 );
and ( n53048 , n53039 , n53046 );
or ( n53049 , n53044 , n53047 , n53048 );
and ( n53050 , n53035 , n53049 );
xor ( n53051 , n52887 , n52891 );
xor ( n53052 , n53051 , n52896 );
and ( n53053 , n53049 , n53052 );
and ( n53054 , n53035 , n53052 );
or ( n53055 , n53050 , n53053 , n53054 );
and ( n53056 , n52037 , n52509 );
and ( n53057 , n52029 , n52507 );
nor ( n53058 , n53056 , n53057 );
xnor ( n53059 , n53058 , n52383 );
and ( n53060 , n52115 , n52432 );
and ( n53061 , n52092 , n52430 );
nor ( n53062 , n53060 , n53061 );
xnor ( n53063 , n53062 , n52255 );
and ( n53064 , n53059 , n53063 );
and ( n53065 , n52304 , n52155 );
and ( n53066 , n52262 , n52153 );
nor ( n53067 , n53065 , n53066 );
xnor ( n53068 , n53067 , n52085 );
and ( n53069 , n53063 , n53068 );
and ( n53070 , n53059 , n53068 );
or ( n53071 , n53064 , n53069 , n53070 );
and ( n53072 , n51946 , n52978 );
and ( n53073 , n51924 , n52976 );
nor ( n53074 , n53072 , n53073 );
xnor ( n53075 , n53074 , n52680 );
and ( n53076 , n53071 , n53075 );
xor ( n53077 , n52961 , n52965 );
xor ( n53078 , n53077 , n52970 );
and ( n53079 , n53075 , n53078 );
and ( n53080 , n53071 , n53078 );
or ( n53081 , n53076 , n53079 , n53080 );
xor ( n53082 , n52933 , n52973 );
xor ( n53083 , n53082 , n52981 );
and ( n53084 , n53081 , n53083 );
xor ( n53085 , n52903 , n52905 );
xor ( n53086 , n53085 , n52908 );
and ( n53087 , n53083 , n53086 );
and ( n53088 , n53081 , n53086 );
or ( n53089 , n53084 , n53087 , n53088 );
and ( n53090 , n53055 , n53089 );
xor ( n53091 , n52899 , n52911 );
xor ( n53092 , n53091 , n52914 );
and ( n53093 , n53089 , n53092 );
and ( n53094 , n53055 , n53092 );
or ( n53095 , n53090 , n53093 , n53094 );
xor ( n53096 , n52858 , n52860 );
xor ( n53097 , n53096 , n52863 );
and ( n53098 , n53095 , n53097 );
xor ( n53099 , n52917 , n52992 );
xor ( n53100 , n53099 , n52995 );
and ( n53101 , n53097 , n53100 );
and ( n53102 , n53095 , n53100 );
or ( n53103 , n53098 , n53101 , n53102 );
and ( n53104 , n53009 , n53103 );
xor ( n53105 , n53095 , n53097 );
xor ( n53106 , n53105 , n53100 );
buf ( n53107 , n578881 );
and ( n53108 , n53107 , n51929 );
buf ( n53109 , n578880 );
and ( n53110 , n53109 , n51927 );
nor ( n53111 , n53108 , n53110 );
not ( n53112 , n53111 );
buf ( n53113 , n53112 );
buf ( n53114 , n579208 );
buf ( n53115 , n579212 );
and ( n53116 , n53114 , n53115 );
not ( n53117 , n53116 );
and ( n53118 , n52942 , n53117 );
not ( n53119 , n53118 );
and ( n53120 , n53113 , n53119 );
and ( n53121 , n53109 , n51929 );
and ( n53122 , n52934 , n51927 );
nor ( n53123 , n53121 , n53122 );
not ( n53124 , n53123 );
and ( n53125 , n53119 , n53124 );
and ( n53126 , n53113 , n53124 );
or ( n53127 , n53120 , n53125 , n53126 );
and ( n53128 , n52816 , n51936 );
and ( n53129 , n52818 , n51934 );
nor ( n53130 , n53128 , n53129 );
xnor ( n53131 , n53130 , n51941 );
and ( n53132 , n53127 , n53131 );
and ( n53133 , n53131 , n52938 );
and ( n53134 , n53127 , n52938 );
or ( n53135 , n53132 , n53133 , n53134 );
and ( n53136 , n52262 , n52273 );
and ( n53137 , n52194 , n52271 );
nor ( n53138 , n53136 , n53137 );
xnor ( n53139 , n53138 , n52137 );
and ( n53140 , n53135 , n53139 );
and ( n53141 , n52533 , n52065 );
and ( n53142 , n52488 , n52063 );
nor ( n53143 , n53141 , n53142 );
xnor ( n53144 , n53143 , n52022 );
and ( n53145 , n53139 , n53144 );
and ( n53146 , n53135 , n53144 );
or ( n53147 , n53140 , n53145 , n53146 );
and ( n53148 , n51967 , n52978 );
and ( n53149 , n51946 , n52976 );
nor ( n53150 , n53148 , n53149 );
xnor ( n53151 , n53150 , n52680 );
and ( n53152 , n53147 , n53151 );
and ( n53153 , n52000 , n52707 );
and ( n53154 , n51965 , n52705 );
nor ( n53155 , n53153 , n53154 );
xnor ( n53156 , n53155 , n52526 );
and ( n53157 , n53151 , n53156 );
and ( n53158 , n53147 , n53156 );
or ( n53159 , n53152 , n53157 , n53158 );
and ( n53160 , n52671 , n51991 );
and ( n53161 , n52626 , n51989 );
nor ( n53162 , n53160 , n53161 );
xnor ( n53163 , n53162 , n51959 );
and ( n53164 , n52818 , n51936 );
and ( n53165 , n52669 , n51934 );
nor ( n53166 , n53164 , n53165 );
xnor ( n53167 , n53166 , n51941 );
and ( n53168 , n53163 , n53167 );
xor ( n53169 , n52940 , n52946 );
xor ( n53170 , n53169 , n52951 );
and ( n53171 , n53167 , n53170 );
and ( n53172 , n53163 , n53170 );
or ( n53173 , n53168 , n53171 , n53172 );
xor ( n53174 , n52677 , n52823 );
xor ( n53175 , n52823 , n52824 );
not ( n53176 , n53175 );
and ( n53177 , n53174 , n53176 );
and ( n53178 , n51924 , n53177 );
not ( n53179 , n53178 );
xnor ( n53180 , n53179 , n52827 );
and ( n53181 , n53173 , n53180 );
xor ( n53182 , n52954 , n52957 );
xor ( n53183 , n53182 , n52820 );
and ( n53184 , n53180 , n53183 );
and ( n53185 , n53173 , n53183 );
or ( n53186 , n53181 , n53184 , n53185 );
and ( n53187 , n53159 , n53186 );
xor ( n53188 , n53039 , n53043 );
xor ( n53189 , n53188 , n53046 );
and ( n53190 , n53186 , n53189 );
and ( n53191 , n53159 , n53189 );
or ( n53192 , n53187 , n53190 , n53191 );
xor ( n53193 , n53035 , n53049 );
xor ( n53194 , n53193 , n53052 );
and ( n53195 , n53192 , n53194 );
xor ( n53196 , n53081 , n53083 );
xor ( n53197 , n53196 , n53086 );
and ( n53198 , n53194 , n53197 );
and ( n53199 , n53192 , n53197 );
or ( n53200 , n53195 , n53198 , n53199 );
xor ( n53201 , n52984 , n52986 );
xor ( n53202 , n53201 , n52989 );
and ( n53203 , n53200 , n53202 );
xor ( n53204 , n53055 , n53089 );
xor ( n53205 , n53204 , n53092 );
and ( n53206 , n53202 , n53205 );
and ( n53207 , n53200 , n53205 );
or ( n53208 , n53203 , n53206 , n53207 );
and ( n53209 , n53106 , n53208 );
xor ( n53210 , n53200 , n53202 );
xor ( n53211 , n53210 , n53205 );
and ( n53212 , n52092 , n52509 );
and ( n53213 , n52037 , n52507 );
nor ( n53214 , n53212 , n53213 );
xnor ( n53215 , n53214 , n52383 );
and ( n53216 , n52144 , n52432 );
and ( n53217 , n52115 , n52430 );
nor ( n53218 , n53216 , n53217 );
xnor ( n53219 , n53218 , n52255 );
and ( n53220 , n53215 , n53219 );
and ( n53221 , n52390 , n52155 );
and ( n53222 , n52304 , n52153 );
nor ( n53223 , n53221 , n53222 );
xnor ( n53224 , n53223 , n52085 );
and ( n53225 , n53219 , n53224 );
and ( n53226 , n53215 , n53224 );
or ( n53227 , n53220 , n53225 , n53226 );
xor ( n53228 , n53013 , n53017 );
xor ( n53229 , n53228 , n53022 );
and ( n53230 , n53227 , n53229 );
xor ( n53231 , n53059 , n53063 );
xor ( n53232 , n53231 , n53068 );
and ( n53233 , n53229 , n53232 );
and ( n53234 , n53227 , n53232 );
or ( n53235 , n53230 , n53233 , n53234 );
xor ( n53236 , n53025 , n53029 );
xor ( n53237 , n53236 , n53032 );
and ( n53238 , n53235 , n53237 );
xor ( n53239 , n53071 , n53075 );
xor ( n53240 , n53239 , n53078 );
and ( n53241 , n53237 , n53240 );
and ( n53242 , n53235 , n53240 );
or ( n53243 , n53238 , n53241 , n53242 );
and ( n53244 , n52037 , n52707 );
and ( n53245 , n52029 , n52705 );
nor ( n53246 , n53244 , n53245 );
xnor ( n53247 , n53246 , n52526 );
and ( n53248 , n52115 , n52509 );
and ( n53249 , n52092 , n52507 );
nor ( n53250 , n53248 , n53249 );
xnor ( n53251 , n53250 , n52383 );
and ( n53252 , n53247 , n53251 );
and ( n53253 , n52626 , n52065 );
and ( n53254 , n52533 , n52063 );
nor ( n53255 , n53253 , n53254 );
xnor ( n53256 , n53255 , n52022 );
and ( n53257 , n53251 , n53256 );
and ( n53258 , n53247 , n53256 );
or ( n53259 , n53252 , n53257 , n53258 );
xor ( n53260 , n53215 , n53219 );
xor ( n53261 , n53260 , n53224 );
and ( n53262 , n53259 , n53261 );
xor ( n53263 , n53135 , n53139 );
xor ( n53264 , n53263 , n53144 );
and ( n53265 , n53261 , n53264 );
and ( n53266 , n53259 , n53264 );
or ( n53267 , n53262 , n53265 , n53266 );
xor ( n53268 , n53147 , n53151 );
xor ( n53269 , n53268 , n53156 );
and ( n53270 , n53267 , n53269 );
xor ( n53271 , n53227 , n53229 );
xor ( n53272 , n53271 , n53232 );
and ( n53273 , n53269 , n53272 );
and ( n53274 , n53267 , n53272 );
or ( n53275 , n53270 , n53273 , n53274 );
and ( n53276 , n52304 , n52273 );
and ( n53277 , n52262 , n52271 );
nor ( n53278 , n53276 , n53277 );
xnor ( n53279 , n53278 , n52137 );
and ( n53280 , n52488 , n52155 );
and ( n580602 , n52390 , n52153 );
nor ( n53281 , n53280 , n580602 );
xnor ( n53282 , n53281 , n52085 );
and ( n53283 , n53279 , n53282 );
xor ( n53284 , n53127 , n53131 );
xor ( n53285 , n53284 , n52938 );
and ( n53286 , n53282 , n53285 );
and ( n53287 , n53279 , n53285 );
or ( n53288 , n53283 , n53286 , n53287 );
and ( n53289 , n51946 , n53177 );
and ( n53290 , n51924 , n53175 );
nor ( n53291 , n53289 , n53290 );
xnor ( n53292 , n53291 , n52827 );
and ( n53293 , n53288 , n53292 );
and ( n53294 , n51965 , n52978 );
and ( n53295 , n51967 , n52976 );
nor ( n53296 , n53294 , n53295 );
xnor ( n53297 , n53296 , n52680 );
and ( n53298 , n53292 , n53297 );
and ( n53299 , n53288 , n53297 );
or ( n53300 , n53293 , n53298 , n53299 );
and ( n53301 , n52818 , n51991 );
and ( n53302 , n52669 , n51989 );
nor ( n53303 , n53301 , n53302 );
xnor ( n53304 , n53303 , n51959 );
and ( n53305 , n52936 , n51936 );
and ( n53306 , n52816 , n51934 );
nor ( n53307 , n53305 , n53306 );
xnor ( n53308 , n53307 , n51941 );
and ( n53309 , n53304 , n53308 );
xor ( n53310 , n53113 , n53119 );
xor ( n53311 , n53310 , n53124 );
and ( n53312 , n53308 , n53311 );
and ( n53313 , n53304 , n53311 );
or ( n53314 , n53309 , n53312 , n53313 );
and ( n53315 , n52194 , n52432 );
and ( n53316 , n52144 , n52430 );
nor ( n53317 , n53315 , n53316 );
xnor ( n53318 , n53317 , n52255 );
and ( n53319 , n53314 , n53318 );
and ( n53320 , n52669 , n51991 );
and ( n53321 , n52671 , n51989 );
nor ( n53322 , n53320 , n53321 );
xnor ( n53323 , n53322 , n51959 );
and ( n53324 , n53318 , n53323 );
and ( n53325 , n53314 , n53323 );
or ( n53326 , n53319 , n53324 , n53325 );
and ( n53327 , n52029 , n52707 );
and ( n53328 , n52000 , n52705 );
nor ( n53329 , n53327 , n53328 );
xnor ( n53330 , n53329 , n52526 );
and ( n53331 , n53326 , n53330 );
xor ( n53332 , n53163 , n53167 );
xor ( n53333 , n53332 , n53170 );
and ( n53334 , n53330 , n53333 );
and ( n53335 , n53326 , n53333 );
or ( n53336 , n53331 , n53334 , n53335 );
and ( n53337 , n53300 , n53336 );
xor ( n53338 , n53173 , n53180 );
xor ( n53339 , n53338 , n53183 );
and ( n53340 , n53336 , n53339 );
and ( n53341 , n53300 , n53339 );
or ( n53342 , n53337 , n53340 , n53341 );
and ( n53343 , n53275 , n53342 );
xor ( n53344 , n53159 , n53186 );
xor ( n53345 , n53344 , n53189 );
and ( n53346 , n53342 , n53345 );
and ( n53347 , n53275 , n53345 );
or ( n53348 , n53343 , n53346 , n53347 );
and ( n53349 , n53243 , n53348 );
xor ( n53350 , n53192 , n53194 );
xor ( n53351 , n53350 , n53197 );
and ( n53352 , n53348 , n53351 );
and ( n53353 , n53243 , n53351 );
or ( n53354 , n53349 , n53352 , n53353 );
and ( n53355 , n53211 , n53354 );
and ( n53356 , n52669 , n52065 );
and ( n53357 , n52671 , n52063 );
nor ( n53358 , n53356 , n53357 );
xnor ( n53359 , n53358 , n52022 );
and ( n53360 , n52816 , n51991 );
and ( n53361 , n52818 , n51989 );
nor ( n53362 , n53360 , n53361 );
xnor ( n53363 , n53362 , n51959 );
and ( n53364 , n53359 , n53363 );
buf ( n53365 , n578883 );
and ( n53366 , n53365 , n51929 );
buf ( n53367 , n578882 );
and ( n53368 , n53367 , n51927 );
nor ( n53369 , n53366 , n53368 );
not ( n53370 , n53369 );
buf ( n53371 , n53370 );
buf ( n53372 , n579216 );
buf ( n53373 , n579220 );
and ( n53374 , n53372 , n53373 );
not ( n53375 , n53374 );
and ( n53376 , n53115 , n53375 );
not ( n53377 , n53376 );
and ( n53378 , n53371 , n53377 );
and ( n53379 , n53109 , n51936 );
and ( n53380 , n52934 , n51934 );
nor ( n53381 , n53379 , n53380 );
xnor ( n53382 , n53381 , n51941 );
and ( n53383 , n53377 , n53382 );
and ( n53384 , n53371 , n53382 );
or ( n53385 , n53378 , n53383 , n53384 );
and ( n53386 , n52934 , n51936 );
and ( n53387 , n52936 , n51934 );
nor ( n53388 , n53386 , n53387 );
xnor ( n53389 , n53388 , n51941 );
xor ( n53390 , n53385 , n53389 );
xor ( n53391 , n53390 , n53111 );
and ( n53392 , n53363 , n53391 );
and ( n53393 , n53359 , n53391 );
or ( n53394 , n53364 , n53392 , n53393 );
and ( n53395 , n52092 , n52707 );
and ( n53396 , n52037 , n52705 );
nor ( n53397 , n53395 , n53396 );
xnor ( n53398 , n53397 , n52526 );
and ( n53399 , n53394 , n53398 );
and ( n53400 , n52144 , n52509 );
and ( n53401 , n52115 , n52507 );
nor ( n53402 , n53400 , n53401 );
xnor ( n53403 , n53402 , n52383 );
and ( n53404 , n53398 , n53403 );
and ( n53405 , n53394 , n53403 );
or ( n53406 , n53399 , n53404 , n53405 );
and ( n53407 , n51967 , n53177 );
and ( n53408 , n51946 , n53175 );
nor ( n53409 , n53407 , n53408 );
xnor ( n53410 , n53409 , n52827 );
and ( n53411 , n53406 , n53410 );
and ( n53412 , n52000 , n52978 );
and ( n580735 , n51965 , n52976 );
nor ( n53413 , n53412 , n580735 );
xnor ( n53414 , n53413 , n52680 );
and ( n53415 , n53410 , n53414 );
and ( n53416 , n53406 , n53414 );
or ( n53417 , n53411 , n53415 , n53416 );
xor ( n53418 , n53247 , n53251 );
xor ( n53419 , n53418 , n53256 );
xor ( n53420 , n53314 , n53318 );
xor ( n53421 , n53420 , n53323 );
and ( n53422 , n53419 , n53421 );
xor ( n53423 , n53279 , n53282 );
xor ( n53424 , n53423 , n53285 );
and ( n53425 , n53421 , n53424 );
and ( n53426 , n53419 , n53424 );
or ( n53427 , n53422 , n53425 , n53426 );
and ( n53428 , n53417 , n53427 );
xor ( n53429 , n53259 , n53261 );
xor ( n53430 , n53429 , n53264 );
and ( n53431 , n53427 , n53430 );
and ( n53432 , n53417 , n53430 );
or ( n53433 , n53428 , n53431 , n53432 );
and ( n53434 , n53385 , n53389 );
and ( n53435 , n53389 , n53111 );
and ( n53436 , n53385 , n53111 );
or ( n53437 , n53434 , n53435 , n53436 );
and ( n53438 , n52262 , n52432 );
and ( n53439 , n52194 , n52430 );
nor ( n53440 , n53438 , n53439 );
xnor ( n53441 , n53440 , n52255 );
and ( n53442 , n53437 , n53441 );
and ( n53443 , n52671 , n52065 );
and ( n53444 , n52626 , n52063 );
nor ( n53445 , n53443 , n53444 );
xnor ( n53446 , n53445 , n52022 );
and ( n53447 , n53441 , n53446 );
and ( n53448 , n53437 , n53446 );
or ( n53449 , n53442 , n53447 , n53448 );
and ( n53450 , n52390 , n52273 );
and ( n53451 , n52304 , n52271 );
nor ( n53452 , n53450 , n53451 );
xnor ( n53453 , n53452 , n52137 );
and ( n53454 , n52533 , n52155 );
and ( n53455 , n52488 , n52153 );
nor ( n53456 , n53454 , n53455 );
xnor ( n53457 , n53456 , n52085 );
and ( n53458 , n53453 , n53457 );
xor ( n53459 , n53304 , n53308 );
xor ( n53460 , n53459 , n53311 );
and ( n53461 , n53457 , n53460 );
and ( n53462 , n53453 , n53460 );
or ( n53463 , n53458 , n53461 , n53462 );
and ( n53464 , n53449 , n53463 );
xor ( n53465 , n52824 , n52941 );
xor ( n53466 , n52941 , n52942 );
not ( n53467 , n53466 );
and ( n53468 , n53465 , n53467 );
and ( n53469 , n51924 , n53468 );
not ( n53470 , n53469 );
xnor ( n53471 , n53470 , n52945 );
and ( n53472 , n53463 , n53471 );
and ( n53473 , n53449 , n53471 );
or ( n53474 , n53464 , n53472 , n53473 );
xor ( n53475 , n53288 , n53292 );
xor ( n53476 , n53475 , n53297 );
and ( n53477 , n53474 , n53476 );
xor ( n53478 , n53326 , n53330 );
xor ( n53479 , n53478 , n53333 );
and ( n53480 , n53476 , n53479 );
and ( n53481 , n53474 , n53479 );
or ( n53482 , n53477 , n53480 , n53481 );
and ( n53483 , n53433 , n53482 );
xor ( n53484 , n53300 , n53336 );
xor ( n53485 , n53484 , n53339 );
and ( n53486 , n53482 , n53485 );
and ( n53487 , n53433 , n53485 );
or ( n53488 , n53483 , n53486 , n53487 );
xor ( n53489 , n53235 , n53237 );
xor ( n53490 , n53489 , n53240 );
and ( n53491 , n53488 , n53490 );
xor ( n53492 , n53275 , n53342 );
xor ( n53493 , n53492 , n53345 );
and ( n53494 , n53490 , n53493 );
and ( n53495 , n53488 , n53493 );
or ( n53496 , n53491 , n53494 , n53495 );
xor ( n53497 , n53243 , n53348 );
xor ( n53498 , n53497 , n53351 );
and ( n53499 , n53496 , n53498 );
and ( n53500 , n52934 , n51991 );
and ( n53501 , n52936 , n51989 );
nor ( n53502 , n53500 , n53501 );
xnor ( n53503 , n53502 , n51959 );
and ( n53504 , n53107 , n51936 );
and ( n53505 , n53109 , n51934 );
nor ( n53506 , n53504 , n53505 );
xnor ( n53507 , n53506 , n51941 );
and ( n53508 , n53503 , n53507 );
and ( n53509 , n53507 , n53369 );
and ( n53510 , n53503 , n53369 );
or ( n53511 , n53508 , n53509 , n53510 );
and ( n53512 , n52936 , n51991 );
and ( n53513 , n52816 , n51989 );
nor ( n53514 , n53512 , n53513 );
xnor ( n53515 , n53514 , n51959 );
and ( n53516 , n53511 , n53515 );
and ( n53517 , n53367 , n51929 );
and ( n53518 , n53107 , n51927 );
nor ( n53519 , n53517 , n53518 );
not ( n53520 , n53519 );
and ( n53521 , n53515 , n53520 );
and ( n53522 , n53511 , n53520 );
or ( n53523 , n53516 , n53521 , n53522 );
and ( n53524 , n52304 , n52432 );
and ( n53525 , n52262 , n52430 );
nor ( n53526 , n53524 , n53525 );
xnor ( n53527 , n53526 , n52255 );
and ( n53528 , n53523 , n53527 );
and ( n53529 , n52488 , n52273 );
and ( n53530 , n52390 , n52271 );
nor ( n53531 , n53529 , n53530 );
xnor ( n53532 , n53531 , n52137 );
and ( n53533 , n53527 , n53532 );
and ( n53534 , n53523 , n53532 );
or ( n53535 , n53528 , n53533 , n53534 );
and ( n53536 , n52194 , n52509 );
and ( n53537 , n52144 , n52507 );
nor ( n53538 , n53536 , n53537 );
xnor ( n53539 , n53538 , n52383 );
and ( n53540 , n52626 , n52155 );
and ( n53541 , n52533 , n52153 );
nor ( n53542 , n53540 , n53541 );
xnor ( n53543 , n53542 , n52085 );
and ( n53544 , n53539 , n53543 );
xor ( n53545 , n53359 , n53363 );
xor ( n53546 , n53545 , n53391 );
and ( n53547 , n53543 , n53546 );
and ( n53548 , n53539 , n53546 );
or ( n53549 , n53544 , n53547 , n53548 );
and ( n53550 , n53535 , n53549 );
and ( n53551 , n51946 , n53468 );
and ( n53552 , n51924 , n53466 );
nor ( n53553 , n53551 , n53552 );
xnor ( n53554 , n53553 , n52945 );
and ( n53555 , n53549 , n53554 );
and ( n53556 , n53535 , n53554 );
or ( n53557 , n53550 , n53555 , n53556 );
and ( n53558 , n51965 , n53177 );
and ( n53559 , n51967 , n53175 );
nor ( n53560 , n53558 , n53559 );
xnor ( n53561 , n53560 , n52827 );
and ( n53562 , n52029 , n52978 );
and ( n53563 , n52000 , n52976 );
nor ( n53564 , n53562 , n53563 );
xnor ( n53565 , n53564 , n52680 );
and ( n53566 , n53561 , n53565 );
xor ( n53567 , n53437 , n53441 );
xor ( n53568 , n53567 , n53446 );
and ( n53569 , n53565 , n53568 );
and ( n53570 , n53561 , n53568 );
or ( n53571 , n53566 , n53569 , n53570 );
and ( n53572 , n53557 , n53571 );
xor ( n53573 , n53449 , n53463 );
xor ( n53574 , n53573 , n53471 );
and ( n53575 , n53571 , n53574 );
and ( n53576 , n53557 , n53574 );
or ( n53577 , n53572 , n53575 , n53576 );
and ( n53578 , n52671 , n52155 );
and ( n53579 , n52626 , n52153 );
nor ( n53580 , n53578 , n53579 );
xnor ( n53581 , n53580 , n52085 );
and ( n53582 , n52818 , n52065 );
and ( n53583 , n52669 , n52063 );
nor ( n53584 , n53582 , n53583 );
xnor ( n53585 , n53584 , n52022 );
and ( n53586 , n53581 , n53585 );
xor ( n53587 , n53371 , n53377 );
xor ( n53588 , n53587 , n53382 );
and ( n53589 , n53585 , n53588 );
and ( n53590 , n53581 , n53588 );
or ( n53591 , n53586 , n53589 , n53590 );
and ( n53592 , n52037 , n52978 );
and ( n53593 , n52029 , n52976 );
nor ( n53594 , n53592 , n53593 );
xnor ( n53595 , n53594 , n52680 );
and ( n53596 , n53591 , n53595 );
and ( n53597 , n52115 , n52707 );
and ( n53598 , n52092 , n52705 );
nor ( n53599 , n53597 , n53598 );
xnor ( n53600 , n53599 , n52526 );
and ( n53601 , n53595 , n53600 );
and ( n53602 , n53591 , n53600 );
or ( n53603 , n53596 , n53601 , n53602 );
xor ( n53604 , n53394 , n53398 );
xor ( n53605 , n53604 , n53403 );
and ( n53606 , n53603 , n53605 );
xor ( n53607 , n53453 , n53457 );
xor ( n53608 , n53607 , n53460 );
and ( n53609 , n53605 , n53608 );
and ( n53610 , n53603 , n53608 );
or ( n53611 , n53606 , n53609 , n53610 );
xor ( n53612 , n53406 , n53410 );
xor ( n53613 , n53612 , n53414 );
and ( n53614 , n53611 , n53613 );
xor ( n53615 , n53419 , n53421 );
xor ( n53616 , n53615 , n53424 );
and ( n53617 , n53613 , n53616 );
and ( n53618 , n53611 , n53616 );
or ( n53619 , n53614 , n53617 , n53618 );
and ( n53620 , n53577 , n53619 );
xor ( n53621 , n53474 , n53476 );
xor ( n53622 , n53621 , n53479 );
and ( n53623 , n53619 , n53622 );
and ( n53624 , n53577 , n53622 );
or ( n53625 , n53620 , n53623 , n53624 );
xor ( n53626 , n53267 , n53269 );
xor ( n53627 , n53626 , n53272 );
and ( n53628 , n53625 , n53627 );
xor ( n53629 , n53433 , n53482 );
xor ( n53630 , n53629 , n53485 );
and ( n53631 , n53627 , n53630 );
and ( n53632 , n53625 , n53630 );
or ( n53633 , n53628 , n53631 , n53632 );
xor ( n53634 , n53488 , n53490 );
xor ( n53635 , n53634 , n53493 );
and ( n53636 , n53633 , n53635 );
xor ( n53637 , n53625 , n53627 );
xor ( n53638 , n53637 , n53630 );
buf ( n53639 , n578885 );
and ( n53640 , n53639 , n51929 );
buf ( n53641 , n578884 );
and ( n53642 , n53641 , n51927 );
nor ( n53643 , n53640 , n53642 );
not ( n53644 , n53643 );
buf ( n53645 , n53644 );
buf ( n53646 , n579224 );
buf ( n53647 , n579228 );
and ( n53648 , n53646 , n53647 );
not ( n53649 , n53648 );
and ( n53650 , n53373 , n53649 );
not ( n53651 , n53650 );
and ( n53652 , n53645 , n53651 );
and ( n53653 , n53641 , n51929 );
and ( n53654 , n53365 , n51927 );
nor ( n53655 , n53653 , n53654 );
not ( n53656 , n53655 );
and ( n53657 , n53651 , n53656 );
and ( n53658 , n53645 , n53656 );
or ( n53659 , n53652 , n53657 , n53658 );
and ( n53660 , n52816 , n52065 );
and ( n53661 , n52818 , n52063 );
nor ( n53662 , n53660 , n53661 );
xnor ( n53663 , n53662 , n52022 );
and ( n53664 , n53659 , n53663 );
xor ( n53665 , n53503 , n53507 );
xor ( n53666 , n53665 , n53369 );
and ( n53667 , n53663 , n53666 );
and ( n53668 , n53659 , n53666 );
or ( n53669 , n53664 , n53667 , n53668 );
and ( n53670 , n52390 , n52432 );
and ( n53671 , n52304 , n52430 );
nor ( n53672 , n53670 , n53671 );
xnor ( n53673 , n53672 , n52255 );
and ( n53674 , n53669 , n53673 );
xor ( n53675 , n53511 , n53515 );
xor ( n53676 , n53675 , n53520 );
and ( n53677 , n53673 , n53676 );
and ( n53678 , n53669 , n53676 );
or ( n53679 , n53674 , n53677 , n53678 );
xor ( n53680 , n52942 , n53114 );
xor ( n53681 , n53114 , n53115 );
not ( n53682 , n53681 );
and ( n53683 , n53680 , n53682 );
and ( n53684 , n51924 , n53683 );
not ( n53685 , n53684 );
xnor ( n53686 , n53685 , n53118 );
and ( n53687 , n53679 , n53686 );
and ( n53688 , n52000 , n53177 );
and ( n53689 , n51965 , n53175 );
nor ( n53690 , n53688 , n53689 );
xnor ( n53691 , n53690 , n52827 );
and ( n53692 , n53686 , n53691 );
and ( n53693 , n53679 , n53691 );
or ( n53694 , n53687 , n53692 , n53693 );
and ( n53695 , n52092 , n52978 );
and ( n53696 , n52037 , n52976 );
nor ( n53697 , n53695 , n53696 );
xnor ( n53698 , n53697 , n52680 );
and ( n53699 , n52262 , n52509 );
and ( n53700 , n52194 , n52507 );
nor ( n53701 , n53699 , n53700 );
xnor ( n53702 , n53701 , n52383 );
and ( n53703 , n53698 , n53702 );
and ( n53704 , n52533 , n52273 );
and ( n53705 , n52488 , n52271 );
nor ( n53706 , n53704 , n53705 );
xnor ( n53707 , n53706 , n52137 );
and ( n53708 , n53702 , n53707 );
and ( n53709 , n53698 , n53707 );
or ( n53710 , n53703 , n53708 , n53709 );
and ( n53711 , n51967 , n53468 );
and ( n53712 , n51946 , n53466 );
nor ( n53713 , n53711 , n53712 );
xnor ( n53714 , n53713 , n52945 );
and ( n53715 , n53710 , n53714 );
xor ( n53716 , n53523 , n53527 );
xor ( n53717 , n53716 , n53532 );
and ( n53718 , n53714 , n53717 );
and ( n53719 , n53710 , n53717 );
or ( n53720 , n53715 , n53718 , n53719 );
and ( n53721 , n53694 , n53720 );
xor ( n53722 , n53561 , n53565 );
xor ( n53723 , n53722 , n53568 );
and ( n53724 , n53720 , n53723 );
and ( n53725 , n53694 , n53723 );
or ( n53726 , n53721 , n53724 , n53725 );
xor ( n53727 , n53557 , n53571 );
xor ( n53728 , n53727 , n53574 );
and ( n53729 , n53726 , n53728 );
xor ( n53730 , n53611 , n53613 );
xor ( n53731 , n53730 , n53616 );
and ( n53732 , n53728 , n53731 );
and ( n53733 , n53726 , n53731 );
or ( n53734 , n53729 , n53732 , n53733 );
xor ( n53735 , n53417 , n53427 );
xor ( n53736 , n53735 , n53430 );
and ( n53737 , n53734 , n53736 );
xor ( n53738 , n53577 , n53619 );
xor ( n53739 , n53738 , n53622 );
and ( n53740 , n53736 , n53739 );
and ( n53741 , n53734 , n53739 );
or ( n53742 , n53737 , n53740 , n53741 );
and ( n53743 , n53638 , n53742 );
xor ( n53744 , n53734 , n53736 );
xor ( n53745 , n53744 , n53739 );
and ( n53746 , n52194 , n52707 );
and ( n53747 , n52144 , n52705 );
nor ( n53748 , n53746 , n53747 );
xnor ( n53749 , n53748 , n52526 );
and ( n53750 , n52304 , n52509 );
and ( n53751 , n52262 , n52507 );
nor ( n53752 , n53750 , n53751 );
xnor ( n53753 , n53752 , n52383 );
and ( n53754 , n53749 , n53753 );
and ( n53755 , n52626 , n52273 );
and ( n53756 , n52533 , n52271 );
nor ( n53757 , n53755 , n53756 );
xnor ( n53758 , n53757 , n52137 );
and ( n53759 , n53753 , n53758 );
and ( n53760 , n53749 , n53758 );
or ( n53761 , n53754 , n53759 , n53760 );
buf ( n53762 , n579236 );
not ( n53763 , n53762 );
buf ( n53764 , n53763 );
buf ( n53765 , n53764 );
buf ( n53766 , n579232 );
and ( n53767 , n53766 , n53762 );
not ( n53768 , n53767 );
and ( n53769 , n53647 , n53768 );
not ( n53770 , n53769 );
and ( n53771 , n53765 , n53770 );
and ( n53772 , n53641 , n51936 );
and ( n53773 , n53365 , n51934 );
nor ( n53774 , n53772 , n53773 );
xnor ( n53775 , n53774 , n51941 );
and ( n53776 , n53770 , n53775 );
and ( n53777 , n53765 , n53775 );
or ( n53778 , n53771 , n53776 , n53777 );
and ( n53779 , n53365 , n51936 );
and ( n53780 , n53367 , n51934 );
nor ( n53781 , n53779 , n53780 );
xnor ( n53782 , n53781 , n51941 );
and ( n53783 , n53778 , n53782 );
and ( n53784 , n53782 , n53643 );
and ( n53785 , n53778 , n53643 );
or ( n53786 , n53783 , n53784 , n53785 );
and ( n53787 , n52818 , n52155 );
and ( n53788 , n52669 , n52153 );
nor ( n53789 , n53787 , n53788 );
xnor ( n53790 , n53789 , n52085 );
and ( n53791 , n53786 , n53790 );
and ( n53792 , n52936 , n52065 );
and ( n53793 , n52816 , n52063 );
nor ( n53794 , n53792 , n53793 );
xnor ( n53795 , n53794 , n52022 );
and ( n53796 , n53790 , n53795 );
and ( n53797 , n53786 , n53795 );
or ( n53798 , n53791 , n53796 , n53797 );
and ( n53799 , n53109 , n51991 );
and ( n53800 , n52934 , n51989 );
nor ( n53801 , n53799 , n53800 );
xnor ( n53802 , n53801 , n51959 );
and ( n53803 , n53367 , n51936 );
and ( n53804 , n53107 , n51934 );
nor ( n53805 , n53803 , n53804 );
xnor ( n53806 , n53805 , n51941 );
and ( n53807 , n53802 , n53806 );
xor ( n53808 , n53645 , n53651 );
xor ( n53809 , n53808 , n53656 );
and ( n53810 , n53806 , n53809 );
and ( n53811 , n53802 , n53809 );
or ( n53812 , n53807 , n53810 , n53811 );
and ( n53813 , n53798 , n53812 );
and ( n53814 , n52669 , n52155 );
and ( n53815 , n52671 , n52153 );
nor ( n53816 , n53814 , n53815 );
xnor ( n53817 , n53816 , n52085 );
and ( n53818 , n53812 , n53817 );
and ( n53819 , n53798 , n53817 );
or ( n53820 , n53813 , n53818 , n53819 );
and ( n53821 , n53761 , n53820 );
and ( n53822 , n51965 , n53468 );
and ( n53823 , n51967 , n53466 );
nor ( n53824 , n53822 , n53823 );
xnor ( n53825 , n53824 , n52945 );
and ( n53826 , n53820 , n53825 );
and ( n53827 , n53761 , n53825 );
or ( n53828 , n53821 , n53826 , n53827 );
not ( n53829 , n53764 );
and ( n53830 , n53639 , n51936 );
and ( n53831 , n53641 , n51934 );
nor ( n53832 , n53830 , n53831 );
xnor ( n53833 , n53832 , n51941 );
and ( n53834 , n53829 , n53833 );
buf ( n53835 , n578887 );
and ( n53836 , n53835 , n51929 );
buf ( n53837 , n578886 );
and ( n53838 , n53837 , n51927 );
nor ( n53839 , n53836 , n53838 );
not ( n53840 , n53839 );
and ( n53841 , n53833 , n53840 );
and ( n53842 , n53829 , n53840 );
or ( n53843 , n53834 , n53841 , n53842 );
and ( n53844 , n53367 , n51991 );
and ( n53845 , n53107 , n51989 );
nor ( n53846 , n53844 , n53845 );
xnor ( n53847 , n53846 , n51959 );
and ( n53848 , n53843 , n53847 );
and ( n53849 , n53837 , n51929 );
and ( n53850 , n53639 , n51927 );
nor ( n53851 , n53849 , n53850 );
not ( n53852 , n53851 );
and ( n53853 , n53847 , n53852 );
and ( n53854 , n53843 , n53852 );
or ( n53855 , n53848 , n53853 , n53854 );
and ( n53856 , n52934 , n52065 );
and ( n53857 , n52936 , n52063 );
nor ( n53858 , n53856 , n53857 );
xnor ( n53859 , n53858 , n52022 );
and ( n53860 , n53855 , n53859 );
and ( n53861 , n53107 , n51991 );
and ( n53862 , n53109 , n51989 );
nor ( n53863 , n53861 , n53862 );
xnor ( n53864 , n53863 , n51959 );
and ( n53865 , n53859 , n53864 );
and ( n53866 , n53855 , n53864 );
or ( n53867 , n53860 , n53865 , n53866 );
and ( n53868 , n52671 , n52273 );
and ( n53869 , n52626 , n52271 );
nor ( n53870 , n53868 , n53869 );
xnor ( n53871 , n53870 , n52137 );
and ( n53872 , n53867 , n53871 );
xor ( n53873 , n53802 , n53806 );
xor ( n53874 , n53873 , n53809 );
and ( n53875 , n53871 , n53874 );
and ( n53876 , n53867 , n53874 );
or ( n53877 , n53872 , n53875 , n53876 );
and ( n53878 , n52488 , n52432 );
and ( n53879 , n52390 , n52430 );
nor ( n53880 , n53878 , n53879 );
xnor ( n53881 , n53880 , n52255 );
and ( n53882 , n53877 , n53881 );
xor ( n53883 , n53659 , n53663 );
xor ( n53884 , n53883 , n53666 );
and ( n53885 , n53881 , n53884 );
and ( n53886 , n53877 , n53884 );
or ( n53887 , n53882 , n53885 , n53886 );
xor ( n53888 , n53698 , n53702 );
xor ( n53889 , n53888 , n53707 );
and ( n53890 , n53887 , n53889 );
xor ( n53891 , n53669 , n53673 );
xor ( n53892 , n53891 , n53676 );
and ( n53893 , n53889 , n53892 );
and ( n53894 , n53887 , n53892 );
or ( n53895 , n53890 , n53893 , n53894 );
and ( n53896 , n53828 , n53895 );
xor ( n53897 , n53679 , n53686 );
xor ( n53898 , n53897 , n53691 );
and ( n53899 , n53895 , n53898 );
and ( n53900 , n53828 , n53898 );
or ( n53901 , n53896 , n53899 , n53900 );
and ( n53902 , n52037 , n53177 );
and ( n53903 , n52029 , n53175 );
nor ( n53904 , n53902 , n53903 );
xnor ( n53905 , n53904 , n52827 );
and ( n53906 , n52115 , n52978 );
and ( n53907 , n52092 , n52976 );
nor ( n53908 , n53906 , n53907 );
xnor ( n53909 , n53908 , n52680 );
and ( n53910 , n53905 , n53909 );
xor ( n53911 , n53798 , n53812 );
xor ( n53912 , n53911 , n53817 );
and ( n53913 , n53909 , n53912 );
and ( n53914 , n53905 , n53912 );
or ( n53915 , n53910 , n53913 , n53914 );
and ( n53916 , n51946 , n53683 );
and ( n53917 , n51924 , n53681 );
nor ( n53918 , n53916 , n53917 );
xnor ( n53919 , n53918 , n53118 );
and ( n53920 , n53915 , n53919 );
and ( n53921 , n52029 , n53177 );
and ( n53922 , n52000 , n53175 );
nor ( n53923 , n53921 , n53922 );
xnor ( n53924 , n53923 , n52827 );
and ( n53925 , n52144 , n52707 );
and ( n53926 , n52115 , n52705 );
nor ( n53927 , n53925 , n53926 );
xnor ( n53928 , n53927 , n52526 );
xor ( n53929 , n53924 , n53928 );
xor ( n53930 , n53581 , n53585 );
xor ( n53931 , n53930 , n53588 );
xor ( n53932 , n53929 , n53931 );
and ( n53933 , n53919 , n53932 );
and ( n53934 , n53915 , n53932 );
or ( n53935 , n53920 , n53933 , n53934 );
xor ( n53936 , n53710 , n53714 );
xor ( n53937 , n53936 , n53717 );
and ( n53938 , n53935 , n53937 );
and ( n53939 , n53924 , n53928 );
and ( n53940 , n53928 , n53931 );
and ( n53941 , n53924 , n53931 );
or ( n53942 , n53939 , n53940 , n53941 );
xor ( n53943 , n53591 , n53595 );
xor ( n53944 , n53943 , n53600 );
xor ( n53945 , n53942 , n53944 );
xor ( n53946 , n53539 , n53543 );
xor ( n53947 , n53946 , n53546 );
xor ( n53948 , n53945 , n53947 );
and ( n53949 , n53937 , n53948 );
and ( n53950 , n53935 , n53948 );
or ( n53951 , n53938 , n53949 , n53950 );
and ( n53952 , n53901 , n53951 );
xor ( n53953 , n53694 , n53720 );
xor ( n53954 , n53953 , n53723 );
and ( n53955 , n53951 , n53954 );
and ( n53956 , n53901 , n53954 );
or ( n53957 , n53952 , n53955 , n53956 );
and ( n53958 , n53942 , n53944 );
and ( n53959 , n53944 , n53947 );
and ( n53960 , n53942 , n53947 );
or ( n53961 , n53958 , n53959 , n53960 );
xor ( n53962 , n53535 , n53549 );
xor ( n53963 , n53962 , n53554 );
and ( n53964 , n53961 , n53963 );
xor ( n53965 , n53603 , n53605 );
xor ( n53966 , n53965 , n53608 );
and ( n53967 , n53963 , n53966 );
and ( n53968 , n53961 , n53966 );
or ( n53969 , n53964 , n53967 , n53968 );
and ( n53970 , n53957 , n53969 );
xor ( n53971 , n53726 , n53728 );
xor ( n53972 , n53971 , n53731 );
and ( n53973 , n53969 , n53972 );
and ( n53974 , n53957 , n53972 );
or ( n53975 , n53970 , n53973 , n53974 );
and ( n53976 , n53745 , n53975 );
xor ( n53977 , n53957 , n53969 );
xor ( n53978 , n53977 , n53972 );
and ( n53979 , n52262 , n52707 );
and ( n53980 , n52194 , n52705 );
nor ( n53981 , n53979 , n53980 );
xnor ( n53982 , n53981 , n52526 );
and ( n53983 , n52533 , n52432 );
and ( n53984 , n52488 , n52430 );
nor ( n53985 , n53983 , n53984 );
xnor ( n53986 , n53985 , n52255 );
and ( n53987 , n53982 , n53986 );
xor ( n53988 , n53786 , n53790 );
xor ( n53989 , n53988 , n53795 );
and ( n53990 , n53986 , n53989 );
and ( n53991 , n53982 , n53989 );
or ( n53992 , n53987 , n53990 , n53991 );
xor ( n53993 , n53115 , n53372 );
xor ( n53994 , n53372 , n53373 );
not ( n53995 , n53994 );
and ( n53996 , n53993 , n53995 );
and ( n53997 , n51924 , n53996 );
not ( n53998 , n53997 );
xnor ( n53999 , n53998 , n53376 );
and ( n54000 , n53992 , n53999 );
and ( n54001 , n52000 , n53468 );
and ( n54002 , n51965 , n53466 );
nor ( n54003 , n54001 , n54002 );
xnor ( n54004 , n54003 , n52945 );
and ( n54005 , n53999 , n54004 );
and ( n54006 , n53992 , n54004 );
or ( n54007 , n54000 , n54005 , n54006 );
and ( n54008 , n52669 , n52273 );
and ( n54009 , n52671 , n52271 );
nor ( n54010 , n54008 , n54009 );
xnor ( n54011 , n54010 , n52137 );
and ( n54012 , n52816 , n52155 );
and ( n54013 , n52818 , n52153 );
nor ( n54014 , n54012 , n54013 );
xnor ( n54015 , n54014 , n52085 );
and ( n54016 , n54011 , n54015 );
xor ( n54017 , n53778 , n53782 );
xor ( n54018 , n54017 , n53643 );
and ( n54019 , n54015 , n54018 );
and ( n54020 , n54011 , n54018 );
or ( n54021 , n54016 , n54019 , n54020 );
and ( n54022 , n52144 , n52978 );
and ( n54023 , n52115 , n52976 );
nor ( n54024 , n54022 , n54023 );
xnor ( n54025 , n54024 , n52680 );
and ( n54026 , n54021 , n54025 );
and ( n54027 , n52390 , n52509 );
and ( n54028 , n52304 , n52507 );
nor ( n54029 , n54027 , n54028 );
xnor ( n54030 , n54029 , n52383 );
and ( n54031 , n54025 , n54030 );
and ( n54032 , n54021 , n54030 );
or ( n54033 , n54026 , n54031 , n54032 );
and ( n54034 , n51967 , n53683 );
and ( n54035 , n51946 , n53681 );
nor ( n54036 , n54034 , n54035 );
xnor ( n54037 , n54036 , n53118 );
and ( n54038 , n54033 , n54037 );
xor ( n54039 , n53877 , n53881 );
xor ( n54040 , n54039 , n53884 );
and ( n54041 , n54037 , n54040 );
and ( n54042 , n54033 , n54040 );
or ( n54043 , n54038 , n54041 , n54042 );
and ( n54044 , n54007 , n54043 );
xor ( n54045 , n53761 , n53820 );
xor ( n54046 , n54045 , n53825 );
and ( n54047 , n54043 , n54046 );
and ( n54048 , n54007 , n54046 );
or ( n54049 , n54044 , n54047 , n54048 );
and ( n54050 , n53837 , n51936 );
and ( n54051 , n53639 , n51934 );
nor ( n54052 , n54050 , n54051 );
xnor ( n54053 , n54052 , n51941 );
and ( n54054 , n53762 , n54053 );
buf ( n54055 , n578888 );
and ( n54056 , n54055 , n51929 );
and ( n54057 , n53835 , n51927 );
nor ( n54058 , n54056 , n54057 );
not ( n54059 , n54058 );
and ( n54060 , n54053 , n54059 );
and ( n54061 , n53762 , n54059 );
or ( n54062 , n54054 , n54060 , n54061 );
and ( n54063 , n53107 , n52065 );
and ( n54064 , n53109 , n52063 );
nor ( n54065 , n54063 , n54064 );
xnor ( n54066 , n54065 , n52022 );
and ( n54067 , n54062 , n54066 );
and ( n54068 , n53365 , n51991 );
and ( n54069 , n53367 , n51989 );
nor ( n54070 , n54068 , n54069 );
xnor ( n54071 , n54070 , n51959 );
and ( n54072 , n54066 , n54071 );
and ( n54073 , n54062 , n54071 );
or ( n54074 , n54067 , n54072 , n54073 );
and ( n54075 , n53109 , n52065 );
and ( n54076 , n52934 , n52063 );
nor ( n54077 , n54075 , n54076 );
xnor ( n54078 , n54077 , n52022 );
and ( n54079 , n54074 , n54078 );
xor ( n54080 , n53765 , n53770 );
xor ( n54081 , n54080 , n53775 );
and ( n54082 , n54078 , n54081 );
and ( n54083 , n54074 , n54081 );
or ( n54084 , n54079 , n54082 , n54083 );
and ( n54085 , n52818 , n52273 );
and ( n54086 , n52669 , n52271 );
nor ( n54087 , n54085 , n54086 );
xnor ( n54088 , n54087 , n52137 );
and ( n54089 , n52936 , n52155 );
and ( n54090 , n52816 , n52153 );
nor ( n54091 , n54089 , n54090 );
xnor ( n54092 , n54091 , n52085 );
and ( n54093 , n54088 , n54092 );
xor ( n54094 , n53843 , n53847 );
xor ( n54095 , n54094 , n53852 );
and ( n54096 , n54092 , n54095 );
and ( n54097 , n54088 , n54095 );
or ( n54098 , n54093 , n54096 , n54097 );
and ( n54099 , n54084 , n54098 );
xor ( n54100 , n53855 , n53859 );
xor ( n54101 , n54100 , n53864 );
and ( n54102 , n54098 , n54101 );
and ( n54103 , n54084 , n54101 );
or ( n54104 , n54099 , n54102 , n54103 );
and ( n54105 , n52029 , n53468 );
and ( n54106 , n52000 , n53466 );
nor ( n54107 , n54105 , n54106 );
xnor ( n54108 , n54107 , n52945 );
and ( n54109 , n54104 , n54108 );
and ( n54110 , n52092 , n53177 );
and ( n54111 , n52037 , n53175 );
nor ( n54112 , n54110 , n54111 );
xnor ( n54113 , n54112 , n52827 );
and ( n54114 , n54108 , n54113 );
and ( n54115 , n54104 , n54113 );
or ( n54116 , n54109 , n54114 , n54115 );
xor ( n54117 , n53749 , n53753 );
xor ( n54118 , n54117 , n53758 );
and ( n54119 , n54116 , n54118 );
xor ( n54120 , n53905 , n53909 );
xor ( n54121 , n54120 , n53912 );
and ( n54122 , n54118 , n54121 );
and ( n54123 , n54116 , n54121 );
or ( n54124 , n54119 , n54122 , n54123 );
xor ( n54125 , n53887 , n53889 );
xor ( n54126 , n54125 , n53892 );
and ( n54127 , n54124 , n54126 );
xor ( n54128 , n53915 , n53919 );
xor ( n54129 , n54128 , n53932 );
and ( n54130 , n54126 , n54129 );
and ( n54131 , n54124 , n54129 );
or ( n54132 , n54127 , n54130 , n54131 );
and ( n54133 , n54049 , n54132 );
xor ( n54134 , n53828 , n53895 );
xor ( n54135 , n54134 , n53898 );
and ( n54136 , n54132 , n54135 );
and ( n54137 , n54049 , n54135 );
or ( n54138 , n54133 , n54136 , n54137 );
xor ( n54139 , n53901 , n53951 );
xor ( n54140 , n54139 , n53954 );
and ( n54141 , n54138 , n54140 );
xor ( n54142 , n53961 , n53963 );
xor ( n54143 , n54142 , n53966 );
and ( n54144 , n54140 , n54143 );
and ( n54145 , n54138 , n54143 );
or ( n54146 , n54141 , n54144 , n54145 );
and ( n54147 , n53978 , n54146 );
xor ( n54148 , n54138 , n54140 );
xor ( n54149 , n54148 , n54143 );
and ( n54150 , n52115 , n53177 );
and ( n54151 , n52092 , n53175 );
nor ( n54152 , n54150 , n54151 );
xnor ( n54153 , n54152 , n52827 );
and ( n54154 , n52626 , n52432 );
and ( n54155 , n52533 , n52430 );
nor ( n54156 , n54154 , n54155 );
xnor ( n54157 , n54156 , n52255 );
and ( n54158 , n54153 , n54157 );
xor ( n54159 , n54011 , n54015 );
xor ( n54160 , n54159 , n54018 );
and ( n54161 , n54157 , n54160 );
and ( n54162 , n54153 , n54160 );
or ( n54163 , n54158 , n54161 , n54162 );
and ( n54164 , n51946 , n53996 );
and ( n54165 , n51924 , n53994 );
nor ( n54166 , n54164 , n54165 );
xnor ( n54167 , n54166 , n53376 );
and ( n54168 , n54163 , n54167 );
xor ( n54169 , n54021 , n54025 );
xor ( n54170 , n54169 , n54030 );
and ( n54171 , n54167 , n54170 );
and ( n54172 , n54163 , n54170 );
or ( n54173 , n54168 , n54171 , n54172 );
and ( n54174 , n52194 , n52978 );
and ( n54175 , n52144 , n52976 );
nor ( n54176 , n54174 , n54175 );
xnor ( n54177 , n54176 , n52680 );
and ( n54178 , n52304 , n52707 );
and ( n54179 , n52262 , n52705 );
nor ( n54180 , n54178 , n54179 );
xnor ( n54181 , n54180 , n52526 );
and ( n54182 , n54177 , n54181 );
and ( n54183 , n52488 , n52509 );
and ( n54184 , n52390 , n52507 );
nor ( n54185 , n54183 , n54184 );
xnor ( n54186 , n54185 , n52383 );
and ( n54187 , n54181 , n54186 );
and ( n54188 , n54177 , n54186 );
or ( n54189 , n54182 , n54187 , n54188 );
and ( n54190 , n51965 , n53683 );
and ( n54191 , n51967 , n53681 );
nor ( n54192 , n54190 , n54191 );
xnor ( n54193 , n54192 , n53118 );
and ( n54194 , n54189 , n54193 );
xor ( n54195 , n53867 , n53871 );
xor ( n54196 , n54195 , n53874 );
and ( n54197 , n54193 , n54196 );
and ( n54198 , n54189 , n54196 );
or ( n54199 , n54194 , n54197 , n54198 );
and ( n54200 , n54173 , n54199 );
xor ( n54201 , n53992 , n53999 );
xor ( n54202 , n54201 , n54004 );
and ( n54203 , n54199 , n54202 );
and ( n54204 , n54173 , n54202 );
or ( n54205 , n54200 , n54203 , n54204 );
and ( n54206 , n53639 , n51991 );
and ( n54207 , n53641 , n51989 );
nor ( n54208 , n54206 , n54207 );
xnor ( n54209 , n54208 , n51959 );
and ( n54210 , n53835 , n51936 );
and ( n54211 , n53837 , n51934 );
nor ( n54212 , n54210 , n54211 );
xnor ( n54213 , n54212 , n51941 );
and ( n54214 , n54209 , n54213 );
buf ( n54215 , n578889 );
and ( n54216 , n54215 , n51929 );
and ( n54217 , n54055 , n51927 );
nor ( n54218 , n54216 , n54217 );
not ( n54219 , n54218 );
and ( n54220 , n54213 , n54219 );
and ( n54221 , n54209 , n54219 );
or ( n54222 , n54214 , n54220 , n54221 );
and ( n54223 , n53367 , n52065 );
and ( n54224 , n53107 , n52063 );
nor ( n54225 , n54223 , n54224 );
xnor ( n54226 , n54225 , n52022 );
and ( n54227 , n54222 , n54226 );
and ( n54228 , n53641 , n51991 );
and ( n54229 , n53365 , n51989 );
nor ( n54230 , n54228 , n54229 );
xnor ( n54231 , n54230 , n51959 );
and ( n54232 , n54226 , n54231 );
and ( n54233 , n54222 , n54231 );
or ( n54234 , n54227 , n54232 , n54233 );
and ( n54235 , n52934 , n52155 );
and ( n54236 , n52936 , n52153 );
nor ( n54237 , n54235 , n54236 );
xnor ( n54238 , n54237 , n52085 );
and ( n54239 , n54234 , n54238 );
xor ( n54240 , n53829 , n53833 );
xor ( n54241 , n54240 , n53840 );
and ( n54242 , n54238 , n54241 );
and ( n54243 , n54234 , n54241 );
or ( n54244 , n54239 , n54242 , n54243 );
and ( n54245 , n52671 , n52432 );
and ( n54246 , n52626 , n52430 );
nor ( n54247 , n54245 , n54246 );
xnor ( n54248 , n54247 , n52255 );
and ( n54249 , n54244 , n54248 );
xor ( n54250 , n54074 , n54078 );
xor ( n54251 , n54250 , n54081 );
and ( n54252 , n54248 , n54251 );
and ( n54253 , n54244 , n54251 );
or ( n54254 , n54249 , n54252 , n54253 );
and ( n54255 , n52037 , n53468 );
and ( n54256 , n52029 , n53466 );
nor ( n54257 , n54255 , n54256 );
xnor ( n54258 , n54257 , n52945 );
and ( n54259 , n54254 , n54258 );
xor ( n54260 , n54084 , n54098 );
xor ( n54261 , n54260 , n54101 );
and ( n54262 , n54258 , n54261 );
and ( n54263 , n54254 , n54261 );
or ( n54264 , n54259 , n54262 , n54263 );
xor ( n54265 , n54104 , n54108 );
xor ( n54266 , n54265 , n54113 );
and ( n54267 , n54264 , n54266 );
xor ( n54268 , n53982 , n53986 );
xor ( n54269 , n54268 , n53989 );
and ( n54270 , n54266 , n54269 );
and ( n54271 , n54264 , n54269 );
or ( n54272 , n54267 , n54270 , n54271 );
xor ( n54273 , n54116 , n54118 );
xor ( n54274 , n54273 , n54121 );
and ( n54275 , n54272 , n54274 );
xor ( n54276 , n54033 , n54037 );
xor ( n54277 , n54276 , n54040 );
and ( n54278 , n54274 , n54277 );
and ( n54279 , n54272 , n54277 );
or ( n54280 , n54275 , n54278 , n54279 );
and ( n54281 , n54205 , n54280 );
xor ( n54282 , n54007 , n54043 );
xor ( n54283 , n54282 , n54046 );
and ( n54284 , n54280 , n54283 );
and ( n54285 , n54205 , n54283 );
or ( n54286 , n54281 , n54284 , n54285 );
xor ( n54287 , n54049 , n54132 );
xor ( n54288 , n54287 , n54135 );
and ( n54289 , n54286 , n54288 );
xor ( n54290 , n53935 , n53937 );
xor ( n54291 , n54290 , n53948 );
and ( n54292 , n54288 , n54291 );
and ( n54293 , n54286 , n54291 );
or ( n54294 , n54289 , n54292 , n54293 );
and ( n54295 , n54149 , n54294 );
xor ( n54296 , n54286 , n54288 );
xor ( n54297 , n54296 , n54291 );
and ( n54298 , n52936 , n52273 );
and ( n54299 , n52816 , n52271 );
nor ( n54300 , n54298 , n54299 );
xnor ( n54301 , n54300 , n52137 );
and ( n54302 , n53109 , n52155 );
and ( n54303 , n52934 , n52153 );
nor ( n54304 , n54302 , n54303 );
xnor ( n54305 , n54304 , n52085 );
and ( n54306 , n54301 , n54305 );
xor ( n54307 , n53762 , n54053 );
xor ( n54308 , n54307 , n54059 );
and ( n54309 , n54305 , n54308 );
and ( n54310 , n54301 , n54308 );
or ( n54311 , n54306 , n54309 , n54310 );
and ( n54312 , n53641 , n52065 );
and ( n54313 , n53365 , n52063 );
nor ( n54314 , n54312 , n54313 );
xnor ( n54315 , n54314 , n52022 );
and ( n54316 , n54055 , n51936 );
and ( n54317 , n53835 , n51934 );
nor ( n54318 , n54316 , n54317 );
xnor ( n54319 , n54318 , n51941 );
and ( n54320 , n54315 , n54319 );
buf ( n54321 , n578890 );
and ( n54322 , n54321 , n51929 );
and ( n54323 , n54215 , n51927 );
nor ( n54324 , n54322 , n54323 );
not ( n54325 , n54324 );
and ( n54326 , n54319 , n54325 );
and ( n54327 , n54315 , n54325 );
or ( n54328 , n54320 , n54326 , n54327 );
and ( n54329 , n53107 , n52155 );
and ( n54330 , n53109 , n52153 );
nor ( n54331 , n54329 , n54330 );
xnor ( n54332 , n54331 , n52085 );
and ( n54333 , n54328 , n54332 );
and ( n54334 , n53365 , n52065 );
and ( n54335 , n53367 , n52063 );
nor ( n54336 , n54334 , n54335 );
xnor ( n54337 , n54336 , n52022 );
and ( n54338 , n54332 , n54337 );
and ( n54339 , n54328 , n54337 );
or ( n54340 , n54333 , n54338 , n54339 );
and ( n54341 , n52818 , n52432 );
and ( n54342 , n52669 , n52430 );
nor ( n54343 , n54341 , n54342 );
xnor ( n54344 , n54343 , n52255 );
and ( n54345 , n54340 , n54344 );
xor ( n54346 , n54222 , n54226 );
xor ( n54347 , n54346 , n54231 );
and ( n54348 , n54344 , n54347 );
and ( n54349 , n54340 , n54347 );
or ( n54350 , n54345 , n54348 , n54349 );
and ( n54351 , n54311 , n54350 );
xor ( n54352 , n54234 , n54238 );
xor ( n54353 , n54352 , n54241 );
and ( n54354 , n54350 , n54353 );
and ( n54355 , n54311 , n54353 );
or ( n54356 , n54351 , n54354 , n54355 );
and ( n54357 , n52029 , n53683 );
and ( n54358 , n52000 , n53681 );
nor ( n54359 , n54357 , n54358 );
xnor ( n54360 , n54359 , n53118 );
and ( n54361 , n54356 , n54360 );
and ( n54362 , n52144 , n53177 );
and ( n54363 , n52115 , n53175 );
nor ( n54364 , n54362 , n54363 );
xnor ( n54365 , n54364 , n52827 );
and ( n54366 , n54360 , n54365 );
and ( n54367 , n54356 , n54365 );
or ( n54368 , n54361 , n54366 , n54367 );
xor ( n54369 , n54177 , n54181 );
xor ( n54370 , n54369 , n54186 );
and ( n54371 , n54368 , n54370 );
xor ( n54372 , n54254 , n54258 );
xor ( n54373 , n54372 , n54261 );
and ( n54374 , n54370 , n54373 );
and ( n54375 , n54368 , n54373 );
or ( n54376 , n54371 , n54374 , n54375 );
xor ( n54377 , n54163 , n54167 );
xor ( n54378 , n54377 , n54170 );
and ( n54379 , n54376 , n54378 );
xor ( n54380 , n54264 , n54266 );
xor ( n54381 , n54380 , n54269 );
and ( n54382 , n54378 , n54381 );
and ( n54383 , n54376 , n54381 );
or ( n54384 , n54379 , n54382 , n54383 );
and ( n54385 , n52669 , n52432 );
and ( n54386 , n52671 , n52430 );
nor ( n54387 , n54385 , n54386 );
xnor ( n54388 , n54387 , n52255 );
and ( n54389 , n52816 , n52273 );
and ( n54390 , n52818 , n52271 );
nor ( n54391 , n54389 , n54390 );
xnor ( n54392 , n54391 , n52137 );
and ( n54393 , n54388 , n54392 );
xor ( n54394 , n54062 , n54066 );
xor ( n54395 , n54394 , n54071 );
and ( n54396 , n54392 , n54395 );
and ( n54397 , n54388 , n54395 );
or ( n54398 , n54393 , n54396 , n54397 );
and ( n54399 , n52262 , n52978 );
and ( n54400 , n52194 , n52976 );
nor ( n54401 , n54399 , n54400 );
xnor ( n54402 , n54401 , n52680 );
and ( n54403 , n54398 , n54402 );
and ( n54404 , n52533 , n52509 );
and ( n54405 , n52488 , n52507 );
nor ( n54406 , n54404 , n54405 );
xnor ( n54407 , n54406 , n52383 );
and ( n54408 , n54402 , n54407 );
and ( n54409 , n54398 , n54407 );
or ( n54410 , n54403 , n54408 , n54409 );
xor ( n54411 , n53373 , n53646 );
xor ( n54412 , n53646 , n53647 );
not ( n54413 , n54412 );
and ( n54414 , n54411 , n54413 );
and ( n54415 , n51924 , n54414 );
not ( n54416 , n54415 );
xnor ( n54417 , n54416 , n53650 );
and ( n54418 , n54410 , n54417 );
and ( n54419 , n52000 , n53683 );
and ( n54420 , n51965 , n53681 );
nor ( n54421 , n54419 , n54420 );
xnor ( n54422 , n54421 , n53118 );
and ( n54423 , n54417 , n54422 );
and ( n54424 , n54410 , n54422 );
or ( n54425 , n54418 , n54423 , n54424 );
and ( n54426 , n52092 , n53468 );
and ( n54427 , n52037 , n53466 );
nor ( n54428 , n54426 , n54427 );
xnor ( n54429 , n54428 , n52945 );
and ( n54430 , n52390 , n52707 );
and ( n54431 , n52304 , n52705 );
nor ( n54432 , n54430 , n54431 );
xnor ( n54433 , n54432 , n52526 );
and ( n54434 , n54429 , n54433 );
xor ( n54435 , n54088 , n54092 );
xor ( n54436 , n54435 , n54095 );
and ( n54437 , n54433 , n54436 );
and ( n54438 , n54429 , n54436 );
or ( n54439 , n54434 , n54437 , n54438 );
and ( n54440 , n51967 , n53996 );
and ( n54441 , n51946 , n53994 );
nor ( n54442 , n54440 , n54441 );
xnor ( n54443 , n54442 , n53376 );
and ( n54444 , n54439 , n54443 );
xor ( n54445 , n54153 , n54157 );
xor ( n54446 , n54445 , n54160 );
and ( n54447 , n54443 , n54446 );
and ( n54448 , n54439 , n54446 );
or ( n54449 , n54444 , n54447 , n54448 );
and ( n54450 , n54425 , n54449 );
xor ( n54451 , n54189 , n54193 );
xor ( n54452 , n54451 , n54196 );
and ( n54453 , n54449 , n54452 );
and ( n54454 , n54425 , n54452 );
or ( n54455 , n54450 , n54453 , n54454 );
and ( n54456 , n54384 , n54455 );
xor ( n54457 , n54173 , n54199 );
xor ( n54458 , n54457 , n54202 );
and ( n54459 , n54455 , n54458 );
and ( n54460 , n54384 , n54458 );
or ( n54461 , n54456 , n54459 , n54460 );
xor ( n54462 , n54205 , n54280 );
xor ( n54463 , n54462 , n54283 );
and ( n54464 , n54461 , n54463 );
xor ( n54465 , n54124 , n54126 );
xor ( n54466 , n54465 , n54129 );
and ( n54467 , n54463 , n54466 );
and ( n54468 , n54461 , n54466 );
or ( n54469 , n54464 , n54467 , n54468 );
and ( n54470 , n54297 , n54469 );
and ( n54471 , n52194 , n53177 );
and ( n54472 , n52144 , n53175 );
nor ( n54473 , n54471 , n54472 );
xnor ( n54474 , n54473 , n52827 );
and ( n54475 , n52304 , n52978 );
and ( n54476 , n52262 , n52976 );
nor ( n54477 , n54475 , n54476 );
xnor ( n54478 , n54477 , n52680 );
and ( n54479 , n54474 , n54478 );
xor ( n54480 , n54388 , n54392 );
xor ( n54481 , n54480 , n54395 );
and ( n54482 , n54478 , n54481 );
and ( n54483 , n54474 , n54481 );
or ( n54484 , n54479 , n54482 , n54483 );
and ( n54485 , n51965 , n53996 );
and ( n54486 , n51967 , n53994 );
nor ( n54487 , n54485 , n54486 );
xnor ( n54488 , n54487 , n53376 );
and ( n54489 , n54484 , n54488 );
xor ( n54490 , n54244 , n54248 );
xor ( n54491 , n54490 , n54251 );
and ( n54492 , n54488 , n54491 );
and ( n54493 , n54484 , n54491 );
or ( n54494 , n54489 , n54492 , n54493 );
and ( n54495 , n51946 , n54414 );
and ( n54496 , n51924 , n54412 );
nor ( n54497 , n54495 , n54496 );
xnor ( n54498 , n54497 , n53650 );
xor ( n54499 , n54398 , n54402 );
xor ( n54500 , n54499 , n54407 );
and ( n54501 , n54498 , n54500 );
xor ( n54502 , n54429 , n54433 );
xor ( n54503 , n54502 , n54436 );
and ( n54504 , n54500 , n54503 );
and ( n54505 , n54498 , n54503 );
or ( n54506 , n54501 , n54504 , n54505 );
and ( n54507 , n54494 , n54506 );
xor ( n54508 , n54410 , n54417 );
xor ( n54509 , n54508 , n54422 );
and ( n54510 , n54506 , n54509 );
and ( n54511 , n54494 , n54509 );
or ( n54512 , n54507 , n54510 , n54511 );
and ( n54513 , n52262 , n53177 );
and ( n54514 , n52194 , n53175 );
nor ( n54515 , n54513 , n54514 );
xnor ( n54516 , n54515 , n52827 );
and ( n54517 , n52390 , n52978 );
and ( n54518 , n52304 , n52976 );
nor ( n54519 , n54517 , n54518 );
xnor ( n54520 , n54519 , n52680 );
and ( n54521 , n54516 , n54520 );
and ( n54522 , n52533 , n52707 );
and ( n54523 , n52488 , n52705 );
nor ( n54524 , n54522 , n54523 );
xnor ( n54525 , n54524 , n52526 );
and ( n54526 , n54520 , n54525 );
and ( n54527 , n54516 , n54525 );
or ( n54528 , n54521 , n54526 , n54527 );
xor ( n54529 , n53647 , n53766 );
xor ( n54530 , n53766 , n53762 );
not ( n54531 , n54530 );
and ( n54532 , n54529 , n54531 );
and ( n54533 , n51924 , n54532 );
not ( n54534 , n54533 );
xnor ( n54535 , n54534 , n53769 );
and ( n54536 , n54528 , n54535 );
and ( n54537 , n52000 , n53996 );
and ( n54538 , n51965 , n53994 );
nor ( n54539 , n54537 , n54538 );
xnor ( n54540 , n54539 , n53376 );
and ( n54541 , n54535 , n54540 );
and ( n54542 , n54528 , n54540 );
or ( n54543 , n54536 , n54541 , n54542 );
and ( n54544 , n53639 , n52065 );
and ( n54545 , n53641 , n52063 );
nor ( n54546 , n54544 , n54545 );
xnor ( n54547 , n54546 , n52022 );
and ( n54548 , n54215 , n51936 );
and ( n54549 , n54055 , n51934 );
nor ( n54550 , n54548 , n54549 );
xnor ( n54551 , n54550 , n51941 );
and ( n54552 , n54547 , n54551 );
buf ( n54553 , n578891 );
and ( n54554 , n54553 , n51929 );
and ( n54555 , n54321 , n51927 );
nor ( n54556 , n54554 , n54555 );
not ( n54557 , n54556 );
and ( n54558 , n54551 , n54557 );
and ( n54559 , n54547 , n54557 );
or ( n54560 , n54552 , n54558 , n54559 );
and ( n54561 , n53367 , n52155 );
and ( n54562 , n53107 , n52153 );
nor ( n54563 , n54561 , n54562 );
xnor ( n54564 , n54563 , n52085 );
and ( n54565 , n54560 , n54564 );
and ( n54566 , n53837 , n51991 );
and ( n54567 , n53639 , n51989 );
nor ( n54568 , n54566 , n54567 );
xnor ( n54569 , n54568 , n51959 );
and ( n54570 , n54564 , n54569 );
and ( n54571 , n54560 , n54569 );
or ( n54572 , n54565 , n54570 , n54571 );
and ( n54573 , n52934 , n52273 );
and ( n54574 , n52936 , n52271 );
nor ( n54575 , n54573 , n54574 );
xnor ( n54576 , n54575 , n52137 );
and ( n54577 , n54572 , n54576 );
xor ( n54578 , n54209 , n54213 );
xor ( n54579 , n54578 , n54219 );
and ( n54580 , n54576 , n54579 );
and ( n54581 , n54572 , n54579 );
or ( n54582 , n54577 , n54580 , n54581 );
and ( n54583 , n52671 , n52509 );
and ( n54584 , n52626 , n52507 );
nor ( n54585 , n54583 , n54584 );
xnor ( n54586 , n54585 , n52383 );
and ( n54587 , n54582 , n54586 );
xor ( n54588 , n54301 , n54305 );
xor ( n54589 , n54588 , n54308 );
and ( n54590 , n54586 , n54589 );
and ( n54591 , n54582 , n54589 );
or ( n54592 , n54587 , n54590 , n54591 );
and ( n54593 , n52488 , n52707 );
and ( n54594 , n52390 , n52705 );
nor ( n54595 , n54593 , n54594 );
xnor ( n54596 , n54595 , n52526 );
and ( n54597 , n54592 , n54596 );
and ( n54598 , n52626 , n52509 );
and ( n54599 , n52533 , n52507 );
nor ( n54600 , n54598 , n54599 );
xnor ( n54601 , n54600 , n52383 );
and ( n54602 , n54596 , n54601 );
and ( n54603 , n54592 , n54601 );
or ( n54604 , n54597 , n54602 , n54603 );
and ( n54605 , n54543 , n54604 );
and ( n54606 , n52037 , n53683 );
and ( n54607 , n52029 , n53681 );
nor ( n54608 , n54606 , n54607 );
xnor ( n54609 , n54608 , n53118 );
and ( n54610 , n52115 , n53468 );
and ( n54611 , n52092 , n53466 );
nor ( n54612 , n54610 , n54611 );
xnor ( n54613 , n54612 , n52945 );
and ( n54614 , n54609 , n54613 );
xor ( n54615 , n54311 , n54350 );
xor ( n54616 , n54615 , n54353 );
and ( n54617 , n54613 , n54616 );
and ( n54618 , n54609 , n54616 );
or ( n54619 , n54614 , n54617 , n54618 );
and ( n54620 , n54604 , n54619 );
and ( n54621 , n54543 , n54619 );
or ( n54622 , n54605 , n54620 , n54621 );
xor ( n54623 , n54439 , n54443 );
xor ( n54624 , n54623 , n54446 );
and ( n54625 , n54622 , n54624 );
xor ( n54626 , n54368 , n54370 );
xor ( n54627 , n54626 , n54373 );
and ( n54628 , n54624 , n54627 );
and ( n54629 , n54622 , n54627 );
or ( n54630 , n54625 , n54628 , n54629 );
and ( n54631 , n54512 , n54630 );
xor ( n54632 , n54425 , n54449 );
xor ( n54633 , n54632 , n54452 );
and ( n54634 , n54630 , n54633 );
and ( n54635 , n54512 , n54633 );
or ( n54636 , n54631 , n54634 , n54635 );
xor ( n54637 , n54384 , n54455 );
xor ( n54638 , n54637 , n54458 );
and ( n54639 , n54636 , n54638 );
xor ( n54640 , n54272 , n54274 );
xor ( n54641 , n54640 , n54277 );
and ( n54642 , n54638 , n54641 );
and ( n54643 , n54636 , n54641 );
or ( n54644 , n54639 , n54642 , n54643 );
xor ( n54645 , n54461 , n54463 );
xor ( n54646 , n54645 , n54466 );
and ( n54647 , n54644 , n54646 );
xor ( n54648 , n54636 , n54638 );
xor ( n54649 , n54648 , n54641 );
and ( n54650 , n52669 , n52509 );
and ( n54651 , n52671 , n52507 );
nor ( n54652 , n54650 , n54651 );
xnor ( n54653 , n54652 , n52383 );
and ( n54654 , n52816 , n52432 );
and ( n54655 , n52818 , n52430 );
nor ( n54656 , n54654 , n54655 );
xnor ( n54657 , n54656 , n52255 );
and ( n54658 , n54653 , n54657 );
xor ( n54659 , n54328 , n54332 );
xor ( n54660 , n54659 , n54337 );
and ( n54661 , n54657 , n54660 );
and ( n54662 , n54653 , n54660 );
or ( n54663 , n54658 , n54661 , n54662 );
and ( n54664 , n52092 , n53683 );
and ( n54665 , n52037 , n53681 );
nor ( n54666 , n54664 , n54665 );
xnor ( n54667 , n54666 , n53118 );
and ( n54668 , n54663 , n54667 );
xor ( n54669 , n54340 , n54344 );
xor ( n54670 , n54669 , n54347 );
and ( n54671 , n54667 , n54670 );
and ( n54672 , n54663 , n54670 );
or ( n54673 , n54668 , n54671 , n54672 );
xor ( n54674 , n54592 , n54596 );
xor ( n54675 , n54674 , n54601 );
and ( n54676 , n54673 , n54675 );
xor ( n54677 , n54474 , n54478 );
xor ( n54678 , n54677 , n54481 );
and ( n54679 , n54675 , n54678 );
and ( n54680 , n54673 , n54678 );
or ( n54681 , n54676 , n54679 , n54680 );
xor ( n54682 , n54356 , n54360 );
xor ( n54683 , n54682 , n54365 );
and ( n54684 , n54681 , n54683 );
xor ( n54685 , n54484 , n54488 );
xor ( n54686 , n54685 , n54491 );
and ( n54687 , n54683 , n54686 );
and ( n54688 , n54681 , n54686 );
or ( n54689 , n54684 , n54687 , n54688 );
and ( n54690 , n52934 , n52432 );
and ( n54691 , n52936 , n52430 );
nor ( n54692 , n54690 , n54691 );
xnor ( n54693 , n54692 , n52255 );
and ( n54694 , n53107 , n52273 );
and ( n54695 , n53109 , n52271 );
nor ( n54696 , n54694 , n54695 );
xnor ( n54697 , n54696 , n52137 );
and ( n54698 , n54693 , n54697 );
xor ( n54699 , n54547 , n54551 );
xor ( n54700 , n54699 , n54557 );
and ( n54701 , n54697 , n54700 );
and ( n54702 , n54693 , n54700 );
or ( n54703 , n54698 , n54701 , n54702 );
and ( n54704 , n52818 , n52509 );
and ( n54705 , n52669 , n52507 );
nor ( n54706 , n54704 , n54705 );
xnor ( n54707 , n54706 , n52383 );
and ( n54708 , n54703 , n54707 );
and ( n54709 , n52936 , n52432 );
and ( n54710 , n52816 , n52430 );
nor ( n54711 , n54709 , n54710 );
xnor ( n54712 , n54711 , n52255 );
and ( n54713 , n54707 , n54712 );
and ( n54714 , n54703 , n54712 );
or ( n54715 , n54708 , n54713 , n54714 );
and ( n54716 , n54055 , n51991 );
and ( n54717 , n53835 , n51989 );
nor ( n54718 , n54716 , n54717 );
xnor ( n54719 , n54718 , n51959 );
and ( n54720 , n54321 , n51936 );
and ( n54721 , n54215 , n51934 );
nor ( n54722 , n54720 , n54721 );
xnor ( n54723 , n54722 , n51941 );
and ( n54724 , n54719 , n54723 );
buf ( n54725 , n578892 );
and ( n54726 , n54725 , n51929 );
and ( n54727 , n54553 , n51927 );
nor ( n54728 , n54726 , n54727 );
not ( n54729 , n54728 );
and ( n54730 , n54723 , n54729 );
and ( n54731 , n54719 , n54729 );
or ( n54732 , n54724 , n54730 , n54731 );
and ( n54733 , n53365 , n52155 );
and ( n54734 , n53367 , n52153 );
nor ( n54735 , n54733 , n54734 );
xnor ( n54736 , n54735 , n52085 );
and ( n54737 , n54732 , n54736 );
and ( n54738 , n53835 , n51991 );
and ( n54739 , n53837 , n51989 );
nor ( n54740 , n54738 , n54739 );
xnor ( n54741 , n54740 , n51959 );
and ( n54742 , n54736 , n54741 );
and ( n54743 , n54732 , n54741 );
or ( n54744 , n54737 , n54742 , n54743 );
and ( n54745 , n53109 , n52273 );
and ( n54746 , n52934 , n52271 );
nor ( n54747 , n54745 , n54746 );
xnor ( n54748 , n54747 , n52137 );
and ( n54749 , n54744 , n54748 );
xor ( n54750 , n54315 , n54319 );
xor ( n54751 , n54750 , n54325 );
and ( n54752 , n54748 , n54751 );
and ( n54753 , n54744 , n54751 );
or ( n54754 , n54749 , n54752 , n54753 );
and ( n54755 , n54715 , n54754 );
xor ( n54756 , n54572 , n54576 );
xor ( n54757 , n54756 , n54579 );
and ( n54758 , n54754 , n54757 );
and ( n54759 , n54715 , n54757 );
or ( n54760 , n54755 , n54758 , n54759 );
and ( n54761 , n52029 , n53996 );
and ( n54762 , n52000 , n53994 );
nor ( n54763 , n54761 , n54762 );
xnor ( n54764 , n54763 , n53376 );
and ( n54765 , n54760 , n54764 );
and ( n54766 , n52144 , n53468 );
and ( n54767 , n52115 , n53466 );
nor ( n54768 , n54766 , n54767 );
xnor ( n54769 , n54768 , n52945 );
and ( n54770 , n54764 , n54769 );
and ( n54771 , n54760 , n54769 );
or ( n54772 , n54765 , n54770 , n54771 );
and ( n54773 , n52194 , n53468 );
and ( n54774 , n52144 , n53466 );
nor ( n54775 , n54773 , n54774 );
xnor ( n54776 , n54775 , n52945 );
and ( n54777 , n52304 , n53177 );
and ( n54778 , n52262 , n53175 );
nor ( n54779 , n54777 , n54778 );
xnor ( n54780 , n54779 , n52827 );
and ( n54781 , n54776 , n54780 );
xor ( n54782 , n54653 , n54657 );
xor ( n54783 , n54782 , n54660 );
and ( n54784 , n54780 , n54783 );
and ( n54785 , n54776 , n54783 );
or ( n54786 , n54781 , n54784 , n54785 );
and ( n54787 , n51965 , n54414 );
and ( n54788 , n51967 , n54412 );
nor ( n54789 , n54787 , n54788 );
xnor ( n54790 , n54789 , n53650 );
and ( n54791 , n54786 , n54790 );
xor ( n54792 , n54582 , n54586 );
xor ( n54793 , n54792 , n54589 );
and ( n54794 , n54790 , n54793 );
and ( n54795 , n54786 , n54793 );
or ( n54796 , n54791 , n54794 , n54795 );
and ( n54797 , n54772 , n54796 );
and ( n54798 , n51967 , n54414 );
and ( n54799 , n51946 , n54412 );
nor ( n54800 , n54798 , n54799 );
xnor ( n54801 , n54800 , n53650 );
and ( n54802 , n54796 , n54801 );
and ( n54803 , n54772 , n54801 );
or ( n54804 , n54797 , n54802 , n54803 );
xor ( n54805 , n54543 , n54604 );
xor ( n54806 , n54805 , n54619 );
and ( n54807 , n54804 , n54806 );
xor ( n54808 , n54498 , n54500 );
xor ( n54809 , n54808 , n54503 );
and ( n54810 , n54806 , n54809 );
and ( n54811 , n54804 , n54809 );
or ( n54812 , n54807 , n54810 , n54811 );
and ( n54813 , n54689 , n54812 );
xor ( n54814 , n54494 , n54506 );
xor ( n54815 , n54814 , n54509 );
and ( n54816 , n54812 , n54815 );
and ( n54817 , n54689 , n54815 );
or ( n54818 , n54813 , n54816 , n54817 );
xor ( n54819 , n54376 , n54378 );
xor ( n54820 , n54819 , n54381 );
and ( n54821 , n54818 , n54820 );
xor ( n54822 , n54512 , n54630 );
xor ( n54823 , n54822 , n54633 );
and ( n54824 , n54820 , n54823 );
and ( n54825 , n54818 , n54823 );
or ( n54826 , n54821 , n54824 , n54825 );
and ( n54827 , n54649 , n54826 );
and ( n54828 , n52671 , n52707 );
and ( n54829 , n52626 , n52705 );
nor ( n54830 , n54828 , n54829 );
xnor ( n54831 , n54830 , n52526 );
xor ( n54832 , n54560 , n54564 );
xor ( n54833 , n54832 , n54569 );
and ( n54834 , n54831 , n54833 );
xor ( n54835 , n54744 , n54748 );
xor ( n54836 , n54835 , n54751 );
and ( n54837 , n54833 , n54836 );
and ( n54838 , n54831 , n54836 );
or ( n54839 , n54834 , n54837 , n54838 );
and ( n54840 , n52488 , n52978 );
and ( n54841 , n52390 , n52976 );
nor ( n54842 , n54840 , n54841 );
xnor ( n54843 , n54842 , n52680 );
and ( n54844 , n54839 , n54843 );
and ( n54845 , n52626 , n52707 );
and ( n54846 , n52533 , n52705 );
nor ( n54847 , n54845 , n54846 );
xnor ( n54848 , n54847 , n52526 );
and ( n54849 , n54843 , n54848 );
and ( n54850 , n54839 , n54848 );
or ( n54851 , n54844 , n54849 , n54850 );
xor ( n54852 , n54516 , n54520 );
xor ( n54853 , n54852 , n54525 );
and ( n54854 , n54851 , n54853 );
xor ( n54855 , n54663 , n54667 );
xor ( n54856 , n54855 , n54670 );
and ( n54857 , n54853 , n54856 );
and ( n54858 , n54851 , n54856 );
or ( n54859 , n54854 , n54857 , n54858 );
xor ( n54860 , n54528 , n54535 );
xor ( n54861 , n54860 , n54540 );
and ( n54862 , n54859 , n54861 );
xor ( n54863 , n54609 , n54613 );
xor ( n54864 , n54863 , n54616 );
and ( n54865 , n54861 , n54864 );
and ( n54866 , n54859 , n54864 );
or ( n54867 , n54862 , n54865 , n54866 );
and ( n54868 , n53109 , n52432 );
and ( n54869 , n52934 , n52430 );
nor ( n54870 , n54868 , n54869 );
xnor ( n54871 , n54870 , n52255 );
and ( n54872 , n53641 , n52155 );
and ( n54873 , n53365 , n52153 );
nor ( n54874 , n54872 , n54873 );
xnor ( n54875 , n54874 , n52085 );
and ( n54876 , n54871 , n54875 );
and ( n54877 , n53837 , n52065 );
and ( n54878 , n53639 , n52063 );
nor ( n54879 , n54877 , n54878 );
xnor ( n54880 , n54879 , n52022 );
and ( n54881 , n54875 , n54880 );
and ( n54882 , n54871 , n54880 );
or ( n54883 , n54876 , n54881 , n54882 );
and ( n54884 , n54215 , n51991 );
and ( n54885 , n54055 , n51989 );
nor ( n54886 , n54884 , n54885 );
xnor ( n54887 , n54886 , n51959 );
and ( n54888 , n54553 , n51936 );
and ( n54889 , n54321 , n51934 );
nor ( n54890 , n54888 , n54889 );
xnor ( n54891 , n54890 , n51941 );
and ( n54892 , n54887 , n54891 );
buf ( n54893 , n578893 );
and ( n54894 , n54893 , n51929 );
and ( n54895 , n54725 , n51927 );
nor ( n54896 , n54894 , n54895 );
not ( n54897 , n54896 );
and ( n54898 , n54891 , n54897 );
and ( n54899 , n54887 , n54897 );
or ( n54900 , n54892 , n54898 , n54899 );
and ( n54901 , n53367 , n52273 );
and ( n54902 , n53107 , n52271 );
nor ( n54903 , n54901 , n54902 );
xnor ( n54904 , n54903 , n52137 );
and ( n54905 , n54900 , n54904 );
xor ( n54906 , n54719 , n54723 );
xor ( n54907 , n54906 , n54729 );
and ( n54908 , n54904 , n54907 );
and ( n54909 , n54900 , n54907 );
or ( n54910 , n54905 , n54908 , n54909 );
and ( n54911 , n54883 , n54910 );
xor ( n54912 , n54732 , n54736 );
xor ( n54913 , n54912 , n54741 );
and ( n54914 , n54910 , n54913 );
and ( n54915 , n54883 , n54913 );
or ( n54916 , n54911 , n54914 , n54915 );
and ( n54917 , n52262 , n53468 );
and ( n54918 , n52194 , n53466 );
nor ( n54919 , n54917 , n54918 );
xnor ( n54920 , n54919 , n52945 );
and ( n54921 , n54916 , n54920 );
and ( n54922 , n52390 , n53177 );
and ( n54923 , n52304 , n53175 );
nor ( n54924 , n54922 , n54923 );
xnor ( n54925 , n54924 , n52827 );
and ( n54926 , n54920 , n54925 );
and ( n54927 , n54916 , n54925 );
or ( n54928 , n54921 , n54926 , n54927 );
and ( n54929 , n52669 , n52707 );
and ( n54930 , n52671 , n52705 );
nor ( n54931 , n54929 , n54930 );
xnor ( n54932 , n54931 , n52526 );
and ( n54933 , n52816 , n52509 );
and ( n54934 , n52818 , n52507 );
nor ( n54935 , n54933 , n54934 );
xnor ( n54936 , n54935 , n52383 );
and ( n54937 , n54932 , n54936 );
xor ( n54938 , n54693 , n54697 );
xor ( n54939 , n54938 , n54700 );
and ( n54940 , n54936 , n54939 );
and ( n54941 , n54932 , n54939 );
or ( n54942 , n54937 , n54940 , n54941 );
and ( n54943 , n52533 , n52978 );
and ( n54944 , n52488 , n52976 );
nor ( n54945 , n54943 , n54944 );
xnor ( n54946 , n54945 , n52680 );
and ( n54947 , n54942 , n54946 );
xor ( n54948 , n54703 , n54707 );
xor ( n54949 , n54948 , n54712 );
and ( n54950 , n54946 , n54949 );
and ( n54951 , n54942 , n54949 );
or ( n54952 , n54947 , n54950 , n54951 );
and ( n54953 , n54928 , n54952 );
and ( n54954 , n52000 , n54414 );
and ( n54955 , n51965 , n54412 );
nor ( n54956 , n54954 , n54955 );
xnor ( n54957 , n54956 , n53650 );
and ( n54958 , n54952 , n54957 );
and ( n54959 , n54928 , n54957 );
or ( n54960 , n54953 , n54958 , n54959 );
and ( n54961 , n52037 , n53996 );
and ( n54962 , n52029 , n53994 );
nor ( n54963 , n54961 , n54962 );
xnor ( n54964 , n54963 , n53376 );
and ( n54965 , n52115 , n53683 );
and ( n54966 , n52092 , n53681 );
nor ( n54967 , n54965 , n54966 );
xnor ( n54968 , n54967 , n53118 );
and ( n54969 , n54964 , n54968 );
xor ( n54970 , n54715 , n54754 );
xor ( n54971 , n54970 , n54757 );
and ( n54972 , n54968 , n54971 );
and ( n54973 , n54964 , n54971 );
or ( n54974 , n54969 , n54972 , n54973 );
and ( n54975 , n54960 , n54974 );
and ( n54976 , n51946 , n54532 );
and ( n54977 , n51924 , n54530 );
nor ( n54978 , n54976 , n54977 );
xnor ( n54979 , n54978 , n53769 );
and ( n54980 , n54974 , n54979 );
and ( n54981 , n54960 , n54979 );
or ( n54982 , n54975 , n54980 , n54981 );
xor ( n54983 , n54772 , n54796 );
xor ( n54984 , n54983 , n54801 );
and ( n54985 , n54982 , n54984 );
xor ( n54986 , n54673 , n54675 );
xor ( n54987 , n54986 , n54678 );
and ( n54988 , n54984 , n54987 );
and ( n54989 , n54982 , n54987 );
or ( n54990 , n54985 , n54988 , n54989 );
and ( n54991 , n54867 , n54990 );
xor ( n54992 , n54681 , n54683 );
xor ( n54993 , n54992 , n54686 );
and ( n54994 , n54990 , n54993 );
and ( n54995 , n54867 , n54993 );
or ( n54996 , n54991 , n54994 , n54995 );
xor ( n54997 , n54689 , n54812 );
xor ( n54998 , n54997 , n54815 );
and ( n54999 , n54996 , n54998 );
xor ( n55000 , n54622 , n54624 );
xor ( n55001 , n55000 , n54627 );
and ( n55002 , n54998 , n55001 );
and ( n55003 , n54996 , n55001 );
or ( n55004 , n54999 , n55002 , n55003 );
xor ( n55005 , n54818 , n54820 );
xor ( n55006 , n55005 , n54823 );
and ( n55007 , n55004 , n55006 );
xor ( n55008 , n54996 , n54998 );
xor ( n55009 , n55008 , n55001 );
buf ( n55010 , n579239 );
xor ( n55011 , n53762 , n55010 );
not ( n55012 , n55010 );
and ( n55013 , n55011 , n55012 );
and ( n55014 , n51924 , n55013 );
not ( n55015 , n55014 );
xnor ( n55016 , n55015 , n53762 );
xor ( n55017 , n54839 , n54843 );
xor ( n55018 , n55017 , n54848 );
and ( n55019 , n55016 , n55018 );
xor ( n55020 , n54776 , n54780 );
xor ( n55021 , n55020 , n54783 );
and ( n55022 , n55018 , n55021 );
and ( n55023 , n55016 , n55021 );
or ( n55024 , n55019 , n55022 , n55023 );
xor ( n55025 , n54760 , n54764 );
xor ( n55026 , n55025 , n54769 );
and ( n55027 , n55024 , n55026 );
xor ( n55028 , n54786 , n54790 );
xor ( n55029 , n55028 , n54793 );
and ( n55030 , n55026 , n55029 );
and ( n55031 , n55024 , n55029 );
or ( n55032 , n55027 , n55030 , n55031 );
and ( n55033 , n53365 , n52273 );
and ( n55034 , n53367 , n52271 );
nor ( n55035 , n55033 , n55034 );
xnor ( n55036 , n55035 , n52137 );
and ( n55037 , n53639 , n52155 );
and ( n55038 , n53641 , n52153 );
nor ( n55039 , n55037 , n55038 );
xnor ( n55040 , n55039 , n52085 );
and ( n55041 , n55036 , n55040 );
and ( n55042 , n53835 , n52065 );
and ( n55043 , n53837 , n52063 );
nor ( n55044 , n55042 , n55043 );
xnor ( n55045 , n55044 , n52022 );
and ( n55046 , n55040 , n55045 );
and ( n55047 , n55036 , n55045 );
or ( n55048 , n55041 , n55046 , n55047 );
and ( n55049 , n54321 , n51991 );
and ( n55050 , n54215 , n51989 );
nor ( n55051 , n55049 , n55050 );
xnor ( n55052 , n55051 , n51959 );
and ( n55053 , n54725 , n51936 );
and ( n55054 , n54553 , n51934 );
nor ( n55055 , n55053 , n55054 );
xnor ( n55056 , n55055 , n51941 );
and ( n55057 , n55052 , n55056 );
buf ( n55058 , n578894 );
and ( n55059 , n55058 , n51929 );
and ( n55060 , n54893 , n51927 );
nor ( n55061 , n55059 , n55060 );
not ( n55062 , n55061 );
and ( n55063 , n55056 , n55062 );
and ( n55064 , n55052 , n55062 );
or ( n55065 , n55057 , n55063 , n55064 );
and ( n55066 , n54553 , n51991 );
and ( n55067 , n54321 , n51989 );
nor ( n55068 , n55066 , n55067 );
xnor ( n55069 , n55068 , n51959 );
and ( n55070 , n54893 , n51936 );
and ( n55071 , n54725 , n51934 );
nor ( n55072 , n55070 , n55071 );
xnor ( n55073 , n55072 , n51941 );
and ( n55074 , n55069 , n55073 );
buf ( n55075 , n578895 );
and ( n55076 , n55075 , n51929 );
and ( n55077 , n55058 , n51927 );
nor ( n55078 , n55076 , n55077 );
not ( n55079 , n55078 );
and ( n55080 , n55073 , n55079 );
and ( n55081 , n55069 , n55079 );
or ( n55082 , n55074 , n55080 , n55081 );
and ( n55083 , n53641 , n52273 );
and ( n55084 , n53365 , n52271 );
nor ( n55085 , n55083 , n55084 );
xnor ( n55086 , n55085 , n52137 );
and ( n55087 , n55082 , n55086 );
and ( n55088 , n54055 , n52065 );
and ( n55089 , n53835 , n52063 );
nor ( n55090 , n55088 , n55089 );
xnor ( n55091 , n55090 , n52022 );
and ( n55092 , n55086 , n55091 );
and ( n55093 , n55082 , n55091 );
or ( n55094 , n55087 , n55092 , n55093 );
and ( n55095 , n55065 , n55094 );
and ( n55096 , n53107 , n52432 );
and ( n55097 , n53109 , n52430 );
nor ( n55098 , n55096 , n55097 );
xnor ( n55099 , n55098 , n52255 );
and ( n55100 , n55094 , n55099 );
and ( n55101 , n55065 , n55099 );
or ( n55102 , n55095 , n55100 , n55101 );
and ( n55103 , n55048 , n55102 );
and ( n55104 , n52936 , n52509 );
and ( n55105 , n52816 , n52507 );
nor ( n55106 , n55104 , n55105 );
xnor ( n55107 , n55106 , n52383 );
and ( n55108 , n55102 , n55107 );
and ( n55109 , n55048 , n55107 );
or ( n55110 , n55103 , n55108 , n55109 );
and ( n55111 , n52818 , n52707 );
and ( n55112 , n52669 , n52705 );
nor ( n55113 , n55111 , n55112 );
xnor ( n55114 , n55113 , n52526 );
xor ( n55115 , n54871 , n54875 );
xor ( n55116 , n55115 , n54880 );
and ( n55117 , n55114 , n55116 );
xor ( n55118 , n54900 , n54904 );
xor ( n55119 , n55118 , n54907 );
and ( n55120 , n55116 , n55119 );
and ( n55121 , n55114 , n55119 );
or ( n55122 , n55117 , n55120 , n55121 );
and ( n55123 , n55110 , n55122 );
xor ( n55124 , n54883 , n54910 );
xor ( n55125 , n55124 , n54913 );
and ( n55126 , n55122 , n55125 );
and ( n55127 , n55110 , n55125 );
or ( n55128 , n55123 , n55126 , n55127 );
and ( n55129 , n52092 , n53996 );
and ( n55130 , n52037 , n53994 );
nor ( n55131 , n55129 , n55130 );
xnor ( n55132 , n55131 , n53376 );
and ( n55133 , n55128 , n55132 );
and ( n55134 , n52144 , n53683 );
and ( n55135 , n52115 , n53681 );
nor ( n55136 , n55134 , n55135 );
xnor ( n55137 , n55136 , n53118 );
and ( n55138 , n55132 , n55137 );
and ( n55139 , n55128 , n55137 );
or ( n55140 , n55133 , n55138 , n55139 );
and ( n55141 , n51965 , n54532 );
and ( n55142 , n51967 , n54530 );
nor ( n55143 , n55141 , n55142 );
xnor ( n55144 , n55143 , n53769 );
and ( n55145 , n52029 , n54414 );
and ( n55146 , n52000 , n54412 );
nor ( n55147 , n55145 , n55146 );
xnor ( n55148 , n55147 , n53650 );
and ( n55149 , n55144 , n55148 );
xor ( n55150 , n54831 , n54833 );
xor ( n55151 , n55150 , n54836 );
and ( n55152 , n55148 , n55151 );
and ( n55153 , n55144 , n55151 );
or ( n55154 , n55149 , n55152 , n55153 );
and ( n55155 , n55140 , n55154 );
and ( n55156 , n51967 , n54532 );
and ( n55157 , n51946 , n54530 );
nor ( n55158 , n55156 , n55157 );
xnor ( n55159 , n55158 , n53769 );
and ( n55160 , n55154 , n55159 );
and ( n55161 , n55140 , n55159 );
or ( n55162 , n55155 , n55160 , n55161 );
xor ( n55163 , n54960 , n54974 );
xor ( n55164 , n55163 , n54979 );
and ( n55165 , n55162 , n55164 );
xor ( n55166 , n54851 , n54853 );
xor ( n55167 , n55166 , n54856 );
and ( n55168 , n55164 , n55167 );
and ( n55169 , n55162 , n55167 );
or ( n55170 , n55165 , n55168 , n55169 );
and ( n55171 , n55032 , n55170 );
xor ( n55172 , n54859 , n54861 );
xor ( n55173 , n55172 , n54864 );
and ( n55174 , n55170 , n55173 );
and ( n55175 , n55032 , n55173 );
or ( n55176 , n55171 , n55174 , n55175 );
xor ( n55177 , n54804 , n54806 );
xor ( n55178 , n55177 , n54809 );
and ( n55179 , n55176 , n55178 );
xor ( n55180 , n54867 , n54990 );
xor ( n55181 , n55180 , n54993 );
and ( n55182 , n55178 , n55181 );
and ( n55183 , n55176 , n55181 );
or ( n55184 , n55179 , n55182 , n55183 );
and ( n55185 , n55009 , n55184 );
xor ( n55186 , n55176 , n55178 );
xor ( n55187 , n55186 , n55181 );
and ( n55188 , n52194 , n53683 );
and ( n55189 , n52144 , n53681 );
nor ( n55190 , n55188 , n55189 );
xnor ( n55191 , n55190 , n53118 );
and ( n55192 , n52488 , n53177 );
and ( n55193 , n52390 , n53175 );
nor ( n55194 , n55192 , n55193 );
xnor ( n55195 , n55194 , n52827 );
and ( n55196 , n55191 , n55195 );
and ( n55197 , n52626 , n52978 );
and ( n55198 , n52533 , n52976 );
nor ( n55199 , n55197 , n55198 );
xnor ( n55200 , n55199 , n52680 );
and ( n55201 , n55195 , n55200 );
and ( n55202 , n55191 , n55200 );
or ( n55203 , n55196 , n55201 , n55202 );
and ( n55204 , n51946 , n55013 );
and ( n55205 , n51924 , n55010 );
nor ( n55206 , n55204 , n55205 );
xnor ( n55207 , n55206 , n53762 );
and ( n55208 , n55203 , n55207 );
xor ( n55209 , n54942 , n54946 );
xor ( n55210 , n55209 , n54949 );
and ( n55211 , n55207 , n55210 );
and ( n55212 , n55203 , n55210 );
or ( n55213 , n55208 , n55211 , n55212 );
xor ( n55214 , n54928 , n54952 );
xor ( n55215 , n55214 , n54957 );
and ( n55216 , n55213 , n55215 );
xor ( n55217 , n54964 , n54968 );
xor ( n55218 , n55217 , n54971 );
and ( n55219 , n55215 , n55218 );
and ( n55220 , n55213 , n55218 );
or ( n55221 , n55216 , n55219 , n55220 );
and ( n55222 , n52115 , n53996 );
and ( n55223 , n52092 , n53994 );
nor ( n55224 , n55222 , n55223 );
xnor ( n55225 , n55224 , n53376 );
and ( n55226 , n52304 , n53468 );
and ( n55227 , n52262 , n53466 );
nor ( n55228 , n55226 , n55227 );
xnor ( n55229 , n55228 , n52945 );
and ( n55230 , n55225 , n55229 );
xor ( n55231 , n54932 , n54936 );
xor ( n55232 , n55231 , n54939 );
and ( n55233 , n55229 , n55232 );
and ( n55234 , n55225 , n55232 );
or ( n55235 , n55230 , n55233 , n55234 );
xor ( n55236 , n54916 , n54920 );
xor ( n55237 , n55236 , n54925 );
and ( n55238 , n55235 , n55237 );
xor ( n55239 , n55128 , n55132 );
xor ( n55240 , n55239 , n55137 );
and ( n55241 , n55237 , n55240 );
and ( n55242 , n55235 , n55240 );
or ( n55243 , n55238 , n55241 , n55242 );
and ( n55244 , n53109 , n52509 );
and ( n55245 , n52934 , n52507 );
nor ( n55246 , n55244 , n55245 );
xnor ( n55247 , n55246 , n52383 );
and ( n55248 , n53837 , n52155 );
and ( n55249 , n53639 , n52153 );
nor ( n55250 , n55248 , n55249 );
xnor ( n55251 , n55250 , n52085 );
and ( n55252 , n55247 , n55251 );
xor ( n55253 , n55052 , n55056 );
xor ( n55254 , n55253 , n55062 );
and ( n55255 , n55251 , n55254 );
and ( n55256 , n55247 , n55254 );
or ( n55257 , n55252 , n55255 , n55256 );
and ( n55258 , n52816 , n52707 );
and ( n55259 , n52818 , n52705 );
nor ( n55260 , n55258 , n55259 );
xnor ( n55261 , n55260 , n52526 );
and ( n55262 , n55257 , n55261 );
xor ( n55263 , n55065 , n55094 );
xor ( n55264 , n55263 , n55099 );
and ( n55265 , n55261 , n55264 );
and ( n55266 , n55257 , n55264 );
or ( n55267 , n55262 , n55265 , n55266 );
and ( n55268 , n53365 , n52432 );
and ( n55269 , n53367 , n52430 );
nor ( n55270 , n55268 , n55269 );
xnor ( n55271 , n55270 , n52255 );
and ( n55272 , n53639 , n52273 );
and ( n55273 , n53641 , n52271 );
nor ( n55274 , n55272 , n55273 );
xnor ( n55275 , n55274 , n52137 );
and ( n55276 , n55271 , n55275 );
and ( n55277 , n53835 , n52155 );
and ( n55278 , n53837 , n52153 );
nor ( n55279 , n55277 , n55278 );
xnor ( n55280 , n55279 , n52085 );
and ( n55281 , n55275 , n55280 );
and ( n55282 , n55271 , n55280 );
or ( n55283 , n55276 , n55281 , n55282 );
and ( n55284 , n54725 , n51991 );
and ( n55285 , n54553 , n51989 );
nor ( n55286 , n55284 , n55285 );
xnor ( n55287 , n55286 , n51959 );
and ( n55288 , n55058 , n51936 );
and ( n55289 , n54893 , n51934 );
nor ( n55290 , n55288 , n55289 );
xnor ( n55291 , n55290 , n51941 );
and ( n55292 , n55287 , n55291 );
buf ( n55293 , n578896 );
and ( n55294 , n55293 , n51929 );
and ( n55295 , n55075 , n51927 );
nor ( n55296 , n55294 , n55295 );
not ( n55297 , n55296 );
and ( n55298 , n55291 , n55297 );
and ( n55299 , n55287 , n55297 );
or ( n55300 , n55292 , n55298 , n55299 );
and ( n55301 , n54215 , n52065 );
and ( n55302 , n54055 , n52063 );
nor ( n55303 , n55301 , n55302 );
xnor ( n55304 , n55303 , n52022 );
and ( n55305 , n55300 , n55304 );
xor ( n55306 , n55069 , n55073 );
xor ( n55307 , n55306 , n55079 );
and ( n55308 , n55304 , n55307 );
and ( n55309 , n55300 , n55307 );
or ( n55310 , n55305 , n55308 , n55309 );
and ( n55311 , n55283 , n55310 );
and ( n55312 , n53367 , n52432 );
and ( n55313 , n53107 , n52430 );
nor ( n55314 , n55312 , n55313 );
xnor ( n55315 , n55314 , n52255 );
and ( n55316 , n55310 , n55315 );
and ( n55317 , n55283 , n55315 );
or ( n55318 , n55311 , n55316 , n55317 );
and ( n55319 , n52669 , n52978 );
and ( n55320 , n52671 , n52976 );
nor ( n55321 , n55319 , n55320 );
xnor ( n55322 , n55321 , n52680 );
and ( n55323 , n55318 , n55322 );
and ( n55324 , n52934 , n52509 );
and ( n55325 , n52936 , n52507 );
nor ( n55326 , n55324 , n55325 );
xnor ( n55327 , n55326 , n52383 );
xor ( n55328 , n54887 , n54891 );
xor ( n55329 , n55328 , n54897 );
xor ( n55330 , n55327 , n55329 );
xor ( n55331 , n55036 , n55040 );
xor ( n55332 , n55331 , n55045 );
xor ( n55333 , n55330 , n55332 );
and ( n55334 , n55322 , n55333 );
and ( n55335 , n55318 , n55333 );
or ( n55336 , n55323 , n55334 , n55335 );
and ( n55337 , n55267 , n55336 );
and ( n55338 , n52262 , n53683 );
and ( n55339 , n52194 , n53681 );
nor ( n55340 , n55338 , n55339 );
xnor ( n55341 , n55340 , n53118 );
and ( n55342 , n55336 , n55341 );
and ( n55343 , n55267 , n55341 );
or ( n55344 , n55337 , n55342 , n55343 );
and ( n55345 , n52390 , n53468 );
and ( n55346 , n52304 , n53466 );
nor ( n55347 , n55345 , n55346 );
xnor ( n55348 , n55347 , n52945 );
and ( n55349 , n52533 , n53177 );
and ( n55350 , n52488 , n53175 );
nor ( n55351 , n55349 , n55350 );
xnor ( n55352 , n55351 , n52827 );
and ( n55353 , n55348 , n55352 );
xor ( n55354 , n55114 , n55116 );
xor ( n55355 , n55354 , n55119 );
and ( n55356 , n55352 , n55355 );
and ( n55357 , n55348 , n55355 );
or ( n55358 , n55353 , n55356 , n55357 );
and ( n55359 , n55344 , n55358 );
and ( n55360 , n52000 , n54532 );
and ( n55361 , n51965 , n54530 );
nor ( n55362 , n55360 , n55361 );
xnor ( n55363 , n55362 , n53769 );
and ( n55364 , n55358 , n55363 );
and ( n55365 , n55344 , n55363 );
or ( n55366 , n55359 , n55364 , n55365 );
and ( n55367 , n55327 , n55329 );
and ( n55368 , n55329 , n55332 );
and ( n55369 , n55327 , n55332 );
or ( n55370 , n55367 , n55368 , n55369 );
and ( n55371 , n52671 , n52978 );
and ( n55372 , n52626 , n52976 );
nor ( n55373 , n55371 , n55372 );
xnor ( n55374 , n55373 , n52680 );
and ( n55375 , n55370 , n55374 );
xor ( n55376 , n55048 , n55102 );
xor ( n55377 , n55376 , n55107 );
and ( n55378 , n55374 , n55377 );
and ( n55379 , n55370 , n55377 );
or ( n55380 , n55375 , n55378 , n55379 );
and ( n55381 , n52037 , n54414 );
and ( n55382 , n52029 , n54412 );
nor ( n55383 , n55381 , n55382 );
xnor ( n55384 , n55383 , n53650 );
and ( n55385 , n55380 , n55384 );
xor ( n55386 , n55110 , n55122 );
xor ( n55387 , n55386 , n55125 );
and ( n55388 , n55384 , n55387 );
and ( n55389 , n55380 , n55387 );
or ( n55390 , n55385 , n55388 , n55389 );
and ( n55391 , n55366 , n55390 );
xor ( n55392 , n55144 , n55148 );
xor ( n55393 , n55392 , n55151 );
and ( n55394 , n55390 , n55393 );
and ( n55395 , n55366 , n55393 );
or ( n55396 , n55391 , n55394 , n55395 );
and ( n55397 , n55243 , n55396 );
xor ( n55398 , n55016 , n55018 );
xor ( n55399 , n55398 , n55021 );
and ( n55400 , n55396 , n55399 );
and ( n55401 , n55243 , n55399 );
or ( n55402 , n55397 , n55400 , n55401 );
and ( n55403 , n55221 , n55402 );
xor ( n55404 , n55024 , n55026 );
xor ( n55405 , n55404 , n55029 );
and ( n55406 , n55402 , n55405 );
and ( n55407 , n55221 , n55405 );
or ( n55408 , n55403 , n55406 , n55407 );
xor ( n55409 , n54982 , n54984 );
xor ( n55410 , n55409 , n54987 );
and ( n55411 , n55408 , n55410 );
xor ( n55412 , n55032 , n55170 );
xor ( n55413 , n55412 , n55173 );
and ( n55414 , n55410 , n55413 );
and ( n55415 , n55408 , n55413 );
or ( n55416 , n55411 , n55414 , n55415 );
and ( n55417 , n55187 , n55416 );
xor ( n55418 , n55408 , n55410 );
xor ( n55419 , n55418 , n55413 );
and ( n55420 , n52092 , n54414 );
and ( n55421 , n52037 , n54412 );
nor ( n55422 , n55420 , n55421 );
xnor ( n55423 , n55422 , n53650 );
and ( n55424 , n52144 , n53996 );
and ( n55425 , n52115 , n53994 );
nor ( n55426 , n55424 , n55425 );
xnor ( n55427 , n55426 , n53376 );
and ( n55428 , n55423 , n55427 );
xor ( n55429 , n55370 , n55374 );
xor ( n55430 , n55429 , n55377 );
and ( n55431 , n55427 , n55430 );
and ( n55432 , n55423 , n55430 );
or ( n55433 , n55428 , n55431 , n55432 );
and ( n55434 , n51967 , n55013 );
and ( n55435 , n51946 , n55010 );
nor ( n55436 , n55434 , n55435 );
xnor ( n55437 , n55436 , n53762 );
and ( n55438 , n55433 , n55437 );
xor ( n55439 , n55191 , n55195 );
xor ( n55440 , n55439 , n55200 );
and ( n55441 , n55437 , n55440 );
and ( n55442 , n55433 , n55440 );
or ( n55443 , n55438 , n55441 , n55442 );
xor ( n55444 , n55235 , n55237 );
xor ( n55445 , n55444 , n55240 );
and ( n55446 , n55443 , n55445 );
xor ( n55447 , n55203 , n55207 );
xor ( n55448 , n55447 , n55210 );
and ( n55449 , n55445 , n55448 );
and ( n55450 , n55443 , n55448 );
or ( n55451 , n55446 , n55449 , n55450 );
xor ( n55452 , n55140 , n55154 );
xor ( n55453 , n55452 , n55159 );
and ( n55454 , n55451 , n55453 );
xor ( n55455 , n55213 , n55215 );
xor ( n55456 , n55455 , n55218 );
and ( n55457 , n55453 , n55456 );
and ( n55458 , n55451 , n55456 );
or ( n55459 , n55454 , n55457 , n55458 );
xor ( n55460 , n55162 , n55164 );
xor ( n55461 , n55460 , n55167 );
and ( n582785 , n55459 , n55461 );
xor ( n582786 , n55221 , n55402 );
xor ( n55464 , n582786 , n55405 );
and ( n582788 , n55461 , n55464 );
and ( n582789 , n55459 , n55464 );
or ( n582790 , n582785 , n582788 , n582789 );
and ( n55468 , n55419 , n582790 );
xor ( n582792 , n55459 , n55461 );
xor ( n55470 , n582792 , n55464 );
and ( n582794 , n52194 , n53996 );
and ( n582795 , n52144 , n53994 );
nor ( n55473 , n582794 , n582795 );
xnor ( n582797 , n55473 , n53376 );
and ( n55475 , n52488 , n53468 );
and ( n582799 , n52390 , n53466 );
nor ( n582800 , n55475 , n582799 );
xnor ( n55478 , n582800 , n52945 );
and ( n582802 , n582797 , n55478 );
and ( n582803 , n52626 , n53177 );
and ( n582804 , n52533 , n53175 );
nor ( n582805 , n582803 , n582804 );
xnor ( n55483 , n582805 , n52827 );
and ( n582807 , n55478 , n55483 );
and ( n582808 , n582797 , n55483 );
or ( n55486 , n582802 , n582807 , n582808 );
xor ( n582810 , n55267 , n55336 );
xor ( n582811 , n582810 , n55341 );
and ( n55489 , n55486 , n582811 );
xor ( n582813 , n55348 , n55352 );
xor ( n582814 , n582813 , n55355 );
and ( n55492 , n582811 , n582814 );
and ( n582816 , n55486 , n582814 );
or ( n582817 , n55489 , n55492 , n582816 );
xor ( n582818 , n55344 , n55358 );
xor ( n55496 , n582818 , n55363 );
and ( n582820 , n582817 , n55496 );
xor ( n582821 , n55433 , n55437 );
xor ( n582822 , n582821 , n55440 );
and ( n55500 , n55496 , n582822 );
and ( n582824 , n582817 , n582822 );
or ( n55502 , n582820 , n55500 , n582824 );
and ( n582826 , n53641 , n52432 );
and ( n582827 , n53365 , n52430 );
nor ( n55505 , n582826 , n582827 );
xnor ( n582829 , n55505 , n52255 );
and ( n55507 , n53837 , n52273 );
and ( n55508 , n53639 , n52271 );
nor ( n55509 , n55507 , n55508 );
xnor ( n55510 , n55509 , n52137 );
and ( n582834 , n582829 , n55510 );
and ( n582835 , n54055 , n52155 );
and ( n582836 , n53835 , n52153 );
nor ( n55514 , n582835 , n582836 );
xnor ( n582838 , n55514 , n52085 );
and ( n582839 , n55510 , n582838 );
and ( n582840 , n582829 , n582838 );
or ( n582841 , n582834 , n582839 , n582840 );
and ( n55519 , n54893 , n51991 );
and ( n582843 , n54725 , n51989 );
nor ( n582844 , n55519 , n582843 );
xnor ( n55522 , n582844 , n51959 );
and ( n582846 , n55075 , n51936 );
and ( n582847 , n55058 , n51934 );
nor ( n55525 , n582846 , n582847 );
xnor ( n582849 , n55525 , n51941 );
and ( n582850 , n55522 , n582849 );
buf ( n55528 , n578897 );
and ( n582852 , n55528 , n51929 );
and ( n582853 , n55293 , n51927 );
nor ( n582854 , n582852 , n582853 );
not ( n582855 , n582854 );
and ( n55533 , n582849 , n582855 );
and ( n582857 , n55522 , n582855 );
or ( n582858 , n582850 , n55533 , n582857 );
and ( n582859 , n54321 , n52065 );
and ( n582860 , n54215 , n52063 );
nor ( n55538 , n582859 , n582860 );
xnor ( n582862 , n55538 , n52022 );
and ( n582863 , n582858 , n582862 );
xor ( n55541 , n55287 , n55291 );
xor ( n582865 , n55541 , n55297 );
and ( n582866 , n582862 , n582865 );
and ( n55544 , n582858 , n582865 );
or ( n582868 , n582863 , n582866 , n55544 );
and ( n582869 , n582841 , n582868 );
and ( n55547 , n53107 , n52509 );
and ( n55548 , n53109 , n52507 );
nor ( n55549 , n55547 , n55548 );
xnor ( n582873 , n55549 , n52383 );
and ( n582874 , n582868 , n582873 );
and ( n55552 , n582841 , n582873 );
or ( n582876 , n582869 , n582874 , n55552 );
and ( n55554 , n52934 , n52707 );
and ( n55555 , n52936 , n52705 );
nor ( n55556 , n55554 , n55555 );
xnor ( n55557 , n55556 , n52526 );
xor ( n55558 , n55271 , n55275 );
xor ( n55559 , n55558 , n55280 );
and ( n582883 , n55557 , n55559 );
xor ( n582884 , n55300 , n55304 );
xor ( n55562 , n582884 , n55307 );
and ( n582886 , n55559 , n55562 );
and ( n582887 , n55557 , n55562 );
or ( n55565 , n582883 , n582886 , n582887 );
and ( n582889 , n582876 , n55565 );
xor ( n582890 , n55283 , n55310 );
xor ( n55568 , n582890 , n55315 );
and ( n582892 , n55565 , n55568 );
and ( n582893 , n582876 , n55568 );
or ( n55571 , n582889 , n582892 , n582893 );
and ( n582895 , n52936 , n52707 );
and ( n55573 , n52816 , n52705 );
nor ( n582897 , n582895 , n55573 );
xnor ( n55575 , n582897 , n52526 );
xor ( n55576 , n55082 , n55086 );
xor ( n55577 , n55576 , n55091 );
and ( n55578 , n55575 , n55577 );
xor ( n582902 , n55247 , n55251 );
xor ( n582903 , n582902 , n55254 );
and ( n55581 , n55577 , n582903 );
and ( n582905 , n55575 , n582903 );
or ( n55583 , n55578 , n55581 , n582905 );
and ( n582907 , n55571 , n55583 );
and ( n55585 , n52304 , n53683 );
and ( n582909 , n52262 , n53681 );
nor ( n582910 , n55585 , n582909 );
xnor ( n55588 , n582910 , n53118 );
and ( n582912 , n55583 , n55588 );
and ( n582913 , n55571 , n55588 );
or ( n582914 , n582907 , n582912 , n582913 );
and ( n582915 , n51965 , n55013 );
and ( n55593 , n51967 , n55010 );
nor ( n582917 , n582915 , n55593 );
xnor ( n582918 , n582917 , n53762 );
and ( n55596 , n582914 , n582918 );
and ( n582920 , n52029 , n54532 );
and ( n582921 , n52000 , n54530 );
nor ( n55599 , n582920 , n582921 );
xnor ( n582923 , n55599 , n53769 );
and ( n582924 , n582918 , n582923 );
and ( n55602 , n582914 , n582923 );
or ( n55603 , n55596 , n582924 , n55602 );
xor ( n55604 , n55225 , n55229 );
xor ( n582928 , n55604 , n55232 );
and ( n582929 , n55603 , n582928 );
xor ( n582930 , n55380 , n55384 );
xor ( n55608 , n582930 , n55387 );
and ( n582932 , n582928 , n55608 );
and ( n55610 , n55603 , n55608 );
or ( n55611 , n582929 , n582932 , n55610 );
and ( n582935 , n55502 , n55611 );
xor ( n582936 , n55366 , n55390 );
xor ( n55614 , n582936 , n55393 );
and ( n582938 , n55611 , n55614 );
and ( n55616 , n55502 , n55614 );
or ( n55617 , n582935 , n582938 , n55616 );
xor ( n55618 , n55243 , n55396 );
xor ( n55619 , n55618 , n55399 );
and ( n55620 , n55617 , n55619 );
xor ( n55621 , n55451 , n55453 );
xor ( n582945 , n55621 , n55456 );
and ( n55623 , n55619 , n582945 );
and ( n582947 , n55617 , n582945 );
or ( n55625 , n55620 , n55623 , n582947 );
and ( n582949 , n55470 , n55625 );
xor ( n582950 , n55617 , n55619 );
xor ( n55628 , n582950 , n582945 );
and ( n582952 , n55058 , n51991 );
and ( n582953 , n54893 , n51989 );
nor ( n582954 , n582952 , n582953 );
xnor ( n582955 , n582954 , n51959 );
and ( n55633 , n55293 , n51936 );
and ( n582957 , n55075 , n51934 );
nor ( n582958 , n55633 , n582957 );
xnor ( n55636 , n582958 , n51941 );
and ( n582960 , n582955 , n55636 );
buf ( n582961 , n578898 );
and ( n55639 , n582961 , n51929 );
and ( n582963 , n55528 , n51927 );
nor ( n582964 , n55639 , n582963 );
not ( n55642 , n582964 );
and ( n55643 , n55636 , n55642 );
and ( n55644 , n582955 , n55642 );
or ( n582968 , n582960 , n55643 , n55644 );
and ( n582969 , n54553 , n52065 );
and ( n582970 , n54321 , n52063 );
nor ( n582971 , n582969 , n582970 );
xnor ( n55649 , n582971 , n52022 );
and ( n582973 , n582968 , n55649 );
xor ( n582974 , n55522 , n582849 );
xor ( n582975 , n582974 , n582855 );
and ( n55653 , n55649 , n582975 );
and ( n582977 , n582968 , n582975 );
or ( n582978 , n582973 , n55653 , n582977 );
and ( n55656 , n53109 , n52707 );
and ( n582980 , n52934 , n52705 );
nor ( n55658 , n55656 , n582980 );
xnor ( n582982 , n55658 , n52526 );
and ( n582983 , n582978 , n582982 );
xor ( n55661 , n582858 , n582862 );
xor ( n582985 , n55661 , n582865 );
and ( n55663 , n582982 , n582985 );
and ( n582987 , n582978 , n582985 );
or ( n55665 , n582983 , n55663 , n582987 );
and ( n55666 , n52816 , n52978 );
and ( n582990 , n52818 , n52976 );
nor ( n582991 , n55666 , n582990 );
xnor ( n55669 , n582991 , n52680 );
and ( n582993 , n55665 , n55669 );
xor ( n582994 , n582841 , n582868 );
xor ( n55672 , n582994 , n582873 );
and ( n582996 , n55669 , n55672 );
and ( n582997 , n55665 , n55672 );
or ( n55675 , n582993 , n582996 , n582997 );
and ( n582999 , n52671 , n53177 );
and ( n583000 , n52626 , n53175 );
nor ( n55678 , n582999 , n583000 );
xnor ( n583002 , n55678 , n52827 );
and ( n583003 , n55675 , n583002 );
and ( n55681 , n52818 , n52978 );
and ( n583005 , n52669 , n52976 );
nor ( n583006 , n55681 , n583005 );
xnor ( n583007 , n583006 , n52680 );
and ( n583008 , n583002 , n583007 );
and ( n55686 , n55675 , n583007 );
or ( n583010 , n583003 , n583008 , n55686 );
and ( n583011 , n52037 , n54532 );
and ( n55689 , n52029 , n54530 );
nor ( n583013 , n583011 , n55689 );
xnor ( n583014 , n583013 , n53769 );
and ( n55692 , n583010 , n583014 );
xor ( n583016 , n55571 , n55583 );
xor ( n583017 , n583016 , n55588 );
and ( n55695 , n583014 , n583017 );
and ( n55696 , n583010 , n583017 );
or ( n55697 , n55692 , n55695 , n55696 );
and ( n583021 , n52115 , n54414 );
and ( n583022 , n52092 , n54412 );
nor ( n55700 , n583021 , n583022 );
xnor ( n55701 , n55700 , n53650 );
xor ( n55702 , n55257 , n55261 );
xor ( n583026 , n55702 , n55264 );
and ( n583027 , n55701 , n583026 );
xor ( n55705 , n55318 , n55322 );
xor ( n583029 , n55705 , n55333 );
and ( n55707 , n583026 , n583029 );
and ( n55708 , n55701 , n583029 );
or ( n55709 , n583027 , n55707 , n55708 );
and ( n55710 , n55697 , n55709 );
xor ( n55711 , n55423 , n55427 );
xor ( n583035 , n55711 , n55430 );
and ( n55713 , n55709 , n583035 );
and ( n583037 , n55697 , n583035 );
or ( n583038 , n55710 , n55713 , n583037 );
and ( n55716 , n55075 , n51991 );
and ( n583040 , n55058 , n51989 );
nor ( n55718 , n55716 , n583040 );
xnor ( n583042 , n55718 , n51959 );
and ( n583043 , n55528 , n51936 );
and ( n55721 , n55293 , n51934 );
nor ( n55722 , n583043 , n55721 );
xnor ( n55723 , n55722 , n51941 );
and ( n55724 , n583042 , n55723 );
buf ( n583048 , n578899 );
and ( n55726 , n583048 , n51929 );
and ( n583050 , n582961 , n51927 );
nor ( n55728 , n55726 , n583050 );
not ( n55729 , n55728 );
and ( n583053 , n55723 , n55729 );
and ( n55731 , n583042 , n55729 );
or ( n583055 , n55724 , n583053 , n55731 );
and ( n583056 , n54725 , n52065 );
and ( n55734 , n54553 , n52063 );
nor ( n583058 , n583056 , n55734 );
xnor ( n55736 , n583058 , n52022 );
and ( n55737 , n583055 , n55736 );
xor ( n583061 , n582955 , n55636 );
xor ( n55739 , n583061 , n55642 );
and ( n55740 , n55736 , n55739 );
and ( n55741 , n583055 , n55739 );
or ( n583065 , n55737 , n55740 , n55741 );
and ( n55743 , n53639 , n52432 );
and ( n55744 , n53641 , n52430 );
nor ( n583068 , n55743 , n55744 );
xnor ( n55746 , n583068 , n52255 );
and ( n55747 , n583065 , n55746 );
and ( n55748 , n54215 , n52155 );
and ( n583072 , n54055 , n52153 );
nor ( n583073 , n55748 , n583072 );
xnor ( n55751 , n583073 , n52085 );
and ( n55752 , n55746 , n55751 );
and ( n55753 , n583065 , n55751 );
or ( n55754 , n55747 , n55752 , n55753 );
and ( n55755 , n53367 , n52509 );
and ( n55756 , n53107 , n52507 );
nor ( n55757 , n55755 , n55756 );
xnor ( n55758 , n55757 , n52383 );
and ( n583082 , n55754 , n55758 );
xor ( n583083 , n582829 , n55510 );
xor ( n583084 , n583083 , n582838 );
and ( n55762 , n55758 , n583084 );
and ( n583086 , n55754 , n583084 );
or ( n583087 , n583082 , n55762 , n583086 );
and ( n583088 , n52669 , n53177 );
and ( n55766 , n52671 , n53175 );
nor ( n583090 , n583088 , n55766 );
xnor ( n583091 , n583090 , n52827 );
and ( n583092 , n583087 , n583091 );
xor ( n55770 , n55557 , n55559 );
xor ( n583094 , n55770 , n55562 );
and ( n583095 , n583091 , n583094 );
and ( n55773 , n583087 , n583094 );
or ( n583097 , n583092 , n583095 , n55773 );
and ( n583098 , n52262 , n53996 );
and ( n55776 , n52194 , n53994 );
nor ( n583100 , n583098 , n55776 );
xnor ( n583101 , n583100 , n53376 );
and ( n583102 , n583097 , n583101 );
and ( n583103 , n52390 , n53683 );
and ( n55781 , n52304 , n53681 );
nor ( n583105 , n583103 , n55781 );
xnor ( n583106 , n583105 , n53118 );
and ( n583107 , n583101 , n583106 );
and ( n583108 , n583097 , n583106 );
or ( n55786 , n583102 , n583107 , n583108 );
and ( n583110 , n52533 , n53468 );
and ( n583111 , n52488 , n53466 );
nor ( n55789 , n583110 , n583111 );
xnor ( n583113 , n55789 , n52945 );
xor ( n583114 , n582876 , n55565 );
xor ( n55792 , n583114 , n55568 );
and ( n583116 , n583113 , n55792 );
xor ( n583117 , n55575 , n55577 );
xor ( n55795 , n583117 , n582903 );
and ( n583119 , n55792 , n55795 );
and ( n583120 , n583113 , n55795 );
or ( n583121 , n583116 , n583119 , n583120 );
and ( n583122 , n55786 , n583121 );
and ( n55800 , n52000 , n55013 );
and ( n583124 , n51965 , n55010 );
nor ( n583125 , n55800 , n583124 );
xnor ( n583126 , n583125 , n53762 );
and ( n583127 , n583121 , n583126 );
and ( n55805 , n55786 , n583126 );
or ( n583129 , n583122 , n583127 , n55805 );
xor ( n583130 , n582914 , n582918 );
xor ( n55808 , n583130 , n582923 );
and ( n583132 , n583129 , n55808 );
xor ( n583133 , n55486 , n582811 );
xor ( n55811 , n583133 , n582814 );
and ( n583135 , n55808 , n55811 );
and ( n583136 , n583129 , n55811 );
or ( n55814 , n583132 , n583135 , n583136 );
and ( n583138 , n583038 , n55814 );
xor ( n583139 , n55603 , n582928 );
xor ( n55817 , n583139 , n55608 );
and ( n583141 , n55814 , n55817 );
and ( n583142 , n583038 , n55817 );
or ( n55820 , n583138 , n583141 , n583142 );
xor ( n55821 , n55443 , n55445 );
xor ( n583145 , n55821 , n55448 );
and ( n55823 , n55820 , n583145 );
xor ( n583147 , n55502 , n55611 );
xor ( n583148 , n583147 , n55614 );
and ( n55826 , n583145 , n583148 );
and ( n55827 , n55820 , n583148 );
or ( n583151 , n55823 , n55826 , n55827 );
and ( n55829 , n55628 , n583151 );
xor ( n583153 , n55820 , n583145 );
xor ( n55831 , n583153 , n583148 );
and ( n583155 , n55293 , n51991 );
and ( n55833 , n55075 , n51989 );
nor ( n583157 , n583155 , n55833 );
xnor ( n583158 , n583157 , n51959 );
and ( n55836 , n582961 , n51936 );
and ( n583160 , n55528 , n51934 );
nor ( n55838 , n55836 , n583160 );
xnor ( n583162 , n55838 , n51941 );
and ( n55840 , n583158 , n583162 );
buf ( n55841 , n578900 );
and ( n55842 , n55841 , n51929 );
and ( n55843 , n583048 , n51927 );
nor ( n55844 , n55842 , n55843 );
not ( n55845 , n55844 );
and ( n55846 , n583162 , n55845 );
and ( n55847 , n583158 , n55845 );
or ( n55848 , n55840 , n55846 , n55847 );
and ( n583172 , n54893 , n52065 );
and ( n583173 , n54725 , n52063 );
nor ( n55851 , n583172 , n583173 );
xnor ( n583175 , n55851 , n52022 );
and ( n583176 , n55848 , n583175 );
xor ( n583177 , n583042 , n55723 );
xor ( n55855 , n583177 , n55729 );
and ( n583179 , n583175 , n55855 );
and ( n583180 , n55848 , n55855 );
or ( n583181 , n583176 , n583179 , n583180 );
and ( n55859 , n53641 , n52509 );
and ( n583183 , n53365 , n52507 );
nor ( n583184 , n55859 , n583183 );
xnor ( n55862 , n583184 , n52383 );
and ( n583186 , n583181 , n55862 );
and ( n55864 , n54321 , n52155 );
and ( n583188 , n54215 , n52153 );
nor ( n583189 , n55864 , n583188 );
xnor ( n55867 , n583189 , n52085 );
and ( n583191 , n55862 , n55867 );
and ( n55869 , n583181 , n55867 );
or ( n583193 , n583186 , n583191 , n55869 );
and ( n55871 , n53837 , n52432 );
and ( n55872 , n53639 , n52430 );
nor ( n583196 , n55871 , n55872 );
xnor ( n583197 , n583196 , n52255 );
and ( n55875 , n54055 , n52273 );
and ( n583199 , n53835 , n52271 );
nor ( n583200 , n55875 , n583199 );
xnor ( n55878 , n583200 , n52137 );
and ( n583202 , n583197 , n55878 );
xor ( n583203 , n583055 , n55736 );
xor ( n55881 , n583203 , n55739 );
and ( n583205 , n55878 , n55881 );
and ( n583206 , n583197 , n55881 );
or ( n583207 , n583202 , n583205 , n583206 );
and ( n55885 , n583193 , n583207 );
and ( n583209 , n53107 , n52707 );
and ( n583210 , n53109 , n52705 );
nor ( n55888 , n583209 , n583210 );
xnor ( n583212 , n55888 , n52526 );
and ( n55890 , n583207 , n583212 );
and ( n583214 , n583193 , n583212 );
or ( n583215 , n55885 , n55890 , n583214 );
and ( n583216 , n52818 , n53177 );
and ( n583217 , n52669 , n53175 );
nor ( n55895 , n583216 , n583217 );
xnor ( n583219 , n55895 , n52827 );
and ( n583220 , n583215 , n583219 );
xor ( n55898 , n55754 , n55758 );
xor ( n583222 , n55898 , n583084 );
and ( n55900 , n583219 , n583222 );
and ( n583224 , n583215 , n583222 );
or ( n55902 , n583220 , n55900 , n583224 );
and ( n55903 , n53365 , n52509 );
and ( n583227 , n53367 , n52507 );
nor ( n583228 , n55903 , n583227 );
xnor ( n55906 , n583228 , n52383 );
and ( n583230 , n53835 , n52273 );
and ( n583231 , n53837 , n52271 );
nor ( n55909 , n583230 , n583231 );
xnor ( n583233 , n55909 , n52137 );
and ( n583234 , n55906 , n583233 );
xor ( n55912 , n582968 , n55649 );
xor ( n583236 , n55912 , n582975 );
and ( n583237 , n583233 , n583236 );
and ( n55915 , n55906 , n583236 );
or ( n583239 , n583234 , n583237 , n55915 );
and ( n583240 , n52936 , n52978 );
and ( n55918 , n52816 , n52976 );
nor ( n583242 , n583240 , n55918 );
xnor ( n583243 , n583242 , n52680 );
and ( n583244 , n583239 , n583243 );
xor ( n55922 , n582978 , n582982 );
xor ( n583246 , n55922 , n582985 );
and ( n55924 , n583243 , n583246 );
and ( n583248 , n583239 , n583246 );
or ( n583249 , n583244 , n55924 , n583248 );
and ( n55927 , n55902 , n583249 );
and ( n583251 , n52194 , n54414 );
and ( n55929 , n52144 , n54412 );
nor ( n55930 , n583251 , n55929 );
xnor ( n55931 , n55930 , n53650 );
and ( n583255 , n583249 , n55931 );
and ( n55933 , n55902 , n55931 );
or ( n55934 , n55927 , n583255 , n55933 );
and ( n55935 , n52304 , n53996 );
and ( n583259 , n52262 , n53994 );
nor ( n583260 , n55935 , n583259 );
xnor ( n55938 , n583260 , n53376 );
and ( n583262 , n52626 , n53468 );
and ( n55940 , n52533 , n53466 );
nor ( n55941 , n583262 , n55940 );
xnor ( n583265 , n55941 , n52945 );
and ( n55943 , n55938 , n583265 );
xor ( n583267 , n55665 , n55669 );
xor ( n583268 , n583267 , n55672 );
and ( n55946 , n583265 , n583268 );
and ( n55947 , n55938 , n583268 );
or ( n55948 , n55943 , n55946 , n55947 );
and ( n583272 , n55934 , n55948 );
xor ( n583273 , n55675 , n583002 );
xor ( n55951 , n583273 , n583007 );
and ( n583275 , n55948 , n55951 );
and ( n583276 , n55934 , n55951 );
or ( n55954 , n583272 , n583275 , n583276 );
and ( n583278 , n52115 , n54532 );
and ( n583279 , n52092 , n54530 );
nor ( n583280 , n583278 , n583279 );
xnor ( n583281 , n583280 , n53769 );
and ( n55959 , n52488 , n53683 );
and ( n583283 , n52390 , n53681 );
nor ( n583284 , n55959 , n583283 );
xnor ( n55962 , n583284 , n53118 );
and ( n583286 , n583281 , n55962 );
xor ( n583287 , n583087 , n583091 );
xor ( n55965 , n583287 , n583094 );
and ( n583289 , n55962 , n55965 );
and ( n583290 , n583281 , n55965 );
or ( n55968 , n583286 , n583289 , n583290 );
xor ( n55969 , n583097 , n583101 );
xor ( n55970 , n55969 , n583106 );
and ( n583294 , n55968 , n55970 );
xor ( n583295 , n583113 , n55792 );
xor ( n55973 , n583295 , n55795 );
and ( n55974 , n55970 , n55973 );
and ( n583298 , n55968 , n55973 );
or ( n583299 , n583294 , n55974 , n583298 );
and ( n55977 , n55954 , n583299 );
xor ( n55978 , n583010 , n583014 );
xor ( n55979 , n55978 , n583017 );
and ( n583303 , n583299 , n55979 );
and ( n583304 , n55954 , n55979 );
or ( n55982 , n55977 , n583303 , n583304 );
and ( n583306 , n52029 , n55013 );
and ( n583307 , n52000 , n55010 );
nor ( n55985 , n583306 , n583307 );
xnor ( n583309 , n55985 , n53762 );
and ( n583310 , n52092 , n54532 );
and ( n55988 , n52037 , n54530 );
nor ( n55989 , n583310 , n55988 );
xnor ( n583313 , n55989 , n53769 );
and ( n583314 , n583309 , n583313 );
and ( n55992 , n52144 , n54414 );
and ( n583316 , n52115 , n54412 );
nor ( n55994 , n55992 , n583316 );
xnor ( n55995 , n55994 , n53650 );
and ( n55996 , n583313 , n55995 );
and ( n55997 , n583309 , n55995 );
or ( n55998 , n583314 , n55996 , n55997 );
xor ( n55999 , n582797 , n55478 );
xor ( n56000 , n55999 , n55483 );
and ( n56001 , n55998 , n56000 );
xor ( n56002 , n55701 , n583026 );
xor ( n56003 , n56002 , n583029 );
and ( n56004 , n56000 , n56003 );
and ( n56005 , n55998 , n56003 );
or ( n56006 , n56001 , n56004 , n56005 );
and ( n56007 , n55982 , n56006 );
xor ( n56008 , n55697 , n55709 );
xor ( n56009 , n56008 , n583035 );
and ( n56010 , n56006 , n56009 );
and ( n56011 , n55982 , n56009 );
or ( n56012 , n56007 , n56010 , n56011 );
xor ( n56013 , n582817 , n55496 );
xor ( n56014 , n56013 , n582822 );
and ( n56015 , n56012 , n56014 );
xor ( n56016 , n583038 , n55814 );
xor ( n56017 , n56016 , n55817 );
and ( n56018 , n56014 , n56017 );
and ( n56019 , n56012 , n56017 );
or ( n56020 , n56015 , n56018 , n56019 );
and ( n56021 , n55831 , n56020 );
xor ( n56022 , n56012 , n56014 );
xor ( n56023 , n56022 , n56017 );
xor ( n56024 , n55786 , n583121 );
xor ( n56025 , n56024 , n583126 );
xor ( n56026 , n55954 , n583299 );
xor ( n56027 , n56026 , n55979 );
and ( n56028 , n56025 , n56027 );
xor ( n56029 , n55998 , n56000 );
xor ( n56030 , n56029 , n56003 );
and ( n56031 , n56027 , n56030 );
and ( n56032 , n56025 , n56030 );
or ( n56033 , n56028 , n56031 , n56032 );
xor ( n56034 , n55982 , n56006 );
xor ( n56035 , n56034 , n56009 );
and ( n56036 , n56033 , n56035 );
xor ( n56037 , n583129 , n55808 );
xor ( n56038 , n56037 , n55811 );
and ( n583362 , n56035 , n56038 );
and ( n583363 , n56033 , n56038 );
or ( n583364 , n56036 , n583362 , n583363 );
and ( n56042 , n56023 , n583364 );
xor ( n583366 , n56033 , n56035 );
xor ( n583367 , n583366 , n56038 );
and ( n583368 , n55528 , n51991 );
and ( n583369 , n55293 , n51989 );
nor ( n56047 , n583368 , n583369 );
xnor ( n583371 , n56047 , n51959 );
and ( n583372 , n583048 , n51936 );
and ( n56050 , n582961 , n51934 );
nor ( n583374 , n583372 , n56050 );
xnor ( n583375 , n583374 , n51941 );
and ( n56053 , n583371 , n583375 );
buf ( n583377 , n578901 );
and ( n583378 , n583377 , n51929 );
and ( n56056 , n55841 , n51927 );
nor ( n583380 , n583378 , n56056 );
not ( n583381 , n583380 );
and ( n583382 , n583375 , n583381 );
and ( n56060 , n583371 , n583381 );
or ( n583384 , n56053 , n583382 , n56060 );
and ( n583385 , n54725 , n52155 );
and ( n583386 , n54553 , n52153 );
nor ( n56064 , n583385 , n583386 );
xnor ( n583388 , n56064 , n52085 );
and ( n56066 , n583384 , n583388 );
and ( n583390 , n55058 , n52065 );
and ( n583391 , n54893 , n52063 );
nor ( n56069 , n583390 , n583391 );
xnor ( n583393 , n56069 , n52022 );
and ( n56071 , n583388 , n583393 );
and ( n56072 , n583384 , n583393 );
or ( n583396 , n56066 , n56071 , n56072 );
and ( n583397 , n54553 , n52155 );
and ( n56075 , n54321 , n52153 );
nor ( n583399 , n583397 , n56075 );
xnor ( n583400 , n583399 , n52085 );
and ( n583401 , n583396 , n583400 );
xor ( n583402 , n55848 , n583175 );
xor ( n56080 , n583402 , n55855 );
and ( n583404 , n583400 , n56080 );
and ( n583405 , n583396 , n56080 );
or ( n56083 , n583401 , n583404 , n583405 );
and ( n583407 , n53109 , n52978 );
and ( n583408 , n52934 , n52976 );
nor ( n56086 , n583407 , n583408 );
xnor ( n583410 , n56086 , n52680 );
and ( n583411 , n56083 , n583410 );
xor ( n56089 , n583181 , n55862 );
xor ( n583413 , n56089 , n55867 );
and ( n56091 , n583410 , n583413 );
and ( n56092 , n56083 , n583413 );
or ( n56093 , n583411 , n56091 , n56092 );
and ( n56094 , n53639 , n52509 );
and ( n56095 , n53641 , n52507 );
nor ( n56096 , n56094 , n56095 );
xnor ( n56097 , n56096 , n52383 );
and ( n56098 , n53835 , n52432 );
and ( n56099 , n53837 , n52430 );
nor ( n583423 , n56098 , n56099 );
xnor ( n583424 , n583423 , n52255 );
and ( n56102 , n56097 , n583424 );
and ( n56103 , n54215 , n52273 );
and ( n56104 , n54055 , n52271 );
nor ( n56105 , n56103 , n56104 );
xnor ( n583429 , n56105 , n52137 );
and ( n583430 , n583424 , n583429 );
and ( n56108 , n56097 , n583429 );
or ( n583432 , n56102 , n583430 , n56108 );
and ( n583433 , n53367 , n52707 );
and ( n56111 , n53107 , n52705 );
nor ( n583435 , n583433 , n56111 );
xnor ( n583436 , n583435 , n52526 );
and ( n583437 , n583432 , n583436 );
xor ( n583438 , n583197 , n55878 );
xor ( n56116 , n583438 , n55881 );
and ( n583440 , n583436 , n56116 );
and ( n583441 , n583432 , n56116 );
or ( n56119 , n583437 , n583440 , n583441 );
and ( n583443 , n56093 , n56119 );
and ( n583444 , n52816 , n53177 );
and ( n56122 , n52818 , n53175 );
nor ( n583446 , n583444 , n56122 );
xnor ( n583447 , n583446 , n52827 );
and ( n56125 , n56119 , n583447 );
and ( n583449 , n56093 , n583447 );
or ( n583450 , n583443 , n56125 , n583449 );
and ( n56128 , n52934 , n52978 );
and ( n583452 , n52936 , n52976 );
nor ( n56130 , n56128 , n583452 );
xnor ( n56131 , n56130 , n52680 );
xor ( n56132 , n583065 , n55746 );
xor ( n56133 , n56132 , n55751 );
and ( n56134 , n56131 , n56133 );
xor ( n56135 , n55906 , n583233 );
xor ( n583459 , n56135 , n583236 );
and ( n56137 , n56133 , n583459 );
and ( n56138 , n56131 , n583459 );
or ( n56139 , n56134 , n56137 , n56138 );
and ( n56140 , n583450 , n56139 );
and ( n583464 , n52671 , n53468 );
and ( n583465 , n52626 , n53466 );
nor ( n56143 , n583464 , n583465 );
xnor ( n583467 , n56143 , n52945 );
and ( n56145 , n56139 , n583467 );
and ( n56146 , n583450 , n583467 );
or ( n56147 , n56140 , n56145 , n56146 );
and ( n56148 , n52669 , n53468 );
and ( n56149 , n52671 , n53466 );
nor ( n56150 , n56148 , n56149 );
xnor ( n56151 , n56150 , n52945 );
xor ( n56152 , n583193 , n583207 );
xor ( n56153 , n56152 , n583212 );
and ( n56154 , n56151 , n56153 );
xor ( n56155 , n56131 , n56133 );
xor ( n56156 , n56155 , n583459 );
and ( n56157 , n56153 , n56156 );
and ( n56158 , n56151 , n56156 );
or ( n56159 , n56154 , n56157 , n56158 );
xor ( n583483 , n583215 , n583219 );
xor ( n56161 , n583483 , n583222 );
and ( n583485 , n56159 , n56161 );
xor ( n583486 , n583239 , n583243 );
xor ( n56164 , n583486 , n583246 );
and ( n583488 , n56161 , n56164 );
and ( n56166 , n56159 , n56164 );
or ( n583490 , n583485 , n583488 , n56166 );
and ( n583491 , n56147 , n583490 );
and ( n56169 , n52037 , n55013 );
and ( n56170 , n52029 , n55010 );
nor ( n56171 , n56169 , n56170 );
xnor ( n583495 , n56171 , n53762 );
and ( n583496 , n583490 , n583495 );
and ( n56174 , n56147 , n583495 );
or ( n56175 , n583491 , n583496 , n56174 );
and ( n56176 , n52262 , n54414 );
and ( n583500 , n52194 , n54412 );
nor ( n583501 , n56176 , n583500 );
xnor ( n56179 , n583501 , n53650 );
and ( n56180 , n52390 , n53996 );
and ( n56181 , n52304 , n53994 );
nor ( n56182 , n56180 , n56181 );
xnor ( n56183 , n56182 , n53376 );
and ( n56184 , n56179 , n56183 );
and ( n56185 , n52533 , n53683 );
and ( n583509 , n52488 , n53681 );
nor ( n583510 , n56185 , n583509 );
xnor ( n56188 , n583510 , n53118 );
and ( n583512 , n56183 , n56188 );
and ( n56190 , n56179 , n56188 );
or ( n583514 , n56184 , n583512 , n56190 );
xor ( n56192 , n55902 , n583249 );
xor ( n583516 , n56192 , n55931 );
and ( n56194 , n583514 , n583516 );
xor ( n583518 , n55938 , n583265 );
xor ( n56196 , n583518 , n583268 );
and ( n56197 , n583516 , n56196 );
and ( n56198 , n583514 , n56196 );
or ( n56199 , n56194 , n56197 , n56198 );
and ( n56200 , n56175 , n56199 );
xor ( n56201 , n583309 , n583313 );
xor ( n56202 , n56201 , n55995 );
and ( n56203 , n56199 , n56202 );
and ( n56204 , n56175 , n56202 );
or ( n56205 , n56200 , n56203 , n56204 );
and ( n56206 , n52092 , n55013 );
and ( n56207 , n52037 , n55010 );
nor ( n56208 , n56206 , n56207 );
xnor ( n56209 , n56208 , n53762 );
and ( n56210 , n52144 , n54532 );
and ( n56211 , n52115 , n54530 );
nor ( n56212 , n56210 , n56211 );
xnor ( n56213 , n56212 , n53769 );
and ( n56214 , n56209 , n56213 );
xor ( n56215 , n583450 , n56139 );
xor ( n56216 , n56215 , n583467 );
and ( n56217 , n56213 , n56216 );
and ( n56218 , n56209 , n56216 );
or ( n56219 , n56214 , n56217 , n56218 );
xor ( n56220 , n56147 , n583490 );
xor ( n56221 , n56220 , n583495 );
and ( n56222 , n56219 , n56221 );
xor ( n56223 , n583281 , n55962 );
xor ( n56224 , n56223 , n55965 );
and ( n56225 , n56221 , n56224 );
and ( n56226 , n56219 , n56224 );
or ( n56227 , n56222 , n56225 , n56226 );
xor ( n56228 , n55934 , n55948 );
xor ( n56229 , n56228 , n55951 );
and ( n56230 , n56227 , n56229 );
xor ( n56231 , n55968 , n55970 );
xor ( n56232 , n56231 , n55973 );
and ( n56233 , n56229 , n56232 );
and ( n56234 , n56227 , n56232 );
or ( n56235 , n56230 , n56233 , n56234 );
and ( n56236 , n56205 , n56235 );
xor ( n56237 , n56025 , n56027 );
xor ( n56238 , n56237 , n56030 );
and ( n56239 , n56235 , n56238 );
and ( n583563 , n56205 , n56238 );
or ( n56241 , n56236 , n56239 , n583563 );
and ( n583565 , n583367 , n56241 );
xor ( n56243 , n56205 , n56235 );
xor ( n56244 , n56243 , n56238 );
and ( n56245 , n53641 , n52707 );
and ( n56246 , n53365 , n52705 );
nor ( n56247 , n56245 , n56246 );
xnor ( n56248 , n56247 , n52526 );
and ( n56249 , n54055 , n52432 );
and ( n56250 , n53835 , n52430 );
nor ( n56251 , n56249 , n56250 );
xnor ( n583575 , n56251 , n52255 );
and ( n583576 , n56248 , n583575 );
and ( n56254 , n54321 , n52273 );
and ( n56255 , n54215 , n52271 );
nor ( n56256 , n56254 , n56255 );
xnor ( n56257 , n56256 , n52137 );
and ( n583581 , n583575 , n56257 );
and ( n56259 , n56248 , n56257 );
or ( n583583 , n583576 , n583581 , n56259 );
and ( n583584 , n52934 , n53177 );
and ( n56262 , n52936 , n53175 );
nor ( n56263 , n583584 , n56262 );
xnor ( n56264 , n56263 , n52827 );
and ( n56265 , n583583 , n56264 );
and ( n583589 , n53107 , n52978 );
and ( n583590 , n53109 , n52976 );
nor ( n56268 , n583589 , n583590 );
xnor ( n583592 , n56268 , n52680 );
and ( n583593 , n56264 , n583592 );
and ( n56271 , n583583 , n583592 );
or ( n56272 , n56265 , n583593 , n56271 );
and ( n56273 , n55293 , n52065 );
and ( n56274 , n55075 , n52063 );
nor ( n583598 , n56273 , n56274 );
xnor ( n583599 , n583598 , n52022 );
and ( n56277 , n55841 , n51936 );
and ( n56278 , n583048 , n51934 );
nor ( n56279 , n56277 , n56278 );
xnor ( n56280 , n56279 , n51941 );
and ( n583604 , n583599 , n56280 );
buf ( n56282 , n578902 );
and ( n583606 , n56282 , n51929 );
and ( n583607 , n583377 , n51927 );
nor ( n56285 , n583606 , n583607 );
not ( n583609 , n56285 );
and ( n583610 , n56280 , n583609 );
and ( n583611 , n583599 , n583609 );
or ( n583612 , n583604 , n583610 , n583611 );
and ( n56290 , n55075 , n52065 );
and ( n583614 , n55058 , n52063 );
nor ( n583615 , n56290 , n583614 );
xnor ( n56293 , n583615 , n52022 );
and ( n583617 , n583612 , n56293 );
xor ( n583618 , n583371 , n583375 );
xor ( n56296 , n583618 , n583381 );
and ( n583620 , n56293 , n56296 );
and ( n583621 , n583612 , n56296 );
or ( n56299 , n583617 , n583620 , n583621 );
xor ( n583623 , n583158 , n583162 );
xor ( n583624 , n583623 , n55845 );
and ( n56302 , n56299 , n583624 );
xor ( n583626 , n583384 , n583388 );
xor ( n583627 , n583626 , n583393 );
and ( n56305 , n583624 , n583627 );
and ( n583629 , n56299 , n583627 );
or ( n583630 , n56302 , n56305 , n583629 );
and ( n56308 , n53365 , n52707 );
and ( n583632 , n53367 , n52705 );
nor ( n583633 , n56308 , n583632 );
xnor ( n56311 , n583633 , n52526 );
and ( n56312 , n583630 , n56311 );
xor ( n583636 , n583396 , n583400 );
xor ( n583637 , n583636 , n56080 );
and ( n56315 , n56311 , n583637 );
and ( n56316 , n583630 , n583637 );
or ( n56317 , n56312 , n56315 , n56316 );
and ( n583641 , n56272 , n56317 );
and ( n56319 , n52936 , n53177 );
and ( n583643 , n52816 , n53175 );
nor ( n583644 , n56319 , n583643 );
xnor ( n56322 , n583644 , n52827 );
and ( n583646 , n56317 , n56322 );
and ( n583647 , n56272 , n56322 );
or ( n56325 , n583641 , n583646 , n583647 );
and ( n583649 , n52818 , n53468 );
and ( n56327 , n52669 , n53466 );
nor ( n56328 , n583649 , n56327 );
xnor ( n583652 , n56328 , n52945 );
xor ( n56330 , n56083 , n583410 );
xor ( n583654 , n56330 , n583413 );
and ( n583655 , n583652 , n583654 );
xor ( n56333 , n583432 , n583436 );
xor ( n56334 , n56333 , n56116 );
and ( n56335 , n583654 , n56334 );
and ( n56336 , n583652 , n56334 );
or ( n583660 , n583655 , n56335 , n56336 );
and ( n583661 , n56325 , n583660 );
and ( n56339 , n52488 , n53996 );
and ( n583663 , n52390 , n53994 );
nor ( n583664 , n56339 , n583663 );
xnor ( n56342 , n583664 , n53376 );
and ( n583666 , n583660 , n56342 );
and ( n56344 , n56325 , n56342 );
or ( n56345 , n583661 , n583666 , n56344 );
and ( n583669 , n52194 , n54532 );
and ( n56347 , n52144 , n54530 );
nor ( n583671 , n583669 , n56347 );
xnor ( n583672 , n583671 , n53769 );
and ( n56350 , n52304 , n54414 );
and ( n583674 , n52262 , n54412 );
nor ( n583675 , n56350 , n583674 );
xnor ( n583676 , n583675 , n53650 );
and ( n56354 , n583672 , n583676 );
xor ( n583678 , n56093 , n56119 );
xor ( n56356 , n583678 , n583447 );
and ( n583680 , n583676 , n56356 );
and ( n583681 , n583672 , n56356 );
or ( n56359 , n56354 , n583680 , n583681 );
and ( n583683 , n56345 , n56359 );
and ( n56361 , n52115 , n55013 );
and ( n56362 , n52092 , n55010 );
nor ( n56363 , n56361 , n56362 );
xnor ( n56364 , n56363 , n53762 );
and ( n56365 , n52626 , n53683 );
and ( n583689 , n52533 , n53681 );
nor ( n583690 , n56365 , n583689 );
xnor ( n583691 , n583690 , n53118 );
and ( n56369 , n56364 , n583691 );
xor ( n583693 , n56151 , n56153 );
xor ( n583694 , n583693 , n56156 );
and ( n583695 , n583691 , n583694 );
and ( n583696 , n56364 , n583694 );
or ( n56374 , n56369 , n583695 , n583696 );
and ( n583698 , n56359 , n56374 );
and ( n583699 , n56345 , n56374 );
or ( n56377 , n583683 , n583698 , n583699 );
xor ( n583701 , n56179 , n56183 );
xor ( n583702 , n583701 , n56188 );
xor ( n56380 , n56209 , n56213 );
xor ( n583704 , n56380 , n56216 );
and ( n583705 , n583702 , n583704 );
xor ( n56383 , n56159 , n56161 );
xor ( n583707 , n56383 , n56164 );
and ( n56385 , n583704 , n583707 );
and ( n56386 , n583702 , n583707 );
or ( n583710 , n583705 , n56385 , n56386 );
and ( n56388 , n56377 , n583710 );
xor ( n56389 , n583514 , n583516 );
xor ( n56390 , n56389 , n56196 );
and ( n56391 , n583710 , n56390 );
and ( n583715 , n56377 , n56390 );
or ( n583716 , n56388 , n56391 , n583715 );
xor ( n56394 , n56175 , n56199 );
xor ( n583718 , n56394 , n56202 );
and ( n583719 , n583716 , n583718 );
xor ( n583720 , n56227 , n56229 );
xor ( n56398 , n583720 , n56232 );
and ( n583722 , n583718 , n56398 );
and ( n583723 , n583716 , n56398 );
or ( n583724 , n583719 , n583722 , n583723 );
and ( n583725 , n56244 , n583724 );
xor ( n56403 , n583716 , n583718 );
xor ( n583727 , n56403 , n56398 );
and ( n583728 , n53639 , n52707 );
and ( n56406 , n53641 , n52705 );
nor ( n583730 , n583728 , n56406 );
xnor ( n583731 , n583730 , n52526 );
and ( n56409 , n53835 , n52509 );
and ( n583733 , n53837 , n52507 );
nor ( n583734 , n56409 , n583733 );
xnor ( n56412 , n583734 , n52383 );
and ( n583736 , n583731 , n56412 );
and ( n583737 , n583048 , n51991 );
and ( n583738 , n582961 , n51989 );
nor ( n56416 , n583737 , n583738 );
xnor ( n583740 , n56416 , n51959 );
and ( n583741 , n583377 , n51936 );
and ( n583742 , n55841 , n51934 );
nor ( n583743 , n583741 , n583742 );
xnor ( n56421 , n583743 , n51941 );
and ( n583745 , n583740 , n56421 );
buf ( n583746 , n578903 );
and ( n56424 , n583746 , n51929 );
and ( n583748 , n56282 , n51927 );
nor ( n583749 , n56424 , n583748 );
not ( n56427 , n583749 );
and ( n583751 , n56421 , n56427 );
and ( n583752 , n583740 , n56427 );
or ( n56430 , n583745 , n583751 , n583752 );
and ( n583754 , n55058 , n52155 );
and ( n56432 , n54893 , n52153 );
nor ( n56433 , n583754 , n56432 );
xnor ( n56434 , n56433 , n52085 );
and ( n56435 , n56430 , n56434 );
and ( n56436 , n582961 , n51991 );
and ( n56437 , n55528 , n51989 );
nor ( n56438 , n56436 , n56437 );
xnor ( n56439 , n56438 , n51959 );
and ( n583763 , n56434 , n56439 );
and ( n56441 , n56430 , n56439 );
or ( n583765 , n56435 , n583763 , n56441 );
and ( n56443 , n54553 , n52273 );
and ( n56444 , n54321 , n52271 );
nor ( n583768 , n56443 , n56444 );
xnor ( n56446 , n583768 , n52137 );
xor ( n583770 , n583765 , n56446 );
and ( n56448 , n54893 , n52155 );
and ( n56449 , n54725 , n52153 );
nor ( n56450 , n56448 , n56449 );
xnor ( n56451 , n56450 , n52085 );
xor ( n56452 , n583770 , n56451 );
and ( n56453 , n56412 , n56452 );
and ( n583777 , n583731 , n56452 );
or ( n56455 , n583736 , n56453 , n583777 );
and ( n583779 , n53109 , n53177 );
and ( n583780 , n52934 , n53175 );
nor ( n56458 , n583779 , n583780 );
xnor ( n56459 , n56458 , n52827 );
and ( n583783 , n56455 , n56459 );
and ( n583784 , n53367 , n52978 );
and ( n56462 , n53107 , n52976 );
nor ( n56463 , n583784 , n56462 );
xnor ( n583787 , n56463 , n52680 );
and ( n583788 , n56459 , n583787 );
and ( n56466 , n56455 , n583787 );
or ( n583790 , n583783 , n583788 , n56466 );
and ( n583791 , n55841 , n51991 );
and ( n56469 , n583048 , n51989 );
nor ( n56470 , n583791 , n56469 );
xnor ( n583794 , n56470 , n51959 );
and ( n583795 , n56282 , n51936 );
and ( n56473 , n583377 , n51934 );
nor ( n583797 , n583795 , n56473 );
xnor ( n583798 , n583797 , n51941 );
and ( n56476 , n583794 , n583798 );
buf ( n583800 , n578904 );
and ( n583801 , n583800 , n51929 );
and ( n56479 , n583746 , n51927 );
nor ( n56480 , n583801 , n56479 );
not ( n56481 , n56480 );
and ( n56482 , n583798 , n56481 );
and ( n56483 , n583794 , n56481 );
or ( n56484 , n56476 , n56482 , n56483 );
and ( n56485 , n55075 , n52155 );
and ( n56486 , n55058 , n52153 );
nor ( n583810 , n56485 , n56486 );
xnor ( n56488 , n583810 , n52085 );
and ( n56489 , n56484 , n56488 );
and ( n56490 , n55528 , n52065 );
and ( n56491 , n55293 , n52063 );
nor ( n583815 , n56490 , n56491 );
xnor ( n56493 , n583815 , n52022 );
and ( n56494 , n56488 , n56493 );
and ( n56495 , n56484 , n56493 );
or ( n56496 , n56489 , n56494 , n56495 );
and ( n56497 , n54725 , n52273 );
and ( n56498 , n54553 , n52271 );
nor ( n56499 , n56497 , n56498 );
xnor ( n56500 , n56499 , n52137 );
and ( n56501 , n56496 , n56500 );
xor ( n56502 , n583599 , n56280 );
xor ( n56503 , n56502 , n583609 );
and ( n56504 , n56500 , n56503 );
and ( n583828 , n56496 , n56503 );
or ( n583829 , n56501 , n56504 , n583828 );
and ( n583830 , n54215 , n52432 );
and ( n56508 , n54055 , n52430 );
nor ( n583832 , n583830 , n56508 );
xnor ( n583833 , n583832 , n52255 );
and ( n56511 , n583829 , n583833 );
xor ( n56512 , n583612 , n56293 );
xor ( n583836 , n56512 , n56296 );
and ( n56514 , n583833 , n583836 );
and ( n56515 , n583829 , n583836 );
or ( n583839 , n56511 , n56514 , n56515 );
xor ( n583840 , n56248 , n583575 );
xor ( n56518 , n583840 , n56257 );
and ( n583842 , n583839 , n56518 );
and ( n583843 , n583765 , n56446 );
and ( n56521 , n56446 , n56451 );
and ( n583845 , n583765 , n56451 );
or ( n583846 , n583843 , n56521 , n583845 );
and ( n56524 , n53837 , n52509 );
and ( n583848 , n53639 , n52507 );
nor ( n583849 , n56524 , n583848 );
xnor ( n56527 , n583849 , n52383 );
xor ( n583851 , n583846 , n56527 );
xor ( n583852 , n56299 , n583624 );
xor ( n583853 , n583852 , n583627 );
xor ( n56531 , n583851 , n583853 );
and ( n583855 , n56518 , n56531 );
and ( n56533 , n583839 , n56531 );
or ( n56534 , n583842 , n583855 , n56533 );
and ( n56535 , n583790 , n56534 );
and ( n56536 , n52816 , n53468 );
and ( n56537 , n52818 , n53466 );
nor ( n56538 , n56536 , n56537 );
xnor ( n56539 , n56538 , n52945 );
and ( n56540 , n56534 , n56539 );
and ( n56541 , n583790 , n56539 );
or ( n56542 , n56535 , n56540 , n56541 );
and ( n56543 , n583846 , n56527 );
and ( n56544 , n56527 , n583853 );
and ( n56545 , n583846 , n583853 );
or ( n56546 , n56543 , n56544 , n56545 );
xor ( n56547 , n56097 , n583424 );
xor ( n583871 , n56547 , n583429 );
and ( n56549 , n56546 , n583871 );
xor ( n583873 , n583630 , n56311 );
xor ( n583874 , n583873 , n583637 );
and ( n56552 , n583871 , n583874 );
and ( n583876 , n56546 , n583874 );
or ( n56554 , n56549 , n56552 , n583876 );
and ( n56555 , n56542 , n56554 );
and ( n56556 , n52671 , n53683 );
and ( n56557 , n52626 , n53681 );
nor ( n56558 , n56556 , n56557 );
xnor ( n56559 , n56558 , n53118 );
and ( n56560 , n56554 , n56559 );
and ( n56561 , n56542 , n56559 );
or ( n56562 , n56555 , n56560 , n56561 );
and ( n56563 , n52533 , n53996 );
and ( n56564 , n52488 , n53994 );
nor ( n583888 , n56563 , n56564 );
xnor ( n56566 , n583888 , n53376 );
xor ( n583890 , n56272 , n56317 );
xor ( n583891 , n583890 , n56322 );
and ( n56569 , n56566 , n583891 );
xor ( n583893 , n583652 , n583654 );
xor ( n583894 , n583893 , n56334 );
and ( n56572 , n583891 , n583894 );
and ( n583896 , n56566 , n583894 );
or ( n583897 , n56569 , n56572 , n583896 );
and ( n56575 , n56562 , n583897 );
xor ( n583899 , n56325 , n583660 );
xor ( n56577 , n583899 , n56342 );
and ( n56578 , n583897 , n56577 );
and ( n56579 , n56562 , n56577 );
or ( n56580 , n56575 , n56578 , n56579 );
and ( n56581 , n52669 , n53683 );
and ( n583905 , n52671 , n53681 );
nor ( n56583 , n56581 , n583905 );
xnor ( n56584 , n56583 , n53118 );
xor ( n583908 , n583583 , n56264 );
xor ( n56586 , n583908 , n583592 );
and ( n56587 , n56584 , n56586 );
xor ( n56588 , n56546 , n583871 );
xor ( n56589 , n56588 , n583874 );
and ( n583913 , n56586 , n56589 );
and ( n583914 , n56584 , n56589 );
or ( n583915 , n56587 , n583913 , n583914 );
and ( n56593 , n52262 , n54532 );
and ( n583917 , n52194 , n54530 );
nor ( n583918 , n56593 , n583917 );
xnor ( n583919 , n583918 , n53769 );
and ( n56597 , n583915 , n583919 );
and ( n583921 , n52390 , n54414 );
and ( n56599 , n52304 , n54412 );
nor ( n583923 , n583921 , n56599 );
xnor ( n583924 , n583923 , n53650 );
and ( n56602 , n583919 , n583924 );
and ( n583926 , n583915 , n583924 );
or ( n56604 , n56597 , n56602 , n583926 );
xor ( n583928 , n583672 , n583676 );
xor ( n583929 , n583928 , n56356 );
and ( n583930 , n56604 , n583929 );
xor ( n56608 , n56364 , n583691 );
xor ( n583932 , n56608 , n583694 );
and ( n583933 , n583929 , n583932 );
and ( n583934 , n56604 , n583932 );
or ( n583935 , n583930 , n583933 , n583934 );
and ( n56613 , n56580 , n583935 );
xor ( n583937 , n56345 , n56359 );
xor ( n583938 , n583937 , n56374 );
and ( n56616 , n583935 , n583938 );
and ( n583940 , n56580 , n583938 );
or ( n583941 , n56613 , n56616 , n583940 );
xor ( n56619 , n56377 , n583710 );
xor ( n583943 , n56619 , n56390 );
and ( n583944 , n583941 , n583943 );
xor ( n56622 , n56219 , n56221 );
xor ( n583946 , n56622 , n56224 );
and ( n583947 , n583943 , n583946 );
and ( n56625 , n583941 , n583946 );
or ( n583949 , n583944 , n583947 , n56625 );
and ( n583950 , n583727 , n583949 );
xor ( n56628 , n583941 , n583943 );
xor ( n583952 , n56628 , n583946 );
and ( n583953 , n52818 , n53683 );
and ( n583954 , n52669 , n53681 );
nor ( n583955 , n583953 , n583954 );
xnor ( n56633 , n583955 , n53118 );
xor ( n583957 , n56455 , n56459 );
xor ( n583958 , n583957 , n583787 );
and ( n56636 , n56633 , n583958 );
xor ( n583960 , n583839 , n56518 );
xor ( n583961 , n583960 , n56531 );
and ( n56639 , n583958 , n583961 );
and ( n583963 , n56633 , n583961 );
or ( n583964 , n56636 , n56639 , n583963 );
and ( n56642 , n52304 , n54532 );
and ( n583966 , n52262 , n54530 );
nor ( n583967 , n56642 , n583966 );
xnor ( n56645 , n583967 , n53769 );
and ( n56646 , n583964 , n56645 );
xor ( n56647 , n583790 , n56534 );
xor ( n583971 , n56647 , n56539 );
and ( n583972 , n56645 , n583971 );
and ( n56650 , n583964 , n583971 );
or ( n583974 , n56646 , n583972 , n56650 );
and ( n583975 , n52144 , n55013 );
and ( n583976 , n52115 , n55010 );
nor ( n583977 , n583975 , n583976 );
xnor ( n56655 , n583977 , n53762 );
and ( n583979 , n583974 , n56655 );
xor ( n56657 , n56542 , n56554 );
xor ( n583981 , n56657 , n56559 );
and ( n583982 , n56655 , n583981 );
and ( n56660 , n583974 , n583981 );
or ( n583984 , n583979 , n583982 , n56660 );
and ( n583985 , n583377 , n51991 );
and ( n583986 , n55841 , n51989 );
nor ( n583987 , n583985 , n583986 );
xnor ( n56665 , n583987 , n51959 );
and ( n583989 , n583746 , n51936 );
and ( n583990 , n56282 , n51934 );
nor ( n56668 , n583989 , n583990 );
xnor ( n583992 , n56668 , n51941 );
and ( n56670 , n56665 , n583992 );
buf ( n56671 , n578905 );
and ( n56672 , n56671 , n51929 );
and ( n56673 , n583800 , n51927 );
nor ( n583997 , n56672 , n56673 );
not ( n583998 , n583997 );
and ( n56676 , n583992 , n583998 );
and ( n584000 , n56665 , n583998 );
or ( n56678 , n56670 , n56676 , n584000 );
and ( n584002 , n55293 , n52155 );
and ( n584003 , n55075 , n52153 );
nor ( n56681 , n584002 , n584003 );
xnor ( n584005 , n56681 , n52085 );
and ( n584006 , n56678 , n584005 );
and ( n584007 , n582961 , n52065 );
and ( n56685 , n55528 , n52063 );
nor ( n584009 , n584007 , n56685 );
xnor ( n584010 , n584009 , n52022 );
and ( n584011 , n584005 , n584010 );
and ( n56689 , n56678 , n584010 );
or ( n584013 , n584006 , n584011 , n56689 );
and ( n584014 , n54893 , n52273 );
and ( n56692 , n54725 , n52271 );
nor ( n584016 , n584014 , n56692 );
xnor ( n56694 , n584016 , n52137 );
and ( n56695 , n584013 , n56694 );
xor ( n56696 , n583740 , n56421 );
xor ( n56697 , n56696 , n56427 );
and ( n56698 , n56694 , n56697 );
and ( n56699 , n584013 , n56697 );
or ( n584023 , n56695 , n56698 , n56699 );
and ( n584024 , n54321 , n52432 );
and ( n56702 , n54215 , n52430 );
nor ( n584026 , n584024 , n56702 );
xnor ( n584027 , n584026 , n52255 );
and ( n56705 , n584023 , n584027 );
xor ( n584029 , n56430 , n56434 );
xor ( n584030 , n584029 , n56439 );
and ( n584031 , n584027 , n584030 );
and ( n56709 , n584023 , n584030 );
or ( n584033 , n56705 , n584031 , n56709 );
and ( n584034 , n53641 , n52978 );
and ( n56712 , n53365 , n52976 );
nor ( n584036 , n584034 , n56712 );
xnor ( n56714 , n584036 , n52680 );
and ( n56715 , n54055 , n52509 );
and ( n584039 , n53835 , n52507 );
nor ( n584040 , n56715 , n584039 );
xnor ( n56718 , n584040 , n52383 );
and ( n584042 , n56714 , n56718 );
xor ( n56720 , n56496 , n56500 );
xor ( n56721 , n56720 , n56503 );
and ( n56722 , n56718 , n56721 );
and ( n56723 , n56714 , n56721 );
or ( n56724 , n584042 , n56722 , n56723 );
and ( n56725 , n584033 , n56724 );
and ( n56726 , n53365 , n52978 );
and ( n56727 , n53367 , n52976 );
nor ( n56728 , n56726 , n56727 );
xnor ( n56729 , n56728 , n52680 );
and ( n56730 , n56724 , n56729 );
and ( n56731 , n584033 , n56729 );
or ( n56732 , n56725 , n56730 , n56731 );
and ( n56733 , n52934 , n53468 );
and ( n584057 , n52936 , n53466 );
nor ( n56735 , n56733 , n584057 );
xnor ( n56736 , n56735 , n52945 );
and ( n584060 , n53107 , n53177 );
and ( n56738 , n53109 , n53175 );
nor ( n56739 , n584060 , n56738 );
xnor ( n584063 , n56739 , n52827 );
and ( n584064 , n56736 , n584063 );
xor ( n56742 , n583829 , n583833 );
xor ( n56743 , n56742 , n583836 );
and ( n584067 , n584063 , n56743 );
and ( n584068 , n56736 , n56743 );
or ( n56746 , n584064 , n584067 , n584068 );
and ( n584070 , n56732 , n56746 );
and ( n584071 , n52936 , n53468 );
and ( n56749 , n52816 , n53466 );
nor ( n56750 , n584071 , n56749 );
xnor ( n584074 , n56750 , n52945 );
and ( n56752 , n56746 , n584074 );
and ( n584076 , n56732 , n584074 );
or ( n584077 , n584070 , n56752 , n584076 );
and ( n56755 , n52194 , n55013 );
and ( n584079 , n52144 , n55010 );
nor ( n584080 , n56755 , n584079 );
xnor ( n56758 , n584080 , n53762 );
and ( n584082 , n584077 , n56758 );
and ( n584083 , n52488 , n54414 );
and ( n56761 , n52390 , n54412 );
nor ( n584085 , n584083 , n56761 );
xnor ( n584086 , n584085 , n53650 );
and ( n584087 , n56758 , n584086 );
and ( n584088 , n584077 , n584086 );
or ( n56766 , n584082 , n584087 , n584088 );
xor ( n584090 , n583915 , n583919 );
xor ( n584091 , n584090 , n583924 );
and ( n56769 , n56766 , n584091 );
xor ( n584093 , n56566 , n583891 );
xor ( n584094 , n584093 , n583894 );
and ( n56772 , n584091 , n584094 );
and ( n584096 , n56766 , n584094 );
or ( n584097 , n56769 , n56772 , n584096 );
and ( n56775 , n583984 , n584097 );
xor ( n584099 , n56562 , n583897 );
xor ( n584100 , n584099 , n56577 );
and ( n584101 , n584097 , n584100 );
and ( n56779 , n583984 , n584100 );
or ( n584103 , n56775 , n584101 , n56779 );
xor ( n584104 , n56580 , n583935 );
xor ( n584105 , n584104 , n583938 );
and ( n56783 , n584103 , n584105 );
xor ( n584107 , n583702 , n583704 );
xor ( n56785 , n584107 , n583707 );
and ( n584109 , n584105 , n56785 );
and ( n584110 , n584103 , n56785 );
or ( n56788 , n56783 , n584109 , n584110 );
and ( n584112 , n583952 , n56788 );
xor ( n56790 , n584103 , n584105 );
xor ( n56791 , n56790 , n56785 );
and ( n56792 , n52816 , n53683 );
and ( n56793 , n52818 , n53681 );
nor ( n584117 , n56792 , n56793 );
xnor ( n584118 , n584117 , n53118 );
xor ( n56796 , n584033 , n56724 );
xor ( n584120 , n56796 , n56729 );
and ( n584121 , n584118 , n584120 );
xor ( n584122 , n56736 , n584063 );
xor ( n56800 , n584122 , n56743 );
and ( n584124 , n584120 , n56800 );
and ( n56802 , n584118 , n56800 );
or ( n584126 , n584121 , n584124 , n56802 );
and ( n584127 , n52390 , n54532 );
and ( n56805 , n52304 , n54530 );
nor ( n584129 , n584127 , n56805 );
xnor ( n56807 , n584129 , n53769 );
and ( n56808 , n584126 , n56807 );
and ( n56809 , n52533 , n54414 );
and ( n56810 , n52488 , n54412 );
nor ( n56811 , n56809 , n56810 );
xnor ( n56812 , n56811 , n53650 );
and ( n56813 , n56807 , n56812 );
and ( n56814 , n584126 , n56812 );
or ( n56815 , n56808 , n56813 , n56814 );
and ( n56816 , n53367 , n53177 );
and ( n56817 , n53107 , n53175 );
nor ( n56818 , n56816 , n56817 );
xnor ( n56819 , n56818 , n52827 );
xor ( n56820 , n56714 , n56718 );
xor ( n584144 , n56820 , n56721 );
and ( n584145 , n56819 , n584144 );
and ( n56823 , n56282 , n51991 );
and ( n584147 , n583377 , n51989 );
nor ( n584148 , n56823 , n584147 );
xnor ( n584149 , n584148 , n51959 );
and ( n56827 , n583800 , n51936 );
and ( n584151 , n583746 , n51934 );
nor ( n56829 , n56827 , n584151 );
xnor ( n584153 , n56829 , n51941 );
and ( n584154 , n584149 , n584153 );
buf ( n56832 , n578906 );
and ( n584156 , n56832 , n51929 );
and ( n56834 , n56671 , n51927 );
nor ( n584158 , n584156 , n56834 );
not ( n584159 , n584158 );
and ( n56837 , n584153 , n584159 );
and ( n584161 , n584149 , n584159 );
or ( n584162 , n584154 , n56837 , n584161 );
and ( n584163 , n583048 , n52065 );
and ( n56841 , n582961 , n52063 );
nor ( n584165 , n584163 , n56841 );
xnor ( n56843 , n584165 , n52022 );
and ( n584167 , n584162 , n56843 );
xor ( n584168 , n56665 , n583992 );
xor ( n56846 , n584168 , n583998 );
and ( n584170 , n56843 , n56846 );
and ( n56848 , n584162 , n56846 );
or ( n56849 , n584167 , n584170 , n56848 );
and ( n56850 , n55058 , n52273 );
and ( n584174 , n54893 , n52271 );
nor ( n584175 , n56850 , n584174 );
xnor ( n56853 , n584175 , n52137 );
and ( n584177 , n56849 , n56853 );
xor ( n584178 , n583794 , n583798 );
xor ( n584179 , n584178 , n56481 );
and ( n584180 , n56853 , n584179 );
and ( n56858 , n56849 , n584179 );
or ( n584182 , n584177 , n584180 , n56858 );
and ( n584183 , n54553 , n52432 );
and ( n56861 , n54321 , n52430 );
nor ( n584185 , n584183 , n56861 );
xnor ( n584186 , n584185 , n52255 );
and ( n56864 , n584182 , n584186 );
xor ( n56865 , n56484 , n56488 );
xor ( n584189 , n56865 , n56493 );
and ( n56867 , n584186 , n584189 );
and ( n56868 , n584182 , n584189 );
or ( n584192 , n56864 , n56867 , n56868 );
and ( n584193 , n53837 , n52707 );
and ( n56871 , n53639 , n52705 );
nor ( n584195 , n584193 , n56871 );
xnor ( n584196 , n584195 , n52526 );
xor ( n56874 , n584192 , n584196 );
xor ( n584198 , n584023 , n584027 );
xor ( n56876 , n584198 , n584030 );
xor ( n56877 , n56874 , n56876 );
and ( n56878 , n584144 , n56877 );
and ( n56879 , n56819 , n56877 );
or ( n56880 , n584145 , n56878 , n56879 );
and ( n56881 , n52669 , n53996 );
and ( n56882 , n52671 , n53994 );
nor ( n56883 , n56881 , n56882 );
xnor ( n584207 , n56883 , n53376 );
and ( n56885 , n56880 , n584207 );
and ( n584209 , n53639 , n52978 );
and ( n584210 , n53641 , n52976 );
nor ( n56888 , n584209 , n584210 );
xnor ( n56889 , n56888 , n52680 );
and ( n584213 , n53835 , n52707 );
and ( n584214 , n53837 , n52705 );
nor ( n56892 , n584213 , n584214 );
xnor ( n56893 , n56892 , n52526 );
and ( n584217 , n56889 , n56893 );
xor ( n56895 , n584182 , n584186 );
xor ( n56896 , n56895 , n584189 );
and ( n584220 , n56893 , n56896 );
and ( n56898 , n56889 , n56896 );
or ( n584222 , n584217 , n584220 , n56898 );
and ( n584223 , n583746 , n51991 );
and ( n56901 , n56282 , n51989 );
nor ( n584225 , n584223 , n56901 );
xnor ( n584226 , n584225 , n51959 );
and ( n584227 , n56671 , n51936 );
and ( n584228 , n583800 , n51934 );
nor ( n56906 , n584227 , n584228 );
xnor ( n584230 , n56906 , n51941 );
and ( n584231 , n584226 , n584230 );
buf ( n56909 , n578907 );
and ( n584233 , n56909 , n51929 );
and ( n584234 , n56832 , n51927 );
nor ( n56912 , n584233 , n584234 );
not ( n584236 , n56912 );
and ( n584237 , n584230 , n584236 );
and ( n56915 , n584226 , n584236 );
or ( n56916 , n584231 , n584237 , n56915 );
and ( n56917 , n55841 , n52065 );
and ( n584241 , n583048 , n52063 );
nor ( n584242 , n56917 , n584241 );
xnor ( n584243 , n584242 , n52022 );
and ( n56921 , n56916 , n584243 );
xor ( n584245 , n584149 , n584153 );
xor ( n584246 , n584245 , n584159 );
and ( n56924 , n584243 , n584246 );
and ( n584248 , n56916 , n584246 );
or ( n584249 , n56921 , n56924 , n584248 );
and ( n56927 , n55075 , n52273 );
and ( n584251 , n55058 , n52271 );
nor ( n584252 , n56927 , n584251 );
xnor ( n56930 , n584252 , n52137 );
and ( n56931 , n584249 , n56930 );
and ( n584255 , n55528 , n52155 );
and ( n584256 , n55293 , n52153 );
nor ( n56934 , n584255 , n584256 );
xnor ( n584258 , n56934 , n52085 );
and ( n584259 , n56930 , n584258 );
and ( n56937 , n584249 , n584258 );
or ( n584261 , n56931 , n584259 , n56937 );
and ( n584262 , n54725 , n52432 );
and ( n56940 , n54553 , n52430 );
nor ( n584264 , n584262 , n56940 );
xnor ( n584265 , n584264 , n52255 );
and ( n56943 , n584261 , n584265 );
xor ( n584267 , n56678 , n584005 );
xor ( n56945 , n584267 , n584010 );
and ( n56946 , n584265 , n56945 );
and ( n56947 , n584261 , n56945 );
or ( n56948 , n56943 , n56946 , n56947 );
and ( n56949 , n54215 , n52509 );
and ( n56950 , n54055 , n52507 );
nor ( n56951 , n56949 , n56950 );
xnor ( n56952 , n56951 , n52383 );
and ( n584276 , n56948 , n56952 );
xor ( n584277 , n584013 , n56694 );
xor ( n56955 , n584277 , n56697 );
and ( n584279 , n56952 , n56955 );
and ( n584280 , n56948 , n56955 );
or ( n584281 , n584276 , n584279 , n584280 );
and ( n584282 , n584222 , n584281 );
and ( n56960 , n53109 , n53468 );
and ( n584284 , n52934 , n53466 );
nor ( n584285 , n56960 , n584284 );
xnor ( n56963 , n584285 , n52945 );
and ( n584287 , n584281 , n56963 );
and ( n584288 , n584222 , n56963 );
or ( n56966 , n584282 , n584287 , n584288 );
and ( n584290 , n584192 , n584196 );
and ( n584291 , n584196 , n56876 );
and ( n56969 , n584192 , n56876 );
or ( n56970 , n584290 , n584291 , n56969 );
xor ( n56971 , n56966 , n56970 );
xor ( n584295 , n583731 , n56412 );
xor ( n584296 , n584295 , n56452 );
xor ( n584297 , n56971 , n584296 );
and ( n584298 , n584207 , n584297 );
and ( n56976 , n56880 , n584297 );
or ( n584300 , n56885 , n584298 , n56976 );
and ( n584301 , n52262 , n55013 );
and ( n584302 , n52194 , n55010 );
nor ( n584303 , n584301 , n584302 );
xnor ( n56981 , n584303 , n53762 );
and ( n584305 , n584300 , n56981 );
xor ( n584306 , n56633 , n583958 );
xor ( n56984 , n584306 , n583961 );
and ( n584308 , n56981 , n56984 );
and ( n584309 , n584300 , n56984 );
or ( n56987 , n584305 , n584308 , n584309 );
and ( n584311 , n56815 , n56987 );
xor ( n584312 , n583964 , n56645 );
xor ( n56990 , n584312 , n583971 );
and ( n56991 , n56987 , n56990 );
and ( n56992 , n56815 , n56990 );
or ( n584316 , n584311 , n56991 , n56992 );
and ( n584317 , n56966 , n56970 );
and ( n56995 , n56970 , n584296 );
and ( n584319 , n56966 , n584296 );
or ( n584320 , n584317 , n56995 , n584319 );
and ( n56998 , n52671 , n53996 );
and ( n584322 , n52626 , n53994 );
nor ( n584323 , n56998 , n584322 );
xnor ( n584324 , n584323 , n53376 );
and ( n584325 , n584320 , n584324 );
xor ( n57003 , n56732 , n56746 );
xor ( n584327 , n57003 , n584074 );
and ( n584328 , n584324 , n584327 );
and ( n57006 , n584320 , n584327 );
or ( n584330 , n584325 , n584328 , n57006 );
and ( n584331 , n52626 , n53996 );
and ( n57009 , n52533 , n53994 );
nor ( n584333 , n584331 , n57009 );
xnor ( n584334 , n584333 , n53376 );
and ( n57012 , n584330 , n584334 );
xor ( n57013 , n56584 , n56586 );
xor ( n57014 , n57013 , n56589 );
and ( n584338 , n584334 , n57014 );
and ( n584339 , n584330 , n57014 );
or ( n57017 , n57012 , n584338 , n584339 );
and ( n584341 , n584316 , n57017 );
xor ( n57019 , n583974 , n56655 );
xor ( n57020 , n57019 , n583981 );
and ( n57021 , n57017 , n57020 );
and ( n57022 , n584316 , n57020 );
or ( n57023 , n584341 , n57021 , n57022 );
xor ( n57024 , n583984 , n584097 );
xor ( n57025 , n57024 , n584100 );
and ( n57026 , n57023 , n57025 );
xor ( n57027 , n56604 , n583929 );
xor ( n584351 , n57027 , n583932 );
and ( n57029 , n57025 , n584351 );
and ( n57030 , n57023 , n584351 );
or ( n57031 , n57026 , n57029 , n57030 );
and ( n57032 , n56791 , n57031 );
xor ( n57033 , n57023 , n57025 );
xor ( n57034 , n57033 , n584351 );
and ( n584358 , n53641 , n53177 );
and ( n584359 , n53365 , n53175 );
nor ( n57037 , n584358 , n584359 );
xnor ( n57038 , n57037 , n52827 );
and ( n57039 , n54055 , n52707 );
and ( n57040 , n53835 , n52705 );
nor ( n584364 , n57039 , n57040 );
xnor ( n57042 , n584364 , n52526 );
and ( n57043 , n57038 , n57042 );
xor ( n57044 , n584261 , n584265 );
xor ( n57045 , n57044 , n56945 );
and ( n584369 , n57042 , n57045 );
and ( n584370 , n57038 , n57045 );
or ( n57048 , n57043 , n584369 , n584370 );
and ( n57049 , n583800 , n51991 );
and ( n57050 , n583746 , n51989 );
nor ( n57051 , n57049 , n57050 );
xnor ( n57052 , n57051 , n51959 );
and ( n584376 , n56832 , n51936 );
and ( n57054 , n56671 , n51934 );
nor ( n584378 , n584376 , n57054 );
xnor ( n584379 , n584378 , n51941 );
and ( n57057 , n57052 , n584379 );
buf ( n57058 , n578908 );
and ( n57059 , n57058 , n51929 );
and ( n57060 , n56909 , n51927 );
nor ( n57061 , n57059 , n57060 );
not ( n584385 , n57061 );
and ( n584386 , n584379 , n584385 );
and ( n57064 , n57052 , n584385 );
or ( n584388 , n57057 , n584386 , n57064 );
and ( n57066 , n583377 , n52065 );
and ( n57067 , n55841 , n52063 );
nor ( n57068 , n57066 , n57067 );
xnor ( n57069 , n57068 , n52022 );
and ( n57070 , n584388 , n57069 );
xor ( n57071 , n584226 , n584230 );
xor ( n57072 , n57071 , n584236 );
and ( n584396 , n57069 , n57072 );
and ( n57074 , n584388 , n57072 );
or ( n584398 , n57070 , n584396 , n57074 );
and ( n584399 , n55293 , n52273 );
and ( n57077 , n55075 , n52271 );
nor ( n584401 , n584399 , n57077 );
xnor ( n57079 , n584401 , n52137 );
and ( n57080 , n584398 , n57079 );
and ( n57081 , n582961 , n52155 );
and ( n584405 , n55528 , n52153 );
nor ( n57083 , n57081 , n584405 );
xnor ( n584407 , n57083 , n52085 );
and ( n584408 , n57079 , n584407 );
and ( n57086 , n584398 , n584407 );
or ( n57087 , n57080 , n584408 , n57086 );
and ( n584411 , n54893 , n52432 );
and ( n57089 , n54725 , n52430 );
nor ( n584413 , n584411 , n57089 );
xnor ( n57091 , n584413 , n52255 );
and ( n584415 , n57087 , n57091 );
xor ( n584416 , n584162 , n56843 );
xor ( n57094 , n584416 , n56846 );
and ( n584418 , n57091 , n57094 );
and ( n584419 , n57087 , n57094 );
or ( n584420 , n584415 , n584418 , n584419 );
and ( n584421 , n54321 , n52509 );
and ( n57099 , n54215 , n52507 );
nor ( n584423 , n584421 , n57099 );
xnor ( n57101 , n584423 , n52383 );
and ( n584425 , n584420 , n57101 );
xor ( n57103 , n56849 , n56853 );
xor ( n57104 , n57103 , n584179 );
and ( n584428 , n57101 , n57104 );
and ( n57106 , n584420 , n57104 );
or ( n584430 , n584425 , n584428 , n57106 );
and ( n584431 , n57048 , n584430 );
and ( n57109 , n53365 , n53177 );
and ( n584433 , n53367 , n53175 );
nor ( n584434 , n57109 , n584433 );
xnor ( n57112 , n584434 , n52827 );
and ( n57113 , n584430 , n57112 );
and ( n57114 , n57048 , n57112 );
or ( n57115 , n584431 , n57113 , n57114 );
and ( n584439 , n52934 , n53683 );
and ( n584440 , n52936 , n53681 );
nor ( n57118 , n584439 , n584440 );
xnor ( n584442 , n57118 , n53118 );
and ( n584443 , n53107 , n53468 );
and ( n57121 , n53109 , n53466 );
nor ( n584445 , n584443 , n57121 );
xnor ( n57123 , n584445 , n52945 );
and ( n584447 , n584442 , n57123 );
xor ( n57125 , n56948 , n56952 );
xor ( n57126 , n57125 , n56955 );
and ( n584450 , n57123 , n57126 );
and ( n57128 , n584442 , n57126 );
or ( n584452 , n584447 , n584450 , n57128 );
and ( n584453 , n57115 , n584452 );
and ( n57131 , n52936 , n53683 );
and ( n584455 , n52816 , n53681 );
nor ( n584456 , n57131 , n584455 );
xnor ( n57134 , n584456 , n53118 );
and ( n584458 , n584452 , n57134 );
and ( n584459 , n57115 , n57134 );
or ( n57137 , n584453 , n584458 , n584459 );
and ( n584461 , n52304 , n55013 );
and ( n57139 , n52262 , n55010 );
nor ( n57140 , n584461 , n57139 );
xnor ( n57141 , n57140 , n53762 );
and ( n57142 , n57137 , n57141 );
and ( n584466 , n52626 , n54414 );
and ( n584467 , n52533 , n54412 );
nor ( n57145 , n584466 , n584467 );
xnor ( n584469 , n57145 , n53650 );
and ( n57147 , n57141 , n584469 );
and ( n57148 , n57137 , n584469 );
or ( n57149 , n57142 , n57147 , n57148 );
and ( n57150 , n52818 , n53996 );
and ( n57151 , n52669 , n53994 );
nor ( n57152 , n57150 , n57151 );
xnor ( n57153 , n57152 , n53376 );
xor ( n57154 , n584222 , n584281 );
xor ( n57155 , n57154 , n56963 );
and ( n57156 , n57153 , n57155 );
xor ( n584480 , n56819 , n584144 );
xor ( n57158 , n584480 , n56877 );
and ( n57159 , n57155 , n57158 );
and ( n57160 , n57153 , n57158 );
or ( n57161 , n57156 , n57159 , n57160 );
and ( n57162 , n52488 , n54532 );
and ( n57163 , n52390 , n54530 );
nor ( n57164 , n57162 , n57163 );
xnor ( n57165 , n57164 , n53769 );
and ( n57166 , n57161 , n57165 );
xor ( n57167 , n584118 , n584120 );
xor ( n57168 , n57167 , n56800 );
and ( n57169 , n57165 , n57168 );
and ( n57170 , n57161 , n57168 );
or ( n57171 , n57166 , n57169 , n57170 );
and ( n57172 , n57149 , n57171 );
xor ( n57173 , n584320 , n584324 );
xor ( n57174 , n57173 , n584327 );
and ( n57175 , n57171 , n57174 );
and ( n57176 , n57149 , n57174 );
or ( n57177 , n57172 , n57175 , n57176 );
xor ( n57178 , n584077 , n56758 );
xor ( n57179 , n57178 , n584086 );
and ( n57180 , n57177 , n57179 );
xor ( n57181 , n584330 , n584334 );
xor ( n57182 , n57181 , n57014 );
and ( n57183 , n57179 , n57182 );
and ( n584507 , n57177 , n57182 );
or ( n57185 , n57180 , n57183 , n584507 );
xor ( n57186 , n584316 , n57017 );
xor ( n584510 , n57186 , n57020 );
and ( n584511 , n57185 , n584510 );
xor ( n57189 , n56766 , n584091 );
xor ( n584513 , n57189 , n584094 );
and ( n57191 , n584510 , n584513 );
and ( n57192 , n57185 , n584513 );
or ( n57193 , n584511 , n57191 , n57192 );
and ( n57194 , n57034 , n57193 );
xor ( n57195 , n57185 , n584510 );
xor ( n57196 , n57195 , n584513 );
and ( n57197 , n583746 , n52065 );
and ( n57198 , n56282 , n52063 );
nor ( n57199 , n57197 , n57198 );
xnor ( n57200 , n57199 , n52022 );
and ( n57201 , n56909 , n51936 );
and ( n57202 , n56832 , n51934 );
nor ( n57203 , n57201 , n57202 );
xnor ( n57204 , n57203 , n51941 );
and ( n57205 , n57200 , n57204 );
buf ( n584529 , n578909 );
and ( n584530 , n584529 , n51929 );
and ( n57208 , n57058 , n51927 );
nor ( n584532 , n584530 , n57208 );
not ( n57210 , n584532 );
and ( n57211 , n57204 , n57210 );
and ( n57212 , n57200 , n57210 );
or ( n57213 , n57205 , n57211 , n57212 );
and ( n57214 , n56282 , n52065 );
and ( n57215 , n583377 , n52063 );
nor ( n57216 , n57214 , n57215 );
xnor ( n584540 , n57216 , n52022 );
and ( n57218 , n57213 , n584540 );
xor ( n57219 , n57052 , n584379 );
xor ( n57220 , n57219 , n584385 );
and ( n584544 , n584540 , n57220 );
and ( n57222 , n57213 , n57220 );
or ( n57223 , n57218 , n584544 , n57222 );
and ( n57224 , n55528 , n52273 );
and ( n57225 , n55293 , n52271 );
nor ( n584549 , n57224 , n57225 );
xnor ( n584550 , n584549 , n52137 );
and ( n57228 , n57223 , n584550 );
and ( n584552 , n583048 , n52155 );
and ( n584553 , n582961 , n52153 );
nor ( n57231 , n584552 , n584553 );
xnor ( n584555 , n57231 , n52085 );
and ( n584556 , n584550 , n584555 );
and ( n57234 , n57223 , n584555 );
or ( n57235 , n57228 , n584556 , n57234 );
and ( n584559 , n55058 , n52432 );
and ( n584560 , n54893 , n52430 );
nor ( n57238 , n584559 , n584560 );
xnor ( n57239 , n57238 , n52255 );
and ( n584563 , n57235 , n57239 );
xor ( n57241 , n56916 , n584243 );
xor ( n57242 , n57241 , n584246 );
and ( n584566 , n57239 , n57242 );
and ( n57244 , n57235 , n57242 );
or ( n584568 , n584563 , n584566 , n57244 );
and ( n584569 , n54553 , n52509 );
and ( n57247 , n54321 , n52507 );
nor ( n57248 , n584569 , n57247 );
xnor ( n57249 , n57248 , n52383 );
and ( n57250 , n584568 , n57249 );
xor ( n57251 , n584249 , n56930 );
xor ( n57252 , n57251 , n584258 );
and ( n57253 , n57249 , n57252 );
and ( n57254 , n584568 , n57252 );
or ( n57255 , n57250 , n57253 , n57254 );
and ( n57256 , n53837 , n52978 );
and ( n57257 , n53639 , n52976 );
nor ( n57258 , n57256 , n57257 );
xnor ( n57259 , n57258 , n52680 );
and ( n57260 , n57255 , n57259 );
xor ( n584584 , n584420 , n57101 );
xor ( n584585 , n584584 , n57104 );
and ( n57263 , n57259 , n584585 );
and ( n584587 , n57255 , n584585 );
or ( n584588 , n57260 , n57263 , n584587 );
xor ( n57266 , n57048 , n584430 );
xor ( n584590 , n57266 , n57112 );
and ( n584591 , n584588 , n584590 );
xor ( n57269 , n56889 , n56893 );
xor ( n57270 , n57269 , n56896 );
and ( n584594 , n584590 , n57270 );
and ( n584595 , n584588 , n57270 );
or ( n57273 , n584591 , n584594 , n584595 );
and ( n57274 , n56832 , n51991 );
and ( n584598 , n56671 , n51989 );
nor ( n57276 , n57274 , n584598 );
xnor ( n57277 , n57276 , n51959 );
and ( n57278 , n57058 , n51936 );
and ( n57279 , n56909 , n51934 );
nor ( n57280 , n57278 , n57279 );
xnor ( n57281 , n57280 , n51941 );
and ( n57282 , n57277 , n57281 );
buf ( n57283 , n578910 );
and ( n57284 , n57283 , n51929 );
and ( n57285 , n584529 , n51927 );
nor ( n57286 , n57284 , n57285 );
not ( n57287 , n57286 );
and ( n57288 , n57281 , n57287 );
and ( n57289 , n57277 , n57287 );
or ( n57290 , n57282 , n57288 , n57289 );
and ( n57291 , n583377 , n52155 );
and ( n57292 , n55841 , n52153 );
nor ( n57293 , n57291 , n57292 );
xnor ( n57294 , n57293 , n52085 );
and ( n57295 , n57290 , n57294 );
and ( n57296 , n56671 , n51991 );
and ( n57297 , n583800 , n51989 );
nor ( n57298 , n57296 , n57297 );
xnor ( n57299 , n57298 , n51959 );
and ( n57300 , n57294 , n57299 );
and ( n57301 , n57290 , n57299 );
or ( n584625 , n57295 , n57300 , n57301 );
and ( n584626 , n582961 , n52273 );
and ( n57304 , n55528 , n52271 );
nor ( n584628 , n584626 , n57304 );
xnor ( n57306 , n584628 , n52137 );
and ( n57307 , n584625 , n57306 );
and ( n57308 , n55841 , n52155 );
and ( n584632 , n583048 , n52153 );
nor ( n584633 , n57308 , n584632 );
xnor ( n57311 , n584633 , n52085 );
and ( n584635 , n57306 , n57311 );
and ( n57313 , n584625 , n57311 );
or ( n57314 , n57307 , n584635 , n57313 );
and ( n57315 , n55075 , n52432 );
and ( n584639 , n55058 , n52430 );
nor ( n57317 , n57315 , n584639 );
xnor ( n584641 , n57317 , n52255 );
and ( n584642 , n57314 , n584641 );
xor ( n57320 , n584388 , n57069 );
xor ( n584644 , n57320 , n57072 );
and ( n584645 , n584641 , n584644 );
and ( n57323 , n57314 , n584644 );
or ( n57324 , n584642 , n584645 , n57323 );
and ( n584648 , n54725 , n52509 );
and ( n584649 , n54553 , n52507 );
nor ( n57327 , n584648 , n584649 );
xnor ( n57328 , n57327 , n52383 );
and ( n584652 , n57324 , n57328 );
xor ( n584653 , n584398 , n57079 );
xor ( n57331 , n584653 , n584407 );
and ( n57332 , n57328 , n57331 );
and ( n57333 , n57324 , n57331 );
or ( n584657 , n584652 , n57332 , n57333 );
and ( n57335 , n53835 , n52978 );
and ( n584659 , n53837 , n52976 );
nor ( n57337 , n57335 , n584659 );
xnor ( n584661 , n57337 , n52680 );
and ( n57339 , n584657 , n584661 );
xor ( n584663 , n584568 , n57249 );
xor ( n57341 , n584663 , n57252 );
and ( n57342 , n584661 , n57341 );
and ( n57343 , n584657 , n57341 );
or ( n584667 , n57339 , n57342 , n57343 );
and ( n57345 , n53639 , n53177 );
and ( n584669 , n53641 , n53175 );
nor ( n57347 , n57345 , n584669 );
xnor ( n584671 , n57347 , n52827 );
and ( n57349 , n54215 , n52707 );
and ( n584673 , n54055 , n52705 );
nor ( n57351 , n57349 , n584673 );
xnor ( n584675 , n57351 , n52526 );
and ( n57353 , n584671 , n584675 );
xor ( n57354 , n57087 , n57091 );
xor ( n57355 , n57354 , n57094 );
and ( n57356 , n584675 , n57355 );
and ( n584680 , n584671 , n57355 );
or ( n57358 , n57353 , n57356 , n584680 );
and ( n584682 , n584667 , n57358 );
and ( n57360 , n53367 , n53468 );
and ( n584684 , n53107 , n53466 );
nor ( n57362 , n57360 , n584684 );
xnor ( n57363 , n57362 , n52945 );
and ( n57364 , n57358 , n57363 );
and ( n57365 , n584667 , n57363 );
or ( n584689 , n584682 , n57364 , n57365 );
and ( n57367 , n52816 , n53996 );
and ( n57368 , n52818 , n53994 );
nor ( n584692 , n57367 , n57368 );
xnor ( n57370 , n584692 , n53376 );
and ( n57371 , n584689 , n57370 );
xor ( n57372 , n584442 , n57123 );
xor ( n57373 , n57372 , n57126 );
and ( n584697 , n57370 , n57373 );
and ( n584698 , n584689 , n57373 );
or ( n584699 , n57371 , n584697 , n584698 );
and ( n57377 , n57273 , n584699 );
and ( n584701 , n52671 , n54414 );
and ( n57379 , n52626 , n54412 );
nor ( n584703 , n584701 , n57379 );
xnor ( n584704 , n584703 , n53650 );
and ( n584705 , n584699 , n584704 );
and ( n584706 , n57273 , n584704 );
or ( n57384 , n57377 , n584705 , n584706 );
and ( n584708 , n52390 , n55013 );
and ( n57386 , n52304 , n55010 );
nor ( n57387 , n584708 , n57386 );
xnor ( n584711 , n57387 , n53762 );
and ( n57389 , n52533 , n54532 );
and ( n57390 , n52488 , n54530 );
nor ( n57391 , n57389 , n57390 );
xnor ( n57392 , n57391 , n53769 );
and ( n584716 , n584711 , n57392 );
xor ( n57394 , n57115 , n584452 );
xor ( n584718 , n57394 , n57134 );
and ( n584719 , n57392 , n584718 );
and ( n57397 , n584711 , n584718 );
or ( n57398 , n584716 , n584719 , n57397 );
and ( n57399 , n57384 , n57398 );
xor ( n57400 , n56880 , n584207 );
xor ( n57401 , n57400 , n584297 );
and ( n57402 , n57398 , n57401 );
and ( n57403 , n57384 , n57401 );
or ( n57404 , n57399 , n57402 , n57403 );
xor ( n57405 , n584126 , n56807 );
xor ( n584729 , n57405 , n56812 );
and ( n57407 , n57404 , n584729 );
xor ( n57408 , n584300 , n56981 );
xor ( n584732 , n57408 , n56984 );
and ( n584733 , n584729 , n584732 );
and ( n57411 , n57404 , n584732 );
or ( n584735 , n57407 , n584733 , n57411 );
xor ( n584736 , n56815 , n56987 );
xor ( n57414 , n584736 , n56990 );
and ( n584738 , n584735 , n57414 );
xor ( n584739 , n57177 , n57179 );
xor ( n57417 , n584739 , n57182 );
and ( n57418 , n57414 , n57417 );
and ( n584742 , n584735 , n57417 );
or ( n584743 , n584738 , n57418 , n584742 );
and ( n57421 , n57196 , n584743 );
xor ( n57422 , n584735 , n57414 );
xor ( n57423 , n57422 , n57417 );
and ( n57424 , n53109 , n53683 );
and ( n57425 , n52934 , n53681 );
nor ( n584749 , n57424 , n57425 );
xnor ( n584750 , n584749 , n53118 );
xor ( n57428 , n57038 , n57042 );
xor ( n584752 , n57428 , n57045 );
and ( n57430 , n584750 , n584752 );
xor ( n57431 , n57255 , n57259 );
xor ( n57432 , n57431 , n584585 );
and ( n57433 , n584752 , n57432 );
and ( n584757 , n584750 , n57432 );
or ( n57435 , n57430 , n57433 , n584757 );
and ( n584759 , n52669 , n54414 );
and ( n584760 , n52671 , n54412 );
nor ( n57438 , n584759 , n584760 );
xnor ( n584762 , n57438 , n53650 );
and ( n584763 , n57435 , n584762 );
xor ( n57441 , n584588 , n584590 );
xor ( n57442 , n57441 , n57270 );
and ( n584766 , n584762 , n57442 );
and ( n584767 , n57435 , n57442 );
or ( n57445 , n584763 , n584766 , n584767 );
xor ( n57446 , n57273 , n584699 );
xor ( n584770 , n57446 , n584704 );
and ( n57448 , n57445 , n584770 );
xor ( n584772 , n57153 , n57155 );
xor ( n584773 , n584772 , n57158 );
and ( n57451 , n584770 , n584773 );
and ( n584775 , n57445 , n584773 );
or ( n57453 , n57448 , n57451 , n584775 );
xor ( n584777 , n57137 , n57141 );
xor ( n57455 , n584777 , n584469 );
and ( n57456 , n57453 , n57455 );
xor ( n57457 , n57161 , n57165 );
xor ( n584781 , n57457 , n57168 );
and ( n584782 , n57455 , n584781 );
and ( n57460 , n57453 , n584781 );
or ( n57461 , n57456 , n584782 , n57460 );
xor ( n584785 , n57149 , n57171 );
xor ( n584786 , n584785 , n57174 );
and ( n57464 , n57461 , n584786 );
xor ( n57465 , n57404 , n584729 );
xor ( n584789 , n57465 , n584732 );
and ( n57467 , n584786 , n584789 );
and ( n57468 , n57461 , n584789 );
or ( n57469 , n57464 , n57467 , n57468 );
and ( n57470 , n57423 , n57469 );
xor ( n584794 , n57461 , n584786 );
xor ( n57472 , n584794 , n584789 );
and ( n584796 , n57058 , n51991 );
and ( n584797 , n56909 , n51989 );
nor ( n57475 , n584796 , n584797 );
xnor ( n584799 , n57475 , n51959 );
and ( n57477 , n57283 , n51936 );
and ( n57478 , n584529 , n51934 );
nor ( n584802 , n57477 , n57478 );
xnor ( n57480 , n584802 , n51941 );
and ( n584804 , n584799 , n57480 );
buf ( n57482 , n578912 );
and ( n584806 , n57482 , n51929 );
buf ( n57484 , n578911 );
and ( n57485 , n57484 , n51927 );
nor ( n584809 , n584806 , n57485 );
not ( n57487 , n584809 );
and ( n584811 , n57480 , n57487 );
and ( n57489 , n584799 , n57487 );
or ( n584813 , n584804 , n584811 , n57489 );
and ( n57491 , n583746 , n52155 );
and ( n57492 , n56282 , n52153 );
nor ( n584816 , n57491 , n57492 );
xnor ( n584817 , n584816 , n52085 );
and ( n57495 , n584813 , n584817 );
and ( n584819 , n56909 , n51991 );
and ( n57497 , n56832 , n51989 );
nor ( n57498 , n584819 , n57497 );
xnor ( n584822 , n57498 , n51959 );
and ( n584823 , n584529 , n51936 );
and ( n584824 , n57058 , n51934 );
nor ( n57502 , n584823 , n584824 );
xnor ( n584826 , n57502 , n51941 );
xor ( n584827 , n584822 , n584826 );
and ( n57505 , n57484 , n51929 );
and ( n57506 , n57283 , n51927 );
nor ( n57507 , n57505 , n57506 );
not ( n57508 , n57507 );
xor ( n57509 , n584827 , n57508 );
and ( n57510 , n584817 , n57509 );
and ( n57511 , n584813 , n57509 );
or ( n584835 , n57495 , n57510 , n57511 );
and ( n57513 , n55841 , n52273 );
and ( n57514 , n583048 , n52271 );
nor ( n584838 , n57513 , n57514 );
xnor ( n584839 , n584838 , n52137 );
and ( n57517 , n584835 , n584839 );
and ( n584841 , n56282 , n52155 );
and ( n584842 , n583377 , n52153 );
nor ( n57520 , n584841 , n584842 );
xnor ( n584844 , n57520 , n52085 );
and ( n584845 , n584839 , n584844 );
and ( n57523 , n584835 , n584844 );
or ( n584847 , n57517 , n584845 , n57523 );
and ( n57525 , n55528 , n52432 );
and ( n57526 , n55293 , n52430 );
nor ( n57527 , n57525 , n57526 );
xnor ( n57528 , n57527 , n52255 );
and ( n57529 , n584847 , n57528 );
xor ( n57530 , n57290 , n57294 );
xor ( n57531 , n57530 , n57299 );
and ( n57532 , n57528 , n57531 );
and ( n584856 , n584847 , n57531 );
or ( n584857 , n57529 , n57532 , n584856 );
and ( n584858 , n55058 , n52509 );
and ( n57536 , n54893 , n52507 );
nor ( n584860 , n584858 , n57536 );
xnor ( n584861 , n584860 , n52383 );
and ( n584862 , n584857 , n584861 );
xor ( n584863 , n584625 , n57306 );
xor ( n57541 , n584863 , n57311 );
and ( n584865 , n584861 , n57541 );
and ( n584866 , n584857 , n57541 );
or ( n57544 , n584862 , n584865 , n584866 );
and ( n584868 , n54553 , n52707 );
and ( n584869 , n54321 , n52705 );
nor ( n57547 , n584868 , n584869 );
xnor ( n584871 , n57547 , n52526 );
and ( n584872 , n57544 , n584871 );
xor ( n57550 , n57314 , n584641 );
xor ( n584874 , n57550 , n584644 );
and ( n584875 , n584871 , n584874 );
and ( n584876 , n57544 , n584874 );
or ( n57554 , n584872 , n584875 , n584876 );
and ( n584878 , n53641 , n53468 );
and ( n584879 , n53365 , n53466 );
nor ( n584880 , n584878 , n584879 );
xnor ( n584881 , n584880 , n52945 );
and ( n57559 , n57554 , n584881 );
and ( n584883 , n54055 , n52978 );
and ( n584884 , n53835 , n52976 );
nor ( n57562 , n584883 , n584884 );
xnor ( n584886 , n57562 , n52680 );
and ( n584887 , n584881 , n584886 );
and ( n57565 , n57554 , n584886 );
or ( n584889 , n57559 , n584887 , n57565 );
and ( n584890 , n584822 , n584826 );
and ( n57568 , n584826 , n57508 );
and ( n584892 , n584822 , n57508 );
or ( n57570 , n584890 , n57568 , n584892 );
and ( n584894 , n583800 , n52065 );
and ( n584895 , n583746 , n52063 );
nor ( n57573 , n584894 , n584895 );
xnor ( n584897 , n57573 , n52022 );
and ( n584898 , n57570 , n584897 );
xor ( n584899 , n57277 , n57281 );
xor ( n584900 , n584899 , n57287 );
and ( n57578 , n584897 , n584900 );
and ( n584902 , n57570 , n584900 );
or ( n584903 , n584898 , n57578 , n584902 );
and ( n57581 , n583048 , n52273 );
and ( n57582 , n582961 , n52271 );
nor ( n57583 , n57581 , n57582 );
xnor ( n57584 , n57583 , n52137 );
and ( n57585 , n584903 , n57584 );
xor ( n584909 , n57200 , n57204 );
xor ( n584910 , n584909 , n57210 );
and ( n57588 , n57584 , n584910 );
and ( n584912 , n584903 , n584910 );
or ( n57590 , n57585 , n57588 , n584912 );
and ( n584914 , n55293 , n52432 );
and ( n57592 , n55075 , n52430 );
nor ( n584916 , n584914 , n57592 );
xnor ( n584917 , n584916 , n52255 );
and ( n57595 , n57590 , n584917 );
xor ( n584919 , n57213 , n584540 );
xor ( n584920 , n584919 , n57220 );
and ( n584921 , n584917 , n584920 );
and ( n57599 , n57590 , n584920 );
or ( n584923 , n57595 , n584921 , n57599 );
and ( n57601 , n54893 , n52509 );
and ( n584925 , n54725 , n52507 );
nor ( n584926 , n57601 , n584925 );
xnor ( n57604 , n584926 , n52383 );
and ( n584928 , n584923 , n57604 );
xor ( n57606 , n57223 , n584550 );
xor ( n584930 , n57606 , n584555 );
and ( n57608 , n57604 , n584930 );
and ( n57609 , n584923 , n584930 );
or ( n57610 , n584928 , n57608 , n57609 );
and ( n57611 , n54321 , n52707 );
and ( n584935 , n54215 , n52705 );
nor ( n57613 , n57611 , n584935 );
xnor ( n57614 , n57613 , n52526 );
and ( n57615 , n57610 , n57614 );
xor ( n57616 , n57235 , n57239 );
xor ( n57617 , n57616 , n57242 );
and ( n57618 , n57614 , n57617 );
and ( n57619 , n57610 , n57617 );
or ( n57620 , n57615 , n57618 , n57619 );
and ( n57621 , n584889 , n57620 );
and ( n57622 , n53365 , n53468 );
and ( n57623 , n53367 , n53466 );
nor ( n584947 , n57622 , n57623 );
xnor ( n57625 , n584947 , n52945 );
and ( n584949 , n57620 , n57625 );
and ( n584950 , n584889 , n57625 );
or ( n57628 , n57621 , n584949 , n584950 );
and ( n584952 , n52936 , n53996 );
and ( n57630 , n52816 , n53994 );
nor ( n57631 , n584952 , n57630 );
xnor ( n57632 , n57631 , n53376 );
and ( n57633 , n57628 , n57632 );
xor ( n57634 , n584667 , n57358 );
xor ( n57635 , n57634 , n57363 );
and ( n57636 , n57632 , n57635 );
and ( n57637 , n57628 , n57635 );
or ( n57638 , n57633 , n57636 , n57637 );
and ( n57639 , n52488 , n55013 );
and ( n57640 , n52390 , n55010 );
nor ( n584964 , n57639 , n57640 );
xnor ( n57642 , n584964 , n53762 );
and ( n584966 , n57638 , n57642 );
and ( n57644 , n52626 , n54532 );
and ( n57645 , n52533 , n54530 );
nor ( n57646 , n57644 , n57645 );
xnor ( n57647 , n57646 , n53769 );
and ( n57648 , n57642 , n57647 );
and ( n57649 , n57638 , n57647 );
or ( n57650 , n584966 , n57648 , n57649 );
and ( n57651 , n52934 , n53996 );
and ( n57652 , n52936 , n53994 );
nor ( n57653 , n57651 , n57652 );
xnor ( n57654 , n57653 , n53376 );
and ( n57655 , n53107 , n53683 );
and ( n57656 , n53109 , n53681 );
nor ( n57657 , n57655 , n57656 );
xnor ( n57658 , n57657 , n53118 );
and ( n57659 , n57654 , n57658 );
xor ( n57660 , n584657 , n584661 );
xor ( n57661 , n57660 , n57341 );
and ( n584985 , n57658 , n57661 );
and ( n57663 , n57654 , n57661 );
or ( n57664 , n57659 , n584985 , n57663 );
and ( n57665 , n52818 , n54414 );
and ( n57666 , n52669 , n54412 );
nor ( n57667 , n57665 , n57666 );
xnor ( n584991 , n57667 , n53650 );
and ( n57669 , n57664 , n584991 );
xor ( n57670 , n584750 , n584752 );
xor ( n57671 , n57670 , n57432 );
and ( n57672 , n584991 , n57671 );
and ( n57673 , n57664 , n57671 );
or ( n57674 , n57669 , n57672 , n57673 );
xor ( n57675 , n57435 , n584762 );
xor ( n57676 , n57675 , n57442 );
and ( n57677 , n57674 , n57676 );
xor ( n57678 , n584689 , n57370 );
xor ( n57679 , n57678 , n57373 );
and ( n57680 , n57676 , n57679 );
and ( n57681 , n57674 , n57679 );
or ( n57682 , n57677 , n57680 , n57681 );
and ( n57683 , n57650 , n57682 );
xor ( n57684 , n584711 , n57392 );
xor ( n57685 , n57684 , n584718 );
and ( n57686 , n57682 , n57685 );
and ( n57687 , n57650 , n57685 );
or ( n57688 , n57683 , n57686 , n57687 );
xor ( n57689 , n57384 , n57398 );
xor ( n57690 , n57689 , n57401 );
and ( n57691 , n57688 , n57690 );
xor ( n57692 , n57453 , n57455 );
xor ( n57693 , n57692 , n584781 );
and ( n57694 , n57690 , n57693 );
and ( n57695 , n57688 , n57693 );
or ( n57696 , n57691 , n57694 , n57695 );
and ( n57697 , n57472 , n57696 );
xor ( n585021 , n57688 , n57690 );
xor ( n585022 , n585021 , n57693 );
and ( n585023 , n53837 , n53177 );
and ( n57701 , n53639 , n53175 );
nor ( n585025 , n585023 , n57701 );
xnor ( n585026 , n585025 , n52827 );
xor ( n57704 , n57324 , n57328 );
xor ( n57705 , n57704 , n57331 );
and ( n57706 , n585026 , n57705 );
xor ( n57707 , n57610 , n57614 );
xor ( n585031 , n57707 , n57617 );
and ( n57709 , n57705 , n585031 );
and ( n585033 , n585026 , n585031 );
or ( n57711 , n57706 , n57709 , n585033 );
xor ( n585035 , n584889 , n57620 );
xor ( n57713 , n585035 , n57625 );
and ( n585037 , n57711 , n57713 );
xor ( n585038 , n584671 , n584675 );
xor ( n57716 , n585038 , n57355 );
and ( n585040 , n57713 , n57716 );
and ( n585041 , n57711 , n57716 );
or ( n585042 , n585037 , n585040 , n585041 );
and ( n57720 , n52671 , n54532 );
and ( n585044 , n52626 , n54530 );
nor ( n585045 , n57720 , n585044 );
xnor ( n57723 , n585045 , n53769 );
and ( n585047 , n585042 , n57723 );
xor ( n57725 , n57628 , n57632 );
xor ( n57726 , n57725 , n57635 );
and ( n57727 , n57723 , n57726 );
and ( n585051 , n585042 , n57726 );
or ( n57729 , n585047 , n57727 , n585051 );
and ( n585053 , n584529 , n51991 );
and ( n585054 , n57058 , n51989 );
nor ( n57732 , n585053 , n585054 );
xnor ( n57733 , n57732 , n51959 );
and ( n57734 , n57484 , n51936 );
and ( n57735 , n57283 , n51934 );
nor ( n585059 , n57734 , n57735 );
xnor ( n585060 , n585059 , n51941 );
and ( n57738 , n57733 , n585060 );
buf ( n585062 , n578913 );
and ( n57740 , n585062 , n51929 );
and ( n57741 , n57482 , n51927 );
nor ( n57742 , n57740 , n57741 );
not ( n57743 , n57742 );
and ( n57744 , n585060 , n57743 );
and ( n57745 , n57733 , n57743 );
or ( n57746 , n57738 , n57744 , n57745 );
and ( n57747 , n56832 , n52065 );
and ( n57748 , n56671 , n52063 );
nor ( n57749 , n57747 , n57748 );
xnor ( n57750 , n57749 , n52022 );
and ( n57751 , n57746 , n57750 );
xor ( n57752 , n584799 , n57480 );
xor ( n57753 , n57752 , n57487 );
and ( n57754 , n57750 , n57753 );
and ( n57755 , n57746 , n57753 );
or ( n57756 , n57751 , n57754 , n57755 );
and ( n57757 , n583377 , n52273 );
and ( n57758 , n55841 , n52271 );
nor ( n57759 , n57757 , n57758 );
xnor ( n57760 , n57759 , n52137 );
and ( n57761 , n57756 , n57760 );
and ( n57762 , n56671 , n52065 );
and ( n585086 , n583800 , n52063 );
nor ( n57764 , n57762 , n585086 );
xnor ( n57765 , n57764 , n52022 );
and ( n57766 , n57760 , n57765 );
and ( n57767 , n57756 , n57765 );
or ( n57768 , n57761 , n57766 , n57767 );
and ( n585092 , n55293 , n52509 );
and ( n57770 , n55075 , n52507 );
nor ( n57771 , n585092 , n57770 );
xnor ( n585095 , n57771 , n52383 );
and ( n57773 , n57768 , n585095 );
xor ( n57774 , n57570 , n584897 );
xor ( n57775 , n57774 , n584900 );
and ( n57776 , n585095 , n57775 );
and ( n585100 , n57768 , n57775 );
or ( n585101 , n57773 , n57776 , n585100 );
and ( n57779 , n55075 , n52509 );
and ( n57780 , n55058 , n52507 );
nor ( n57781 , n57779 , n57780 );
xnor ( n57782 , n57781 , n52383 );
and ( n57783 , n585101 , n57782 );
xor ( n57784 , n584903 , n57584 );
xor ( n585108 , n57784 , n584910 );
and ( n57786 , n57782 , n585108 );
and ( n57787 , n585101 , n585108 );
or ( n585111 , n57783 , n57786 , n57787 );
and ( n57789 , n54725 , n52707 );
and ( n57790 , n54553 , n52705 );
nor ( n57791 , n57789 , n57790 );
xnor ( n57792 , n57791 , n52526 );
and ( n57793 , n585111 , n57792 );
xor ( n585117 , n57590 , n584917 );
xor ( n57795 , n585117 , n584920 );
and ( n57796 , n57792 , n57795 );
and ( n585120 , n585111 , n57795 );
or ( n585121 , n57793 , n57796 , n585120 );
and ( n57799 , n53639 , n53468 );
and ( n57800 , n53641 , n53466 );
nor ( n585124 , n57799 , n57800 );
xnor ( n57802 , n585124 , n52945 );
and ( n57803 , n585121 , n57802 );
xor ( n57804 , n584923 , n57604 );
xor ( n57805 , n57804 , n584930 );
and ( n57806 , n57802 , n57805 );
and ( n585130 , n585121 , n57805 );
or ( n57808 , n57803 , n57806 , n585130 );
and ( n57809 , n53109 , n53996 );
and ( n57810 , n52934 , n53994 );
nor ( n57811 , n57809 , n57810 );
xnor ( n57812 , n57811 , n53376 );
and ( n57813 , n57808 , n57812 );
and ( n585137 , n53367 , n53683 );
and ( n585138 , n53107 , n53681 );
nor ( n585139 , n585137 , n585138 );
xnor ( n57817 , n585139 , n53118 );
and ( n585141 , n57812 , n57817 );
and ( n585142 , n57808 , n57817 );
or ( n57820 , n57813 , n585141 , n585142 );
and ( n585144 , n53365 , n53683 );
and ( n585145 , n53367 , n53681 );
nor ( n57823 , n585144 , n585145 );
xnor ( n585147 , n57823 , n53118 );
and ( n585148 , n53835 , n53177 );
and ( n57826 , n53837 , n53175 );
nor ( n57827 , n585148 , n57826 );
xnor ( n585151 , n57827 , n52827 );
and ( n585152 , n585147 , n585151 );
and ( n57830 , n54215 , n52978 );
and ( n585154 , n54055 , n52976 );
nor ( n585155 , n57830 , n585154 );
xnor ( n57833 , n585155 , n52680 );
and ( n585157 , n585151 , n57833 );
and ( n585158 , n585147 , n57833 );
or ( n57836 , n585152 , n585157 , n585158 );
xor ( n585160 , n57554 , n584881 );
xor ( n585161 , n585160 , n584886 );
and ( n57839 , n57836 , n585161 );
xor ( n585163 , n585026 , n57705 );
xor ( n585164 , n585163 , n585031 );
and ( n585165 , n585161 , n585164 );
and ( n585166 , n57836 , n585164 );
or ( n57844 , n57839 , n585165 , n585166 );
and ( n585168 , n57820 , n57844 );
and ( n585169 , n52816 , n54414 );
and ( n585170 , n52818 , n54412 );
nor ( n585171 , n585169 , n585170 );
xnor ( n57849 , n585171 , n53650 );
and ( n585173 , n57844 , n57849 );
and ( n585174 , n57820 , n57849 );
or ( n57852 , n585168 , n585173 , n585174 );
and ( n585176 , n52533 , n55013 );
and ( n585177 , n52488 , n55010 );
nor ( n57855 , n585176 , n585177 );
xnor ( n585179 , n57855 , n53762 );
and ( n57857 , n57852 , n585179 );
xor ( n585181 , n57664 , n584991 );
xor ( n57859 , n585181 , n57671 );
and ( n57860 , n585179 , n57859 );
and ( n585184 , n57852 , n57859 );
or ( n585185 , n57857 , n57860 , n585184 );
and ( n57863 , n57729 , n585185 );
xor ( n585187 , n57638 , n57642 );
xor ( n585188 , n585187 , n57647 );
and ( n57866 , n585185 , n585188 );
and ( n585190 , n57729 , n585188 );
or ( n585191 , n57863 , n57866 , n585190 );
xor ( n57869 , n57650 , n57682 );
xor ( n585193 , n57869 , n57685 );
and ( n585194 , n585191 , n585193 );
xor ( n57872 , n57445 , n584770 );
xor ( n585196 , n57872 , n584773 );
and ( n585197 , n585193 , n585196 );
and ( n57875 , n585191 , n585196 );
or ( n585199 , n585194 , n585197 , n57875 );
and ( n585200 , n585022 , n585199 );
xor ( n585201 , n585191 , n585193 );
xor ( n57879 , n585201 , n585196 );
and ( n585203 , n57058 , n52065 );
and ( n585204 , n56909 , n52063 );
nor ( n57882 , n585203 , n585204 );
xnor ( n585206 , n57882 , n52022 );
and ( n57884 , n57283 , n51991 );
and ( n585208 , n584529 , n51989 );
nor ( n585209 , n57884 , n585208 );
xnor ( n57887 , n585209 , n51959 );
and ( n57888 , n585206 , n57887 );
and ( n585212 , n57484 , n51991 );
and ( n585213 , n57283 , n51989 );
nor ( n57891 , n585212 , n585213 );
xnor ( n585215 , n57891 , n51959 );
and ( n585216 , n585062 , n51936 );
and ( n57894 , n57482 , n51934 );
nor ( n585218 , n585216 , n57894 );
xnor ( n585219 , n585218 , n51941 );
and ( n57897 , n585215 , n585219 );
buf ( n585221 , n578915 );
and ( n585222 , n585221 , n51929 );
buf ( n57900 , n578914 );
and ( n585224 , n57900 , n51927 );
nor ( n585225 , n585222 , n585224 );
not ( n585226 , n585225 );
and ( n57904 , n585219 , n585226 );
and ( n585228 , n585215 , n585226 );
or ( n585229 , n57897 , n57904 , n585228 );
and ( n57907 , n57482 , n51936 );
and ( n585231 , n57484 , n51934 );
nor ( n585232 , n57907 , n585231 );
xnor ( n57910 , n585232 , n51941 );
xor ( n57911 , n585229 , n57910 );
and ( n585235 , n57900 , n51929 );
and ( n57913 , n585062 , n51927 );
nor ( n585237 , n585235 , n57913 );
not ( n585238 , n585237 );
xor ( n57916 , n57911 , n585238 );
and ( n57917 , n57887 , n57916 );
and ( n585241 , n585206 , n57916 );
or ( n585242 , n57888 , n57917 , n585241 );
and ( n57920 , n583746 , n52273 );
and ( n57921 , n56282 , n52271 );
nor ( n57922 , n57920 , n57921 );
xnor ( n585246 , n57922 , n52137 );
and ( n585247 , n585242 , n585246 );
and ( n57925 , n585229 , n57910 );
and ( n57926 , n57910 , n585238 );
and ( n57927 , n585229 , n585238 );
or ( n57928 , n57925 , n57926 , n57927 );
and ( n57929 , n56909 , n52065 );
and ( n585253 , n56832 , n52063 );
nor ( n57931 , n57929 , n585253 );
xnor ( n57932 , n57931 , n52022 );
xor ( n57933 , n57928 , n57932 );
xor ( n585257 , n57733 , n585060 );
xor ( n57935 , n585257 , n57743 );
xor ( n585259 , n57933 , n57935 );
and ( n585260 , n585246 , n585259 );
and ( n57938 , n585242 , n585259 );
or ( n585262 , n585247 , n585260 , n57938 );
and ( n57940 , n55841 , n52432 );
and ( n57941 , n583048 , n52430 );
nor ( n57942 , n57940 , n57941 );
xnor ( n585266 , n57942 , n52255 );
and ( n57944 , n585262 , n585266 );
and ( n585268 , n56282 , n52273 );
and ( n585269 , n583377 , n52271 );
nor ( n57947 , n585268 , n585269 );
xnor ( n585271 , n57947 , n52137 );
and ( n57949 , n585266 , n585271 );
and ( n585273 , n585262 , n585271 );
or ( n585274 , n57944 , n57949 , n585273 );
and ( n57952 , n55528 , n52509 );
and ( n585276 , n55293 , n52507 );
nor ( n585277 , n57952 , n585276 );
xnor ( n57955 , n585277 , n52383 );
and ( n57956 , n585274 , n57955 );
xor ( n585280 , n57756 , n57760 );
xor ( n585281 , n585280 , n57765 );
and ( n57959 , n57955 , n585281 );
and ( n57960 , n585274 , n585281 );
or ( n585284 , n57956 , n57959 , n57960 );
and ( n585285 , n55058 , n52707 );
and ( n585286 , n54893 , n52705 );
nor ( n57964 , n585285 , n585286 );
xnor ( n585288 , n57964 , n52526 );
and ( n585289 , n585284 , n585288 );
xor ( n57967 , n57768 , n585095 );
xor ( n585291 , n57967 , n57775 );
and ( n585292 , n585288 , n585291 );
and ( n57970 , n585284 , n585291 );
or ( n57971 , n585289 , n585292 , n57970 );
and ( n585295 , n54553 , n52978 );
and ( n585296 , n54321 , n52976 );
nor ( n57974 , n585295 , n585296 );
xnor ( n57975 , n57974 , n52680 );
and ( n585299 , n57971 , n57975 );
xor ( n585300 , n585101 , n57782 );
xor ( n57978 , n585300 , n585108 );
and ( n585302 , n57975 , n57978 );
and ( n57980 , n57971 , n57978 );
or ( n585304 , n585299 , n585302 , n57980 );
and ( n585305 , n53641 , n53683 );
and ( n57983 , n53365 , n53681 );
nor ( n585307 , n585305 , n57983 );
xnor ( n585308 , n585307 , n53118 );
and ( n57986 , n585304 , n585308 );
and ( n57987 , n53837 , n53468 );
and ( n585311 , n53639 , n53466 );
nor ( n585312 , n57987 , n585311 );
xnor ( n57990 , n585312 , n52945 );
and ( n57991 , n585308 , n57990 );
and ( n585315 , n585304 , n57990 );
or ( n585316 , n57986 , n57991 , n585315 );
and ( n57994 , n57928 , n57932 );
and ( n57995 , n57932 , n57935 );
and ( n57996 , n57928 , n57935 );
or ( n585320 , n57994 , n57995 , n57996 );
and ( n57998 , n583800 , n52155 );
and ( n57999 , n583746 , n52153 );
nor ( n58000 , n57998 , n57999 );
xnor ( n585324 , n58000 , n52085 );
and ( n585325 , n585320 , n585324 );
xor ( n58003 , n57746 , n57750 );
xor ( n585327 , n58003 , n57753 );
and ( n58005 , n585324 , n585327 );
and ( n58006 , n585320 , n585327 );
or ( n58007 , n585325 , n58005 , n58006 );
and ( n58008 , n583048 , n52432 );
and ( n58009 , n582961 , n52430 );
nor ( n58010 , n58008 , n58009 );
xnor ( n58011 , n58010 , n52255 );
and ( n58012 , n58007 , n58011 );
xor ( n58013 , n584813 , n584817 );
xor ( n58014 , n58013 , n57509 );
and ( n58015 , n58011 , n58014 );
and ( n58016 , n58007 , n58014 );
or ( n58017 , n58012 , n58015 , n58016 );
and ( n58018 , n582961 , n52432 );
and ( n58019 , n55528 , n52430 );
nor ( n585343 , n58018 , n58019 );
xnor ( n585344 , n585343 , n52255 );
and ( n58022 , n58017 , n585344 );
xor ( n585346 , n584835 , n584839 );
xor ( n585347 , n585346 , n584844 );
and ( n58025 , n585344 , n585347 );
and ( n585349 , n58017 , n585347 );
or ( n585350 , n58022 , n58025 , n585349 );
and ( n58028 , n54893 , n52707 );
and ( n585352 , n54725 , n52705 );
nor ( n585353 , n58028 , n585352 );
xnor ( n58031 , n585353 , n52526 );
and ( n58032 , n585350 , n58031 );
xor ( n585356 , n584847 , n57528 );
xor ( n585357 , n585356 , n57531 );
and ( n58035 , n58031 , n585357 );
and ( n585359 , n585350 , n585357 );
or ( n585360 , n58032 , n58035 , n585359 );
and ( n58038 , n54321 , n52978 );
and ( n585362 , n54215 , n52976 );
nor ( n585363 , n58038 , n585362 );
xnor ( n58041 , n585363 , n52680 );
and ( n585365 , n585360 , n58041 );
xor ( n585366 , n584857 , n584861 );
xor ( n58044 , n585366 , n57541 );
and ( n585368 , n58041 , n58044 );
and ( n585369 , n585360 , n58044 );
or ( n585370 , n585365 , n585368 , n585369 );
and ( n585371 , n585316 , n585370 );
xor ( n58049 , n57544 , n584871 );
xor ( n585373 , n58049 , n584874 );
and ( n585374 , n585370 , n585373 );
and ( n585375 , n585316 , n585373 );
or ( n585376 , n585371 , n585374 , n585375 );
and ( n58054 , n52936 , n54414 );
and ( n585378 , n52816 , n54412 );
nor ( n585379 , n58054 , n585378 );
xnor ( n58057 , n585379 , n53650 );
and ( n585381 , n585376 , n58057 );
xor ( n585382 , n57808 , n57812 );
xor ( n58060 , n585382 , n57817 );
and ( n585384 , n58057 , n58060 );
and ( n58062 , n585376 , n58060 );
or ( n585386 , n585381 , n585384 , n58062 );
and ( n58064 , n53107 , n53996 );
and ( n58065 , n53109 , n53994 );
nor ( n585389 , n58064 , n58065 );
xnor ( n585390 , n585389 , n53376 );
xor ( n58068 , n585147 , n585151 );
xor ( n585392 , n58068 , n57833 );
and ( n585393 , n585390 , n585392 );
xor ( n58071 , n585121 , n57802 );
xor ( n585395 , n58071 , n57805 );
and ( n585396 , n585392 , n585395 );
and ( n58074 , n585390 , n585395 );
or ( n585398 , n585393 , n585396 , n58074 );
and ( n585399 , n52818 , n54532 );
and ( n58077 , n52669 , n54530 );
nor ( n585401 , n585399 , n58077 );
xnor ( n585402 , n585401 , n53769 );
and ( n58080 , n585398 , n585402 );
xor ( n585404 , n57836 , n585161 );
xor ( n585405 , n585404 , n585164 );
and ( n58083 , n585402 , n585405 );
and ( n585407 , n585398 , n585405 );
or ( n585408 , n58080 , n58083 , n585407 );
and ( n58086 , n585386 , n585408 );
and ( n585410 , n52626 , n55013 );
and ( n585411 , n52533 , n55010 );
nor ( n58089 , n585410 , n585411 );
xnor ( n58090 , n58089 , n53762 );
and ( n585414 , n585408 , n58090 );
and ( n585415 , n585386 , n58090 );
or ( n58093 , n58086 , n585414 , n585415 );
and ( n585417 , n52669 , n54532 );
and ( n585418 , n52671 , n54530 );
nor ( n58096 , n585417 , n585418 );
xnor ( n585420 , n58096 , n53769 );
xor ( n585421 , n57654 , n57658 );
xor ( n58099 , n585421 , n57661 );
and ( n585423 , n585420 , n58099 );
xor ( n585424 , n57711 , n57713 );
xor ( n58102 , n585424 , n57716 );
and ( n585426 , n58099 , n58102 );
and ( n585427 , n585420 , n58102 );
or ( n58105 , n585423 , n585426 , n585427 );
and ( n58106 , n58093 , n58105 );
xor ( n58107 , n585042 , n57723 );
xor ( n585431 , n58107 , n57726 );
and ( n585432 , n58105 , n585431 );
and ( n58110 , n58093 , n585431 );
or ( n58111 , n58106 , n585432 , n58110 );
xor ( n585435 , n57729 , n585185 );
xor ( n585436 , n585435 , n585188 );
and ( n58114 , n58111 , n585436 );
xor ( n585438 , n57674 , n57676 );
xor ( n585439 , n585438 , n57679 );
and ( n58117 , n585436 , n585439 );
and ( n58118 , n58111 , n585439 );
or ( n58119 , n58114 , n58117 , n58118 );
and ( n58120 , n57879 , n58119 );
xor ( n58121 , n58111 , n585436 );
xor ( n58122 , n58121 , n585439 );
and ( n58123 , n54055 , n53177 );
and ( n58124 , n53835 , n53175 );
nor ( n58125 , n58123 , n58124 );
xnor ( n585449 , n58125 , n52827 );
xor ( n585450 , n585360 , n58041 );
xor ( n58128 , n585450 , n58044 );
and ( n585452 , n585449 , n58128 );
xor ( n58130 , n585111 , n57792 );
xor ( n585454 , n58130 , n57795 );
and ( n585455 , n58128 , n585454 );
and ( n58133 , n585449 , n585454 );
or ( n585457 , n585452 , n585455 , n58133 );
and ( n58135 , n52934 , n54414 );
and ( n58136 , n52936 , n54412 );
nor ( n585460 , n58135 , n58136 );
xnor ( n585461 , n585460 , n53650 );
and ( n58139 , n585457 , n585461 );
xor ( n585463 , n585316 , n585370 );
xor ( n585464 , n585463 , n585373 );
and ( n58142 , n585461 , n585464 );
and ( n585466 , n585457 , n585464 );
or ( n585467 , n58139 , n58142 , n585466 );
and ( n58145 , n52671 , n55013 );
and ( n585469 , n52626 , n55010 );
nor ( n58147 , n58145 , n585469 );
xnor ( n58148 , n58147 , n53762 );
and ( n58149 , n585467 , n58148 );
xor ( n58150 , n585376 , n58057 );
xor ( n585474 , n58150 , n58060 );
and ( n58152 , n58148 , n585474 );
and ( n58153 , n585467 , n585474 );
or ( n585477 , n58149 , n58152 , n58153 );
xor ( n58155 , n57820 , n57844 );
xor ( n585479 , n58155 , n57849 );
and ( n58157 , n585477 , n585479 );
xor ( n585481 , n585420 , n58099 );
xor ( n585482 , n585481 , n58102 );
and ( n58160 , n585479 , n585482 );
and ( n585484 , n585477 , n585482 );
or ( n585485 , n58157 , n58160 , n585484 );
xor ( n58163 , n58093 , n58105 );
xor ( n585487 , n58163 , n585431 );
and ( n58165 , n585485 , n585487 );
xor ( n58166 , n57852 , n585179 );
xor ( n58167 , n58166 , n57859 );
and ( n58168 , n585487 , n58167 );
and ( n58169 , n585485 , n58167 );
or ( n58170 , n58165 , n58168 , n58169 );
and ( n58171 , n58122 , n58170 );
xor ( n58172 , n585485 , n585487 );
xor ( n58173 , n58172 , n58167 );
and ( n585497 , n53639 , n53683 );
and ( n58175 , n53641 , n53681 );
nor ( n585499 , n585497 , n58175 );
xnor ( n58177 , n585499 , n53118 );
and ( n58178 , n54215 , n53177 );
and ( n58179 , n54055 , n53175 );
nor ( n585503 , n58178 , n58179 );
xnor ( n585504 , n585503 , n52827 );
and ( n58182 , n58177 , n585504 );
xor ( n585506 , n585350 , n58031 );
xor ( n58184 , n585506 , n585357 );
and ( n585508 , n585504 , n58184 );
and ( n58186 , n58177 , n58184 );
or ( n585510 , n58182 , n585508 , n58186 );
and ( n585511 , n53109 , n54414 );
and ( n58189 , n52934 , n54412 );
nor ( n58190 , n585511 , n58189 );
xnor ( n585514 , n58190 , n53650 );
and ( n585515 , n585510 , n585514 );
and ( n58193 , n53367 , n53996 );
and ( n58194 , n53107 , n53994 );
nor ( n58195 , n58193 , n58194 );
xnor ( n58196 , n58195 , n53376 );
and ( n58197 , n585514 , n58196 );
and ( n58198 , n585510 , n58196 );
or ( n58199 , n585515 , n58197 , n58198 );
and ( n58200 , n52816 , n54532 );
and ( n58201 , n52818 , n54530 );
nor ( n58202 , n58200 , n58201 );
xnor ( n58203 , n58202 , n53769 );
and ( n58204 , n58199 , n58203 );
xor ( n58205 , n585390 , n585392 );
xor ( n58206 , n58205 , n585395 );
and ( n58207 , n58203 , n58206 );
and ( n585531 , n58199 , n58206 );
or ( n58209 , n58204 , n58207 , n585531 );
and ( n585533 , n57482 , n51991 );
and ( n585534 , n57484 , n51989 );
nor ( n58212 , n585533 , n585534 );
xnor ( n58213 , n58212 , n51959 );
and ( n58214 , n57900 , n51936 );
and ( n585538 , n585062 , n51934 );
nor ( n58216 , n58214 , n585538 );
xnor ( n58217 , n58216 , n51941 );
and ( n58218 , n58213 , n58217 );
buf ( n58219 , n578916 );
and ( n58220 , n58219 , n51929 );
and ( n58221 , n585221 , n51927 );
nor ( n58222 , n58220 , n58221 );
not ( n585546 , n58222 );
and ( n58224 , n58217 , n585546 );
and ( n585548 , n58213 , n585546 );
or ( n58226 , n58218 , n58224 , n585548 );
and ( n58227 , n584529 , n52065 );
and ( n585551 , n57058 , n52063 );
nor ( n58229 , n58227 , n585551 );
xnor ( n585553 , n58229 , n52022 );
and ( n585554 , n58226 , n585553 );
xor ( n585555 , n585215 , n585219 );
xor ( n58233 , n585555 , n585226 );
and ( n585557 , n585553 , n58233 );
and ( n58235 , n58226 , n58233 );
or ( n58236 , n585554 , n585557 , n58235 );
and ( n585560 , n585062 , n51991 );
and ( n58238 , n57482 , n51989 );
nor ( n585562 , n585560 , n58238 );
xnor ( n58240 , n585562 , n51959 );
and ( n58241 , n585221 , n51936 );
and ( n58242 , n57900 , n51934 );
nor ( n58243 , n58241 , n58242 );
xnor ( n58244 , n58243 , n51941 );
and ( n58245 , n58240 , n58244 );
buf ( n58246 , n578917 );
and ( n58247 , n58246 , n51929 );
and ( n58248 , n58219 , n51927 );
nor ( n58249 , n58247 , n58248 );
not ( n58250 , n58249 );
and ( n58251 , n58244 , n58250 );
and ( n58252 , n58240 , n58250 );
or ( n58253 , n58245 , n58251 , n58252 );
and ( n58254 , n57900 , n51991 );
and ( n585578 , n585062 , n51989 );
nor ( n58256 , n58254 , n585578 );
xnor ( n585580 , n58256 , n51959 );
and ( n58258 , n58219 , n51936 );
and ( n585582 , n585221 , n51934 );
nor ( n58260 , n58258 , n585582 );
xnor ( n585584 , n58260 , n51941 );
and ( n58262 , n585580 , n585584 );
buf ( n585586 , n578918 );
and ( n58264 , n585586 , n51929 );
and ( n585588 , n58246 , n51927 );
nor ( n585589 , n58264 , n585588 );
not ( n58267 , n585589 );
and ( n585591 , n585584 , n58267 );
and ( n58269 , n585580 , n58267 );
or ( n585593 , n58262 , n585591 , n58269 );
and ( n585594 , n57484 , n52065 );
and ( n58272 , n57283 , n52063 );
nor ( n58273 , n585594 , n58272 );
xnor ( n58274 , n58273 , n52022 );
and ( n58275 , n585593 , n58274 );
xor ( n585599 , n58240 , n58244 );
xor ( n58277 , n585599 , n58250 );
and ( n585601 , n58274 , n58277 );
and ( n58279 , n585593 , n58277 );
or ( n58280 , n58275 , n585601 , n58279 );
and ( n58281 , n58253 , n58280 );
xor ( n58282 , n58213 , n58217 );
xor ( n585606 , n58282 , n585546 );
and ( n58284 , n58280 , n585606 );
and ( n58285 , n58253 , n585606 );
or ( n585609 , n58281 , n58284 , n58285 );
and ( n58287 , n56909 , n52155 );
and ( n58288 , n56832 , n52153 );
nor ( n585612 , n58287 , n58288 );
xnor ( n58290 , n585612 , n52085 );
and ( n585614 , n585609 , n58290 );
xor ( n585615 , n58226 , n585553 );
xor ( n58293 , n585615 , n58233 );
and ( n585617 , n58290 , n58293 );
and ( n585618 , n585609 , n58293 );
or ( n58296 , n585614 , n585617 , n585618 );
and ( n58297 , n58236 , n58296 );
xor ( n585621 , n585206 , n57887 );
xor ( n58299 , n585621 , n57916 );
and ( n58300 , n58296 , n58299 );
and ( n58301 , n58236 , n58299 );
or ( n58302 , n58297 , n58300 , n58301 );
and ( n585626 , n583377 , n52432 );
and ( n58304 , n55841 , n52430 );
nor ( n58305 , n585626 , n58304 );
xnor ( n58306 , n58305 , n52255 );
and ( n58307 , n58302 , n58306 );
and ( n585631 , n56671 , n52155 );
and ( n585632 , n583800 , n52153 );
nor ( n585633 , n585631 , n585632 );
xnor ( n58311 , n585633 , n52085 );
and ( n585635 , n58306 , n58311 );
and ( n585636 , n58302 , n58311 );
or ( n58314 , n58307 , n585635 , n585636 );
and ( n585638 , n55293 , n52707 );
and ( n58316 , n55075 , n52705 );
nor ( n58317 , n585638 , n58316 );
xnor ( n585641 , n58317 , n52526 );
and ( n585642 , n58314 , n585641 );
xor ( n58320 , n585320 , n585324 );
xor ( n585644 , n58320 , n585327 );
and ( n585645 , n585641 , n585644 );
and ( n58323 , n58314 , n585644 );
or ( n585647 , n585642 , n585645 , n58323 );
and ( n585648 , n55075 , n52707 );
and ( n58326 , n55058 , n52705 );
nor ( n58327 , n585648 , n58326 );
xnor ( n58328 , n58327 , n52526 );
and ( n58329 , n585647 , n58328 );
xor ( n585653 , n58007 , n58011 );
xor ( n58331 , n585653 , n58014 );
and ( n58332 , n58328 , n58331 );
and ( n58333 , n585647 , n58331 );
or ( n58334 , n58329 , n58332 , n58333 );
and ( n585658 , n54725 , n52978 );
and ( n585659 , n54553 , n52976 );
nor ( n58337 , n585658 , n585659 );
xnor ( n585661 , n58337 , n52680 );
and ( n585662 , n58334 , n585661 );
xor ( n58340 , n58017 , n585344 );
xor ( n585664 , n58340 , n585347 );
and ( n585665 , n585661 , n585664 );
and ( n585666 , n58334 , n585664 );
or ( n58344 , n585662 , n585665 , n585666 );
and ( n585668 , n53835 , n53468 );
and ( n58346 , n53837 , n53466 );
nor ( n58347 , n585668 , n58346 );
xnor ( n58348 , n58347 , n52945 );
and ( n58349 , n58344 , n58348 );
xor ( n58350 , n57971 , n57975 );
xor ( n58351 , n58350 , n57978 );
and ( n58352 , n58348 , n58351 );
and ( n58353 , n58344 , n58351 );
or ( n58354 , n58349 , n58352 , n58353 );
xor ( n58355 , n585304 , n585308 );
xor ( n58356 , n58355 , n57990 );
and ( n58357 , n58354 , n58356 );
xor ( n58358 , n585449 , n58128 );
xor ( n58359 , n58358 , n585454 );
and ( n58360 , n58356 , n58359 );
and ( n58361 , n58354 , n58359 );
or ( n58362 , n58357 , n58360 , n58361 );
and ( n58363 , n52669 , n55013 );
and ( n58364 , n52671 , n55010 );
nor ( n58365 , n58363 , n58364 );
xnor ( n58366 , n58365 , n53762 );
and ( n58367 , n58362 , n58366 );
xor ( n58368 , n585457 , n585461 );
xor ( n58369 , n58368 , n585464 );
and ( n58370 , n58366 , n58369 );
and ( n58371 , n58362 , n58369 );
or ( n58372 , n58367 , n58370 , n58371 );
and ( n58373 , n58209 , n58372 );
xor ( n58374 , n585398 , n585402 );
xor ( n58375 , n58374 , n585405 );
and ( n58376 , n58372 , n58375 );
and ( n585700 , n58209 , n58375 );
or ( n58378 , n58373 , n58376 , n585700 );
xor ( n585702 , n585386 , n585408 );
xor ( n585703 , n585702 , n58090 );
and ( n585704 , n58378 , n585703 );
xor ( n585705 , n585477 , n585479 );
xor ( n58383 , n585705 , n585482 );
and ( n585707 , n585703 , n58383 );
and ( n58385 , n58378 , n58383 );
or ( n585709 , n585704 , n585707 , n58385 );
and ( n58387 , n58173 , n585709 );
xor ( n585711 , n58378 , n585703 );
xor ( n58389 , n585711 , n58383 );
and ( n58390 , n57058 , n52155 );
and ( n58391 , n56909 , n52153 );
nor ( n58392 , n58390 , n58391 );
xnor ( n58393 , n58392 , n52085 );
and ( n58394 , n57283 , n52065 );
and ( n58395 , n584529 , n52063 );
nor ( n58396 , n58394 , n58395 );
xnor ( n585720 , n58396 , n52022 );
and ( n585721 , n58393 , n585720 );
xor ( n58399 , n58253 , n58280 );
xor ( n58400 , n58399 , n585606 );
and ( n58401 , n585720 , n58400 );
and ( n58402 , n58393 , n58400 );
or ( n585726 , n585721 , n58401 , n58402 );
and ( n585727 , n56671 , n52273 );
and ( n58405 , n583800 , n52271 );
nor ( n585729 , n585727 , n58405 );
xnor ( n585730 , n585729 , n52137 );
and ( n58408 , n585726 , n585730 );
xor ( n585732 , n585609 , n58290 );
xor ( n585733 , n585732 , n58293 );
and ( n585734 , n585730 , n585733 );
and ( n585735 , n585726 , n585733 );
or ( n58413 , n58408 , n585734 , n585735 );
and ( n585737 , n55841 , n52509 );
and ( n585738 , n583048 , n52507 );
nor ( n58416 , n585737 , n585738 );
xnor ( n585740 , n58416 , n52383 );
and ( n585741 , n58413 , n585740 );
and ( n58419 , n56282 , n52432 );
and ( n585743 , n583377 , n52430 );
nor ( n585744 , n58419 , n585743 );
xnor ( n58422 , n585744 , n52255 );
and ( n585746 , n585740 , n58422 );
and ( n585747 , n58413 , n58422 );
or ( n58425 , n585741 , n585746 , n585747 );
and ( n585749 , n55528 , n52707 );
and ( n585750 , n55293 , n52705 );
nor ( n585751 , n585749 , n585750 );
xnor ( n585752 , n585751 , n52526 );
and ( n58430 , n58425 , n585752 );
xor ( n585754 , n58302 , n58306 );
xor ( n585755 , n585754 , n58311 );
and ( n585756 , n585752 , n585755 );
and ( n58434 , n58425 , n585755 );
or ( n585758 , n58430 , n585756 , n58434 );
and ( n58436 , n55058 , n52978 );
and ( n585760 , n54893 , n52976 );
nor ( n585761 , n58436 , n585760 );
xnor ( n58439 , n585761 , n52680 );
and ( n585763 , n585758 , n58439 );
xor ( n58441 , n58314 , n585641 );
xor ( n585765 , n58441 , n585644 );
and ( n585766 , n58439 , n585765 );
and ( n58444 , n585758 , n585765 );
or ( n585768 , n585763 , n585766 , n58444 );
and ( n585769 , n54553 , n53177 );
and ( n585770 , n54321 , n53175 );
nor ( n585771 , n585769 , n585770 );
xnor ( n58449 , n585771 , n52827 );
and ( n585773 , n585768 , n58449 );
xor ( n585774 , n585647 , n58328 );
xor ( n58452 , n585774 , n58331 );
and ( n585776 , n58449 , n58452 );
and ( n585777 , n585768 , n58452 );
or ( n58455 , n585773 , n585776 , n585777 );
and ( n585779 , n53837 , n53683 );
and ( n585780 , n53639 , n53681 );
nor ( n58458 , n585779 , n585780 );
xnor ( n585782 , n58458 , n53118 );
and ( n585783 , n58455 , n585782 );
xor ( n585784 , n58334 , n585661 );
xor ( n58462 , n585784 , n585664 );
and ( n585786 , n585782 , n58462 );
and ( n585787 , n58455 , n58462 );
or ( n585788 , n585783 , n585786 , n585787 );
and ( n585789 , n583800 , n52273 );
and ( n58467 , n583746 , n52271 );
nor ( n585791 , n585789 , n58467 );
xnor ( n585792 , n585791 , n52137 );
and ( n58470 , n56832 , n52155 );
and ( n585794 , n56671 , n52153 );
nor ( n585795 , n58470 , n585794 );
xnor ( n58473 , n585795 , n52085 );
and ( n585797 , n585792 , n58473 );
xor ( n585798 , n58236 , n58296 );
xor ( n58476 , n585798 , n58299 );
and ( n585800 , n58473 , n58476 );
and ( n58478 , n585792 , n58476 );
or ( n58479 , n585797 , n585800 , n58478 );
and ( n585803 , n583048 , n52509 );
and ( n58481 , n582961 , n52507 );
nor ( n585805 , n585803 , n58481 );
xnor ( n58483 , n585805 , n52383 );
and ( n58484 , n58479 , n58483 );
xor ( n58485 , n585242 , n585246 );
xor ( n58486 , n58485 , n585259 );
and ( n58487 , n58483 , n58486 );
and ( n585811 , n58479 , n58486 );
or ( n58489 , n58484 , n58487 , n585811 );
and ( n58490 , n582961 , n52509 );
and ( n585814 , n55528 , n52507 );
nor ( n58492 , n58490 , n585814 );
xnor ( n585816 , n58492 , n52383 );
and ( n585817 , n58489 , n585816 );
xor ( n585818 , n585262 , n585266 );
xor ( n585819 , n585818 , n585271 );
and ( n58497 , n585816 , n585819 );
and ( n585821 , n58489 , n585819 );
or ( n585822 , n585817 , n58497 , n585821 );
and ( n58500 , n54893 , n52978 );
and ( n585824 , n54725 , n52976 );
nor ( n585825 , n58500 , n585824 );
xnor ( n58503 , n585825 , n52680 );
and ( n585827 , n585822 , n58503 );
xor ( n58505 , n585274 , n57955 );
xor ( n58506 , n58505 , n585281 );
and ( n585830 , n58503 , n58506 );
and ( n58508 , n585822 , n58506 );
or ( n585832 , n585827 , n585830 , n58508 );
and ( n58510 , n54321 , n53177 );
and ( n58511 , n54215 , n53175 );
nor ( n585835 , n58510 , n58511 );
xnor ( n58513 , n585835 , n52827 );
and ( n585837 , n585832 , n58513 );
xor ( n585838 , n585284 , n585288 );
xor ( n58516 , n585838 , n585291 );
and ( n585840 , n58513 , n58516 );
and ( n58518 , n585832 , n58516 );
or ( n585842 , n585837 , n585840 , n58518 );
and ( n58520 , n585788 , n585842 );
and ( n58521 , n53365 , n53996 );
and ( n585845 , n53367 , n53994 );
nor ( n58523 , n58521 , n585845 );
xnor ( n585847 , n58523 , n53376 );
and ( n585848 , n585842 , n585847 );
and ( n58526 , n585788 , n585847 );
or ( n585850 , n58520 , n585848 , n58526 );
and ( n585851 , n52818 , n55013 );
and ( n585852 , n52669 , n55010 );
nor ( n585853 , n585851 , n585852 );
xnor ( n58531 , n585853 , n53762 );
and ( n585855 , n585850 , n58531 );
and ( n585856 , n52936 , n54532 );
and ( n58534 , n52816 , n54530 );
nor ( n585858 , n585856 , n58534 );
xnor ( n585859 , n585858 , n53769 );
and ( n58537 , n58531 , n585859 );
and ( n585861 , n585850 , n585859 );
or ( n585862 , n585855 , n58537 , n585861 );
and ( n58540 , n53107 , n54414 );
and ( n58541 , n53109 , n54412 );
nor ( n585865 , n58540 , n58541 );
xnor ( n585866 , n585865 , n53650 );
xor ( n58544 , n58177 , n585504 );
xor ( n585868 , n58544 , n58184 );
and ( n585869 , n585866 , n585868 );
xor ( n58547 , n58344 , n58348 );
xor ( n585871 , n58547 , n58351 );
and ( n585872 , n585868 , n585871 );
and ( n585873 , n585866 , n585871 );
or ( n58551 , n585869 , n585872 , n585873 );
xor ( n585875 , n585510 , n585514 );
xor ( n585876 , n585875 , n58196 );
and ( n585877 , n58551 , n585876 );
xor ( n58555 , n58354 , n58356 );
xor ( n585879 , n58555 , n58359 );
and ( n585880 , n585876 , n585879 );
and ( n58558 , n58551 , n585879 );
or ( n585882 , n585877 , n585880 , n58558 );
and ( n58560 , n585862 , n585882 );
xor ( n58561 , n58199 , n58203 );
xor ( n585885 , n58561 , n58206 );
and ( n58563 , n585882 , n585885 );
and ( n585887 , n585862 , n585885 );
or ( n58565 , n58560 , n58563 , n585887 );
xor ( n585889 , n585467 , n58148 );
xor ( n585890 , n585889 , n585474 );
and ( n58568 , n58565 , n585890 );
xor ( n585892 , n58209 , n58372 );
xor ( n585893 , n585892 , n58375 );
and ( n58571 , n585890 , n585893 );
and ( n58572 , n58565 , n585893 );
or ( n585896 , n58568 , n58571 , n58572 );
and ( n58574 , n58389 , n585896 );
xor ( n58575 , n58565 , n585890 );
xor ( n58576 , n58575 , n585893 );
and ( n58577 , n585221 , n51991 );
and ( n585901 , n57900 , n51989 );
nor ( n58579 , n58577 , n585901 );
xnor ( n58580 , n58579 , n51959 );
and ( n585904 , n58246 , n51936 );
and ( n585905 , n58219 , n51934 );
nor ( n585906 , n585904 , n585905 );
xnor ( n58584 , n585906 , n51941 );
and ( n585908 , n58580 , n58584 );
buf ( n585909 , n578919 );
and ( n585910 , n585909 , n51929 );
and ( n58588 , n585586 , n51927 );
nor ( n585912 , n585910 , n58588 );
not ( n585913 , n585912 );
and ( n58591 , n58584 , n585913 );
and ( n585915 , n58580 , n585913 );
or ( n58593 , n585908 , n58591 , n585915 );
and ( n58594 , n57482 , n52065 );
and ( n58595 , n57484 , n52063 );
nor ( n58596 , n58594 , n58595 );
xnor ( n585920 , n58596 , n52022 );
and ( n58598 , n58593 , n585920 );
xor ( n585922 , n585580 , n585584 );
xor ( n585923 , n585922 , n58267 );
and ( n58601 , n585920 , n585923 );
and ( n58602 , n58593 , n585923 );
or ( n585926 , n58598 , n58601 , n58602 );
and ( n585927 , n584529 , n52155 );
and ( n58605 , n57058 , n52153 );
nor ( n58606 , n585927 , n58605 );
xnor ( n585930 , n58606 , n52085 );
and ( n58608 , n585926 , n585930 );
xor ( n58609 , n585593 , n58274 );
xor ( n58610 , n58609 , n58277 );
and ( n58611 , n585930 , n58610 );
and ( n585935 , n585926 , n58610 );
or ( n585936 , n58608 , n58611 , n585935 );
and ( n585937 , n58219 , n51991 );
and ( n58615 , n585221 , n51989 );
nor ( n585939 , n585937 , n58615 );
xnor ( n585940 , n585939 , n51959 );
and ( n585941 , n585586 , n51936 );
and ( n585942 , n58246 , n51934 );
nor ( n58620 , n585941 , n585942 );
xnor ( n585944 , n58620 , n51941 );
and ( n585945 , n585940 , n585944 );
buf ( n58623 , n578920 );
and ( n585947 , n58623 , n51929 );
and ( n585948 , n585909 , n51927 );
nor ( n58626 , n585947 , n585948 );
not ( n585950 , n58626 );
and ( n585951 , n585944 , n585950 );
and ( n58629 , n585940 , n585950 );
or ( n585953 , n585945 , n585951 , n58629 );
and ( n585954 , n585062 , n52065 );
and ( n58632 , n57482 , n52063 );
nor ( n585956 , n585954 , n58632 );
xnor ( n585957 , n585956 , n52022 );
and ( n58635 , n585953 , n585957 );
xor ( n585959 , n58580 , n58584 );
xor ( n585960 , n585959 , n585913 );
and ( n585961 , n585957 , n585960 );
and ( n585962 , n585953 , n585960 );
or ( n58640 , n58635 , n585961 , n585962 );
and ( n585964 , n58246 , n51991 );
and ( n585965 , n58219 , n51989 );
nor ( n58643 , n585964 , n585965 );
xnor ( n585967 , n58643 , n51959 );
and ( n585968 , n585909 , n51936 );
and ( n58646 , n585586 , n51934 );
nor ( n585970 , n585968 , n58646 );
xnor ( n585971 , n585970 , n51941 );
and ( n58649 , n585967 , n585971 );
buf ( n585973 , n578921 );
and ( n585974 , n585973 , n51929 );
and ( n585975 , n58623 , n51927 );
nor ( n585976 , n585974 , n585975 );
not ( n58654 , n585976 );
and ( n585978 , n585971 , n58654 );
and ( n585979 , n585967 , n58654 );
or ( n585980 , n58649 , n585978 , n585979 );
and ( n585981 , n57900 , n52065 );
and ( n58659 , n585062 , n52063 );
nor ( n585983 , n585981 , n58659 );
xnor ( n585984 , n585983 , n52022 );
and ( n58662 , n585980 , n585984 );
xor ( n585986 , n585940 , n585944 );
xor ( n585987 , n585986 , n585950 );
and ( n58665 , n585984 , n585987 );
and ( n585989 , n585980 , n585987 );
or ( n585990 , n58662 , n58665 , n585989 );
and ( n58668 , n57484 , n52155 );
and ( n58669 , n57283 , n52153 );
nor ( n58670 , n58668 , n58669 );
xnor ( n585994 , n58670 , n52085 );
and ( n585995 , n585990 , n585994 );
xor ( n58673 , n585953 , n585957 );
xor ( n585997 , n58673 , n585960 );
and ( n585998 , n585994 , n585997 );
and ( n58676 , n585990 , n585997 );
or ( n58677 , n585995 , n585998 , n58676 );
and ( n586001 , n58640 , n58677 );
xor ( n586002 , n58593 , n585920 );
xor ( n58680 , n586002 , n585923 );
and ( n58681 , n58677 , n58680 );
and ( n586005 , n58640 , n58680 );
or ( n586006 , n586001 , n58681 , n586005 );
and ( n586007 , n56909 , n52273 );
and ( n586008 , n56832 , n52271 );
nor ( n58686 , n586007 , n586008 );
xnor ( n586010 , n58686 , n52137 );
and ( n586011 , n586006 , n586010 );
xor ( n58689 , n585926 , n585930 );
xor ( n586013 , n58689 , n58610 );
and ( n586014 , n586010 , n586013 );
and ( n58692 , n586006 , n586013 );
or ( n586016 , n586011 , n586014 , n58692 );
and ( n586017 , n585936 , n586016 );
xor ( n58695 , n58393 , n585720 );
xor ( n58696 , n58695 , n58400 );
and ( n586020 , n586016 , n58696 );
and ( n586021 , n585936 , n58696 );
or ( n58699 , n586017 , n586020 , n586021 );
and ( n58700 , n583377 , n52509 );
and ( n586024 , n55841 , n52507 );
nor ( n586025 , n58700 , n586024 );
xnor ( n58703 , n586025 , n52383 );
and ( n58704 , n58699 , n58703 );
and ( n58705 , n583746 , n52432 );
and ( n58706 , n56282 , n52430 );
nor ( n58707 , n58705 , n58706 );
xnor ( n58708 , n58707 , n52255 );
and ( n58709 , n58703 , n58708 );
and ( n58710 , n58699 , n58708 );
or ( n586034 , n58704 , n58709 , n58710 );
xor ( n58712 , n58413 , n585740 );
xor ( n586036 , n58712 , n58422 );
and ( n586037 , n586034 , n586036 );
xor ( n58715 , n585792 , n58473 );
xor ( n58716 , n58715 , n58476 );
and ( n586040 , n586036 , n58716 );
and ( n58718 , n586034 , n58716 );
or ( n586042 , n586037 , n586040 , n58718 );
and ( n58720 , n55075 , n52978 );
and ( n586044 , n55058 , n52976 );
nor ( n586045 , n58720 , n586044 );
xnor ( n58723 , n586045 , n52680 );
and ( n586047 , n586042 , n58723 );
xor ( n58725 , n58479 , n58483 );
xor ( n58726 , n58725 , n58486 );
and ( n586050 , n58723 , n58726 );
and ( n58728 , n586042 , n58726 );
or ( n586052 , n586047 , n586050 , n58728 );
and ( n586053 , n54725 , n53177 );
and ( n58731 , n54553 , n53175 );
nor ( n586055 , n586053 , n58731 );
xnor ( n586056 , n586055 , n52827 );
and ( n58734 , n586052 , n586056 );
xor ( n586058 , n58489 , n585816 );
xor ( n586059 , n586058 , n585819 );
and ( n58737 , n586056 , n586059 );
and ( n58738 , n586052 , n586059 );
or ( n586062 , n58734 , n58737 , n58738 );
and ( n586063 , n53835 , n53683 );
and ( n58741 , n53837 , n53681 );
nor ( n58742 , n586063 , n58741 );
xnor ( n586066 , n58742 , n53118 );
and ( n586067 , n586062 , n586066 );
xor ( n58745 , n585822 , n58503 );
xor ( n58746 , n58745 , n58506 );
and ( n586070 , n586066 , n58746 );
and ( n58748 , n586062 , n58746 );
or ( n58749 , n586067 , n586070 , n58748 );
and ( n586073 , n53109 , n54532 );
and ( n586074 , n52934 , n54530 );
nor ( n58752 , n586073 , n586074 );
xnor ( n58753 , n58752 , n53769 );
and ( n586077 , n58749 , n58753 );
and ( n586078 , n53367 , n54414 );
and ( n58756 , n53107 , n54412 );
nor ( n58757 , n586078 , n58756 );
xnor ( n586081 , n58757 , n53650 );
and ( n586082 , n58753 , n586081 );
and ( n58760 , n58749 , n586081 );
or ( n586084 , n586077 , n586082 , n58760 );
and ( n58762 , n53639 , n53996 );
and ( n58763 , n53641 , n53994 );
nor ( n586087 , n58762 , n58763 );
xnor ( n586088 , n586087 , n53376 );
and ( n58766 , n54215 , n53468 );
and ( n586090 , n54055 , n53466 );
nor ( n58768 , n58766 , n586090 );
xnor ( n586092 , n58768 , n52945 );
and ( n58770 , n586088 , n586092 );
xor ( n58771 , n585768 , n58449 );
xor ( n58772 , n58771 , n58452 );
and ( n58773 , n586092 , n58772 );
and ( n58774 , n586088 , n58772 );
or ( n58775 , n58770 , n58773 , n58774 );
xor ( n58776 , n58455 , n585782 );
xor ( n58777 , n58776 , n58462 );
and ( n58778 , n58775 , n58777 );
and ( n58779 , n53641 , n53996 );
and ( n58780 , n53365 , n53994 );
nor ( n58781 , n58779 , n58780 );
xnor ( n58782 , n58781 , n53376 );
and ( n58783 , n54055 , n53468 );
and ( n58784 , n53835 , n53466 );
nor ( n58785 , n58783 , n58784 );
xnor ( n58786 , n58785 , n52945 );
xor ( n58787 , n58782 , n58786 );
xor ( n58788 , n585832 , n58513 );
xor ( n58789 , n58788 , n58516 );
xor ( n58790 , n58787 , n58789 );
and ( n58791 , n58777 , n58790 );
and ( n58792 , n58775 , n58790 );
or ( n58793 , n58778 , n58791 , n58792 );
and ( n586117 , n586084 , n58793 );
and ( n58795 , n52816 , n55013 );
and ( n586119 , n52818 , n55010 );
nor ( n586120 , n58795 , n586119 );
xnor ( n586121 , n586120 , n53762 );
and ( n58799 , n58793 , n586121 );
and ( n586123 , n586084 , n586121 );
or ( n586124 , n586117 , n58799 , n586123 );
and ( n586125 , n58782 , n58786 );
and ( n58803 , n58786 , n58789 );
and ( n586127 , n58782 , n58789 );
or ( n586128 , n586125 , n58803 , n586127 );
and ( n586129 , n52934 , n54532 );
and ( n58807 , n52936 , n54530 );
nor ( n586131 , n586129 , n58807 );
xnor ( n586132 , n586131 , n53769 );
and ( n58810 , n586128 , n586132 );
xor ( n586134 , n585788 , n585842 );
xor ( n58812 , n586134 , n585847 );
and ( n586136 , n586132 , n58812 );
and ( n586137 , n586128 , n58812 );
or ( n58815 , n58810 , n586136 , n586137 );
and ( n586139 , n586124 , n58815 );
xor ( n586140 , n585850 , n58531 );
xor ( n58818 , n586140 , n585859 );
and ( n586142 , n58815 , n58818 );
and ( n586143 , n586124 , n58818 );
or ( n58821 , n586139 , n586142 , n586143 );
xor ( n58822 , n585862 , n585882 );
xor ( n58823 , n58822 , n585885 );
and ( n586147 , n58821 , n58823 );
xor ( n586148 , n58362 , n58366 );
xor ( n586149 , n586148 , n58369 );
and ( n58827 , n58823 , n586149 );
and ( n586151 , n58821 , n586149 );
or ( n586152 , n586147 , n58827 , n586151 );
and ( n586153 , n58576 , n586152 );
xor ( n58831 , n58821 , n58823 );
xor ( n586155 , n58831 , n586149 );
and ( n58833 , n57058 , n52273 );
and ( n586157 , n56909 , n52271 );
nor ( n586158 , n58833 , n586157 );
xnor ( n58836 , n586158 , n52137 );
and ( n586160 , n57283 , n52155 );
and ( n586161 , n584529 , n52153 );
nor ( n58839 , n586160 , n586161 );
xnor ( n586163 , n58839 , n52085 );
and ( n586164 , n58836 , n586163 );
xor ( n58842 , n58640 , n58677 );
xor ( n58843 , n58842 , n58680 );
and ( n58844 , n586163 , n58843 );
and ( n586168 , n58836 , n58843 );
or ( n58846 , n586164 , n58844 , n586168 );
and ( n58847 , n583746 , n52509 );
and ( n58848 , n56282 , n52507 );
nor ( n58849 , n58847 , n58848 );
xnor ( n58850 , n58849 , n52383 );
and ( n58851 , n58846 , n58850 );
xor ( n58852 , n586006 , n586010 );
xor ( n58853 , n58852 , n586013 );
and ( n58854 , n58850 , n58853 );
and ( n586178 , n58846 , n58853 );
or ( n586179 , n58851 , n58854 , n586178 );
and ( n58857 , n56282 , n52509 );
and ( n586181 , n583377 , n52507 );
nor ( n58859 , n58857 , n586181 );
xnor ( n58860 , n58859 , n52383 );
and ( n58861 , n586179 , n58860 );
and ( n58862 , n583800 , n52432 );
and ( n58863 , n583746 , n52430 );
nor ( n586187 , n58862 , n58863 );
xnor ( n586188 , n586187 , n52255 );
and ( n58866 , n56832 , n52273 );
and ( n586190 , n56671 , n52271 );
nor ( n586191 , n58866 , n586190 );
xnor ( n58869 , n586191 , n52137 );
xor ( n586193 , n586188 , n58869 );
xor ( n586194 , n585936 , n586016 );
xor ( n58872 , n586194 , n58696 );
xor ( n586196 , n586193 , n58872 );
and ( n586197 , n58860 , n586196 );
and ( n586198 , n586179 , n586196 );
or ( n586199 , n58861 , n586197 , n586198 );
and ( n58877 , n55528 , n52978 );
and ( n586201 , n55293 , n52976 );
nor ( n586202 , n58877 , n586201 );
xnor ( n58880 , n586202 , n52680 );
and ( n586204 , n586199 , n58880 );
xor ( n586205 , n58699 , n58703 );
xor ( n58883 , n586205 , n58708 );
and ( n58884 , n58880 , n58883 );
and ( n586208 , n586199 , n58883 );
or ( n586209 , n586204 , n58884 , n586208 );
and ( n58887 , n55058 , n53177 );
and ( n58888 , n54893 , n53175 );
nor ( n586212 , n58887 , n58888 );
xnor ( n586213 , n586212 , n52827 );
and ( n586214 , n586209 , n586213 );
xor ( n58892 , n586034 , n586036 );
xor ( n586216 , n58892 , n58716 );
and ( n586217 , n586213 , n586216 );
and ( n586218 , n586209 , n586216 );
or ( n58896 , n586214 , n586217 , n586218 );
and ( n586220 , n54553 , n53468 );
and ( n586221 , n54321 , n53466 );
nor ( n58899 , n586220 , n586221 );
xnor ( n586223 , n58899 , n52945 );
and ( n586224 , n58896 , n586223 );
xor ( n586225 , n586042 , n58723 );
xor ( n586226 , n586225 , n58726 );
and ( n58904 , n586223 , n586226 );
and ( n586228 , n58896 , n586226 );
or ( n586229 , n586224 , n58904 , n586228 );
and ( n58907 , n54055 , n53683 );
and ( n586231 , n53835 , n53681 );
nor ( n586232 , n58907 , n586231 );
xnor ( n58910 , n586232 , n53118 );
and ( n586234 , n586229 , n58910 );
xor ( n586235 , n586052 , n586056 );
xor ( n58913 , n586235 , n586059 );
and ( n58914 , n58910 , n58913 );
and ( n58915 , n586229 , n58913 );
or ( n586239 , n586234 , n58914 , n58915 );
and ( n586240 , n586188 , n58869 );
and ( n58918 , n58869 , n58872 );
and ( n586242 , n586188 , n58872 );
or ( n586243 , n586240 , n58918 , n586242 );
and ( n58921 , n583048 , n52707 );
and ( n586245 , n582961 , n52705 );
nor ( n586246 , n58921 , n586245 );
xnor ( n58924 , n586246 , n52526 );
and ( n586248 , n586243 , n58924 );
xor ( n586249 , n585726 , n585730 );
xor ( n58927 , n586249 , n585733 );
and ( n586251 , n58924 , n58927 );
and ( n586252 , n586243 , n58927 );
or ( n586253 , n586248 , n586251 , n586252 );
and ( n586254 , n55293 , n52978 );
and ( n58932 , n55075 , n52976 );
nor ( n586256 , n586254 , n58932 );
xnor ( n586257 , n586256 , n52680 );
and ( n58935 , n586253 , n586257 );
and ( n586259 , n582961 , n52707 );
and ( n586260 , n55528 , n52705 );
nor ( n58938 , n586259 , n586260 );
xnor ( n58939 , n58938 , n52526 );
and ( n586263 , n586257 , n58939 );
and ( n586264 , n586253 , n58939 );
or ( n58942 , n58935 , n586263 , n586264 );
and ( n58943 , n54893 , n53177 );
and ( n586267 , n54725 , n53175 );
nor ( n586268 , n58943 , n586267 );
xnor ( n58946 , n586268 , n52827 );
and ( n58947 , n58942 , n58946 );
xor ( n58948 , n58425 , n585752 );
xor ( n586272 , n58948 , n585755 );
and ( n58950 , n58946 , n586272 );
and ( n58951 , n58942 , n586272 );
or ( n58952 , n58947 , n58950 , n58951 );
and ( n586276 , n54321 , n53468 );
and ( n586277 , n54215 , n53466 );
nor ( n58955 , n586276 , n586277 );
xnor ( n586279 , n58955 , n52945 );
and ( n586280 , n58952 , n586279 );
xor ( n586281 , n585758 , n58439 );
xor ( n58959 , n586281 , n585765 );
and ( n586283 , n586279 , n58959 );
and ( n58961 , n58952 , n58959 );
or ( n58962 , n586280 , n586283 , n58961 );
and ( n58963 , n586239 , n58962 );
and ( n58964 , n53365 , n54414 );
and ( n58965 , n53367 , n54412 );
nor ( n58966 , n58964 , n58965 );
xnor ( n586290 , n58966 , n53650 );
and ( n586291 , n58962 , n586290 );
and ( n58969 , n586239 , n586290 );
or ( n586293 , n58963 , n586291 , n58969 );
and ( n58971 , n52934 , n55013 );
and ( n586295 , n52936 , n55010 );
nor ( n58973 , n58971 , n586295 );
xnor ( n58974 , n58973 , n53762 );
and ( n586298 , n53107 , n54532 );
and ( n58976 , n53109 , n54530 );
nor ( n586300 , n586298 , n58976 );
xnor ( n586301 , n586300 , n53769 );
and ( n58979 , n58974 , n586301 );
xor ( n586303 , n586088 , n586092 );
xor ( n586304 , n586303 , n58772 );
and ( n586305 , n586301 , n586304 );
and ( n586306 , n58974 , n586304 );
or ( n58984 , n58979 , n586305 , n586306 );
and ( n586308 , n586293 , n58984 );
and ( n586309 , n52936 , n55013 );
and ( n58987 , n52816 , n55010 );
nor ( n586311 , n586309 , n58987 );
xnor ( n586312 , n586311 , n53762 );
and ( n58990 , n58984 , n586312 );
and ( n586314 , n586293 , n586312 );
or ( n586315 , n586308 , n58990 , n586314 );
xor ( n58993 , n586128 , n586132 );
xor ( n58994 , n58993 , n58812 );
and ( n586318 , n586315 , n58994 );
xor ( n586319 , n585866 , n585868 );
xor ( n58997 , n586319 , n585871 );
and ( n586321 , n58994 , n58997 );
and ( n586322 , n586315 , n58997 );
or ( n59000 , n586318 , n586321 , n586322 );
xor ( n586324 , n586124 , n58815 );
xor ( n586325 , n586324 , n58818 );
and ( n59003 , n59000 , n586325 );
xor ( n586327 , n58551 , n585876 );
xor ( n586328 , n586327 , n585879 );
and ( n59006 , n586325 , n586328 );
and ( n586330 , n59000 , n586328 );
or ( n586331 , n59003 , n59006 , n586330 );
and ( n59009 , n586155 , n586331 );
xor ( n586333 , n59000 , n586325 );
xor ( n59011 , n586333 , n586328 );
and ( n59012 , n53641 , n54414 );
and ( n59013 , n53365 , n54412 );
nor ( n59014 , n59012 , n59013 );
xnor ( n59015 , n59014 , n53650 );
and ( n59016 , n53837 , n53996 );
and ( n59017 , n53639 , n53994 );
nor ( n59018 , n59016 , n59017 );
xnor ( n59019 , n59018 , n53376 );
and ( n586343 , n59015 , n59019 );
xor ( n586344 , n58952 , n586279 );
xor ( n586345 , n586344 , n58959 );
and ( n59023 , n59019 , n586345 );
and ( n586347 , n59015 , n586345 );
or ( n586348 , n586343 , n59023 , n586347 );
xor ( n586349 , n586239 , n58962 );
xor ( n586350 , n586349 , n586290 );
and ( n59028 , n586348 , n586350 );
xor ( n586352 , n586062 , n586066 );
xor ( n586353 , n586352 , n58746 );
and ( n59031 , n586350 , n586353 );
and ( n586355 , n586348 , n586353 );
or ( n586356 , n59028 , n59031 , n586355 );
xor ( n59034 , n58749 , n58753 );
xor ( n586358 , n59034 , n586081 );
and ( n586359 , n586356 , n586358 );
xor ( n59037 , n58775 , n58777 );
xor ( n586361 , n59037 , n58790 );
and ( n586362 , n586358 , n586361 );
and ( n586363 , n586356 , n586361 );
or ( n586364 , n586359 , n586362 , n586363 );
xor ( n59042 , n586084 , n58793 );
xor ( n586366 , n59042 , n586121 );
and ( n586367 , n586364 , n586366 );
xor ( n59045 , n586315 , n58994 );
xor ( n586369 , n59045 , n58997 );
and ( n586370 , n586366 , n586369 );
and ( n59048 , n586364 , n586369 );
or ( n586372 , n586367 , n586370 , n59048 );
and ( n586373 , n59011 , n586372 );
xor ( n59051 , n586364 , n586366 );
xor ( n59052 , n59051 , n586369 );
and ( n59053 , n585586 , n51991 );
and ( n586377 , n58246 , n51989 );
nor ( n586378 , n59053 , n586377 );
xnor ( n59056 , n586378 , n51959 );
and ( n59057 , n58623 , n51936 );
and ( n586381 , n585909 , n51934 );
nor ( n586382 , n59057 , n586381 );
xnor ( n59060 , n586382 , n51941 );
and ( n59061 , n59056 , n59060 );
and ( n586385 , n585973 , n51927 );
nor ( n586386 , n51929 , n586385 );
not ( n586387 , n586386 );
and ( n586388 , n59060 , n586387 );
and ( n59066 , n59056 , n586387 );
or ( n586390 , n59061 , n586388 , n59066 );
and ( n59068 , n585221 , n52065 );
and ( n59069 , n57900 , n52063 );
nor ( n59070 , n59068 , n59069 );
xnor ( n586394 , n59070 , n52022 );
and ( n586395 , n586390 , n586394 );
xor ( n59073 , n585967 , n585971 );
xor ( n586397 , n59073 , n58654 );
and ( n59075 , n586394 , n586397 );
and ( n586399 , n586390 , n586397 );
or ( n59077 , n586395 , n59075 , n586399 );
and ( n59078 , n57482 , n52155 );
and ( n59079 , n57484 , n52153 );
nor ( n59080 , n59078 , n59079 );
xnor ( n59081 , n59080 , n52085 );
and ( n586405 , n59077 , n59081 );
xor ( n586406 , n585980 , n585984 );
xor ( n59084 , n586406 , n585987 );
and ( n586408 , n59081 , n59084 );
and ( n59086 , n59077 , n59084 );
or ( n59087 , n586405 , n586408 , n59086 );
and ( n586411 , n584529 , n52273 );
and ( n59089 , n57058 , n52271 );
nor ( n586413 , n586411 , n59089 );
xnor ( n59091 , n586413 , n52137 );
and ( n59092 , n59087 , n59091 );
xor ( n586416 , n585990 , n585994 );
xor ( n586417 , n586416 , n585997 );
and ( n59095 , n59091 , n586417 );
and ( n586419 , n59087 , n586417 );
or ( n59097 , n59092 , n59095 , n586419 );
and ( n586421 , n585909 , n51991 );
and ( n586422 , n585586 , n51989 );
nor ( n59100 , n586421 , n586422 );
xnor ( n586424 , n59100 , n51959 );
and ( n59102 , n585973 , n51936 );
and ( n59103 , n58623 , n51934 );
nor ( n59104 , n59102 , n59103 );
xnor ( n59105 , n59104 , n51941 );
and ( n59106 , n586424 , n59105 );
nor ( n59107 , n51929 , n51927 );
not ( n59108 , n59107 );
and ( n59109 , n59105 , n59108 );
and ( n59110 , n586424 , n59108 );
or ( n59111 , n59106 , n59109 , n59110 );
and ( n59112 , n58219 , n52065 );
and ( n59113 , n585221 , n52063 );
nor ( n59114 , n59112 , n59113 );
xnor ( n586438 , n59114 , n52022 );
and ( n59116 , n59111 , n586438 );
xor ( n586440 , n59056 , n59060 );
xor ( n586441 , n586440 , n586387 );
and ( n59119 , n586438 , n586441 );
and ( n586443 , n59111 , n586441 );
or ( n586444 , n59116 , n59119 , n586443 );
and ( n59122 , n585062 , n52155 );
and ( n586446 , n57482 , n52153 );
nor ( n586447 , n59122 , n586446 );
xnor ( n586448 , n586447 , n52085 );
and ( n586449 , n586444 , n586448 );
xor ( n59127 , n586390 , n586394 );
xor ( n586451 , n59127 , n586397 );
and ( n586452 , n586448 , n586451 );
and ( n59130 , n586444 , n586451 );
or ( n586454 , n586449 , n586452 , n59130 );
and ( n586455 , n58623 , n51991 );
and ( n59133 , n585909 , n51989 );
nor ( n586457 , n586455 , n59133 );
xnor ( n586458 , n586457 , n51959 );
and ( n59136 , n585973 , n51934 );
nor ( n586460 , n51936 , n59136 );
xnor ( n586461 , n586460 , n51941 );
and ( n586462 , n586458 , n586461 );
nor ( n586463 , n51929 , n51927 );
not ( n59141 , n586463 );
and ( n586465 , n586461 , n59141 );
and ( n586466 , n586458 , n59141 );
or ( n586467 , n586462 , n586465 , n586466 );
and ( n586468 , n58246 , n52065 );
and ( n59146 , n58219 , n52063 );
nor ( n586470 , n586468 , n59146 );
xnor ( n586471 , n586470 , n52022 );
and ( n59149 , n586467 , n586471 );
xor ( n586473 , n586424 , n59105 );
xor ( n586474 , n586473 , n59108 );
and ( n59152 , n586471 , n586474 );
and ( n586476 , n586467 , n586474 );
or ( n586477 , n59149 , n59152 , n586476 );
and ( n59155 , n57900 , n52155 );
and ( n586479 , n585062 , n52153 );
nor ( n586480 , n59155 , n586479 );
xnor ( n59158 , n586480 , n52085 );
and ( n59159 , n586477 , n59158 );
xor ( n59160 , n59111 , n586438 );
xor ( n586484 , n59160 , n586441 );
and ( n586485 , n59158 , n586484 );
and ( n59163 , n586477 , n586484 );
or ( n59164 , n59159 , n586485 , n59163 );
and ( n59165 , n57484 , n52273 );
and ( n586489 , n57283 , n52271 );
nor ( n586490 , n59165 , n586489 );
xnor ( n59168 , n586490 , n52137 );
and ( n586492 , n59164 , n59168 );
xor ( n586493 , n586444 , n586448 );
xor ( n59171 , n586493 , n586451 );
and ( n59172 , n59168 , n59171 );
and ( n59173 , n59164 , n59171 );
or ( n59174 , n586492 , n59172 , n59173 );
and ( n586498 , n586454 , n59174 );
xor ( n59176 , n59077 , n59081 );
xor ( n59177 , n59176 , n59084 );
and ( n59178 , n59174 , n59177 );
and ( n59179 , n586454 , n59177 );
or ( n586503 , n586498 , n59178 , n59179 );
and ( n59181 , n56909 , n52432 );
and ( n59182 , n56832 , n52430 );
nor ( n59183 , n59181 , n59182 );
xnor ( n59184 , n59183 , n52255 );
and ( n59185 , n586503 , n59184 );
xor ( n59186 , n59087 , n59091 );
xor ( n59187 , n59186 , n586417 );
and ( n59188 , n59184 , n59187 );
and ( n59189 , n586503 , n59187 );
or ( n59190 , n59185 , n59188 , n59189 );
and ( n586514 , n59097 , n59190 );
xor ( n59192 , n58836 , n586163 );
xor ( n586516 , n59192 , n58843 );
and ( n586517 , n59190 , n586516 );
and ( n59195 , n59097 , n586516 );
or ( n586519 , n586514 , n586517 , n59195 );
and ( n586520 , n56671 , n52432 );
and ( n59198 , n583800 , n52430 );
nor ( n586522 , n586520 , n59198 );
xnor ( n59200 , n586522 , n52255 );
and ( n59201 , n586519 , n59200 );
xor ( n586525 , n58846 , n58850 );
xor ( n59203 , n586525 , n58853 );
and ( n586527 , n59200 , n59203 );
and ( n59205 , n586519 , n59203 );
or ( n586529 , n59201 , n586527 , n59205 );
and ( n59207 , n55293 , n53177 );
and ( n586531 , n55075 , n53175 );
nor ( n586532 , n59207 , n586531 );
xnor ( n59210 , n586532 , n52827 );
and ( n59211 , n586529 , n59210 );
and ( n59212 , n55841 , n52707 );
and ( n586536 , n583048 , n52705 );
nor ( n586537 , n59212 , n586536 );
xnor ( n586538 , n586537 , n52526 );
and ( n586539 , n59210 , n586538 );
and ( n59217 , n586529 , n586538 );
or ( n586541 , n59211 , n586539 , n59217 );
and ( n59219 , n55075 , n53177 );
and ( n586543 , n55058 , n53175 );
nor ( n59221 , n59219 , n586543 );
xnor ( n59222 , n59221 , n52827 );
and ( n586546 , n586541 , n59222 );
xor ( n59224 , n586243 , n58924 );
xor ( n586548 , n59224 , n58927 );
and ( n586549 , n59222 , n586548 );
and ( n59227 , n586541 , n586548 );
or ( n586551 , n586546 , n586549 , n59227 );
and ( n586552 , n54725 , n53468 );
and ( n59230 , n54553 , n53466 );
nor ( n586554 , n586552 , n59230 );
xnor ( n586555 , n586554 , n52945 );
and ( n59233 , n586551 , n586555 );
xor ( n586557 , n586253 , n586257 );
xor ( n586558 , n586557 , n58939 );
and ( n59236 , n586555 , n586558 );
and ( n586560 , n586551 , n586558 );
or ( n586561 , n59233 , n59236 , n586560 );
and ( n59239 , n54215 , n53683 );
and ( n586563 , n54055 , n53681 );
nor ( n586564 , n59239 , n586563 );
xnor ( n586565 , n586564 , n53118 );
and ( n586566 , n586561 , n586565 );
xor ( n59244 , n58942 , n58946 );
xor ( n586568 , n59244 , n586272 );
and ( n586569 , n586565 , n586568 );
and ( n59247 , n586561 , n586568 );
or ( n586571 , n586566 , n586569 , n59247 );
and ( n586572 , n53109 , n55013 );
and ( n59250 , n52934 , n55010 );
nor ( n59251 , n586572 , n59250 );
xnor ( n586575 , n59251 , n53762 );
and ( n586576 , n586571 , n586575 );
and ( n59254 , n53367 , n54532 );
and ( n59255 , n53107 , n54530 );
nor ( n586579 , n59254 , n59255 );
xnor ( n586580 , n586579 , n53769 );
and ( n59258 , n586575 , n586580 );
and ( n59259 , n586571 , n586580 );
or ( n586583 , n586576 , n59258 , n59259 );
and ( n586584 , n53639 , n54414 );
and ( n59262 , n53641 , n54412 );
nor ( n59263 , n586584 , n59262 );
xnor ( n586587 , n59263 , n53650 );
and ( n586588 , n53835 , n53996 );
and ( n586589 , n53837 , n53994 );
nor ( n59267 , n586588 , n586589 );
xnor ( n586591 , n59267 , n53376 );
and ( n59269 , n586587 , n586591 );
xor ( n59270 , n58896 , n586223 );
xor ( n59271 , n59270 , n586226 );
and ( n59272 , n586591 , n59271 );
and ( n586596 , n586587 , n59271 );
or ( n59274 , n59269 , n59272 , n586596 );
xor ( n59275 , n586229 , n58910 );
xor ( n586599 , n59275 , n58913 );
and ( n59277 , n59274 , n586599 );
xor ( n586601 , n59015 , n59019 );
xor ( n586602 , n586601 , n586345 );
and ( n59280 , n586599 , n586602 );
and ( n59281 , n59274 , n586602 );
or ( n586605 , n59277 , n59280 , n59281 );
and ( n586606 , n586583 , n586605 );
xor ( n59284 , n58974 , n586301 );
xor ( n59285 , n59284 , n586304 );
and ( n59286 , n586605 , n59285 );
and ( n59287 , n586583 , n59285 );
or ( n586611 , n586606 , n59286 , n59287 );
xor ( n586612 , n586293 , n58984 );
xor ( n59290 , n586612 , n586312 );
and ( n59291 , n586611 , n59290 );
xor ( n59292 , n586356 , n586358 );
xor ( n59293 , n59292 , n586361 );
and ( n59294 , n59290 , n59293 );
and ( n586618 , n586611 , n59293 );
or ( n586619 , n59291 , n59294 , n586618 );
and ( n59297 , n59052 , n586619 );
and ( n586621 , n57058 , n52432 );
and ( n586622 , n56909 , n52430 );
nor ( n59300 , n586621 , n586622 );
xnor ( n59301 , n59300 , n52255 );
and ( n586625 , n57283 , n52273 );
and ( n59303 , n584529 , n52271 );
nor ( n59304 , n586625 , n59303 );
xnor ( n59305 , n59304 , n52137 );
and ( n59306 , n59301 , n59305 );
xor ( n586630 , n586454 , n59174 );
xor ( n59308 , n586630 , n59177 );
and ( n59309 , n59305 , n59308 );
and ( n59310 , n59301 , n59308 );
or ( n59311 , n59306 , n59309 , n59310 );
and ( n59312 , n583746 , n52707 );
and ( n59313 , n56282 , n52705 );
nor ( n59314 , n59312 , n59313 );
xnor ( n59315 , n59314 , n52526 );
and ( n59316 , n59311 , n59315 );
xor ( n586640 , n586503 , n59184 );
xor ( n59318 , n586640 , n59187 );
and ( n586642 , n59315 , n59318 );
and ( n59320 , n59311 , n59318 );
or ( n586644 , n59316 , n586642 , n59320 );
and ( n59322 , n55841 , n52978 );
and ( n59323 , n583048 , n52976 );
nor ( n586647 , n59322 , n59323 );
xnor ( n59325 , n586647 , n52680 );
and ( n586649 , n586644 , n59325 );
and ( n586650 , n56282 , n52707 );
and ( n59328 , n583377 , n52705 );
nor ( n586652 , n586650 , n59328 );
xnor ( n586653 , n586652 , n52526 );
and ( n59331 , n59325 , n586653 );
and ( n59332 , n586644 , n586653 );
or ( n586656 , n586649 , n59331 , n59332 );
and ( n586657 , n55528 , n53177 );
and ( n59335 , n55293 , n53175 );
nor ( n59336 , n586657 , n59335 );
xnor ( n586660 , n59336 , n52827 );
and ( n59338 , n586656 , n586660 );
xor ( n586662 , n586519 , n59200 );
xor ( n586663 , n586662 , n59203 );
and ( n59341 , n586660 , n586663 );
and ( n586665 , n586656 , n586663 );
or ( n586666 , n59338 , n59341 , n586665 );
and ( n59344 , n55058 , n53468 );
and ( n586668 , n54893 , n53466 );
nor ( n586669 , n59344 , n586668 );
xnor ( n59347 , n586669 , n52945 );
and ( n586671 , n586666 , n59347 );
xor ( n586672 , n586529 , n59210 );
xor ( n59350 , n586672 , n586538 );
and ( n59351 , n59347 , n59350 );
and ( n586675 , n586666 , n59350 );
or ( n586676 , n586671 , n59351 , n586675 );
and ( n59354 , n54553 , n53683 );
and ( n586678 , n54321 , n53681 );
nor ( n586679 , n59354 , n586678 );
xnor ( n59357 , n586679 , n53118 );
and ( n586681 , n586676 , n59357 );
xor ( n586682 , n586541 , n59222 );
xor ( n59360 , n586682 , n586548 );
and ( n586684 , n59357 , n59360 );
and ( n586685 , n586676 , n59360 );
or ( n59363 , n586681 , n586684 , n586685 );
and ( n586687 , n53837 , n54414 );
and ( n586688 , n53639 , n54412 );
nor ( n586689 , n586687 , n586688 );
xnor ( n586690 , n586689 , n53650 );
and ( n59368 , n59363 , n586690 );
and ( n586692 , n54055 , n53996 );
and ( n586693 , n53835 , n53994 );
nor ( n586694 , n586692 , n586693 );
xnor ( n586695 , n586694 , n53376 );
and ( n59373 , n586690 , n586695 );
and ( n586697 , n59363 , n586695 );
or ( n586698 , n59368 , n59373 , n586697 );
and ( n59376 , n583800 , n52509 );
and ( n586700 , n583746 , n52507 );
nor ( n586701 , n59376 , n586700 );
xnor ( n59379 , n586701 , n52383 );
and ( n586703 , n56832 , n52432 );
and ( n586704 , n56671 , n52430 );
nor ( n59382 , n586703 , n586704 );
xnor ( n59383 , n59382 , n52255 );
and ( n586707 , n59379 , n59383 );
xor ( n59385 , n59097 , n59190 );
xor ( n59386 , n59385 , n586516 );
and ( n59387 , n59383 , n59386 );
and ( n59388 , n59379 , n59386 );
or ( n59389 , n586707 , n59387 , n59388 );
and ( n59390 , n583048 , n52978 );
and ( n59391 , n582961 , n52976 );
nor ( n59392 , n59390 , n59391 );
xnor ( n59393 , n59392 , n52680 );
and ( n59394 , n59389 , n59393 );
and ( n59395 , n583377 , n52707 );
and ( n59396 , n55841 , n52705 );
nor ( n59397 , n59395 , n59396 );
xnor ( n59398 , n59397 , n52526 );
and ( n586722 , n59393 , n59398 );
and ( n59400 , n59389 , n59398 );
or ( n586724 , n59394 , n586722 , n59400 );
and ( n59402 , n582961 , n52978 );
and ( n586726 , n55528 , n52976 );
nor ( n59404 , n59402 , n586726 );
xnor ( n59405 , n59404 , n52680 );
and ( n586729 , n586724 , n59405 );
xor ( n586730 , n586179 , n58860 );
xor ( n59408 , n586730 , n586196 );
and ( n59409 , n59405 , n59408 );
and ( n59410 , n586724 , n59408 );
or ( n59411 , n586729 , n59409 , n59410 );
and ( n59412 , n54893 , n53468 );
and ( n59413 , n54725 , n53466 );
nor ( n586737 , n59412 , n59413 );
xnor ( n59415 , n586737 , n52945 );
and ( n586739 , n59411 , n59415 );
xor ( n59417 , n586199 , n58880 );
xor ( n59418 , n59417 , n58883 );
and ( n59419 , n59415 , n59418 );
and ( n59420 , n59411 , n59418 );
or ( n59421 , n586739 , n59419 , n59420 );
and ( n59422 , n54321 , n53683 );
and ( n59423 , n54215 , n53681 );
nor ( n586747 , n59422 , n59423 );
xnor ( n586748 , n586747 , n53118 );
and ( n59426 , n59421 , n586748 );
xor ( n586750 , n586209 , n586213 );
xor ( n586751 , n586750 , n586216 );
and ( n586752 , n586748 , n586751 );
and ( n586753 , n59421 , n586751 );
or ( n59431 , n59426 , n586752 , n586753 );
and ( n586755 , n586698 , n59431 );
and ( n586756 , n53365 , n54532 );
and ( n59434 , n53367 , n54530 );
nor ( n586758 , n586756 , n59434 );
xnor ( n59436 , n586758 , n53769 );
and ( n586760 , n59431 , n59436 );
and ( n59438 , n586698 , n59436 );
or ( n59439 , n586755 , n586760 , n59438 );
and ( n586763 , n53107 , n55013 );
and ( n586764 , n53109 , n55010 );
nor ( n59442 , n586763 , n586764 );
xnor ( n586766 , n59442 , n53762 );
xor ( n586767 , n586561 , n586565 );
xor ( n59445 , n586767 , n586568 );
and ( n586769 , n586766 , n59445 );
xor ( n586770 , n586587 , n586591 );
xor ( n59448 , n586770 , n59271 );
and ( n586772 , n59445 , n59448 );
and ( n586773 , n586766 , n59448 );
or ( n586774 , n586769 , n586772 , n586773 );
and ( n59452 , n59439 , n586774 );
xor ( n586776 , n586571 , n586575 );
xor ( n586777 , n586776 , n586580 );
and ( n59455 , n586774 , n586777 );
and ( n586779 , n59439 , n586777 );
or ( n586780 , n59452 , n59455 , n586779 );
xor ( n59458 , n586348 , n586350 );
xor ( n586782 , n59458 , n586353 );
and ( n586783 , n586780 , n586782 );
xor ( n59461 , n586583 , n586605 );
xor ( n59462 , n59461 , n59285 );
and ( n586786 , n586782 , n59462 );
and ( n586787 , n586780 , n59462 );
or ( n59465 , n586783 , n586786 , n586787 );
xor ( n586789 , n586611 , n59290 );
xor ( n586790 , n586789 , n59293 );
and ( n59468 , n59465 , n586790 );
xor ( n586792 , n586780 , n586782 );
xor ( n586793 , n586792 , n59462 );
and ( n59471 , n585973 , n51991 );
and ( n586795 , n58623 , n51989 );
nor ( n586796 , n59471 , n586795 );
xnor ( n59474 , n586796 , n51959 );
nor ( n586798 , n51936 , n51934 );
xnor ( n59476 , n586798 , n51941 );
and ( n59477 , n59474 , n59476 );
nor ( n59478 , n51929 , n51927 );
not ( n59479 , n59478 );
and ( n59480 , n59476 , n59479 );
and ( n59481 , n59474 , n59479 );
or ( n59482 , n59477 , n59480 , n59481 );
and ( n59483 , n585586 , n52065 );
and ( n586807 , n58246 , n52063 );
nor ( n59485 , n59483 , n586807 );
xnor ( n586809 , n59485 , n52022 );
and ( n586810 , n59482 , n586809 );
xor ( n586811 , n586458 , n586461 );
xor ( n59489 , n586811 , n59141 );
and ( n586813 , n586809 , n59489 );
and ( n59491 , n59482 , n59489 );
or ( n59492 , n586810 , n586813 , n59491 );
and ( n59493 , n585221 , n52155 );
and ( n59494 , n57900 , n52153 );
nor ( n59495 , n59493 , n59494 );
xnor ( n59496 , n59495 , n52085 );
and ( n59497 , n59492 , n59496 );
xor ( n586821 , n586467 , n586471 );
xor ( n59499 , n586821 , n586474 );
and ( n59500 , n59496 , n59499 );
and ( n586824 , n59492 , n59499 );
or ( n59502 , n59497 , n59500 , n586824 );
and ( n59503 , n57482 , n52273 );
and ( n59504 , n57484 , n52271 );
nor ( n586828 , n59503 , n59504 );
xnor ( n59506 , n586828 , n52137 );
and ( n59507 , n59502 , n59506 );
xor ( n59508 , n586477 , n59158 );
xor ( n586832 , n59508 , n586484 );
and ( n586833 , n59506 , n586832 );
and ( n59511 , n59502 , n586832 );
or ( n586835 , n59507 , n586833 , n59511 );
and ( n586836 , n584529 , n52432 );
and ( n586837 , n57058 , n52430 );
nor ( n59515 , n586836 , n586837 );
xnor ( n586839 , n59515 , n52255 );
and ( n59517 , n586835 , n586839 );
xor ( n59518 , n59164 , n59168 );
xor ( n59519 , n59518 , n59171 );
and ( n59520 , n586839 , n59519 );
and ( n59521 , n586835 , n59519 );
or ( n59522 , n59517 , n59520 , n59521 );
and ( n59523 , n56832 , n52509 );
and ( n59524 , n56671 , n52507 );
nor ( n59525 , n59523 , n59524 );
xnor ( n59526 , n59525 , n52383 );
and ( n586850 , n59522 , n59526 );
xor ( n59528 , n59301 , n59305 );
xor ( n59529 , n59528 , n59308 );
and ( n586853 , n59526 , n59529 );
and ( n59531 , n59522 , n59529 );
or ( n586855 , n586850 , n586853 , n59531 );
and ( n59533 , n583377 , n52978 );
and ( n586857 , n55841 , n52976 );
nor ( n59535 , n59533 , n586857 );
xnor ( n586859 , n59535 , n52680 );
and ( n586860 , n586855 , n586859 );
and ( n59538 , n56671 , n52509 );
and ( n586862 , n583800 , n52507 );
nor ( n59540 , n59538 , n586862 );
xnor ( n586864 , n59540 , n52383 );
and ( n586865 , n586859 , n586864 );
and ( n59543 , n586855 , n586864 );
or ( n586867 , n586860 , n586865 , n59543 );
and ( n586868 , n55293 , n53468 );
and ( n59546 , n55075 , n53466 );
nor ( n59547 , n586868 , n59546 );
xnor ( n586871 , n59547 , n52945 );
and ( n59549 , n586867 , n586871 );
xor ( n586873 , n59379 , n59383 );
xor ( n59551 , n586873 , n59386 );
and ( n586875 , n586871 , n59551 );
and ( n586876 , n586867 , n59551 );
or ( n59554 , n59549 , n586875 , n586876 );
and ( n586878 , n55075 , n53468 );
and ( n586879 , n55058 , n53466 );
nor ( n59557 , n586878 , n586879 );
xnor ( n59558 , n59557 , n52945 );
and ( n586882 , n59554 , n59558 );
xor ( n59560 , n59389 , n59393 );
xor ( n59561 , n59560 , n59398 );
and ( n59562 , n59558 , n59561 );
and ( n59563 , n59554 , n59561 );
or ( n586887 , n586882 , n59562 , n59563 );
and ( n586888 , n54725 , n53683 );
and ( n59566 , n54553 , n53681 );
nor ( n586890 , n586888 , n59566 );
xnor ( n59568 , n586890 , n53118 );
and ( n586892 , n586887 , n59568 );
xor ( n59570 , n586724 , n59405 );
xor ( n59571 , n59570 , n59408 );
and ( n586895 , n59568 , n59571 );
and ( n586896 , n586887 , n59571 );
or ( n59574 , n586892 , n586895 , n586896 );
and ( n59575 , n53835 , n54414 );
and ( n586899 , n53837 , n54412 );
nor ( n586900 , n59575 , n586899 );
xnor ( n59578 , n586900 , n53650 );
and ( n59579 , n59574 , n59578 );
xor ( n586903 , n59411 , n59415 );
xor ( n586904 , n586903 , n59418 );
and ( n59582 , n59578 , n586904 );
and ( n59583 , n59574 , n586904 );
or ( n586907 , n59579 , n59582 , n59583 );
and ( n586908 , n53639 , n54532 );
and ( n59586 , n53641 , n54530 );
nor ( n59587 , n586908 , n59586 );
xnor ( n586911 , n59587 , n53769 );
and ( n59589 , n54215 , n53996 );
and ( n59590 , n54055 , n53994 );
nor ( n59591 , n59589 , n59590 );
xnor ( n59592 , n59591 , n53376 );
and ( n586916 , n586911 , n59592 );
xor ( n586917 , n586676 , n59357 );
xor ( n59595 , n586917 , n59360 );
and ( n586919 , n59592 , n59595 );
and ( n586920 , n586911 , n59595 );
or ( n59598 , n586916 , n586919 , n586920 );
and ( n59599 , n586907 , n59598 );
and ( n586923 , n53367 , n55013 );
and ( n59601 , n53107 , n55010 );
nor ( n59602 , n586923 , n59601 );
xnor ( n586926 , n59602 , n53762 );
and ( n586927 , n59598 , n586926 );
and ( n586928 , n586907 , n586926 );
or ( n59606 , n59599 , n586927 , n586928 );
and ( n586930 , n53641 , n54532 );
and ( n586931 , n53365 , n54530 );
nor ( n586932 , n586930 , n586931 );
xnor ( n59610 , n586932 , n53769 );
xor ( n586934 , n586551 , n586555 );
xor ( n586935 , n586934 , n586558 );
and ( n59613 , n59610 , n586935 );
xor ( n586937 , n59421 , n586748 );
xor ( n586938 , n586937 , n586751 );
and ( n59616 , n586935 , n586938 );
and ( n59617 , n59610 , n586938 );
or ( n59618 , n59613 , n59616 , n59617 );
and ( n59619 , n59606 , n59618 );
xor ( n586943 , n586698 , n59431 );
xor ( n586944 , n586943 , n59436 );
and ( n59622 , n59618 , n586944 );
and ( n586946 , n59606 , n586944 );
or ( n586947 , n59619 , n59622 , n586946 );
xor ( n586948 , n59439 , n586774 );
xor ( n59626 , n586948 , n586777 );
and ( n586950 , n586947 , n59626 );
xor ( n586951 , n59274 , n586599 );
xor ( n586952 , n586951 , n586602 );
and ( n59630 , n59626 , n586952 );
and ( n59631 , n586947 , n586952 );
or ( n586955 , n586950 , n59630 , n59631 );
and ( n59633 , n586793 , n586955 );
xor ( n59634 , n586947 , n59626 );
xor ( n59635 , n59634 , n586952 );
and ( n59636 , n585973 , n51989 );
nor ( n59637 , n51991 , n59636 );
xnor ( n59638 , n59637 , n51959 );
nor ( n59639 , n51936 , n51934 );
xnor ( n59640 , n59639 , n51941 );
and ( n59641 , n59638 , n59640 );
nor ( n59642 , n51929 , n51927 );
not ( n59643 , n59642 );
and ( n59644 , n59640 , n59643 );
and ( n59645 , n59638 , n59643 );
or ( n59646 , n59641 , n59644 , n59645 );
and ( n586970 , n585909 , n52065 );
and ( n59648 , n585586 , n52063 );
nor ( n586972 , n586970 , n59648 );
xnor ( n59650 , n586972 , n52022 );
and ( n59651 , n59646 , n59650 );
xor ( n586975 , n59474 , n59476 );
xor ( n586976 , n586975 , n59479 );
and ( n59654 , n59650 , n586976 );
and ( n59655 , n59646 , n586976 );
or ( n586979 , n59651 , n59654 , n59655 );
nor ( n59657 , n51991 , n51989 );
xnor ( n59658 , n59657 , n51959 );
nor ( n59659 , n51936 , n51934 );
xnor ( n59660 , n59659 , n51941 );
and ( n59661 , n59658 , n59660 );
nor ( n59662 , n51929 , n51927 );
not ( n586986 , n59662 );
and ( n586987 , n59660 , n586986 );
and ( n59665 , n59658 , n586986 );
or ( n586989 , n59661 , n586987 , n59665 );
and ( n586990 , n58623 , n52065 );
and ( n59668 , n585909 , n52063 );
nor ( n586992 , n586990 , n59668 );
xnor ( n586993 , n586992 , n52022 );
and ( n59671 , n586989 , n586993 );
xor ( n586995 , n59638 , n59640 );
xor ( n586996 , n586995 , n59643 );
and ( n59674 , n586993 , n586996 );
and ( n59675 , n586989 , n586996 );
or ( n586999 , n59671 , n59674 , n59675 );
and ( n587000 , n585973 , n52063 );
nor ( n59678 , n52065 , n587000 );
xnor ( n587002 , n59678 , n52022 );
nor ( n587003 , n51936 , n51934 );
xnor ( n59681 , n587003 , n51941 );
and ( n587005 , n587002 , n59681 );
nor ( n587006 , n51929 , n51927 );
not ( n59684 , n587006 );
and ( n587008 , n59681 , n59684 );
and ( n587009 , n587002 , n59684 );
or ( n59687 , n587005 , n587008 , n587009 );
and ( n587011 , n585973 , n52065 );
and ( n587012 , n58623 , n52063 );
nor ( n587013 , n587011 , n587012 );
xnor ( n587014 , n587013 , n52022 );
and ( n59692 , n59687 , n587014 );
xor ( n587016 , n59658 , n59660 );
xor ( n587017 , n587016 , n586986 );
and ( n59695 , n587014 , n587017 );
and ( n587019 , n59687 , n587017 );
or ( n587020 , n59692 , n59695 , n587019 );
and ( n59698 , n585586 , n52155 );
and ( n587022 , n58246 , n52153 );
nor ( n587023 , n59698 , n587022 );
xnor ( n59701 , n587023 , n52085 );
and ( n59702 , n587020 , n59701 );
xor ( n587026 , n586989 , n586993 );
xor ( n587027 , n587026 , n586996 );
and ( n59705 , n59701 , n587027 );
and ( n587029 , n587020 , n587027 );
or ( n587030 , n59702 , n59705 , n587029 );
and ( n59708 , n586999 , n587030 );
xor ( n587032 , n59646 , n59650 );
xor ( n587033 , n587032 , n586976 );
and ( n59711 , n587030 , n587033 );
and ( n587035 , n586999 , n587033 );
or ( n587036 , n59708 , n59711 , n587035 );
and ( n59714 , n586979 , n587036 );
xor ( n587038 , n59482 , n586809 );
xor ( n587039 , n587038 , n59489 );
and ( n59717 , n587036 , n587039 );
and ( n587041 , n586979 , n587039 );
or ( n587042 , n59714 , n59717 , n587041 );
and ( n59720 , n585062 , n52273 );
and ( n587044 , n57482 , n52271 );
nor ( n587045 , n59720 , n587044 );
xnor ( n59723 , n587045 , n52137 );
and ( n587047 , n587042 , n59723 );
xor ( n587048 , n59492 , n59496 );
xor ( n59726 , n587048 , n59499 );
and ( n587050 , n59723 , n59726 );
and ( n587051 , n587042 , n59726 );
or ( n59729 , n587047 , n587050 , n587051 );
and ( n59730 , n57900 , n52273 );
and ( n587054 , n585062 , n52271 );
nor ( n587055 , n59730 , n587054 );
xnor ( n59733 , n587055 , n52137 );
and ( n587057 , n58219 , n52155 );
and ( n587058 , n585221 , n52153 );
nor ( n59736 , n587057 , n587058 );
xnor ( n587060 , n59736 , n52085 );
and ( n587061 , n59733 , n587060 );
xor ( n59739 , n586979 , n587036 );
xor ( n587063 , n59739 , n587039 );
and ( n587064 , n587060 , n587063 );
and ( n59742 , n59733 , n587063 );
or ( n587066 , n587061 , n587064 , n59742 );
and ( n587067 , n57484 , n52432 );
and ( n59745 , n57283 , n52430 );
nor ( n59746 , n587067 , n59745 );
xnor ( n59747 , n59746 , n52255 );
and ( n587071 , n587066 , n59747 );
xor ( n587072 , n587042 , n59723 );
xor ( n59750 , n587072 , n59726 );
and ( n587074 , n59747 , n59750 );
and ( n587075 , n587066 , n59750 );
or ( n59753 , n587071 , n587074 , n587075 );
and ( n59754 , n59729 , n59753 );
xor ( n587078 , n59502 , n59506 );
xor ( n587079 , n587078 , n586832 );
and ( n59757 , n59753 , n587079 );
and ( n587081 , n59729 , n587079 );
or ( n587082 , n59754 , n59757 , n587081 );
and ( n59760 , n56909 , n52509 );
and ( n587084 , n56832 , n52507 );
nor ( n59762 , n59760 , n587084 );
xnor ( n587086 , n59762 , n52383 );
and ( n587087 , n587082 , n587086 );
xor ( n59765 , n586835 , n586839 );
xor ( n587089 , n59765 , n59519 );
and ( n587090 , n587086 , n587089 );
and ( n59768 , n587082 , n587089 );
or ( n59769 , n587087 , n587090 , n59768 );
and ( n587093 , n583800 , n52707 );
and ( n587094 , n583746 , n52705 );
nor ( n59772 , n587093 , n587094 );
xnor ( n59773 , n59772 , n52526 );
and ( n587097 , n59769 , n59773 );
xor ( n587098 , n59522 , n59526 );
xor ( n587099 , n587098 , n59529 );
and ( n59777 , n59773 , n587099 );
and ( n587101 , n59769 , n587099 );
or ( n587102 , n587097 , n59777 , n587101 );
and ( n59780 , n583048 , n53177 );
and ( n587104 , n582961 , n53175 );
nor ( n587105 , n59780 , n587104 );
xnor ( n59783 , n587105 , n52827 );
and ( n59784 , n587102 , n59783 );
xor ( n587108 , n59311 , n59315 );
xor ( n587109 , n587108 , n59318 );
and ( n59787 , n59783 , n587109 );
and ( n59788 , n587102 , n587109 );
or ( n587112 , n59784 , n59787 , n59788 );
and ( n587113 , n582961 , n53177 );
and ( n59791 , n55528 , n53175 );
nor ( n587115 , n587113 , n59791 );
xnor ( n587116 , n587115 , n52827 );
and ( n59794 , n587112 , n587116 );
xor ( n587118 , n586644 , n59325 );
xor ( n587119 , n587118 , n586653 );
and ( n59797 , n587116 , n587119 );
and ( n59798 , n587112 , n587119 );
or ( n59799 , n59794 , n59797 , n59798 );
and ( n59800 , n54893 , n53683 );
and ( n59801 , n54725 , n53681 );
nor ( n587125 , n59800 , n59801 );
xnor ( n59803 , n587125 , n53118 );
and ( n59804 , n59799 , n59803 );
xor ( n587128 , n586656 , n586660 );
xor ( n587129 , n587128 , n586663 );
and ( n59807 , n59803 , n587129 );
and ( n587131 , n59799 , n587129 );
or ( n587132 , n59804 , n59807 , n587131 );
and ( n59810 , n54321 , n53996 );
and ( n587134 , n54215 , n53994 );
nor ( n587135 , n59810 , n587134 );
xnor ( n587136 , n587135 , n53376 );
and ( n59814 , n587132 , n587136 );
xor ( n587138 , n586666 , n59347 );
xor ( n59816 , n587138 , n59350 );
and ( n587140 , n587136 , n59816 );
and ( n587141 , n587132 , n59816 );
or ( n59819 , n59814 , n587140 , n587141 );
and ( n587143 , n53641 , n55013 );
and ( n587144 , n53365 , n55010 );
nor ( n59822 , n587143 , n587144 );
xnor ( n587146 , n59822 , n53762 );
and ( n587147 , n53837 , n54532 );
and ( n59825 , n53639 , n54530 );
nor ( n59826 , n587147 , n59825 );
xnor ( n59827 , n59826 , n53769 );
and ( n587151 , n587146 , n59827 );
xor ( n587152 , n586887 , n59568 );
xor ( n59830 , n587152 , n59571 );
and ( n59831 , n59827 , n59830 );
and ( n59832 , n587146 , n59830 );
or ( n587156 , n587151 , n59831 , n59832 );
and ( n59834 , n59819 , n587156 );
and ( n59835 , n53365 , n55013 );
and ( n59836 , n53367 , n55010 );
nor ( n59837 , n59835 , n59836 );
xnor ( n59838 , n59837 , n53762 );
and ( n59839 , n587156 , n59838 );
and ( n59840 , n59819 , n59838 );
or ( n59841 , n59834 , n59839 , n59840 );
xor ( n59842 , n59363 , n586690 );
xor ( n59843 , n59842 , n586695 );
and ( n59844 , n59841 , n59843 );
xor ( n59845 , n59610 , n586935 );
xor ( n59846 , n59845 , n586938 );
and ( n59847 , n59843 , n59846 );
and ( n59848 , n59841 , n59846 );
or ( n59849 , n59844 , n59847 , n59848 );
xor ( n59850 , n59606 , n59618 );
xor ( n587174 , n59850 , n586944 );
and ( n587175 , n59849 , n587174 );
xor ( n587176 , n586766 , n59445 );
xor ( n59854 , n587176 , n59448 );
and ( n587178 , n587174 , n59854 );
and ( n587179 , n59849 , n59854 );
or ( n59857 , n587175 , n587178 , n587179 );
and ( n587181 , n59635 , n59857 );
xor ( n587182 , n59849 , n587174 );
xor ( n59860 , n587182 , n59854 );
and ( n59861 , n57058 , n52509 );
and ( n587185 , n56909 , n52507 );
nor ( n587186 , n59861 , n587185 );
xnor ( n59864 , n587186 , n52383 );
and ( n59865 , n57283 , n52432 );
and ( n587189 , n584529 , n52430 );
nor ( n587190 , n59865 , n587189 );
xnor ( n587191 , n587190 , n52255 );
and ( n59869 , n59864 , n587191 );
xor ( n587193 , n59729 , n59753 );
xor ( n587194 , n587193 , n587079 );
and ( n59872 , n587191 , n587194 );
and ( n587196 , n59864 , n587194 );
or ( n587197 , n59869 , n59872 , n587196 );
and ( n59875 , n583746 , n52978 );
and ( n59876 , n56282 , n52976 );
nor ( n587200 , n59875 , n59876 );
xnor ( n587201 , n587200 , n52680 );
and ( n59879 , n587197 , n587201 );
xor ( n59880 , n587082 , n587086 );
xor ( n587204 , n59880 , n587089 );
and ( n587205 , n587201 , n587204 );
and ( n59883 , n587197 , n587204 );
or ( n59884 , n59879 , n587205 , n59883 );
and ( n59885 , n55841 , n53177 );
and ( n587209 , n583048 , n53175 );
nor ( n59887 , n59885 , n587209 );
xnor ( n59888 , n59887 , n52827 );
and ( n59889 , n59884 , n59888 );
and ( n587213 , n56282 , n52978 );
and ( n587214 , n583377 , n52976 );
nor ( n59892 , n587213 , n587214 );
xnor ( n587216 , n59892 , n52680 );
and ( n587217 , n59888 , n587216 );
and ( n59895 , n59884 , n587216 );
or ( n587219 , n59889 , n587217 , n59895 );
and ( n59897 , n55528 , n53468 );
and ( n587221 , n55293 , n53466 );
nor ( n587222 , n59897 , n587221 );
xnor ( n59900 , n587222 , n52945 );
and ( n59901 , n587219 , n59900 );
xor ( n59902 , n586855 , n586859 );
xor ( n587226 , n59902 , n586864 );
and ( n59904 , n59900 , n587226 );
and ( n59905 , n587219 , n587226 );
or ( n59906 , n59901 , n59904 , n59905 );
and ( n59907 , n55058 , n53683 );
and ( n59908 , n54893 , n53681 );
nor ( n587232 , n59907 , n59908 );
xnor ( n59910 , n587232 , n53118 );
and ( n587234 , n59906 , n59910 );
xor ( n59912 , n586867 , n586871 );
xor ( n587236 , n59912 , n59551 );
and ( n59914 , n59910 , n587236 );
and ( n59915 , n59906 , n587236 );
or ( n587239 , n587234 , n59914 , n59915 );
and ( n587240 , n54553 , n53996 );
and ( n59918 , n54321 , n53994 );
nor ( n587242 , n587240 , n59918 );
xnor ( n587243 , n587242 , n53376 );
and ( n59921 , n587239 , n587243 );
xor ( n59922 , n59554 , n59558 );
xor ( n587246 , n59922 , n59561 );
and ( n587247 , n587243 , n587246 );
and ( n59925 , n587239 , n587246 );
or ( n587249 , n59921 , n587247 , n59925 );
and ( n587250 , n54055 , n54414 );
and ( n587251 , n53835 , n54412 );
nor ( n587252 , n587250 , n587251 );
xnor ( n59930 , n587252 , n53650 );
and ( n587254 , n587249 , n59930 );
xor ( n587255 , n587132 , n587136 );
xor ( n59933 , n587255 , n59816 );
and ( n587257 , n59930 , n59933 );
and ( n59935 , n587249 , n59933 );
or ( n587259 , n587254 , n587257 , n59935 );
xor ( n59937 , n59574 , n59578 );
xor ( n59938 , n59937 , n586904 );
and ( n587262 , n587259 , n59938 );
xor ( n587263 , n586911 , n59592 );
xor ( n59941 , n587263 , n59595 );
and ( n587265 , n59938 , n59941 );
and ( n587266 , n587259 , n59941 );
or ( n59944 , n587262 , n587265 , n587266 );
xor ( n587268 , n586907 , n59598 );
xor ( n587269 , n587268 , n586926 );
and ( n59947 , n59944 , n587269 );
xor ( n587271 , n59841 , n59843 );
xor ( n59949 , n587271 , n59846 );
and ( n587273 , n587269 , n59949 );
and ( n587274 , n59944 , n59949 );
or ( n59952 , n59947 , n587273 , n587274 );
and ( n587276 , n59860 , n59952 );
xor ( n587277 , n59944 , n587269 );
xor ( n587278 , n587277 , n59949 );
and ( n59956 , n585221 , n52273 );
and ( n587280 , n57900 , n52271 );
nor ( n587281 , n59956 , n587280 );
xnor ( n587282 , n587281 , n52137 );
and ( n59960 , n58246 , n52155 );
and ( n587284 , n58219 , n52153 );
nor ( n587285 , n59960 , n587284 );
xnor ( n59963 , n587285 , n52085 );
and ( n587287 , n587282 , n59963 );
xor ( n587288 , n586999 , n587030 );
xor ( n59966 , n587288 , n587033 );
and ( n587290 , n59963 , n59966 );
and ( n587291 , n587282 , n59966 );
or ( n59969 , n587287 , n587290 , n587291 );
and ( n59970 , n57482 , n52432 );
and ( n59971 , n57484 , n52430 );
nor ( n587295 , n59970 , n59971 );
xnor ( n59973 , n587295 , n52255 );
and ( n59974 , n59969 , n59973 );
xor ( n59975 , n59733 , n587060 );
xor ( n59976 , n59975 , n587063 );
and ( n59977 , n59973 , n59976 );
and ( n59978 , n59969 , n59976 );
or ( n59979 , n59974 , n59977 , n59978 );
and ( n59980 , n584529 , n52509 );
and ( n59981 , n57058 , n52507 );
nor ( n59982 , n59980 , n59981 );
xnor ( n59983 , n59982 , n52383 );
and ( n59984 , n59979 , n59983 );
xor ( n59985 , n587066 , n59747 );
xor ( n587309 , n59985 , n59750 );
and ( n59987 , n59983 , n587309 );
and ( n587311 , n59979 , n587309 );
or ( n587312 , n59984 , n59987 , n587311 );
nor ( n59990 , n52065 , n52063 );
xnor ( n587314 , n59990 , n52022 );
nor ( n587315 , n51936 , n51934 );
xnor ( n587316 , n587315 , n51941 );
and ( n587317 , n587314 , n587316 );
nor ( n59995 , n51929 , n51927 );
not ( n587319 , n59995 );
and ( n587320 , n587316 , n587319 );
and ( n59998 , n587314 , n587319 );
or ( n587322 , n587317 , n587320 , n59998 );
nor ( n60000 , n51991 , n51989 );
xnor ( n587324 , n60000 , n51959 );
and ( n60002 , n587322 , n587324 );
xor ( n60003 , n587002 , n59681 );
xor ( n587327 , n60003 , n59684 );
and ( n587328 , n587324 , n587327 );
and ( n60006 , n587322 , n587327 );
or ( n587330 , n60002 , n587328 , n60006 );
and ( n587331 , n585909 , n52155 );
and ( n60009 , n585586 , n52153 );
nor ( n587333 , n587331 , n60009 );
xnor ( n587334 , n587333 , n52085 );
and ( n60012 , n587330 , n587334 );
xor ( n587336 , n59687 , n587014 );
xor ( n587337 , n587336 , n587017 );
and ( n587338 , n587334 , n587337 );
and ( n587339 , n587330 , n587337 );
or ( n60017 , n60012 , n587338 , n587339 );
nor ( n587341 , n52065 , n52063 );
xnor ( n587342 , n587341 , n52022 );
nor ( n587343 , n51936 , n51934 );
xnor ( n587344 , n587343 , n51941 );
and ( n60022 , n587342 , n587344 );
and ( n587346 , n587344 , n51927 );
and ( n587347 , n587342 , n51927 );
or ( n60025 , n60022 , n587346 , n587347 );
and ( n587349 , n585973 , n52155 );
and ( n60027 , n58623 , n52153 );
nor ( n587351 , n587349 , n60027 );
xnor ( n60029 , n587351 , n52085 );
and ( n60030 , n60025 , n60029 );
nor ( n587354 , n51991 , n51989 );
xnor ( n587355 , n587354 , n51959 );
and ( n60033 , n60029 , n587355 );
and ( n587357 , n60025 , n587355 );
or ( n587358 , n60030 , n60033 , n587357 );
and ( n60036 , n58623 , n52155 );
and ( n587360 , n585909 , n52153 );
nor ( n587361 , n60036 , n587360 );
xnor ( n60039 , n587361 , n52085 );
and ( n587363 , n587358 , n60039 );
xor ( n587364 , n587322 , n587324 );
xor ( n60042 , n587364 , n587327 );
and ( n60043 , n60039 , n60042 );
and ( n587367 , n587358 , n60042 );
or ( n60045 , n587363 , n60043 , n587367 );
nor ( n60046 , n52065 , n52063 );
xnor ( n60047 , n60046 , n52022 );
and ( n587371 , n51935 , n51941 );
and ( n587372 , n60047 , n587371 );
and ( n60050 , n585973 , n52153 );
nor ( n60051 , n52155 , n60050 );
xnor ( n60052 , n60051 , n52085 );
and ( n587376 , n587372 , n60052 );
nor ( n587377 , n51991 , n51989 );
xnor ( n60055 , n587377 , n51959 );
and ( n60056 , n60052 , n60055 );
and ( n587380 , n587372 , n60055 );
or ( n587381 , n587376 , n60056 , n587380 );
xor ( n60059 , n587314 , n587316 );
xor ( n587383 , n60059 , n587319 );
and ( n60061 , n587381 , n587383 );
xor ( n587385 , n60025 , n60029 );
xor ( n587386 , n587385 , n587355 );
and ( n60064 , n587383 , n587386 );
and ( n587388 , n587381 , n587386 );
or ( n587389 , n60061 , n60064 , n587388 );
and ( n60067 , n585586 , n52273 );
and ( n60068 , n58246 , n52271 );
nor ( n587392 , n60067 , n60068 );
xnor ( n587393 , n587392 , n52137 );
and ( n60071 , n587389 , n587393 );
xor ( n60072 , n587358 , n60039 );
xor ( n587396 , n60072 , n60042 );
and ( n587397 , n587393 , n587396 );
and ( n587398 , n587389 , n587396 );
or ( n60076 , n60071 , n587397 , n587398 );
and ( n587400 , n60045 , n60076 );
xor ( n587401 , n587330 , n587334 );
xor ( n60079 , n587401 , n587337 );
and ( n587403 , n60076 , n60079 );
and ( n587404 , n60045 , n60079 );
or ( n60082 , n587400 , n587403 , n587404 );
and ( n60083 , n60017 , n60082 );
xor ( n587407 , n587020 , n59701 );
xor ( n587408 , n587407 , n587027 );
and ( n60086 , n60082 , n587408 );
and ( n60087 , n60017 , n587408 );
or ( n587411 , n60083 , n60086 , n60087 );
and ( n587412 , n585062 , n52432 );
and ( n60090 , n57482 , n52430 );
nor ( n587414 , n587412 , n60090 );
xnor ( n60092 , n587414 , n52255 );
and ( n587416 , n587411 , n60092 );
xor ( n587417 , n587282 , n59963 );
xor ( n60095 , n587417 , n59966 );
and ( n587419 , n60092 , n60095 );
and ( n587420 , n587411 , n60095 );
or ( n60098 , n587416 , n587419 , n587420 );
and ( n60099 , n57900 , n52432 );
and ( n587423 , n585062 , n52430 );
nor ( n587424 , n60099 , n587423 );
xnor ( n60102 , n587424 , n52255 );
and ( n60103 , n58219 , n52273 );
and ( n587427 , n585221 , n52271 );
nor ( n587428 , n60103 , n587427 );
xnor ( n60106 , n587428 , n52137 );
and ( n60107 , n60102 , n60106 );
xor ( n60108 , n60017 , n60082 );
xor ( n587432 , n60108 , n587408 );
and ( n587433 , n60106 , n587432 );
and ( n60111 , n60102 , n587432 );
or ( n60112 , n60107 , n587433 , n60111 );
and ( n587436 , n57484 , n52509 );
and ( n587437 , n57283 , n52507 );
nor ( n60115 , n587436 , n587437 );
xnor ( n60116 , n60115 , n52383 );
and ( n60117 , n60112 , n60116 );
xor ( n587441 , n587411 , n60092 );
xor ( n587442 , n587441 , n60095 );
and ( n60120 , n60116 , n587442 );
and ( n60121 , n60112 , n587442 );
or ( n60122 , n60117 , n60120 , n60121 );
and ( n587446 , n60098 , n60122 );
xor ( n587447 , n59969 , n59973 );
xor ( n60125 , n587447 , n59976 );
and ( n60126 , n60122 , n60125 );
and ( n60127 , n60098 , n60125 );
or ( n587451 , n587446 , n60126 , n60127 );
and ( n587452 , n56909 , n52707 );
and ( n60130 , n56832 , n52705 );
nor ( n60131 , n587452 , n60130 );
xnor ( n587455 , n60131 , n52526 );
and ( n60133 , n587451 , n587455 );
xor ( n60134 , n59979 , n59983 );
xor ( n60135 , n60134 , n587309 );
and ( n60136 , n587455 , n60135 );
and ( n60137 , n587451 , n60135 );
or ( n60138 , n60133 , n60136 , n60137 );
and ( n60139 , n587312 , n60138 );
xor ( n60140 , n59864 , n587191 );
xor ( n60141 , n60140 , n587194 );
and ( n60142 , n60138 , n60141 );
and ( n587466 , n587312 , n60141 );
or ( n60144 , n60139 , n60142 , n587466 );
and ( n60145 , n583377 , n53177 );
and ( n587469 , n55841 , n53175 );
nor ( n60147 , n60145 , n587469 );
xnor ( n60148 , n60147 , n52827 );
and ( n60149 , n60144 , n60148 );
and ( n60150 , n56671 , n52707 );
and ( n587474 , n583800 , n52705 );
nor ( n587475 , n60150 , n587474 );
xnor ( n60153 , n587475 , n52526 );
and ( n587477 , n60148 , n60153 );
and ( n60155 , n60144 , n60153 );
or ( n60156 , n60149 , n587477 , n60155 );
xor ( n587480 , n59884 , n59888 );
xor ( n587481 , n587480 , n587216 );
and ( n60159 , n60156 , n587481 );
xor ( n60160 , n59769 , n59773 );
xor ( n587484 , n60160 , n587099 );
and ( n587485 , n587481 , n587484 );
and ( n60163 , n60156 , n587484 );
or ( n587487 , n60159 , n587485 , n60163 );
and ( n60165 , n55075 , n53683 );
and ( n60166 , n55058 , n53681 );
nor ( n587490 , n60165 , n60166 );
xnor ( n587491 , n587490 , n53118 );
and ( n60169 , n587487 , n587491 );
xor ( n60170 , n587102 , n59783 );
xor ( n587494 , n60170 , n587109 );
and ( n587495 , n587491 , n587494 );
and ( n60173 , n587487 , n587494 );
or ( n587497 , n60169 , n587495 , n60173 );
and ( n60175 , n54725 , n53996 );
and ( n587499 , n54553 , n53994 );
nor ( n60177 , n60175 , n587499 );
xnor ( n60178 , n60177 , n53376 );
and ( n587502 , n587497 , n60178 );
xor ( n587503 , n587112 , n587116 );
xor ( n60181 , n587503 , n587119 );
and ( n60182 , n60178 , n60181 );
and ( n587506 , n587497 , n60181 );
or ( n587507 , n587502 , n60182 , n587506 );
and ( n60185 , n53835 , n54532 );
and ( n587509 , n53837 , n54530 );
nor ( n60187 , n60185 , n587509 );
xnor ( n60188 , n60187 , n53769 );
and ( n587512 , n587507 , n60188 );
xor ( n587513 , n587239 , n587243 );
xor ( n60191 , n587513 , n587246 );
and ( n60192 , n60188 , n60191 );
and ( n587516 , n587507 , n60191 );
or ( n587517 , n587512 , n60192 , n587516 );
and ( n60195 , n53639 , n55013 );
and ( n60196 , n53641 , n55010 );
nor ( n587520 , n60195 , n60196 );
xnor ( n587521 , n587520 , n53762 );
and ( n60199 , n54215 , n54414 );
and ( n60200 , n54055 , n54412 );
nor ( n60201 , n60199 , n60200 );
xnor ( n587525 , n60201 , n53650 );
and ( n587526 , n587521 , n587525 );
xor ( n60204 , n59799 , n59803 );
xor ( n587528 , n60204 , n587129 );
and ( n587529 , n587525 , n587528 );
and ( n60207 , n587521 , n587528 );
or ( n587531 , n587526 , n587529 , n60207 );
and ( n587532 , n587517 , n587531 );
xor ( n60210 , n587146 , n59827 );
xor ( n587534 , n60210 , n59830 );
and ( n587535 , n587531 , n587534 );
and ( n60213 , n587517 , n587534 );
or ( n587537 , n587532 , n587535 , n60213 );
xor ( n587538 , n59819 , n587156 );
xor ( n60216 , n587538 , n59838 );
and ( n587540 , n587537 , n60216 );
xor ( n587541 , n587259 , n59938 );
xor ( n60219 , n587541 , n59941 );
and ( n587543 , n60216 , n60219 );
and ( n60221 , n587537 , n60219 );
or ( n60222 , n587540 , n587543 , n60221 );
and ( n60223 , n587278 , n60222 );
xor ( n60224 , n587537 , n60216 );
xor ( n60225 , n60224 , n60219 );
and ( n60226 , n57058 , n52707 );
and ( n60227 , n56909 , n52705 );
nor ( n60228 , n60226 , n60227 );
xnor ( n60229 , n60228 , n52526 );
and ( n60230 , n57283 , n52509 );
and ( n60231 , n584529 , n52507 );
nor ( n60232 , n60230 , n60231 );
xnor ( n60233 , n60232 , n52383 );
and ( n60234 , n60229 , n60233 );
xor ( n60235 , n60098 , n60122 );
xor ( n587559 , n60235 , n60125 );
and ( n587560 , n60233 , n587559 );
and ( n60238 , n60229 , n587559 );
or ( n587562 , n60234 , n587560 , n60238 );
and ( n587563 , n56671 , n52978 );
and ( n60241 , n583800 , n52976 );
nor ( n587565 , n587563 , n60241 );
xnor ( n587566 , n587565 , n52680 );
and ( n60244 , n587562 , n587566 );
xor ( n587568 , n587451 , n587455 );
xor ( n587569 , n587568 , n60135 );
and ( n60247 , n587566 , n587569 );
and ( n60248 , n587562 , n587569 );
or ( n587572 , n60244 , n60247 , n60248 );
and ( n587573 , n56282 , n53177 );
and ( n60251 , n583377 , n53175 );
nor ( n587575 , n587573 , n60251 );
xnor ( n587576 , n587575 , n52827 );
and ( n60254 , n587572 , n587576 );
and ( n587578 , n583800 , n52978 );
and ( n587579 , n583746 , n52976 );
nor ( n60257 , n587578 , n587579 );
xnor ( n587581 , n60257 , n52680 );
and ( n587582 , n56832 , n52707 );
and ( n60260 , n56671 , n52705 );
nor ( n587584 , n587582 , n60260 );
xnor ( n587585 , n587584 , n52526 );
xor ( n60263 , n587581 , n587585 );
xor ( n587587 , n587312 , n60138 );
xor ( n60265 , n587587 , n60141 );
xor ( n60266 , n60263 , n60265 );
and ( n587590 , n587576 , n60266 );
and ( n60268 , n587572 , n60266 );
or ( n60269 , n60254 , n587590 , n60268 );
and ( n60270 , n55528 , n53683 );
and ( n60271 , n55293 , n53681 );
nor ( n60272 , n60270 , n60271 );
xnor ( n60273 , n60272 , n53118 );
and ( n60274 , n60269 , n60273 );
xor ( n60275 , n60144 , n60148 );
xor ( n60276 , n60275 , n60153 );
and ( n60277 , n60273 , n60276 );
and ( n60278 , n60269 , n60276 );
or ( n60279 , n60274 , n60277 , n60278 );
and ( n60280 , n55058 , n53996 );
and ( n60281 , n54893 , n53994 );
nor ( n60282 , n60280 , n60281 );
xnor ( n60283 , n60282 , n53376 );
and ( n60284 , n60279 , n60283 );
xor ( n587608 , n60156 , n587481 );
xor ( n60286 , n587608 , n587484 );
and ( n60287 , n60283 , n60286 );
and ( n60288 , n60279 , n60286 );
or ( n587612 , n60284 , n60287 , n60288 );
and ( n587613 , n54553 , n54414 );
and ( n587614 , n54321 , n54412 );
nor ( n60292 , n587613 , n587614 );
xnor ( n587616 , n60292 , n53650 );
and ( n587617 , n587612 , n587616 );
xor ( n60295 , n587487 , n587491 );
xor ( n587619 , n60295 , n587494 );
and ( n587620 , n587616 , n587619 );
and ( n60298 , n587612 , n587619 );
or ( n587622 , n587617 , n587620 , n60298 );
and ( n587623 , n53837 , n55013 );
and ( n60301 , n53639 , n55010 );
nor ( n60302 , n587623 , n60301 );
xnor ( n587626 , n60302 , n53762 );
and ( n587627 , n587622 , n587626 );
and ( n60305 , n54055 , n54532 );
and ( n587629 , n53835 , n54530 );
nor ( n587630 , n60305 , n587629 );
xnor ( n60308 , n587630 , n53769 );
and ( n587632 , n587626 , n60308 );
and ( n587633 , n587622 , n60308 );
or ( n60311 , n587627 , n587632 , n587633 );
and ( n587635 , n587581 , n587585 );
and ( n587636 , n587585 , n60265 );
and ( n60314 , n587581 , n60265 );
or ( n587638 , n587635 , n587636 , n60314 );
and ( n587639 , n583048 , n53468 );
and ( n587640 , n582961 , n53466 );
nor ( n587641 , n587639 , n587640 );
xnor ( n60319 , n587641 , n52945 );
and ( n587643 , n587638 , n60319 );
xor ( n587644 , n587197 , n587201 );
xor ( n60322 , n587644 , n587204 );
and ( n587646 , n60319 , n60322 );
and ( n587647 , n587638 , n60322 );
or ( n60325 , n587643 , n587646 , n587647 );
and ( n587649 , n55293 , n53683 );
and ( n587650 , n55075 , n53681 );
nor ( n60328 , n587649 , n587650 );
xnor ( n60329 , n60328 , n53118 );
and ( n587653 , n60325 , n60329 );
and ( n587654 , n582961 , n53468 );
and ( n60332 , n55528 , n53466 );
nor ( n587656 , n587654 , n60332 );
xnor ( n587657 , n587656 , n52945 );
and ( n60335 , n60329 , n587657 );
and ( n587659 , n60325 , n587657 );
or ( n587660 , n587653 , n60335 , n587659 );
and ( n60338 , n54893 , n53996 );
and ( n587662 , n54725 , n53994 );
nor ( n587663 , n60338 , n587662 );
xnor ( n60341 , n587663 , n53376 );
and ( n587665 , n587660 , n60341 );
xor ( n587666 , n587219 , n59900 );
xor ( n60344 , n587666 , n587226 );
and ( n587668 , n60341 , n60344 );
and ( n587669 , n587660 , n60344 );
or ( n60347 , n587665 , n587668 , n587669 );
and ( n587671 , n54321 , n54414 );
and ( n60349 , n54215 , n54412 );
nor ( n587673 , n587671 , n60349 );
xnor ( n60351 , n587673 , n53650 );
and ( n60352 , n60347 , n60351 );
xor ( n587676 , n59906 , n59910 );
xor ( n587677 , n587676 , n587236 );
and ( n60355 , n60351 , n587677 );
and ( n60356 , n60347 , n587677 );
or ( n587680 , n60352 , n60355 , n60356 );
and ( n587681 , n60311 , n587680 );
xor ( n60359 , n587507 , n60188 );
xor ( n587683 , n60359 , n60191 );
and ( n60361 , n587680 , n587683 );
and ( n60362 , n60311 , n587683 );
or ( n587686 , n587681 , n60361 , n60362 );
xor ( n587687 , n587249 , n59930 );
xor ( n60365 , n587687 , n59933 );
and ( n60366 , n587686 , n60365 );
xor ( n587690 , n587517 , n587531 );
xor ( n587691 , n587690 , n587534 );
and ( n60369 , n60365 , n587691 );
and ( n60370 , n587686 , n587691 );
or ( n60371 , n60366 , n60369 , n60370 );
and ( n587695 , n60225 , n60371 );
xor ( n587696 , n587686 , n60365 );
xor ( n60374 , n587696 , n587691 );
and ( n587698 , n585221 , n52432 );
and ( n587699 , n57900 , n52430 );
nor ( n60377 , n587698 , n587699 );
xnor ( n60378 , n60377 , n52255 );
and ( n587702 , n58246 , n52273 );
and ( n587703 , n58219 , n52271 );
nor ( n60381 , n587702 , n587703 );
xnor ( n60382 , n60381 , n52137 );
and ( n60383 , n60378 , n60382 );
xor ( n587707 , n60045 , n60076 );
xor ( n587708 , n587707 , n60079 );
and ( n60386 , n60382 , n587708 );
and ( n60387 , n60378 , n587708 );
or ( n60388 , n60383 , n60386 , n60387 );
and ( n587712 , n57482 , n52509 );
and ( n60390 , n57484 , n52507 );
nor ( n60391 , n587712 , n60390 );
xnor ( n60392 , n60391 , n52383 );
and ( n587716 , n60388 , n60392 );
xor ( n60394 , n60102 , n60106 );
xor ( n60395 , n60394 , n587432 );
and ( n60396 , n60392 , n60395 );
and ( n587720 , n60388 , n60395 );
or ( n60398 , n587716 , n60396 , n587720 );
and ( n60399 , n584529 , n52707 );
and ( n587723 , n57058 , n52705 );
nor ( n587724 , n60399 , n587723 );
xnor ( n60402 , n587724 , n52526 );
and ( n60403 , n60398 , n60402 );
xor ( n587727 , n60112 , n60116 );
xor ( n587728 , n587727 , n587442 );
and ( n60406 , n60402 , n587728 );
and ( n60407 , n60398 , n587728 );
or ( n587731 , n60403 , n60406 , n60407 );
and ( n60409 , n56832 , n52978 );
and ( n60410 , n56671 , n52976 );
nor ( n60411 , n60409 , n60410 );
xnor ( n60412 , n60411 , n52680 );
and ( n587736 , n587731 , n60412 );
xor ( n60414 , n60229 , n60233 );
xor ( n587738 , n60414 , n587559 );
and ( n60416 , n60412 , n587738 );
and ( n60417 , n587731 , n587738 );
or ( n587741 , n587736 , n60416 , n60417 );
and ( n60419 , n583377 , n53468 );
and ( n587743 , n55841 , n53466 );
nor ( n587744 , n60419 , n587743 );
xnor ( n60422 , n587744 , n52945 );
and ( n60423 , n587741 , n60422 );
and ( n60424 , n583746 , n53177 );
and ( n60425 , n56282 , n53175 );
nor ( n60426 , n60424 , n60425 );
xnor ( n60427 , n60426 , n52827 );
and ( n60428 , n60422 , n60427 );
and ( n60429 , n587741 , n60427 );
or ( n60430 , n60423 , n60428 , n60429 );
and ( n60431 , n55293 , n53996 );
and ( n60432 , n55075 , n53994 );
nor ( n60433 , n60431 , n60432 );
xnor ( n60434 , n60433 , n53376 );
and ( n60435 , n60430 , n60434 );
and ( n587759 , n55841 , n53468 );
and ( n60437 , n583048 , n53466 );
nor ( n60438 , n587759 , n60437 );
xnor ( n587762 , n60438 , n52945 );
and ( n60440 , n60434 , n587762 );
and ( n587764 , n60430 , n587762 );
or ( n60442 , n60435 , n60440 , n587764 );
and ( n587766 , n55075 , n53996 );
and ( n587767 , n55058 , n53994 );
nor ( n60445 , n587766 , n587767 );
xnor ( n587769 , n60445 , n53376 );
and ( n587770 , n60442 , n587769 );
xor ( n587771 , n587638 , n60319 );
xor ( n60449 , n587771 , n60322 );
and ( n587773 , n587769 , n60449 );
and ( n587774 , n60442 , n60449 );
or ( n587775 , n587770 , n587773 , n587774 );
and ( n587776 , n54725 , n54414 );
and ( n60454 , n54553 , n54412 );
nor ( n587778 , n587776 , n60454 );
xnor ( n587779 , n587778 , n53650 );
and ( n60457 , n587775 , n587779 );
xor ( n587781 , n60325 , n60329 );
xor ( n587782 , n587781 , n587657 );
and ( n60460 , n587779 , n587782 );
and ( n587784 , n587775 , n587782 );
or ( n587785 , n60457 , n60460 , n587784 );
and ( n60463 , n53835 , n55013 );
and ( n60464 , n53837 , n55010 );
nor ( n60465 , n60463 , n60464 );
xnor ( n587789 , n60465 , n53762 );
and ( n587790 , n587785 , n587789 );
xor ( n587791 , n587660 , n60341 );
xor ( n587792 , n587791 , n60344 );
and ( n60470 , n587789 , n587792 );
and ( n587794 , n587785 , n587792 );
or ( n587795 , n587790 , n60470 , n587794 );
xor ( n587796 , n587497 , n60178 );
xor ( n587797 , n587796 , n60181 );
and ( n60475 , n587795 , n587797 );
xor ( n587799 , n60347 , n60351 );
xor ( n587800 , n587799 , n587677 );
and ( n60478 , n587797 , n587800 );
and ( n587802 , n587795 , n587800 );
or ( n587803 , n60475 , n60478 , n587802 );
xor ( n60481 , n60311 , n587680 );
xor ( n587805 , n60481 , n587683 );
and ( n587806 , n587803 , n587805 );
xor ( n60484 , n587521 , n587525 );
xor ( n60485 , n60484 , n587528 );
and ( n60486 , n587805 , n60485 );
and ( n587810 , n587803 , n60485 );
or ( n587811 , n587806 , n60486 , n587810 );
and ( n60489 , n60374 , n587811 );
nor ( n60490 , n52155 , n52153 );
xnor ( n587814 , n60490 , n52085 );
nor ( n587815 , n51991 , n51989 );
xnor ( n60493 , n587815 , n51959 );
and ( n587817 , n587814 , n60493 );
nor ( n587818 , n51936 , n51934 );
xnor ( n60496 , n587818 , n51941 );
and ( n587820 , n60493 , n60496 );
and ( n60498 , n587814 , n60496 );
or ( n60499 , n587817 , n587820 , n60498 );
xor ( n60500 , n587342 , n587344 );
xor ( n60501 , n60500 , n51927 );
and ( n60502 , n60499 , n60501 );
xor ( n60503 , n587372 , n60052 );
xor ( n60504 , n60503 , n60055 );
and ( n60505 , n60501 , n60504 );
and ( n60506 , n60499 , n60504 );
or ( n60507 , n60502 , n60505 , n60506 );
and ( n60508 , n585909 , n52273 );
and ( n60509 , n585586 , n52271 );
nor ( n60510 , n60508 , n60509 );
xnor ( n60511 , n60510 , n52137 );
and ( n60512 , n60507 , n60511 );
xor ( n60513 , n587381 , n587383 );
xor ( n60514 , n60513 , n587386 );
and ( n587838 , n60511 , n60514 );
and ( n587839 , n60507 , n60514 );
or ( n60517 , n60512 , n587838 , n587839 );
xor ( n587841 , n60047 , n587371 );
nor ( n587842 , n52065 , n52063 );
xnor ( n587843 , n587842 , n52022 );
nor ( n60521 , n51991 , n51989 );
xnor ( n587845 , n60521 , n51959 );
and ( n60523 , n587843 , n587845 );
and ( n587847 , n587845 , n51934 );
and ( n587848 , n587843 , n51934 );
or ( n60526 , n60523 , n587847 , n587848 );
and ( n587850 , n587841 , n60526 );
and ( n60528 , n585973 , n52273 );
and ( n60529 , n58623 , n52271 );
nor ( n60530 , n60528 , n60529 );
xnor ( n60531 , n60530 , n52137 );
and ( n60532 , n60526 , n60531 );
and ( n60533 , n587841 , n60531 );
or ( n60534 , n587850 , n60532 , n60533 );
and ( n587858 , n58623 , n52273 );
and ( n587859 , n585909 , n52271 );
nor ( n587860 , n587858 , n587859 );
xnor ( n60538 , n587860 , n52137 );
and ( n587862 , n60534 , n60538 );
xor ( n60540 , n60499 , n60501 );
xor ( n587864 , n60540 , n60504 );
and ( n60542 , n60538 , n587864 );
and ( n60543 , n60534 , n587864 );
or ( n587867 , n587862 , n60542 , n60543 );
and ( n60545 , n58246 , n52432 );
and ( n587869 , n58219 , n52430 );
nor ( n587870 , n60545 , n587869 );
xnor ( n60548 , n587870 , n52255 );
and ( n587872 , n587867 , n60548 );
xor ( n587873 , n60507 , n60511 );
xor ( n60551 , n587873 , n60514 );
and ( n60552 , n60548 , n60551 );
and ( n60553 , n587867 , n60551 );
or ( n60554 , n587872 , n60552 , n60553 );
and ( n587878 , n60517 , n60554 );
xor ( n587879 , n587389 , n587393 );
xor ( n60557 , n587879 , n587396 );
and ( n60558 , n60554 , n60557 );
and ( n60559 , n60517 , n60557 );
or ( n587883 , n587878 , n60558 , n60559 );
and ( n60561 , n585062 , n52509 );
and ( n60562 , n57482 , n52507 );
nor ( n60563 , n60561 , n60562 );
xnor ( n587887 , n60563 , n52383 );
and ( n587888 , n587883 , n587887 );
xor ( n60566 , n60378 , n60382 );
xor ( n587890 , n60566 , n587708 );
and ( n60568 , n587887 , n587890 );
and ( n60569 , n587883 , n587890 );
or ( n60570 , n587888 , n60568 , n60569 );
and ( n60571 , n57900 , n52509 );
and ( n60572 , n585062 , n52507 );
nor ( n60573 , n60571 , n60572 );
xnor ( n60574 , n60573 , n52383 );
and ( n60575 , n58219 , n52432 );
and ( n60576 , n585221 , n52430 );
nor ( n60577 , n60575 , n60576 );
xnor ( n60578 , n60577 , n52255 );
and ( n60579 , n60574 , n60578 );
xor ( n60580 , n60517 , n60554 );
xor ( n60581 , n60580 , n60557 );
and ( n60582 , n60578 , n60581 );
and ( n60583 , n60574 , n60581 );
or ( n60584 , n60579 , n60582 , n60583 );
and ( n60585 , n57484 , n52707 );
and ( n60586 , n57283 , n52705 );
nor ( n60587 , n60585 , n60586 );
xnor ( n587911 , n60587 , n52526 );
and ( n60589 , n60584 , n587911 );
xor ( n60590 , n587883 , n587887 );
xor ( n587914 , n60590 , n587890 );
and ( n60592 , n587911 , n587914 );
and ( n60593 , n60584 , n587914 );
or ( n587917 , n60589 , n60592 , n60593 );
and ( n587918 , n60570 , n587917 );
xor ( n60596 , n60388 , n60392 );
xor ( n587920 , n60596 , n60395 );
and ( n60598 , n587917 , n587920 );
and ( n60599 , n60570 , n587920 );
or ( n587923 , n587918 , n60598 , n60599 );
and ( n587924 , n56909 , n52978 );
and ( n60602 , n56832 , n52976 );
nor ( n587926 , n587924 , n60602 );
xnor ( n60604 , n587926 , n52680 );
and ( n587928 , n587923 , n60604 );
xor ( n587929 , n60398 , n60402 );
xor ( n60607 , n587929 , n587728 );
and ( n587931 , n60604 , n60607 );
and ( n60609 , n587923 , n60607 );
or ( n60610 , n587928 , n587931 , n60609 );
and ( n587934 , n583800 , n53177 );
and ( n60612 , n583746 , n53175 );
nor ( n587936 , n587934 , n60612 );
xnor ( n60614 , n587936 , n52827 );
and ( n60615 , n60610 , n60614 );
xor ( n60616 , n587731 , n60412 );
xor ( n60617 , n60616 , n587738 );
and ( n60618 , n60614 , n60617 );
and ( n60619 , n60610 , n60617 );
or ( n587943 , n60615 , n60618 , n60619 );
and ( n587944 , n583048 , n53683 );
and ( n60622 , n582961 , n53681 );
nor ( n587946 , n587944 , n60622 );
xnor ( n587947 , n587946 , n53118 );
and ( n60625 , n587943 , n587947 );
xor ( n587949 , n587562 , n587566 );
xor ( n60627 , n587949 , n587569 );
and ( n60628 , n587947 , n60627 );
and ( n60629 , n587943 , n60627 );
or ( n60630 , n60625 , n60628 , n60629 );
and ( n60631 , n582961 , n53683 );
and ( n60632 , n55528 , n53681 );
nor ( n60633 , n60631 , n60632 );
xnor ( n60634 , n60633 , n53118 );
and ( n60635 , n60630 , n60634 );
xor ( n60636 , n587572 , n587576 );
xor ( n587960 , n60636 , n60266 );
and ( n587961 , n60634 , n587960 );
and ( n60639 , n60630 , n587960 );
or ( n587963 , n60635 , n587961 , n60639 );
and ( n587964 , n54893 , n54414 );
and ( n587965 , n54725 , n54412 );
nor ( n60643 , n587964 , n587965 );
xnor ( n587967 , n60643 , n53650 );
and ( n60645 , n587963 , n587967 );
xor ( n60646 , n60269 , n60273 );
xor ( n60647 , n60646 , n60276 );
and ( n60648 , n587967 , n60647 );
and ( n60649 , n587963 , n60647 );
or ( n60650 , n60645 , n60648 , n60649 );
and ( n587974 , n54321 , n54532 );
and ( n587975 , n54215 , n54530 );
nor ( n60653 , n587974 , n587975 );
xnor ( n587977 , n60653 , n53769 );
and ( n60655 , n60650 , n587977 );
xor ( n587979 , n60279 , n60283 );
xor ( n587980 , n587979 , n60286 );
and ( n60658 , n587977 , n587980 );
and ( n587982 , n60650 , n587980 );
or ( n60660 , n60655 , n60658 , n587982 );
and ( n60661 , n54215 , n54532 );
and ( n60662 , n54055 , n54530 );
nor ( n60663 , n60661 , n60662 );
xnor ( n60664 , n60663 , n53769 );
and ( n60665 , n60660 , n60664 );
xor ( n60666 , n587612 , n587616 );
xor ( n60667 , n60666 , n587619 );
and ( n60668 , n60664 , n60667 );
and ( n60669 , n60660 , n60667 );
or ( n60670 , n60665 , n60668 , n60669 );
xor ( n587994 , n587622 , n587626 );
xor ( n60672 , n587994 , n60308 );
and ( n60673 , n60670 , n60672 );
xor ( n60674 , n587795 , n587797 );
xor ( n60675 , n60674 , n587800 );
and ( n60676 , n60672 , n60675 );
and ( n60677 , n60670 , n60675 );
or ( n60678 , n60673 , n60676 , n60677 );
xor ( n60679 , n587803 , n587805 );
xor ( n60680 , n60679 , n60485 );
and ( n60681 , n60678 , n60680 );
xor ( n60682 , n60670 , n60672 );
xor ( n60683 , n60682 , n60675 );
and ( n60684 , n57058 , n52978 );
and ( n60685 , n56909 , n52976 );
nor ( n60686 , n60684 , n60685 );
xnor ( n60687 , n60686 , n52680 );
and ( n60688 , n57283 , n52707 );
and ( n60689 , n584529 , n52705 );
nor ( n60690 , n60688 , n60689 );
xnor ( n60691 , n60690 , n52526 );
and ( n60692 , n60687 , n60691 );
xor ( n60693 , n60570 , n587917 );
xor ( n60694 , n60693 , n587920 );
and ( n60695 , n60691 , n60694 );
and ( n60696 , n60687 , n60694 );
or ( n60697 , n60692 , n60695 , n60696 );
and ( n60698 , n56671 , n53177 );
and ( n60699 , n583800 , n53175 );
nor ( n60700 , n60698 , n60699 );
xnor ( n60701 , n60700 , n52827 );
and ( n60702 , n60697 , n60701 );
xor ( n60703 , n587923 , n60604 );
xor ( n60704 , n60703 , n60607 );
and ( n588028 , n60701 , n60704 );
and ( n588029 , n60697 , n60704 );
or ( n60707 , n60702 , n588028 , n588029 );
and ( n588031 , n55841 , n53683 );
and ( n588032 , n583048 , n53681 );
nor ( n588033 , n588031 , n588032 );
xnor ( n60711 , n588033 , n53118 );
and ( n588035 , n60707 , n60711 );
and ( n60713 , n56282 , n53468 );
and ( n60714 , n583377 , n53466 );
nor ( n588038 , n60713 , n60714 );
xnor ( n588039 , n588038 , n52945 );
and ( n60717 , n60711 , n588039 );
and ( n588041 , n60707 , n588039 );
or ( n60719 , n588035 , n60717 , n588041 );
and ( n588043 , n55528 , n53996 );
and ( n588044 , n55293 , n53994 );
nor ( n60722 , n588043 , n588044 );
xnor ( n588046 , n60722 , n53376 );
and ( n588047 , n60719 , n588046 );
xor ( n60725 , n587741 , n60422 );
xor ( n588049 , n60725 , n60427 );
and ( n588050 , n588046 , n588049 );
and ( n60728 , n60719 , n588049 );
or ( n588052 , n588047 , n588050 , n60728 );
and ( n588053 , n55058 , n54414 );
and ( n60731 , n54893 , n54412 );
nor ( n588055 , n588053 , n60731 );
xnor ( n60733 , n588055 , n53650 );
and ( n588057 , n588052 , n60733 );
xor ( n588058 , n60430 , n60434 );
xor ( n60736 , n588058 , n587762 );
and ( n60737 , n60733 , n60736 );
and ( n60738 , n588052 , n60736 );
or ( n588062 , n588057 , n60737 , n60738 );
and ( n60740 , n54553 , n54532 );
and ( n60741 , n54321 , n54530 );
nor ( n60742 , n60740 , n60741 );
xnor ( n588066 , n60742 , n53769 );
and ( n60744 , n588062 , n588066 );
xor ( n60745 , n60442 , n587769 );
xor ( n588069 , n60745 , n60449 );
and ( n60747 , n588066 , n588069 );
and ( n60748 , n588062 , n588069 );
or ( n60749 , n60744 , n60747 , n60748 );
and ( n60750 , n54055 , n55013 );
and ( n588074 , n53835 , n55010 );
nor ( n588075 , n60750 , n588074 );
xnor ( n588076 , n588075 , n53762 );
and ( n60754 , n60749 , n588076 );
xor ( n588078 , n587775 , n587779 );
xor ( n588079 , n588078 , n587782 );
and ( n588080 , n588076 , n588079 );
and ( n588081 , n60749 , n588079 );
or ( n60759 , n60754 , n588080 , n588081 );
xor ( n588083 , n587785 , n587789 );
xor ( n588084 , n588083 , n587792 );
and ( n60762 , n60759 , n588084 );
xor ( n588086 , n60660 , n60664 );
xor ( n588087 , n588086 , n60667 );
and ( n60765 , n588084 , n588087 );
and ( n588089 , n60759 , n588087 );
or ( n588090 , n60762 , n60765 , n588089 );
and ( n588091 , n60683 , n588090 );
nor ( n588092 , n52065 , n52063 );
xnor ( n60770 , n588092 , n52022 );
and ( n588094 , n51990 , n51959 );
and ( n588095 , n60770 , n588094 );
and ( n60773 , n585973 , n52271 );
nor ( n588097 , n52273 , n60773 );
xnor ( n60775 , n588097 , n52137 );
and ( n588099 , n588095 , n60775 );
nor ( n60777 , n52155 , n52153 );
xnor ( n60778 , n60777 , n52085 );
and ( n588102 , n60775 , n60778 );
and ( n588103 , n588095 , n60778 );
or ( n60781 , n588099 , n588102 , n588103 );
xor ( n588105 , n587814 , n60493 );
xor ( n588106 , n588105 , n60496 );
and ( n60784 , n60781 , n588106 );
xor ( n588108 , n587841 , n60526 );
xor ( n588109 , n588108 , n60531 );
and ( n60787 , n588106 , n588109 );
and ( n588111 , n60781 , n588109 );
or ( n588112 , n60784 , n60787 , n588111 );
and ( n60790 , n585586 , n52432 );
and ( n588114 , n58246 , n52430 );
nor ( n588115 , n60790 , n588114 );
xnor ( n588116 , n588115 , n52255 );
and ( n588117 , n588112 , n588116 );
xor ( n60795 , n60534 , n60538 );
xor ( n588119 , n60795 , n587864 );
and ( n588120 , n588116 , n588119 );
and ( n60798 , n588112 , n588119 );
or ( n588122 , n588117 , n588120 , n60798 );
and ( n588123 , n585221 , n52509 );
and ( n60801 , n57900 , n52507 );
nor ( n588125 , n588123 , n60801 );
xnor ( n588126 , n588125 , n52383 );
and ( n60804 , n588122 , n588126 );
xor ( n60805 , n587867 , n60548 );
xor ( n588129 , n60805 , n60551 );
and ( n588130 , n588126 , n588129 );
and ( n60808 , n588122 , n588129 );
or ( n60809 , n60804 , n588130 , n60808 );
and ( n588133 , n57482 , n52707 );
and ( n588134 , n57484 , n52705 );
nor ( n60812 , n588133 , n588134 );
xnor ( n588136 , n60812 , n52526 );
and ( n588137 , n60809 , n588136 );
xor ( n60815 , n60574 , n60578 );
xor ( n588139 , n60815 , n60581 );
and ( n588140 , n588136 , n588139 );
and ( n60818 , n60809 , n588139 );
or ( n60819 , n588137 , n588140 , n60818 );
and ( n588143 , n584529 , n52978 );
and ( n588144 , n57058 , n52976 );
nor ( n60822 , n588143 , n588144 );
xnor ( n60823 , n60822 , n52680 );
and ( n588147 , n60819 , n60823 );
xor ( n588148 , n60584 , n587911 );
xor ( n60826 , n588148 , n587914 );
and ( n588150 , n60823 , n60826 );
and ( n60828 , n60819 , n60826 );
or ( n588152 , n588147 , n588150 , n60828 );
nor ( n588153 , n52273 , n52271 );
xnor ( n60831 , n588153 , n52137 );
nor ( n588155 , n52155 , n52153 );
xnor ( n60833 , n588155 , n52085 );
and ( n60834 , n60831 , n60833 );
nor ( n60835 , n51991 , n51989 );
xnor ( n60836 , n60835 , n51959 );
and ( n60837 , n60833 , n60836 );
and ( n60838 , n60831 , n60836 );
or ( n60839 , n60834 , n60837 , n60838 );
xor ( n60840 , n587843 , n587845 );
xor ( n60841 , n60840 , n51934 );
and ( n60842 , n60839 , n60841 );
xor ( n60843 , n588095 , n60775 );
xor ( n60844 , n60843 , n60778 );
and ( n60845 , n60841 , n60844 );
and ( n60846 , n60839 , n60844 );
or ( n60847 , n60842 , n60845 , n60846 );
and ( n60848 , n585909 , n52432 );
and ( n60849 , n585586 , n52430 );
nor ( n60850 , n60848 , n60849 );
xnor ( n60851 , n60850 , n52255 );
and ( n60852 , n60847 , n60851 );
xor ( n60853 , n60781 , n588106 );
xor ( n60854 , n60853 , n588109 );
and ( n588178 , n60851 , n60854 );
and ( n60856 , n60847 , n60854 );
or ( n60857 , n60852 , n588178 , n60856 );
and ( n60858 , n58219 , n52509 );
and ( n60859 , n585221 , n52507 );
nor ( n60860 , n60858 , n60859 );
xnor ( n60861 , n60860 , n52383 );
and ( n60862 , n60857 , n60861 );
xor ( n588186 , n588112 , n588116 );
xor ( n588187 , n588186 , n588119 );
and ( n60865 , n60861 , n588187 );
and ( n588189 , n60857 , n588187 );
or ( n588190 , n60862 , n60865 , n588189 );
and ( n588191 , n585062 , n52707 );
and ( n588192 , n57482 , n52705 );
nor ( n60870 , n588191 , n588192 );
xnor ( n588194 , n60870 , n52526 );
and ( n588195 , n588190 , n588194 );
xor ( n60873 , n588122 , n588126 );
xor ( n588197 , n60873 , n588129 );
and ( n588198 , n588194 , n588197 );
and ( n60876 , n588190 , n588197 );
or ( n588200 , n588195 , n588198 , n60876 );
xor ( n588201 , n60770 , n588094 );
and ( n60879 , n585973 , n52430 );
nor ( n588203 , n52432 , n60879 );
xnor ( n588204 , n588203 , n52255 );
nor ( n60882 , n52065 , n52063 );
xnor ( n588206 , n60882 , n52022 );
and ( n588207 , n588204 , n588206 );
and ( n60885 , n588206 , n51989 );
and ( n588209 , n588204 , n51989 );
or ( n588210 , n588207 , n60885 , n588209 );
and ( n60888 , n588201 , n588210 );
and ( n588212 , n585973 , n52432 );
and ( n60890 , n58623 , n52430 );
nor ( n60891 , n588212 , n60890 );
xnor ( n60892 , n60891 , n52255 );
and ( n60893 , n588210 , n60892 );
and ( n60894 , n588201 , n60892 );
or ( n60895 , n60888 , n60893 , n60894 );
and ( n60896 , n58623 , n52432 );
and ( n60897 , n585909 , n52430 );
nor ( n60898 , n60896 , n60897 );
xnor ( n60899 , n60898 , n52255 );
and ( n60900 , n60895 , n60899 );
xor ( n60901 , n60839 , n60841 );
xor ( n60902 , n60901 , n60844 );
and ( n60903 , n60899 , n60902 );
and ( n60904 , n60895 , n60902 );
or ( n60905 , n60900 , n60903 , n60904 );
and ( n588229 , n58246 , n52509 );
and ( n588230 , n58219 , n52507 );
nor ( n60908 , n588229 , n588230 );
xnor ( n588232 , n60908 , n52383 );
and ( n60910 , n60905 , n588232 );
xor ( n588234 , n60847 , n60851 );
xor ( n60912 , n588234 , n60854 );
and ( n60913 , n588232 , n60912 );
and ( n588237 , n60905 , n60912 );
or ( n60915 , n60910 , n60913 , n588237 );
and ( n588239 , n57900 , n52707 );
and ( n588240 , n585062 , n52705 );
nor ( n60918 , n588239 , n588240 );
xnor ( n588242 , n60918 , n52526 );
and ( n588243 , n60915 , n588242 );
xor ( n588244 , n60857 , n60861 );
xor ( n588245 , n588244 , n588187 );
and ( n60923 , n588242 , n588245 );
and ( n588247 , n60915 , n588245 );
or ( n60925 , n588243 , n60923 , n588247 );
and ( n588249 , n57484 , n52978 );
and ( n60927 , n57283 , n52976 );
nor ( n60928 , n588249 , n60927 );
xnor ( n588252 , n60928 , n52680 );
and ( n60930 , n60925 , n588252 );
xor ( n588254 , n588190 , n588194 );
xor ( n588255 , n588254 , n588197 );
and ( n60933 , n588252 , n588255 );
and ( n588257 , n60925 , n588255 );
or ( n588258 , n60930 , n60933 , n588257 );
and ( n60936 , n588200 , n588258 );
xor ( n588260 , n60809 , n588136 );
xor ( n588261 , n588260 , n588139 );
and ( n60939 , n588258 , n588261 );
and ( n588263 , n588200 , n588261 );
or ( n588264 , n60936 , n60939 , n588263 );
and ( n60942 , n56909 , n53177 );
and ( n588266 , n56832 , n53175 );
nor ( n60944 , n60942 , n588266 );
xnor ( n60945 , n60944 , n52827 );
and ( n588269 , n588264 , n60945 );
xor ( n588270 , n60819 , n60823 );
xor ( n60948 , n588270 , n60826 );
and ( n60949 , n60945 , n60948 );
and ( n588273 , n588264 , n60948 );
or ( n588274 , n588269 , n60949 , n588273 );
and ( n60952 , n588152 , n588274 );
xor ( n60953 , n60687 , n60691 );
xor ( n60954 , n60953 , n60694 );
and ( n588278 , n588274 , n60954 );
and ( n60956 , n588152 , n60954 );
or ( n60957 , n60952 , n588278 , n60956 );
and ( n60958 , n583377 , n53683 );
and ( n60959 , n55841 , n53681 );
nor ( n60960 , n60958 , n60959 );
xnor ( n60961 , n60960 , n53118 );
and ( n60962 , n60957 , n60961 );
and ( n60963 , n583746 , n53468 );
and ( n60964 , n56282 , n53466 );
nor ( n60965 , n60963 , n60964 );
xnor ( n60966 , n60965 , n52945 );
and ( n60967 , n60961 , n60966 );
and ( n60968 , n60957 , n60966 );
or ( n60969 , n60962 , n60967 , n60968 );
and ( n60970 , n55293 , n54414 );
and ( n60971 , n55075 , n54412 );
nor ( n60972 , n60970 , n60971 );
xnor ( n60973 , n60972 , n53650 );
and ( n588297 , n60969 , n60973 );
xor ( n60975 , n60610 , n60614 );
xor ( n60976 , n60975 , n60617 );
and ( n60977 , n60973 , n60976 );
and ( n60978 , n60969 , n60976 );
or ( n60979 , n588297 , n60977 , n60978 );
and ( n60980 , n55075 , n54414 );
and ( n60981 , n55058 , n54412 );
nor ( n60982 , n60980 , n60981 );
xnor ( n60983 , n60982 , n53650 );
and ( n60984 , n60979 , n60983 );
xor ( n60985 , n587943 , n587947 );
xor ( n60986 , n60985 , n60627 );
and ( n588310 , n60983 , n60986 );
and ( n60988 , n60979 , n60986 );
or ( n60989 , n60984 , n588310 , n60988 );
and ( n588313 , n54725 , n54532 );
and ( n60991 , n54553 , n54530 );
nor ( n588315 , n588313 , n60991 );
xnor ( n60993 , n588315 , n53769 );
and ( n588317 , n60989 , n60993 );
xor ( n60995 , n60630 , n60634 );
xor ( n60996 , n60995 , n587960 );
and ( n60997 , n60993 , n60996 );
and ( n60998 , n60989 , n60996 );
or ( n588322 , n588317 , n60997 , n60998 );
and ( n588323 , n54215 , n55013 );
and ( n61001 , n54055 , n55010 );
nor ( n588325 , n588323 , n61001 );
xnor ( n588326 , n588325 , n53762 );
and ( n588327 , n588322 , n588326 );
xor ( n588328 , n587963 , n587967 );
xor ( n61006 , n588328 , n60647 );
and ( n588330 , n588326 , n61006 );
and ( n588331 , n588322 , n61006 );
or ( n588332 , n588327 , n588330 , n588331 );
xor ( n588333 , n60749 , n588076 );
xor ( n61011 , n588333 , n588079 );
and ( n588335 , n588332 , n61011 );
xor ( n588336 , n60650 , n587977 );
xor ( n61014 , n588336 , n587980 );
and ( n588338 , n61011 , n61014 );
and ( n588339 , n588332 , n61014 );
or ( n61017 , n588335 , n588338 , n588339 );
xor ( n588341 , n60759 , n588084 );
xor ( n588342 , n588341 , n588087 );
and ( n61020 , n61017 , n588342 );
xor ( n588344 , n588332 , n61011 );
xor ( n588345 , n588344 , n61014 );
and ( n61023 , n583800 , n53468 );
and ( n588347 , n583746 , n53466 );
nor ( n588348 , n61023 , n588347 );
xnor ( n61026 , n588348 , n52945 );
and ( n588350 , n56832 , n53177 );
and ( n588351 , n56671 , n53175 );
nor ( n61029 , n588350 , n588351 );
xnor ( n588353 , n61029 , n52827 );
and ( n588354 , n61026 , n588353 );
xor ( n61032 , n588152 , n588274 );
xor ( n588356 , n61032 , n60954 );
and ( n588357 , n588353 , n588356 );
and ( n588358 , n61026 , n588356 );
or ( n588359 , n588354 , n588357 , n588358 );
and ( n61037 , n583048 , n53996 );
and ( n588361 , n582961 , n53994 );
nor ( n588362 , n61037 , n588361 );
xnor ( n61040 , n588362 , n53376 );
and ( n588364 , n588359 , n61040 );
xor ( n588365 , n60697 , n60701 );
xor ( n61043 , n588365 , n60704 );
and ( n61044 , n61040 , n61043 );
and ( n588368 , n588359 , n61043 );
or ( n588369 , n588364 , n61044 , n588368 );
and ( n61047 , n582961 , n53996 );
and ( n61048 , n55528 , n53994 );
nor ( n588372 , n61047 , n61048 );
xnor ( n588373 , n588372 , n53376 );
and ( n61051 , n588369 , n588373 );
xor ( n588375 , n60707 , n60711 );
xor ( n588376 , n588375 , n588039 );
and ( n588377 , n588373 , n588376 );
and ( n61055 , n588369 , n588376 );
or ( n61056 , n61051 , n588377 , n61055 );
and ( n61057 , n54893 , n54532 );
and ( n588381 , n54725 , n54530 );
nor ( n61059 , n61057 , n588381 );
xnor ( n61060 , n61059 , n53769 );
and ( n588384 , n61056 , n61060 );
xor ( n61062 , n60719 , n588046 );
xor ( n588386 , n61062 , n588049 );
and ( n61064 , n61060 , n588386 );
and ( n588388 , n61056 , n588386 );
or ( n588389 , n588384 , n61064 , n588388 );
and ( n61067 , n54321 , n55013 );
and ( n588391 , n54215 , n55010 );
nor ( n588392 , n61067 , n588391 );
xnor ( n61070 , n588392 , n53762 );
and ( n588394 , n588389 , n61070 );
xor ( n588395 , n588052 , n60733 );
xor ( n61073 , n588395 , n60736 );
and ( n588397 , n61070 , n61073 );
and ( n61075 , n588389 , n61073 );
or ( n588399 , n588394 , n588397 , n61075 );
xor ( n61077 , n588322 , n588326 );
xor ( n61078 , n61077 , n61006 );
and ( n588402 , n588399 , n61078 );
xor ( n61080 , n588062 , n588066 );
xor ( n588404 , n61080 , n588069 );
and ( n588405 , n61078 , n588404 );
and ( n61083 , n588399 , n588404 );
or ( n588407 , n588402 , n588405 , n61083 );
and ( n588408 , n588345 , n588407 );
xor ( n61086 , n588399 , n61078 );
xor ( n61087 , n61086 , n588404 );
and ( n61088 , n57058 , n53177 );
and ( n61089 , n56909 , n53175 );
nor ( n61090 , n61088 , n61089 );
xnor ( n588414 , n61090 , n52827 );
and ( n61092 , n57283 , n52978 );
and ( n61093 , n584529 , n52976 );
nor ( n61094 , n61092 , n61093 );
xnor ( n61095 , n61094 , n52680 );
and ( n61096 , n588414 , n61095 );
xor ( n61097 , n588200 , n588258 );
xor ( n588421 , n61097 , n588261 );
and ( n61099 , n61095 , n588421 );
and ( n588423 , n588414 , n588421 );
or ( n588424 , n61096 , n61099 , n588423 );
and ( n61102 , n583746 , n53683 );
and ( n588426 , n56282 , n53681 );
nor ( n588427 , n61102 , n588426 );
xnor ( n61105 , n588427 , n53118 );
and ( n61106 , n588424 , n61105 );
xor ( n588430 , n588264 , n60945 );
xor ( n61108 , n588430 , n60948 );
and ( n61109 , n61105 , n61108 );
and ( n61110 , n588424 , n61108 );
or ( n61111 , n61106 , n61109 , n61110 );
and ( n588435 , n55841 , n53996 );
and ( n588436 , n583048 , n53994 );
nor ( n588437 , n588435 , n588436 );
xnor ( n61115 , n588437 , n53376 );
and ( n588439 , n61111 , n61115 );
and ( n588440 , n56282 , n53683 );
and ( n588441 , n583377 , n53681 );
nor ( n61119 , n588440 , n588441 );
xnor ( n588443 , n61119 , n53118 );
and ( n61121 , n61115 , n588443 );
and ( n588445 , n61111 , n588443 );
or ( n588446 , n588439 , n61121 , n588445 );
and ( n61124 , n55528 , n54414 );
and ( n588448 , n55293 , n54412 );
nor ( n61126 , n61124 , n588448 );
xnor ( n588450 , n61126 , n53650 );
and ( n588451 , n588446 , n588450 );
xor ( n61129 , n60957 , n60961 );
xor ( n588453 , n61129 , n60966 );
and ( n588454 , n588450 , n588453 );
and ( n588455 , n588446 , n588453 );
or ( n61133 , n588451 , n588454 , n588455 );
and ( n588457 , n55058 , n54532 );
and ( n61135 , n54893 , n54530 );
nor ( n588459 , n588457 , n61135 );
xnor ( n588460 , n588459 , n53769 );
and ( n61138 , n61133 , n588460 );
xor ( n588462 , n60969 , n60973 );
xor ( n61140 , n588462 , n60976 );
and ( n61141 , n588460 , n61140 );
and ( n61142 , n61133 , n61140 );
or ( n588466 , n61138 , n61141 , n61142 );
and ( n588467 , n54553 , n55013 );
and ( n61145 , n54321 , n55010 );
nor ( n588469 , n588467 , n61145 );
xnor ( n588470 , n588469 , n53762 );
and ( n588471 , n588466 , n588470 );
xor ( n588472 , n60979 , n60983 );
xor ( n61150 , n588472 , n60986 );
and ( n588474 , n588470 , n61150 );
and ( n588475 , n588466 , n61150 );
or ( n61153 , n588471 , n588474 , n588475 );
xor ( n588477 , n588389 , n61070 );
xor ( n588478 , n588477 , n61073 );
and ( n61156 , n61153 , n588478 );
xor ( n588480 , n60989 , n60993 );
xor ( n588481 , n588480 , n60996 );
and ( n61159 , n588478 , n588481 );
and ( n588483 , n61153 , n588481 );
or ( n61161 , n61156 , n61159 , n588483 );
and ( n61162 , n61087 , n61161 );
xor ( n588486 , n61056 , n61060 );
xor ( n588487 , n588486 , n588386 );
xor ( n588488 , n588466 , n588470 );
xor ( n61166 , n588488 , n61150 );
and ( n588490 , n588487 , n61166 );
and ( n588491 , n54725 , n55013 );
and ( n588492 , n54553 , n55010 );
nor ( n588493 , n588491 , n588492 );
xnor ( n61171 , n588493 , n53762 );
xor ( n588495 , n588369 , n588373 );
xor ( n588496 , n588495 , n588376 );
and ( n61174 , n61171 , n588496 );
and ( n588498 , n61166 , n61174 );
and ( n588499 , n588487 , n61174 );
or ( n61177 , n588490 , n588498 , n588499 );
xor ( n588501 , n61153 , n588478 );
xor ( n588502 , n588501 , n588481 );
and ( n61180 , n61177 , n588502 );
and ( n61181 , n55058 , n55013 );
and ( n61182 , n54893 , n55010 );
nor ( n588506 , n61181 , n61182 );
xnor ( n61184 , n588506 , n53762 );
and ( n61185 , n582961 , n54414 );
and ( n61186 , n55528 , n54412 );
nor ( n588510 , n61185 , n61186 );
xnor ( n588511 , n588510 , n53650 );
and ( n61189 , n61184 , n588511 );
and ( n588513 , n55075 , n55013 );
and ( n588514 , n55058 , n55010 );
nor ( n588515 , n588513 , n588514 );
xnor ( n588516 , n588515 , n53762 );
and ( n61194 , n55528 , n54532 );
and ( n588518 , n55293 , n54530 );
nor ( n588519 , n61194 , n588518 );
xnor ( n61197 , n588519 , n53769 );
and ( n588521 , n588516 , n61197 );
and ( n588522 , n583048 , n54414 );
and ( n61200 , n582961 , n54412 );
nor ( n588524 , n588522 , n61200 );
xnor ( n588525 , n588524 , n53650 );
and ( n61203 , n61197 , n588525 );
and ( n588527 , n588516 , n588525 );
or ( n61205 , n588521 , n61203 , n588527 );
and ( n61206 , n588511 , n61205 );
and ( n61207 , n61184 , n61205 );
or ( n61208 , n61189 , n61206 , n61207 );
and ( n61209 , n583377 , n53996 );
and ( n588533 , n55841 , n53994 );
nor ( n61211 , n61209 , n588533 );
xnor ( n588535 , n61211 , n53376 );
and ( n588536 , n56671 , n53468 );
and ( n61214 , n583800 , n53466 );
nor ( n588538 , n588536 , n61214 );
xnor ( n588539 , n588538 , n52945 );
and ( n61217 , n588535 , n588539 );
and ( n588541 , n583800 , n53683 );
and ( n588542 , n583746 , n53681 );
nor ( n588543 , n588541 , n588542 );
xnor ( n588544 , n588543 , n53118 );
and ( n61222 , n56832 , n53468 );
and ( n588546 , n56671 , n53466 );
nor ( n588547 , n61222 , n588546 );
xnor ( n61225 , n588547 , n52945 );
and ( n588549 , n588544 , n61225 );
and ( n61227 , n588539 , n588549 );
and ( n588551 , n588535 , n588549 );
or ( n61229 , n61217 , n61227 , n588551 );
xor ( n61230 , n61184 , n588511 );
xor ( n588554 , n61230 , n61205 );
and ( n61232 , n61229 , n588554 );
and ( n588556 , n55293 , n55013 );
and ( n588557 , n55075 , n55010 );
nor ( n588558 , n588556 , n588557 );
xnor ( n61236 , n588558 , n53762 );
and ( n588560 , n582961 , n54532 );
and ( n588561 , n55528 , n54530 );
nor ( n61239 , n588560 , n588561 );
xnor ( n588563 , n61239 , n53769 );
and ( n588564 , n61236 , n588563 );
xor ( n61242 , n588516 , n61197 );
xor ( n588566 , n61242 , n588525 );
and ( n588567 , n588564 , n588566 );
and ( n588568 , n55841 , n54414 );
and ( n61246 , n583048 , n54412 );
nor ( n61247 , n588568 , n61246 );
xnor ( n588571 , n61247 , n53650 );
and ( n61249 , n56282 , n53996 );
and ( n588573 , n583377 , n53994 );
nor ( n588574 , n61249 , n588573 );
xnor ( n61252 , n588574 , n53376 );
and ( n588576 , n588571 , n61252 );
xor ( n61254 , n588544 , n61225 );
and ( n588578 , n61252 , n61254 );
and ( n61256 , n588571 , n61254 );
or ( n588580 , n588576 , n588578 , n61256 );
and ( n588581 , n588566 , n588580 );
and ( n61259 , n588564 , n588580 );
or ( n61260 , n588567 , n588581 , n61259 );
and ( n588584 , n588554 , n61260 );
and ( n588585 , n61229 , n61260 );
or ( n61263 , n61232 , n588584 , n588585 );
and ( n588587 , n61208 , n61263 );
xor ( n588588 , n61236 , n588563 );
and ( n61266 , n55528 , n55013 );
and ( n588590 , n55293 , n55010 );
nor ( n588591 , n61266 , n588590 );
xnor ( n61269 , n588591 , n53762 );
and ( n588593 , n583048 , n54532 );
and ( n588594 , n582961 , n54530 );
nor ( n61272 , n588593 , n588594 );
xnor ( n61273 , n61272 , n53769 );
and ( n588597 , n61269 , n61273 );
and ( n588598 , n583377 , n54414 );
and ( n61276 , n55841 , n54412 );
nor ( n588600 , n588598 , n61276 );
xnor ( n61278 , n588600 , n53650 );
and ( n588602 , n61273 , n61278 );
and ( n588603 , n61269 , n61278 );
or ( n61281 , n588597 , n588602 , n588603 );
and ( n588605 , n588588 , n61281 );
and ( n61283 , n583746 , n53996 );
and ( n61284 , n56282 , n53994 );
nor ( n61285 , n61283 , n61284 );
xnor ( n61286 , n61285 , n53376 );
and ( n61287 , n56671 , n53683 );
and ( n61288 , n583800 , n53681 );
nor ( n61289 , n61287 , n61288 );
xnor ( n61290 , n61289 , n53118 );
and ( n61291 , n61286 , n61290 );
and ( n61292 , n56909 , n53468 );
and ( n61293 , n56832 , n53466 );
nor ( n61294 , n61292 , n61293 );
xnor ( n61295 , n61294 , n52945 );
and ( n61296 , n61290 , n61295 );
and ( n61297 , n61286 , n61295 );
or ( n61298 , n61291 , n61296 , n61297 );
and ( n61299 , n61281 , n61298 );
and ( n61300 , n588588 , n61298 );
or ( n61301 , n588605 , n61299 , n61300 );
xor ( n61302 , n588535 , n588539 );
xor ( n61303 , n61302 , n588549 );
and ( n61304 , n61301 , n61303 );
and ( n61305 , n583800 , n53996 );
and ( n588629 , n583746 , n53994 );
nor ( n61307 , n61305 , n588629 );
xnor ( n61308 , n61307 , n53376 );
and ( n588632 , n56832 , n53683 );
and ( n61310 , n56671 , n53681 );
nor ( n588634 , n588632 , n61310 );
xnor ( n61312 , n588634 , n53118 );
and ( n588636 , n61308 , n61312 );
and ( n588637 , n582961 , n55013 );
and ( n61315 , n55528 , n55010 );
nor ( n588639 , n588637 , n61315 );
xnor ( n588640 , n588639 , n53762 );
and ( n61318 , n55841 , n54532 );
and ( n61319 , n583048 , n54530 );
nor ( n588643 , n61318 , n61319 );
xnor ( n588644 , n588643 , n53769 );
and ( n61322 , n588640 , n588644 );
and ( n588646 , n56282 , n54414 );
and ( n588647 , n583377 , n54412 );
nor ( n61325 , n588646 , n588647 );
xnor ( n588649 , n61325 , n53650 );
and ( n588650 , n588644 , n588649 );
and ( n61328 , n588640 , n588649 );
or ( n61329 , n61322 , n588650 , n61328 );
and ( n61330 , n588636 , n61329 );
xor ( n61331 , n61269 , n61273 );
xor ( n61332 , n61331 , n61278 );
and ( n61333 , n61329 , n61332 );
and ( n61334 , n588636 , n61332 );
or ( n61335 , n61330 , n61333 , n61334 );
xor ( n61336 , n588571 , n61252 );
xor ( n61337 , n61336 , n61254 );
and ( n61338 , n61335 , n61337 );
xor ( n61339 , n588588 , n61281 );
xor ( n61340 , n61339 , n61298 );
and ( n61341 , n61337 , n61340 );
and ( n588665 , n61335 , n61340 );
or ( n61343 , n61338 , n61341 , n588665 );
and ( n61344 , n61303 , n61343 );
and ( n588668 , n61301 , n61343 );
or ( n588669 , n61304 , n61344 , n588668 );
xor ( n61347 , n61229 , n588554 );
xor ( n588671 , n61347 , n61260 );
and ( n588672 , n588669 , n588671 );
xor ( n588673 , n588564 , n588566 );
xor ( n61351 , n588673 , n588580 );
xor ( n588675 , n61301 , n61303 );
xor ( n61353 , n588675 , n61343 );
and ( n588677 , n61351 , n61353 );
xor ( n61355 , n61286 , n61290 );
xor ( n61356 , n61355 , n61295 );
and ( n588680 , n57058 , n53468 );
and ( n61358 , n56909 , n53466 );
nor ( n588682 , n588680 , n61358 );
xnor ( n588683 , n588682 , n52945 );
and ( n61361 , n57283 , n53177 );
and ( n588685 , n584529 , n53175 );
nor ( n61363 , n61361 , n588685 );
xnor ( n61364 , n61363 , n52827 );
and ( n61365 , n588683 , n61364 );
xor ( n588689 , n61308 , n61312 );
and ( n588690 , n61364 , n588689 );
and ( n61368 , n588683 , n588689 );
or ( n588692 , n61365 , n588690 , n61368 );
and ( n588693 , n61356 , n588692 );
and ( n588694 , n583048 , n55013 );
and ( n588695 , n582961 , n55010 );
nor ( n61373 , n588694 , n588695 );
xnor ( n588697 , n61373 , n53762 );
and ( n588698 , n583377 , n54532 );
and ( n61376 , n55841 , n54530 );
nor ( n588700 , n588698 , n61376 );
xnor ( n588701 , n588700 , n53769 );
and ( n61379 , n588697 , n588701 );
and ( n588703 , n583746 , n54414 );
and ( n588704 , n56282 , n54412 );
nor ( n61382 , n588703 , n588704 );
xnor ( n588706 , n61382 , n53650 );
and ( n61384 , n588701 , n588706 );
and ( n61385 , n588697 , n588706 );
or ( n61386 , n61379 , n61384 , n61385 );
and ( n61387 , n56671 , n53996 );
and ( n588711 , n583800 , n53994 );
nor ( n61389 , n61387 , n588711 );
xnor ( n61390 , n61389 , n53376 );
and ( n61391 , n56909 , n53683 );
and ( n61392 , n56832 , n53681 );
nor ( n61393 , n61391 , n61392 );
xnor ( n61394 , n61393 , n53118 );
and ( n61395 , n61390 , n61394 );
and ( n61396 , n584529 , n53468 );
and ( n61397 , n57058 , n53466 );
nor ( n61398 , n61396 , n61397 );
xnor ( n61399 , n61398 , n52945 );
and ( n588723 , n61394 , n61399 );
and ( n588724 , n61390 , n61399 );
or ( n61402 , n61395 , n588723 , n588724 );
and ( n588726 , n61386 , n61402 );
xor ( n61404 , n588640 , n588644 );
xor ( n61405 , n61404 , n588649 );
and ( n61406 , n61402 , n61405 );
and ( n61407 , n61386 , n61405 );
or ( n61408 , n588726 , n61406 , n61407 );
and ( n61409 , n588692 , n61408 );
and ( n61410 , n61356 , n61408 );
or ( n588734 , n588693 , n61409 , n61410 );
xor ( n61412 , n61335 , n61337 );
xor ( n588736 , n61412 , n61340 );
and ( n61414 , n588734 , n588736 );
xor ( n61415 , n588636 , n61329 );
xor ( n588739 , n61415 , n61332 );
and ( n61417 , n57484 , n53177 );
and ( n588741 , n57283 , n53175 );
nor ( n61419 , n61417 , n588741 );
xnor ( n61420 , n61419 , n52827 );
and ( n588744 , n585062 , n52978 );
and ( n61422 , n57482 , n52976 );
nor ( n61423 , n588744 , n61422 );
xnor ( n61424 , n61423 , n52680 );
and ( n61425 , n61420 , n61424 );
and ( n61426 , n55841 , n55013 );
and ( n61427 , n583048 , n55010 );
nor ( n61428 , n61426 , n61427 );
xnor ( n61429 , n61428 , n53762 );
and ( n61430 , n56282 , n54532 );
and ( n588754 , n583377 , n54530 );
nor ( n588755 , n61430 , n588754 );
xnor ( n61433 , n588755 , n53769 );
and ( n588757 , n61429 , n61433 );
and ( n61435 , n583800 , n54414 );
and ( n588759 , n583746 , n54412 );
nor ( n588760 , n61435 , n588759 );
xnor ( n588761 , n588760 , n53650 );
and ( n61439 , n61433 , n588761 );
and ( n588763 , n61429 , n588761 );
or ( n61441 , n588757 , n61439 , n588763 );
and ( n588765 , n61424 , n61441 );
and ( n588766 , n61420 , n61441 );
or ( n61444 , n61425 , n588765 , n588766 );
and ( n588768 , n56832 , n53996 );
and ( n61446 , n56671 , n53994 );
nor ( n61447 , n588768 , n61446 );
xnor ( n61448 , n61447 , n53376 );
and ( n61449 , n57058 , n53683 );
and ( n588773 , n56909 , n53681 );
nor ( n588774 , n61449 , n588773 );
xnor ( n61452 , n588774 , n53118 );
and ( n588776 , n61448 , n61452 );
and ( n588777 , n57283 , n53468 );
and ( n588778 , n584529 , n53466 );
nor ( n588779 , n588777 , n588778 );
xnor ( n61457 , n588779 , n52945 );
and ( n588781 , n61452 , n61457 );
and ( n588782 , n61448 , n61457 );
or ( n61460 , n588776 , n588781 , n588782 );
and ( n588784 , n57482 , n53177 );
and ( n588785 , n57484 , n53175 );
nor ( n61463 , n588784 , n588785 );
xnor ( n588787 , n61463 , n52827 );
and ( n588788 , n57900 , n52978 );
and ( n61466 , n585062 , n52976 );
nor ( n588790 , n588788 , n61466 );
xnor ( n588791 , n588790 , n52680 );
and ( n588792 , n588787 , n588791 );
and ( n588793 , n58219 , n52707 );
and ( n61471 , n585221 , n52705 );
nor ( n588795 , n588793 , n61471 );
xnor ( n588796 , n588795 , n52526 );
and ( n588797 , n588791 , n588796 );
and ( n588798 , n588787 , n588796 );
or ( n61476 , n588792 , n588797 , n588798 );
and ( n588800 , n61460 , n61476 );
xor ( n588801 , n588697 , n588701 );
xor ( n61479 , n588801 , n588706 );
and ( n588803 , n61476 , n61479 );
and ( n588804 , n61460 , n61479 );
or ( n61482 , n588800 , n588803 , n588804 );
and ( n588806 , n61444 , n61482 );
xor ( n588807 , n588683 , n61364 );
xor ( n61485 , n588807 , n588689 );
and ( n588809 , n61482 , n61485 );
and ( n588810 , n61444 , n61485 );
or ( n61488 , n588806 , n588809 , n588810 );
and ( n588812 , n588739 , n61488 );
xor ( n61490 , n61356 , n588692 );
xor ( n588814 , n61490 , n61408 );
and ( n61492 , n61488 , n588814 );
and ( n588816 , n588739 , n588814 );
or ( n61494 , n588812 , n61492 , n588816 );
and ( n588818 , n588736 , n61494 );
and ( n61496 , n588734 , n61494 );
or ( n61497 , n61414 , n588818 , n61496 );
and ( n588821 , n61353 , n61497 );
and ( n588822 , n61351 , n61497 );
or ( n61500 , n588677 , n588821 , n588822 );
and ( n61501 , n588671 , n61500 );
and ( n588825 , n588669 , n61500 );
or ( n588826 , n588672 , n61501 , n588825 );
and ( n61504 , n61263 , n588826 );
and ( n588828 , n61208 , n588826 );
or ( n588829 , n588587 , n61504 , n588828 );
xor ( n61507 , n61133 , n588460 );
xor ( n588831 , n61507 , n61140 );
and ( n588832 , n588829 , n588831 );
and ( n61510 , n55075 , n54532 );
and ( n61511 , n55058 , n54530 );
nor ( n588835 , n61510 , n61511 );
xnor ( n588836 , n588835 , n53769 );
xor ( n61514 , n588359 , n61040 );
xor ( n61515 , n61514 , n61043 );
and ( n588839 , n588836 , n61515 );
and ( n588840 , n588831 , n588839 );
and ( n61518 , n588829 , n588839 );
or ( n61519 , n588832 , n588840 , n61518 );
and ( n61520 , n54893 , n55013 );
and ( n61521 , n54725 , n55010 );
nor ( n588845 , n61520 , n61521 );
xnor ( n588846 , n588845 , n53762 );
xor ( n61524 , n588446 , n588450 );
xor ( n588848 , n61524 , n588453 );
and ( n61526 , n588846 , n588848 );
xor ( n588850 , n61208 , n61263 );
xor ( n61528 , n588850 , n588826 );
and ( n61529 , n55293 , n54532 );
and ( n588853 , n55075 , n54530 );
nor ( n588854 , n61529 , n588853 );
xnor ( n61532 , n588854 , n53769 );
xor ( n61533 , n61111 , n61115 );
xor ( n588857 , n61533 , n588443 );
and ( n61535 , n61532 , n588857 );
and ( n61536 , n61528 , n61535 );
xor ( n61537 , n588669 , n588671 );
xor ( n61538 , n61537 , n61500 );
xor ( n61539 , n61026 , n588353 );
xor ( n588863 , n61539 , n588356 );
and ( n61541 , n61538 , n588863 );
xor ( n61542 , n61351 , n61353 );
xor ( n61543 , n61542 , n61497 );
xor ( n588867 , n588424 , n61105 );
xor ( n588868 , n588867 , n61108 );
and ( n61546 , n61543 , n588868 );
nor ( n588870 , n52273 , n52271 );
xnor ( n588871 , n588870 , n52137 );
nor ( n61549 , n52155 , n52153 );
xnor ( n61550 , n61549 , n52085 );
and ( n588874 , n588871 , n61550 );
xor ( n61552 , n60831 , n60833 );
xor ( n61553 , n61552 , n60836 );
and ( n61554 , n588874 , n61553 );
xor ( n61555 , n588201 , n588210 );
xor ( n588879 , n61555 , n60892 );
and ( n61557 , n61553 , n588879 );
and ( n61558 , n588874 , n588879 );
or ( n61559 , n61554 , n61557 , n61558 );
and ( n61560 , n585586 , n52509 );
and ( n588884 , n58246 , n52507 );
nor ( n588885 , n61560 , n588884 );
xnor ( n588886 , n588885 , n52383 );
and ( n61564 , n61559 , n588886 );
xor ( n588888 , n60895 , n60899 );
xor ( n61566 , n588888 , n60902 );
and ( n61567 , n588886 , n61566 );
and ( n588891 , n61559 , n61566 );
or ( n588892 , n61564 , n61567 , n588891 );
and ( n61570 , n585221 , n52707 );
and ( n61571 , n57900 , n52705 );
nor ( n588895 , n61570 , n61571 );
xnor ( n588896 , n588895 , n52526 );
and ( n61574 , n588892 , n588896 );
xor ( n588898 , n60905 , n588232 );
xor ( n588899 , n588898 , n60912 );
and ( n588900 , n588896 , n588899 );
and ( n588901 , n588892 , n588899 );
or ( n61579 , n61574 , n588900 , n588901 );
and ( n588903 , n57482 , n52978 );
and ( n61581 , n57484 , n52976 );
nor ( n588905 , n588903 , n61581 );
xnor ( n588906 , n588905 , n52680 );
and ( n61584 , n61579 , n588906 );
xor ( n61585 , n60915 , n588242 );
xor ( n61586 , n61585 , n588245 );
and ( n61587 , n588906 , n61586 );
and ( n588911 , n61579 , n61586 );
or ( n61589 , n61584 , n61587 , n588911 );
and ( n61590 , n584529 , n53177 );
and ( n61591 , n57058 , n53175 );
nor ( n61592 , n61590 , n61591 );
xnor ( n588916 , n61592 , n52827 );
and ( n588917 , n61589 , n588916 );
xor ( n61595 , n60925 , n588252 );
xor ( n61596 , n61595 , n588255 );
and ( n61597 , n588916 , n61596 );
and ( n61598 , n61589 , n61596 );
or ( n61599 , n588917 , n61597 , n61598 );
xor ( n588923 , n588414 , n61095 );
xor ( n588924 , n588923 , n588421 );
and ( n588925 , n61599 , n588924 );
and ( n61603 , n588868 , n588925 );
and ( n588927 , n61543 , n588925 );
or ( n588928 , n61546 , n61603 , n588927 );
and ( n61606 , n588863 , n588928 );
and ( n588930 , n61538 , n588928 );
or ( n588931 , n61541 , n61606 , n588930 );
and ( n61609 , n61535 , n588931 );
and ( n61610 , n61528 , n588931 );
or ( n588934 , n61536 , n61609 , n61610 );
and ( n588935 , n61526 , n588934 );
xor ( n61613 , n61171 , n588496 );
and ( n61614 , n588934 , n61613 );
and ( n588938 , n61526 , n61613 );
or ( n588939 , n588935 , n61614 , n588938 );
and ( n61617 , n61519 , n588939 );
xor ( n61618 , n588487 , n61166 );
xor ( n61619 , n61618 , n61174 );
and ( n61620 , n588939 , n61619 );
and ( n588944 , n61519 , n61619 );
or ( n588945 , n61617 , n61620 , n588944 );
and ( n61623 , n588502 , n588945 );
and ( n588947 , n61177 , n588945 );
or ( n588948 , n61180 , n61623 , n588947 );
and ( n61626 , n61161 , n588948 );
and ( n588950 , n61087 , n588948 );
or ( n588951 , n61162 , n61626 , n588950 );
and ( n61629 , n588407 , n588951 );
and ( n588953 , n588345 , n588951 );
or ( n61631 , n588408 , n61629 , n588953 );
and ( n61632 , n588342 , n61631 );
and ( n61633 , n61017 , n61631 );
or ( n61634 , n61020 , n61632 , n61633 );
and ( n61635 , n588090 , n61634 );
and ( n588959 , n60683 , n61634 );
or ( n588960 , n588091 , n61635 , n588959 );
and ( n61638 , n60680 , n588960 );
and ( n61639 , n60678 , n588960 );
or ( n61640 , n60681 , n61638 , n61639 );
and ( n61641 , n587811 , n61640 );
and ( n588965 , n60374 , n61640 );
or ( n588966 , n60489 , n61641 , n588965 );
and ( n61644 , n60371 , n588966 );
and ( n588968 , n60225 , n588966 );
or ( n61646 , n587695 , n61644 , n588968 );
and ( n588970 , n60222 , n61646 );
and ( n61648 , n587278 , n61646 );
or ( n588972 , n60223 , n588970 , n61648 );
and ( n588973 , n59952 , n588972 );
and ( n61651 , n59860 , n588972 );
or ( n588975 , n587276 , n588973 , n61651 );
and ( n588976 , n59857 , n588975 );
and ( n61654 , n59635 , n588975 );
or ( n588978 , n587181 , n588976 , n61654 );
and ( n61656 , n586955 , n588978 );
and ( n61657 , n586793 , n588978 );
or ( n61658 , n59633 , n61656 , n61657 );
and ( n61659 , n586790 , n61658 );
and ( n61660 , n59465 , n61658 );
or ( n588984 , n59468 , n61659 , n61660 );
and ( n61662 , n586619 , n588984 );
and ( n588986 , n59052 , n588984 );
or ( n588987 , n59297 , n61662 , n588986 );
and ( n61665 , n586372 , n588987 );
and ( n588989 , n59011 , n588987 );
or ( n588990 , n586373 , n61665 , n588989 );
and ( n61668 , n586331 , n588990 );
and ( n61669 , n586155 , n588990 );
or ( n61670 , n59009 , n61668 , n61669 );
and ( n61671 , n586152 , n61670 );
and ( n588995 , n58576 , n61670 );
or ( n588996 , n586153 , n61671 , n588995 );
and ( n588997 , n585896 , n588996 );
and ( n588998 , n58389 , n588996 );
or ( n61676 , n58574 , n588997 , n588998 );
and ( n589000 , n585709 , n61676 );
and ( n589001 , n58173 , n61676 );
or ( n61679 , n58387 , n589000 , n589001 );
and ( n61680 , n58170 , n61679 );
and ( n61681 , n58122 , n61679 );
or ( n61682 , n58171 , n61680 , n61681 );
and ( n589006 , n58119 , n61682 );
and ( n61684 , n57879 , n61682 );
or ( n61685 , n58120 , n589006 , n61684 );
and ( n61686 , n585199 , n61685 );
and ( n61687 , n585022 , n61685 );
or ( n61688 , n585200 , n61686 , n61687 );
and ( n589012 , n57696 , n61688 );
and ( n589013 , n57472 , n61688 );
or ( n61691 , n57697 , n589012 , n589013 );
and ( n589015 , n57469 , n61691 );
and ( n589016 , n57423 , n61691 );
or ( n589017 , n57470 , n589015 , n589016 );
and ( n589018 , n584743 , n589017 );
and ( n61696 , n57196 , n589017 );
or ( n589020 , n57421 , n589018 , n61696 );
and ( n589021 , n57193 , n589020 );
and ( n61699 , n57034 , n589020 );
or ( n589023 , n57194 , n589021 , n61699 );
and ( n61701 , n57031 , n589023 );
and ( n589025 , n56791 , n589023 );
or ( n61703 , n57032 , n61701 , n589025 );
and ( n61704 , n56788 , n61703 );
and ( n589028 , n583952 , n61703 );
or ( n589029 , n584112 , n61704 , n589028 );
and ( n61707 , n583949 , n589029 );
and ( n589031 , n583727 , n589029 );
or ( n589032 , n583950 , n61707 , n589031 );
and ( n61710 , n583724 , n589032 );
and ( n589034 , n56244 , n589032 );
or ( n589035 , n583725 , n61710 , n589034 );
and ( n61713 , n56241 , n589035 );
and ( n589037 , n583367 , n589035 );
or ( n589038 , n583565 , n61713 , n589037 );
and ( n589039 , n583364 , n589038 );
and ( n589040 , n56023 , n589038 );
or ( n61718 , n56042 , n589039 , n589040 );
and ( n589042 , n56020 , n61718 );
and ( n589043 , n55831 , n61718 );
or ( n589044 , n56021 , n589042 , n589043 );
and ( n589045 , n583151 , n589044 );
and ( n61723 , n55628 , n589044 );
or ( n589047 , n55829 , n589045 , n61723 );
and ( n589048 , n55625 , n589047 );
and ( n61726 , n55470 , n589047 );
or ( n589050 , n582949 , n589048 , n61726 );
and ( n589051 , n582790 , n589050 );
and ( n61729 , n55419 , n589050 );
or ( n589053 , n55468 , n589051 , n61729 );
and ( n589054 , n55416 , n589053 );
and ( n61732 , n55187 , n589053 );
or ( n61733 , n55417 , n589054 , n61732 );
and ( n61734 , n55184 , n61733 );
and ( n589058 , n55009 , n61733 );
or ( n589059 , n55185 , n61734 , n589058 );
and ( n61737 , n55006 , n589059 );
and ( n589061 , n55004 , n589059 );
or ( n589062 , n55007 , n61737 , n589061 );
and ( n61740 , n54826 , n589062 );
and ( n589064 , n54649 , n589062 );
or ( n589065 , n54827 , n61740 , n589064 );
and ( n589066 , n54646 , n589065 );
and ( n61744 , n54644 , n589065 );
or ( n589068 , n54647 , n589066 , n61744 );
and ( n61746 , n54469 , n589068 );
and ( n589070 , n54297 , n589068 );
or ( n589071 , n54470 , n61746 , n589070 );
and ( n61749 , n54294 , n589071 );
and ( n589073 , n54149 , n589071 );
or ( n61751 , n54295 , n61749 , n589073 );
and ( n61752 , n54146 , n61751 );
and ( n61753 , n53978 , n61751 );
or ( n589077 , n54147 , n61752 , n61753 );
and ( n61755 , n53975 , n589077 );
and ( n61756 , n53745 , n589077 );
or ( n61757 , n53976 , n61755 , n61756 );
and ( n589081 , n53742 , n61757 );
and ( n589082 , n53638 , n61757 );
or ( n589083 , n53743 , n589081 , n589082 );
and ( n61761 , n53635 , n589083 );
and ( n589085 , n53633 , n589083 );
or ( n589086 , n53636 , n61761 , n589085 );
and ( n61764 , n53498 , n589086 );
and ( n589088 , n53496 , n589086 );
or ( n61766 , n53499 , n61764 , n589088 );
and ( n589090 , n53354 , n61766 );
and ( n61768 , n53211 , n61766 );
or ( n589092 , n53355 , n589090 , n61768 );
and ( n589093 , n53208 , n589092 );
and ( n61771 , n53106 , n589092 );
or ( n589095 , n53209 , n589093 , n61771 );
and ( n61773 , n53103 , n589095 );
and ( n61774 , n53009 , n589095 );
or ( n61775 , n53104 , n61773 , n61774 );
and ( n61776 , n53006 , n61775 );
and ( n61777 , n52883 , n61775 );
or ( n61778 , n53007 , n61776 , n61777 );
and ( n61779 , n52880 , n61778 );
and ( n61780 , n52771 , n61778 );
or ( n61781 , n52881 , n61779 , n61780 );
and ( n61782 , n52768 , n61781 );
and ( n61783 , n52668 , n61781 );
or ( n589107 , n52769 , n61782 , n61783 );
and ( n61785 , n52665 , n589107 );
and ( n589109 , n52575 , n589107 );
or ( n61787 , n52666 , n61785 , n589109 );
and ( n589111 , n52572 , n61787 );
and ( n61789 , n52570 , n61787 );
or ( n589113 , n52573 , n589111 , n61789 );
and ( n61791 , n52477 , n589113 );
and ( n589115 , n52362 , n589113 );
or ( n61793 , n52478 , n61791 , n589115 );
and ( n61794 , n52359 , n61793 );
and ( n61795 , n52303 , n61793 );
or ( n589119 , n52360 , n61794 , n61795 );
and ( n589120 , n52300 , n589119 );
and ( n61798 , n52250 , n589119 );
or ( n589122 , n52301 , n589120 , n61798 );
and ( n589123 , n52247 , n589122 );
and ( n61801 , n52193 , n589122 );
or ( n589125 , n52248 , n589123 , n61801 );
and ( n61803 , n52190 , n589125 );
and ( n589127 , n52114 , n589125 );
or ( n61805 , n52191 , n61803 , n589127 );
and ( n61806 , n52111 , n61805 );
and ( n589130 , n52061 , n61805 );
or ( n589131 , n52112 , n61806 , n589130 );
and ( n61809 , n52058 , n589131 );
and ( n589133 , n52017 , n589131 );
or ( n589134 , n52059 , n61809 , n589133 );
and ( n589135 , n52014 , n589134 );
and ( n61813 , n51987 , n589134 );
or ( n589137 , n52015 , n589135 , n61813 );
and ( n61815 , n51984 , n589137 );
and ( n589139 , n51982 , n589137 );
or ( n61817 , n51985 , n61815 , n589139 );
xor ( n61818 , n51954 , n61817 );
not ( n589142 , n61818 );
xor ( n589143 , n51982 , n51984 );
xor ( n61821 , n589143 , n589137 );
xor ( n61822 , n51987 , n52014 );
xor ( n589146 , n61822 , n589134 );
xor ( n589147 , n52017 , n52058 );
xor ( n61825 , n589147 , n589131 );
xor ( n61826 , n52061 , n52111 );
xor ( n589150 , n61826 , n61805 );
xor ( n589151 , n52114 , n52190 );
xor ( n61829 , n589151 , n589125 );
xor ( n61830 , n52193 , n52247 );
xor ( n589154 , n61830 , n589122 );
xor ( n589155 , n52250 , n52300 );
xor ( n61833 , n589155 , n589119 );
xor ( n589157 , n52303 , n52359 );
xor ( n61835 , n589157 , n61793 );
xor ( n589159 , n52362 , n52477 );
xor ( n61837 , n589159 , n589113 );
xor ( n589161 , n52570 , n52572 );
xor ( n61839 , n589161 , n61787 );
xor ( n61840 , n52575 , n52665 );
xor ( n589164 , n61840 , n589107 );
xor ( n589165 , n52668 , n52768 );
xor ( n61843 , n589165 , n61781 );
xor ( n61844 , n52771 , n52880 );
xor ( n589168 , n61844 , n61778 );
xor ( n589169 , n52883 , n53006 );
xor ( n61847 , n589169 , n61775 );
xor ( n61848 , n53009 , n53103 );
xor ( n589172 , n61848 , n589095 );
xor ( n589173 , n53106 , n53208 );
xor ( n61851 , n589173 , n589092 );
xor ( n61852 , n53211 , n53354 );
xor ( n589176 , n61852 , n61766 );
xor ( n589177 , n53496 , n53498 );
xor ( n589178 , n589177 , n589086 );
xor ( n61856 , n53633 , n53635 );
xor ( n589180 , n61856 , n589083 );
xor ( n589181 , n53638 , n53742 );
xor ( n61859 , n589181 , n61757 );
xor ( n589183 , n53745 , n53975 );
xor ( n589184 , n589183 , n589077 );
xor ( n61862 , n53978 , n54146 );
xor ( n61863 , n61862 , n61751 );
xor ( n589187 , n54149 , n54294 );
xor ( n589188 , n589187 , n589071 );
xor ( n61866 , n54297 , n54469 );
xor ( n61867 , n61866 , n589068 );
xor ( n589191 , n54644 , n54646 );
xor ( n589192 , n589191 , n589065 );
xor ( n61870 , n54649 , n54826 );
xor ( n589194 , n61870 , n589062 );
xor ( n589195 , n55004 , n55006 );
xor ( n61873 , n589195 , n589059 );
xor ( n589197 , n55009 , n55184 );
xor ( n589198 , n589197 , n61733 );
xor ( n589199 , n55187 , n55416 );
xor ( n589200 , n589199 , n589053 );
xor ( n61878 , n55419 , n582790 );
xor ( n589202 , n61878 , n589050 );
xor ( n589203 , n55470 , n55625 );
xor ( n61881 , n589203 , n589047 );
xor ( n589205 , n55628 , n583151 );
xor ( n589206 , n589205 , n589044 );
xor ( n61884 , n55831 , n56020 );
xor ( n61885 , n61884 , n61718 );
xor ( n589209 , n56023 , n583364 );
xor ( n61887 , n589209 , n589038 );
xor ( n61888 , n583367 , n56241 );
xor ( n589212 , n61888 , n589035 );
xor ( n589213 , n56244 , n583724 );
xor ( n61891 , n589213 , n589032 );
xor ( n589215 , n583727 , n583949 );
xor ( n589216 , n589215 , n589029 );
xor ( n61894 , n583952 , n56788 );
xor ( n589218 , n61894 , n61703 );
xor ( n589219 , n56791 , n57031 );
xor ( n61897 , n589219 , n589023 );
xor ( n61898 , n57034 , n57193 );
xor ( n61899 , n61898 , n589020 );
xor ( n589223 , n57196 , n584743 );
xor ( n589224 , n589223 , n589017 );
xor ( n61902 , n57423 , n57469 );
xor ( n61903 , n61902 , n61691 );
xor ( n61904 , n57472 , n57696 );
xor ( n589228 , n61904 , n61688 );
xor ( n589229 , n585022 , n585199 );
xor ( n61907 , n589229 , n61685 );
xor ( n61908 , n57879 , n58119 );
xor ( n589232 , n61908 , n61682 );
xor ( n589233 , n58122 , n58170 );
xor ( n61911 , n589233 , n61679 );
xor ( n61912 , n58173 , n585709 );
xor ( n589236 , n61912 , n61676 );
xor ( n61914 , n58389 , n585896 );
xor ( n61915 , n61914 , n588996 );
xor ( n61916 , n58576 , n586152 );
xor ( n61917 , n61916 , n61670 );
xor ( n589241 , n586155 , n586331 );
xor ( n61919 , n589241 , n588990 );
xor ( n61920 , n59011 , n586372 );
xor ( n61921 , n61920 , n588987 );
xor ( n61922 , n59052 , n586619 );
xor ( n589246 , n61922 , n588984 );
xor ( n589247 , n59465 , n586790 );
xor ( n589248 , n589247 , n61658 );
xor ( n61926 , n586793 , n586955 );
xor ( n589250 , n61926 , n588978 );
xor ( n589251 , n59635 , n59857 );
xor ( n589252 , n589251 , n588975 );
xor ( n589253 , n59860 , n59952 );
xor ( n61931 , n589253 , n588972 );
xor ( n589255 , n587278 , n60222 );
xor ( n589256 , n589255 , n61646 );
xor ( n61934 , n60225 , n60371 );
xor ( n589258 , n61934 , n588966 );
xor ( n61936 , n60374 , n587811 );
xor ( n589260 , n61936 , n61640 );
xor ( n61938 , n60678 , n60680 );
xor ( n61939 , n61938 , n588960 );
xor ( n589263 , n60683 , n588090 );
xor ( n589264 , n589263 , n61634 );
xor ( n61942 , n61017 , n588342 );
xor ( n589266 , n61942 , n61631 );
xor ( n589267 , n588345 , n588407 );
xor ( n61945 , n589267 , n588951 );
xor ( n589269 , n61087 , n61161 );
xor ( n589270 , n589269 , n588948 );
xor ( n61948 , n61177 , n588502 );
xor ( n589272 , n61948 , n588945 );
xor ( n589273 , n588836 , n61515 );
xor ( n589274 , n588846 , n588848 );
and ( n589275 , n589273 , n589274 );
xor ( n61953 , n61528 , n61535 );
xor ( n589277 , n61953 , n588931 );
and ( n589278 , n589274 , n589277 );
and ( n589279 , n589273 , n589277 );
or ( n589280 , n589275 , n589278 , n589279 );
xor ( n61958 , n588829 , n588831 );
xor ( n589282 , n61958 , n588839 );
and ( n589283 , n589280 , n589282 );
xor ( n61961 , n61526 , n588934 );
xor ( n589285 , n61961 , n61613 );
and ( n589286 , n589282 , n589285 );
and ( n61964 , n589280 , n589285 );
or ( n589288 , n589283 , n589286 , n61964 );
xor ( n589289 , n61519 , n588939 );
xor ( n61967 , n589289 , n61619 );
and ( n61968 , n589288 , n61967 );
xor ( n61969 , n589288 , n61967 );
xor ( n589293 , n589280 , n589282 );
xor ( n589294 , n589293 , n589285 );
xor ( n61972 , n589273 , n589274 );
xor ( n589296 , n61972 , n589277 );
xor ( n61974 , n61532 , n588857 );
xor ( n589298 , n61538 , n588863 );
xor ( n61976 , n589298 , n588928 );
and ( n61977 , n61974 , n61976 );
xor ( n589301 , n61974 , n61976 );
xor ( n589302 , n588734 , n588736 );
xor ( n61980 , n589302 , n61494 );
xor ( n61981 , n61386 , n61402 );
xor ( n589305 , n61981 , n61405 );
xor ( n589306 , n61390 , n61394 );
xor ( n61984 , n589306 , n61399 );
and ( n589308 , n583377 , n55013 );
and ( n61986 , n55841 , n55010 );
nor ( n61987 , n589308 , n61986 );
xnor ( n589311 , n61987 , n53762 );
and ( n589312 , n583746 , n54532 );
and ( n61990 , n56282 , n54530 );
nor ( n61991 , n589312 , n61990 );
xnor ( n589315 , n61991 , n53769 );
and ( n589316 , n589311 , n589315 );
and ( n61994 , n56671 , n54414 );
and ( n61995 , n583800 , n54412 );
nor ( n61996 , n61994 , n61995 );
xnor ( n589320 , n61996 , n53650 );
and ( n589321 , n589315 , n589320 );
and ( n61999 , n589311 , n589320 );
or ( n589323 , n589316 , n589321 , n61999 );
and ( n589324 , n56909 , n53996 );
and ( n62002 , n56832 , n53994 );
nor ( n589326 , n589324 , n62002 );
xnor ( n589327 , n589326 , n53376 );
and ( n62005 , n584529 , n53683 );
and ( n589329 , n57058 , n53681 );
nor ( n589330 , n62005 , n589329 );
xnor ( n62008 , n589330 , n53118 );
and ( n589332 , n589327 , n62008 );
and ( n589333 , n57484 , n53468 );
and ( n62011 , n57283 , n53466 );
nor ( n589335 , n589333 , n62011 );
xnor ( n589336 , n589335 , n52945 );
and ( n62014 , n62008 , n589336 );
and ( n589338 , n589327 , n589336 );
or ( n589339 , n589332 , n62014 , n589338 );
and ( n62017 , n589323 , n589339 );
and ( n589341 , n585062 , n53177 );
and ( n62019 , n57482 , n53175 );
nor ( n589343 , n589341 , n62019 );
xnor ( n62021 , n589343 , n52827 );
and ( n589345 , n585221 , n52978 );
and ( n589346 , n57900 , n52976 );
nor ( n62024 , n589345 , n589346 );
xnor ( n62025 , n62024 , n52680 );
and ( n589349 , n62021 , n62025 );
and ( n62027 , n58246 , n52707 );
and ( n589351 , n58219 , n52705 );
nor ( n62029 , n62027 , n589351 );
xnor ( n589353 , n62029 , n52526 );
and ( n589354 , n62025 , n589353 );
and ( n62032 , n62021 , n589353 );
or ( n589356 , n589349 , n589354 , n62032 );
and ( n589357 , n589339 , n589356 );
and ( n62035 , n589323 , n589356 );
or ( n62036 , n62017 , n589357 , n62035 );
and ( n589360 , n61984 , n62036 );
xor ( n62038 , n61429 , n61433 );
xor ( n589362 , n62038 , n588761 );
xor ( n62040 , n61448 , n61452 );
xor ( n589364 , n62040 , n61457 );
and ( n589365 , n589362 , n589364 );
xor ( n62043 , n588787 , n588791 );
xor ( n589367 , n62043 , n588796 );
and ( n589368 , n589364 , n589367 );
and ( n62046 , n589362 , n589367 );
or ( n589370 , n589365 , n589368 , n62046 );
and ( n589371 , n62036 , n589370 );
and ( n62049 , n61984 , n589370 );
or ( n62050 , n589360 , n589371 , n62049 );
and ( n589374 , n589305 , n62050 );
xor ( n589375 , n61444 , n61482 );
xor ( n62053 , n589375 , n61485 );
and ( n589377 , n62050 , n62053 );
and ( n589378 , n589305 , n62053 );
or ( n62056 , n589374 , n589377 , n589378 );
xor ( n589380 , n588739 , n61488 );
xor ( n589381 , n589380 , n588814 );
and ( n62059 , n62056 , n589381 );
xor ( n62060 , n61420 , n61424 );
xor ( n589384 , n62060 , n61441 );
xor ( n62062 , n61460 , n61476 );
xor ( n62063 , n62062 , n61479 );
and ( n589387 , n589384 , n62063 );
and ( n589388 , n583800 , n54532 );
and ( n589389 , n583746 , n54530 );
nor ( n62067 , n589388 , n589389 );
xnor ( n589391 , n62067 , n53769 );
and ( n589392 , n56832 , n54414 );
and ( n62070 , n56671 , n54412 );
nor ( n62071 , n589392 , n62070 );
xnor ( n589395 , n62071 , n53650 );
and ( n589396 , n589391 , n589395 );
and ( n62074 , n56282 , n55013 );
and ( n589398 , n583377 , n55010 );
nor ( n589399 , n62074 , n589398 );
xnor ( n62077 , n589399 , n53762 );
and ( n589401 , n57058 , n53996 );
and ( n589402 , n56909 , n53994 );
nor ( n62080 , n589401 , n589402 );
xnor ( n589404 , n62080 , n53376 );
and ( n589405 , n62077 , n589404 );
and ( n62083 , n57283 , n53683 );
and ( n62084 , n584529 , n53681 );
nor ( n589408 , n62083 , n62084 );
xnor ( n589409 , n589408 , n53118 );
and ( n62087 , n589404 , n589409 );
and ( n589411 , n62077 , n589409 );
or ( n589412 , n589405 , n62087 , n589411 );
and ( n62090 , n589396 , n589412 );
and ( n589414 , n57482 , n53468 );
and ( n589415 , n57484 , n53466 );
nor ( n62093 , n589414 , n589415 );
xnor ( n62094 , n62093 , n52945 );
and ( n589418 , n57900 , n53177 );
and ( n589419 , n585062 , n53175 );
nor ( n589420 , n589418 , n589419 );
xnor ( n589421 , n589420 , n52827 );
and ( n589422 , n62094 , n589421 );
and ( n62100 , n58219 , n52978 );
and ( n589424 , n585221 , n52976 );
nor ( n589425 , n62100 , n589424 );
xnor ( n62103 , n589425 , n52680 );
and ( n62104 , n589421 , n62103 );
and ( n589428 , n62094 , n62103 );
or ( n62106 , n589422 , n62104 , n589428 );
and ( n589430 , n589412 , n62106 );
and ( n589431 , n589396 , n62106 );
or ( n62109 , n62090 , n589430 , n589431 );
xor ( n62110 , n589311 , n589315 );
xor ( n589434 , n62110 , n589320 );
xor ( n589435 , n589327 , n62008 );
xor ( n62113 , n589435 , n589336 );
and ( n62114 , n589434 , n62113 );
xor ( n589438 , n62021 , n62025 );
xor ( n62116 , n589438 , n589353 );
and ( n62117 , n62113 , n62116 );
and ( n62118 , n589434 , n62116 );
or ( n62119 , n62114 , n62117 , n62118 );
and ( n589443 , n62109 , n62119 );
xor ( n589444 , n589323 , n589339 );
xor ( n589445 , n589444 , n589356 );
and ( n62123 , n62119 , n589445 );
and ( n589447 , n62109 , n589445 );
or ( n589448 , n589443 , n62123 , n589447 );
and ( n589449 , n62063 , n589448 );
and ( n62127 , n589384 , n589448 );
or ( n589451 , n589387 , n589449 , n62127 );
xor ( n62129 , n589305 , n62050 );
xor ( n589453 , n62129 , n62053 );
and ( n589454 , n589451 , n589453 );
xor ( n62132 , n61984 , n62036 );
xor ( n589456 , n62132 , n589370 );
xor ( n62134 , n589362 , n589364 );
xor ( n62135 , n62134 , n589367 );
and ( n62136 , n585586 , n52707 );
and ( n62137 , n58246 , n52705 );
nor ( n62138 , n62136 , n62137 );
xnor ( n62139 , n62138 , n52526 );
and ( n62140 , n58623 , n52509 );
and ( n62141 , n585909 , n52507 );
nor ( n62142 , n62140 , n62141 );
xnor ( n62143 , n62142 , n52383 );
and ( n589467 , n62139 , n62143 );
xor ( n62145 , n589391 , n589395 );
and ( n589469 , n62143 , n62145 );
and ( n589470 , n62139 , n62145 );
or ( n62148 , n589467 , n589469 , n589470 );
and ( n589472 , n583746 , n55013 );
and ( n589473 , n56282 , n55010 );
nor ( n62151 , n589472 , n589473 );
xnor ( n62152 , n62151 , n53762 );
and ( n589476 , n56671 , n54532 );
and ( n589477 , n583800 , n54530 );
nor ( n62155 , n589476 , n589477 );
xnor ( n62156 , n62155 , n53769 );
and ( n589480 , n62152 , n62156 );
and ( n589481 , n56909 , n54414 );
and ( n62159 , n56832 , n54412 );
nor ( n62160 , n589481 , n62159 );
xnor ( n589484 , n62160 , n53650 );
and ( n62162 , n62156 , n589484 );
and ( n62163 , n62152 , n589484 );
or ( n589487 , n589480 , n62162 , n62163 );
and ( n589488 , n584529 , n53996 );
and ( n62166 , n57058 , n53994 );
nor ( n62167 , n589488 , n62166 );
xnor ( n589491 , n62167 , n53376 );
and ( n62169 , n57484 , n53683 );
and ( n62170 , n57283 , n53681 );
nor ( n62171 , n62169 , n62170 );
xnor ( n62172 , n62171 , n53118 );
and ( n62173 , n589491 , n62172 );
and ( n62174 , n585062 , n53468 );
and ( n589498 , n57482 , n53466 );
nor ( n62176 , n62174 , n589498 );
xnor ( n62177 , n62176 , n52945 );
and ( n62178 , n62172 , n62177 );
and ( n589502 , n589491 , n62177 );
or ( n62180 , n62173 , n62178 , n589502 );
and ( n62181 , n589487 , n62180 );
and ( n62182 , n585221 , n53177 );
and ( n62183 , n57900 , n53175 );
nor ( n62184 , n62182 , n62183 );
xnor ( n62185 , n62184 , n52827 );
and ( n589509 , n58246 , n52978 );
and ( n62187 , n58219 , n52976 );
nor ( n62188 , n589509 , n62187 );
xnor ( n62189 , n62188 , n52680 );
and ( n62190 , n62185 , n62189 );
and ( n62191 , n585909 , n52707 );
and ( n589515 , n585586 , n52705 );
nor ( n62193 , n62191 , n589515 );
xnor ( n62194 , n62193 , n52526 );
and ( n589518 , n62189 , n62194 );
and ( n589519 , n62185 , n62194 );
or ( n62197 , n62190 , n589518 , n589519 );
and ( n62198 , n62180 , n62197 );
and ( n589522 , n589487 , n62197 );
or ( n589523 , n62181 , n62198 , n589522 );
and ( n62201 , n62148 , n589523 );
and ( n589525 , n585973 , n52509 );
and ( n589526 , n58623 , n52507 );
nor ( n62204 , n589525 , n589526 );
xnor ( n589528 , n62204 , n52383 );
nor ( n589529 , n52065 , n52063 );
xnor ( n62207 , n589529 , n52022 );
and ( n589531 , n589528 , n62207 );
and ( n589532 , n52064 , n52022 );
and ( n589533 , n62207 , n589532 );
and ( n589534 , n589528 , n589532 );
or ( n62212 , n589531 , n589533 , n589534 );
xor ( n589536 , n62077 , n589404 );
xor ( n589537 , n589536 , n589409 );
and ( n62215 , n62212 , n589537 );
xor ( n589539 , n62094 , n589421 );
xor ( n62217 , n589539 , n62103 );
and ( n589541 , n589537 , n62217 );
and ( n62219 , n62212 , n62217 );
or ( n62220 , n62215 , n589541 , n62219 );
and ( n589544 , n589523 , n62220 );
and ( n589545 , n62148 , n62220 );
or ( n62223 , n62201 , n589544 , n589545 );
and ( n589547 , n62135 , n62223 );
xor ( n589548 , n62109 , n62119 );
xor ( n62226 , n589548 , n589445 );
and ( n589550 , n62223 , n62226 );
and ( n589551 , n62135 , n62226 );
or ( n62229 , n589547 , n589550 , n589551 );
and ( n589553 , n589456 , n62229 );
xor ( n589554 , n589384 , n62063 );
xor ( n589555 , n589554 , n589448 );
and ( n589556 , n62229 , n589555 );
and ( n62234 , n589456 , n589555 );
or ( n589558 , n589553 , n589556 , n62234 );
and ( n589559 , n589453 , n589558 );
and ( n62237 , n589451 , n589558 );
or ( n62238 , n589454 , n589559 , n62237 );
and ( n589562 , n589381 , n62238 );
and ( n62240 , n62056 , n62238 );
or ( n62241 , n62059 , n589562 , n62240 );
and ( n62242 , n61980 , n62241 );
xor ( n589566 , n62056 , n589381 );
xor ( n589567 , n589566 , n62238 );
xor ( n62245 , n61589 , n588916 );
xor ( n62246 , n62245 , n61596 );
and ( n62247 , n589567 , n62246 );
xor ( n589571 , n589451 , n589453 );
xor ( n589572 , n589571 , n589558 );
xor ( n589573 , n589456 , n62229 );
xor ( n589574 , n589573 , n589555 );
xor ( n62252 , n588892 , n588896 );
xor ( n589576 , n62252 , n588899 );
and ( n62254 , n589574 , n589576 );
xor ( n62255 , n588871 , n61550 );
nor ( n589579 , n52432 , n52430 );
xnor ( n589580 , n589579 , n52255 );
nor ( n62258 , n52273 , n52271 );
xnor ( n62259 , n62258 , n52137 );
and ( n589583 , n589580 , n62259 );
nor ( n589584 , n52155 , n52153 );
xnor ( n62262 , n589584 , n52085 );
and ( n62263 , n62259 , n62262 );
and ( n589587 , n589580 , n62262 );
or ( n62265 , n589583 , n62263 , n589587 );
and ( n589589 , n62255 , n62265 );
xor ( n589590 , n588204 , n588206 );
xor ( n62268 , n589590 , n51989 );
and ( n62269 , n62265 , n62268 );
and ( n589593 , n62255 , n62268 );
or ( n62271 , n589589 , n62269 , n589593 );
and ( n589595 , n585909 , n52509 );
and ( n62273 , n585586 , n52507 );
nor ( n589597 , n589595 , n62273 );
xnor ( n589598 , n589597 , n52383 );
and ( n62276 , n62271 , n589598 );
xor ( n589600 , n588874 , n61553 );
xor ( n589601 , n589600 , n588879 );
and ( n62279 , n589598 , n589601 );
and ( n62280 , n62271 , n589601 );
or ( n589604 , n62276 , n62279 , n62280 );
xor ( n589605 , n61559 , n588886 );
xor ( n62283 , n589605 , n61566 );
and ( n62284 , n589604 , n62283 );
and ( n589608 , n589576 , n62284 );
and ( n589609 , n589574 , n62284 );
or ( n62287 , n62254 , n589608 , n589609 );
and ( n62288 , n589572 , n62287 );
xor ( n62289 , n61579 , n588906 );
xor ( n589613 , n62289 , n61586 );
and ( n589614 , n62287 , n589613 );
and ( n62292 , n589572 , n589613 );
or ( n589616 , n62288 , n589614 , n62292 );
and ( n62294 , n62246 , n589616 );
and ( n62295 , n589567 , n589616 );
or ( n589619 , n62247 , n62294 , n62295 );
and ( n62297 , n62241 , n589619 );
and ( n589621 , n61980 , n589619 );
or ( n62299 , n62242 , n62297 , n589621 );
xor ( n589623 , n61543 , n588868 );
xor ( n62301 , n589623 , n588925 );
and ( n62302 , n62299 , n62301 );
xor ( n62303 , n62299 , n62301 );
xor ( n62304 , n61599 , n588924 );
xor ( n62305 , n61980 , n62241 );
xor ( n62306 , n62305 , n589619 );
and ( n62307 , n62304 , n62306 );
xor ( n62308 , n62304 , n62306 );
xor ( n589632 , n589567 , n62246 );
xor ( n62310 , n589632 , n589616 );
xor ( n589634 , n589396 , n589412 );
xor ( n62312 , n589634 , n62106 );
xor ( n62313 , n589434 , n62113 );
xor ( n589637 , n62313 , n62116 );
and ( n62315 , n62312 , n589637 );
xor ( n62316 , n62255 , n62265 );
xor ( n589640 , n62316 , n62268 );
xor ( n62318 , n589580 , n62259 );
xor ( n62319 , n62318 , n62262 );
nor ( n589643 , n52432 , n52430 );
xnor ( n62321 , n589643 , n52255 );
nor ( n62322 , n52273 , n52271 );
xnor ( n589646 , n62322 , n52137 );
and ( n62324 , n62321 , n589646 );
and ( n62325 , n589646 , n52063 );
and ( n62326 , n62321 , n52063 );
or ( n62327 , n62324 , n62325 , n62326 );
and ( n589651 , n62319 , n62327 );
and ( n62329 , n585973 , n52507 );
nor ( n62330 , n52509 , n62329 );
xnor ( n589654 , n62330 , n52383 );
nor ( n589655 , n52155 , n52153 );
xnor ( n62333 , n589655 , n52085 );
and ( n589657 , n589654 , n62333 );
and ( n589658 , n62327 , n589657 );
and ( n62336 , n62319 , n589657 );
or ( n62337 , n589651 , n589658 , n62336 );
and ( n589661 , n589640 , n62337 );
and ( n62339 , n583800 , n55013 );
and ( n62340 , n583746 , n55010 );
nor ( n62341 , n62339 , n62340 );
xnor ( n62342 , n62341 , n53762 );
and ( n62343 , n56832 , n54532 );
and ( n62344 , n56671 , n54530 );
nor ( n589668 , n62343 , n62344 );
xnor ( n62346 , n589668 , n53769 );
and ( n62347 , n62342 , n62346 );
and ( n589671 , n57058 , n54414 );
and ( n62349 , n56909 , n54412 );
nor ( n62350 , n589671 , n62349 );
xnor ( n62351 , n62350 , n53650 );
and ( n62352 , n57283 , n53996 );
and ( n589676 , n584529 , n53994 );
nor ( n589677 , n62352 , n589676 );
xnor ( n62355 , n589677 , n53376 );
and ( n589679 , n62351 , n62355 );
and ( n62357 , n57482 , n53683 );
and ( n62358 , n57484 , n53681 );
nor ( n62359 , n62357 , n62358 );
xnor ( n589683 , n62359 , n53118 );
and ( n589684 , n62355 , n589683 );
and ( n589685 , n62351 , n589683 );
or ( n62363 , n589679 , n589684 , n589685 );
and ( n589687 , n62347 , n62363 );
and ( n589688 , n57900 , n53468 );
and ( n62366 , n585062 , n53466 );
nor ( n62367 , n589688 , n62366 );
xnor ( n589691 , n62367 , n52945 );
and ( n589692 , n58219 , n53177 );
and ( n589693 , n585221 , n53175 );
nor ( n62371 , n589692 , n589693 );
xnor ( n589695 , n62371 , n52827 );
and ( n589696 , n589691 , n589695 );
and ( n589697 , n585586 , n52978 );
and ( n589698 , n58246 , n52976 );
nor ( n62376 , n589697 , n589698 );
xnor ( n589700 , n62376 , n52680 );
and ( n589701 , n589695 , n589700 );
and ( n62379 , n589691 , n589700 );
or ( n589703 , n589696 , n589701 , n62379 );
and ( n589704 , n62363 , n589703 );
and ( n62382 , n62347 , n589703 );
or ( n589706 , n589687 , n589704 , n62382 );
and ( n589707 , n62337 , n589706 );
and ( n62385 , n589640 , n589706 );
or ( n589709 , n589661 , n589707 , n62385 );
and ( n589710 , n589637 , n589709 );
and ( n62388 , n62312 , n589709 );
or ( n589712 , n62315 , n589710 , n62388 );
xor ( n589713 , n62135 , n62223 );
xor ( n62391 , n589713 , n62226 );
and ( n589715 , n589712 , n62391 );
xor ( n589716 , n62152 , n62156 );
xor ( n62394 , n589716 , n589484 );
xor ( n589718 , n589491 , n62172 );
xor ( n589719 , n589718 , n62177 );
and ( n62397 , n62394 , n589719 );
xor ( n589721 , n62185 , n62189 );
xor ( n589722 , n589721 , n62194 );
and ( n589723 , n589719 , n589722 );
and ( n589724 , n62394 , n589722 );
or ( n62402 , n62397 , n589723 , n589724 );
xor ( n589726 , n62139 , n62143 );
xor ( n589727 , n589726 , n62145 );
and ( n62405 , n62402 , n589727 );
xor ( n589729 , n589487 , n62180 );
xor ( n589730 , n589729 , n62197 );
and ( n62408 , n589727 , n589730 );
and ( n62409 , n62402 , n589730 );
or ( n589733 , n62405 , n62408 , n62409 );
xor ( n589734 , n62148 , n589523 );
xor ( n62412 , n589734 , n62220 );
and ( n62413 , n589733 , n62412 );
xor ( n589737 , n62271 , n589598 );
xor ( n589738 , n589737 , n589601 );
and ( n62416 , n62412 , n589738 );
and ( n62417 , n589733 , n589738 );
or ( n589741 , n62413 , n62416 , n62417 );
and ( n589742 , n62391 , n589741 );
and ( n62420 , n589712 , n589741 );
or ( n62421 , n589715 , n589742 , n62420 );
xor ( n589745 , n589604 , n62283 );
xor ( n589746 , n62212 , n589537 );
xor ( n62424 , n589746 , n62217 );
xor ( n589748 , n589528 , n62207 );
xor ( n589749 , n589748 , n589532 );
and ( n62427 , n58623 , n52707 );
and ( n62428 , n585909 , n52705 );
nor ( n62429 , n62427 , n62428 );
xnor ( n62430 , n62429 , n52526 );
xor ( n62431 , n62321 , n589646 );
xor ( n589755 , n62431 , n52063 );
and ( n62433 , n62430 , n589755 );
xor ( n589757 , n589654 , n62333 );
and ( n589758 , n589755 , n589757 );
and ( n62436 , n62430 , n589757 );
or ( n62437 , n62433 , n589758 , n62436 );
and ( n589761 , n589749 , n62437 );
xor ( n589762 , n62342 , n62346 );
nor ( n62440 , n52509 , n52507 );
xnor ( n589764 , n62440 , n52383 );
nor ( n589765 , n52432 , n52430 );
xnor ( n62443 , n589765 , n52255 );
and ( n589767 , n589764 , n62443 );
nor ( n62445 , n52273 , n52271 );
xnor ( n62446 , n62445 , n52137 );
and ( n62447 , n62443 , n62446 );
and ( n62448 , n589764 , n62446 );
or ( n62449 , n589767 , n62447 , n62448 );
and ( n62450 , n589762 , n62449 );
and ( n62451 , n56671 , n55013 );
and ( n62452 , n583800 , n55010 );
nor ( n589776 , n62451 , n62452 );
xnor ( n589777 , n589776 , n53762 );
and ( n62455 , n56909 , n54532 );
and ( n589779 , n56832 , n54530 );
nor ( n62457 , n62455 , n589779 );
xnor ( n62458 , n62457 , n53769 );
and ( n62459 , n589777 , n62458 );
and ( n62460 , n584529 , n54414 );
and ( n62461 , n57058 , n54412 );
nor ( n62462 , n62460 , n62461 );
xnor ( n62463 , n62462 , n53650 );
and ( n62464 , n62458 , n62463 );
and ( n62465 , n589777 , n62463 );
or ( n62466 , n62459 , n62464 , n62465 );
and ( n62467 , n62449 , n62466 );
and ( n62468 , n589762 , n62466 );
or ( n62469 , n62450 , n62467 , n62468 );
and ( n62470 , n62437 , n62469 );
and ( n589794 , n589749 , n62469 );
or ( n62472 , n589761 , n62470 , n589794 );
and ( n62473 , n62424 , n62472 );
and ( n62474 , n57484 , n53996 );
and ( n62475 , n57283 , n53994 );
nor ( n589799 , n62474 , n62475 );
xnor ( n62477 , n589799 , n53376 );
and ( n589801 , n585062 , n53683 );
and ( n589802 , n57482 , n53681 );
nor ( n62480 , n589801 , n589802 );
xnor ( n589804 , n62480 , n53118 );
and ( n589805 , n62477 , n589804 );
and ( n589806 , n585221 , n53468 );
and ( n589807 , n57900 , n53466 );
nor ( n62485 , n589806 , n589807 );
xnor ( n589809 , n62485 , n52945 );
and ( n589810 , n589804 , n589809 );
and ( n62488 , n62477 , n589809 );
or ( n589812 , n589805 , n589810 , n62488 );
and ( n589813 , n58246 , n53177 );
and ( n62491 , n58219 , n53175 );
nor ( n589815 , n589813 , n62491 );
xnor ( n589816 , n589815 , n52827 );
and ( n62494 , n585909 , n52978 );
and ( n589818 , n585586 , n52976 );
nor ( n62496 , n62494 , n589818 );
xnor ( n589820 , n62496 , n52680 );
and ( n62498 , n589816 , n589820 );
and ( n589822 , n585973 , n52707 );
and ( n62500 , n58623 , n52705 );
nor ( n62501 , n589822 , n62500 );
xnor ( n589825 , n62501 , n52526 );
and ( n589826 , n589820 , n589825 );
and ( n62504 , n589816 , n589825 );
or ( n589828 , n62498 , n589826 , n62504 );
and ( n62506 , n589812 , n589828 );
xor ( n589830 , n62351 , n62355 );
xor ( n589831 , n589830 , n589683 );
and ( n62509 , n589828 , n589831 );
and ( n589833 , n589812 , n589831 );
or ( n62511 , n62506 , n62509 , n589833 );
xor ( n62512 , n62319 , n62327 );
xor ( n62513 , n62512 , n589657 );
and ( n62514 , n62511 , n62513 );
xor ( n62515 , n62347 , n62363 );
xor ( n62516 , n62515 , n589703 );
and ( n589840 , n62513 , n62516 );
and ( n62518 , n62511 , n62516 );
or ( n62519 , n62514 , n589840 , n62518 );
and ( n589843 , n62472 , n62519 );
and ( n62521 , n62424 , n62519 );
or ( n589845 , n62473 , n589843 , n62521 );
xor ( n62523 , n62312 , n589637 );
xor ( n62524 , n62523 , n589709 );
and ( n589848 , n589845 , n62524 );
xor ( n589849 , n589640 , n62337 );
xor ( n62527 , n589849 , n589706 );
xor ( n589851 , n62402 , n589727 );
xor ( n62529 , n589851 , n589730 );
and ( n62530 , n62527 , n62529 );
xor ( n62531 , n62394 , n589719 );
xor ( n62532 , n62531 , n589722 );
xor ( n62533 , n589691 , n589695 );
xor ( n62534 , n62533 , n589700 );
nor ( n62535 , n52155 , n52153 );
xnor ( n62536 , n62535 , n52085 );
and ( n62537 , n52154 , n52085 );
and ( n62538 , n62536 , n62537 );
xor ( n62539 , n589764 , n62443 );
xor ( n62540 , n62539 , n62446 );
and ( n62541 , n62537 , n62540 );
and ( n62542 , n62536 , n62540 );
or ( n62543 , n62538 , n62541 , n62542 );
and ( n62544 , n62534 , n62543 );
nor ( n62545 , n52509 , n52507 );
xnor ( n62546 , n62545 , n52383 );
nor ( n62547 , n52432 , n52430 );
xnor ( n589871 , n62547 , n52255 );
and ( n62549 , n62546 , n589871 );
nor ( n62550 , n52273 , n52271 );
xnor ( n589874 , n62550 , n52137 );
and ( n589875 , n589871 , n589874 );
and ( n62553 , n62546 , n589874 );
or ( n589877 , n62549 , n589875 , n62553 );
and ( n62555 , n585973 , n52705 );
nor ( n589879 , n52707 , n62555 );
xnor ( n589880 , n589879 , n52526 );
and ( n62558 , n589880 , n52153 );
and ( n589882 , n589877 , n62558 );
and ( n589883 , n56832 , n55013 );
and ( n589884 , n56671 , n55010 );
nor ( n62562 , n589883 , n589884 );
xnor ( n589886 , n62562 , n53762 );
and ( n589887 , n57058 , n54532 );
and ( n62565 , n56909 , n54530 );
nor ( n589889 , n589887 , n62565 );
xnor ( n62567 , n589889 , n53769 );
and ( n62568 , n589886 , n62567 );
and ( n589892 , n57283 , n54414 );
and ( n589893 , n584529 , n54412 );
nor ( n62571 , n589892 , n589893 );
xnor ( n589895 , n62571 , n53650 );
and ( n589896 , n62567 , n589895 );
and ( n62574 , n589886 , n589895 );
or ( n589898 , n62568 , n589896 , n62574 );
and ( n62576 , n62558 , n589898 );
and ( n62577 , n589877 , n589898 );
or ( n62578 , n589882 , n62576 , n62577 );
and ( n62579 , n62543 , n62578 );
and ( n62580 , n62534 , n62578 );
or ( n589904 , n62544 , n62579 , n62580 );
and ( n589905 , n62532 , n589904 );
and ( n62583 , n57482 , n53996 );
and ( n589907 , n57484 , n53994 );
nor ( n62585 , n62583 , n589907 );
xnor ( n589909 , n62585 , n53376 );
and ( n62587 , n57900 , n53683 );
and ( n62588 , n585062 , n53681 );
nor ( n589912 , n62587 , n62588 );
xnor ( n62590 , n589912 , n53118 );
and ( n589914 , n589909 , n62590 );
and ( n589915 , n58219 , n53468 );
and ( n62593 , n585221 , n53466 );
nor ( n589917 , n589915 , n62593 );
xnor ( n62595 , n589917 , n52945 );
and ( n62596 , n62590 , n62595 );
and ( n62597 , n589909 , n62595 );
or ( n62598 , n589914 , n62596 , n62597 );
xor ( n589922 , n589777 , n62458 );
xor ( n62600 , n589922 , n62463 );
and ( n62601 , n62598 , n62600 );
xor ( n589925 , n62477 , n589804 );
xor ( n589926 , n589925 , n589809 );
and ( n62604 , n62600 , n589926 );
and ( n589928 , n62598 , n589926 );
or ( n62606 , n62601 , n62604 , n589928 );
xor ( n62607 , n62430 , n589755 );
xor ( n589931 , n62607 , n589757 );
and ( n62609 , n62606 , n589931 );
xor ( n589933 , n589762 , n62449 );
xor ( n62611 , n589933 , n62466 );
and ( n589935 , n589931 , n62611 );
and ( n589936 , n62606 , n62611 );
or ( n62614 , n62609 , n589935 , n589936 );
and ( n589938 , n589904 , n62614 );
and ( n62616 , n62532 , n62614 );
or ( n62617 , n589905 , n589938 , n62616 );
and ( n589941 , n62529 , n62617 );
and ( n62619 , n62527 , n62617 );
or ( n589943 , n62530 , n589941 , n62619 );
and ( n62621 , n62524 , n589943 );
and ( n589945 , n589845 , n589943 );
or ( n589946 , n589848 , n62621 , n589945 );
and ( n62624 , n589745 , n589946 );
xor ( n589948 , n589712 , n62391 );
xor ( n62626 , n589948 , n589741 );
and ( n62627 , n589946 , n62626 );
and ( n62628 , n589745 , n62626 );
or ( n62629 , n62624 , n62627 , n62628 );
and ( n62630 , n62421 , n62629 );
xor ( n589954 , n589574 , n589576 );
xor ( n62632 , n589954 , n62284 );
and ( n589956 , n62629 , n62632 );
and ( n62634 , n62421 , n62632 );
or ( n589958 , n62630 , n589956 , n62634 );
xor ( n62636 , n589572 , n62287 );
xor ( n62637 , n62636 , n589613 );
and ( n62638 , n589958 , n62637 );
xor ( n62639 , n589958 , n62637 );
xor ( n62640 , n62421 , n62629 );
xor ( n62641 , n62640 , n62632 );
xor ( n589965 , n589733 , n62412 );
xor ( n62643 , n589965 , n589738 );
xor ( n62644 , n62424 , n62472 );
xor ( n589968 , n62644 , n62519 );
xor ( n62646 , n589749 , n62437 );
xor ( n62647 , n62646 , n62469 );
xor ( n589971 , n62511 , n62513 );
xor ( n62649 , n589971 , n62516 );
and ( n62650 , n62647 , n62649 );
xor ( n62651 , n589812 , n589828 );
xor ( n62652 , n62651 , n589831 );
xor ( n589976 , n589816 , n589820 );
xor ( n62654 , n589976 , n589825 );
and ( n589978 , n585586 , n53177 );
and ( n62656 , n58246 , n53175 );
nor ( n589980 , n589978 , n62656 );
xnor ( n589981 , n589980 , n52827 );
and ( n62659 , n58623 , n52978 );
and ( n589983 , n585909 , n52976 );
nor ( n589984 , n62659 , n589983 );
xnor ( n62662 , n589984 , n52680 );
and ( n62663 , n589981 , n62662 );
xor ( n589987 , n62546 , n589871 );
xor ( n589988 , n589987 , n589874 );
and ( n62666 , n62662 , n589988 );
and ( n62667 , n589981 , n589988 );
or ( n589991 , n62663 , n62666 , n62667 );
and ( n589992 , n62654 , n589991 );
xor ( n589993 , n589880 , n52153 );
nor ( n589994 , n52707 , n52705 );
xnor ( n589995 , n589994 , n52526 );
nor ( n62673 , n52509 , n52507 );
xnor ( n589997 , n62673 , n52383 );
and ( n589998 , n589995 , n589997 );
nor ( n62676 , n52432 , n52430 );
xnor ( n590000 , n62676 , n52255 );
and ( n62678 , n589997 , n590000 );
and ( n590002 , n589995 , n590000 );
or ( n590003 , n589998 , n62678 , n590002 );
and ( n62681 , n589993 , n590003 );
and ( n62682 , n56909 , n55013 );
and ( n62683 , n56832 , n55010 );
nor ( n62684 , n62682 , n62683 );
xnor ( n62685 , n62684 , n53762 );
and ( n62686 , n584529 , n54532 );
and ( n62687 , n57058 , n54530 );
nor ( n590011 , n62686 , n62687 );
xnor ( n62689 , n590011 , n53769 );
and ( n590013 , n62685 , n62689 );
and ( n590014 , n57484 , n54414 );
and ( n62692 , n57283 , n54412 );
nor ( n590016 , n590014 , n62692 );
xnor ( n590017 , n590016 , n53650 );
and ( n62695 , n62689 , n590017 );
and ( n590019 , n62685 , n590017 );
or ( n590020 , n590013 , n62695 , n590019 );
and ( n590021 , n590003 , n590020 );
and ( n62699 , n589993 , n590020 );
or ( n590023 , n62681 , n590021 , n62699 );
and ( n62701 , n589991 , n590023 );
and ( n590025 , n62654 , n590023 );
or ( n590026 , n589992 , n62701 , n590025 );
and ( n62704 , n62652 , n590026 );
and ( n62705 , n585062 , n53996 );
and ( n62706 , n57482 , n53994 );
nor ( n62707 , n62705 , n62706 );
xnor ( n590031 , n62707 , n53376 );
and ( n62709 , n585221 , n53683 );
and ( n62710 , n57900 , n53681 );
nor ( n62711 , n62709 , n62710 );
xnor ( n62712 , n62711 , n53118 );
and ( n590036 , n590031 , n62712 );
and ( n590037 , n58246 , n53468 );
and ( n62715 , n58219 , n53466 );
nor ( n62716 , n590037 , n62715 );
xnor ( n590040 , n62716 , n52945 );
and ( n62718 , n62712 , n590040 );
and ( n590042 , n590031 , n590040 );
or ( n62720 , n590036 , n62718 , n590042 );
and ( n62721 , n585909 , n53177 );
and ( n62722 , n585586 , n53175 );
nor ( n590046 , n62721 , n62722 );
xnor ( n62724 , n590046 , n52827 );
and ( n590048 , n585973 , n52978 );
and ( n590049 , n58623 , n52976 );
nor ( n590050 , n590048 , n590049 );
xnor ( n62728 , n590050 , n52680 );
and ( n590052 , n62724 , n62728 );
nor ( n590053 , n52273 , n52271 );
xnor ( n62731 , n590053 , n52137 );
and ( n590055 , n62728 , n62731 );
and ( n590056 , n62724 , n62731 );
or ( n62734 , n590052 , n590055 , n590056 );
and ( n62735 , n62720 , n62734 );
xor ( n590059 , n589886 , n62567 );
xor ( n590060 , n590059 , n589895 );
and ( n62738 , n62734 , n590060 );
and ( n62739 , n62720 , n590060 );
or ( n590063 , n62735 , n62738 , n62739 );
xor ( n62741 , n62536 , n62537 );
xor ( n62742 , n62741 , n62540 );
and ( n62743 , n590063 , n62742 );
xor ( n62744 , n589877 , n62558 );
xor ( n62745 , n62744 , n589898 );
and ( n590069 , n62742 , n62745 );
and ( n62747 , n590063 , n62745 );
or ( n590071 , n62743 , n590069 , n62747 );
and ( n590072 , n590026 , n590071 );
and ( n62750 , n62652 , n590071 );
or ( n590074 , n62704 , n590072 , n62750 );
and ( n590075 , n62649 , n590074 );
and ( n62753 , n62647 , n590074 );
or ( n62754 , n62650 , n590075 , n62753 );
and ( n590078 , n589968 , n62754 );
xor ( n590079 , n62527 , n62529 );
xor ( n62757 , n590079 , n62617 );
and ( n62758 , n62754 , n62757 );
and ( n590082 , n589968 , n62757 );
or ( n62760 , n590078 , n62758 , n590082 );
and ( n62761 , n62643 , n62760 );
xor ( n62762 , n589845 , n62524 );
xor ( n62763 , n62762 , n589943 );
and ( n62764 , n62760 , n62763 );
and ( n62765 , n62643 , n62763 );
or ( n62766 , n62761 , n62764 , n62765 );
xor ( n62767 , n589745 , n589946 );
xor ( n62768 , n62767 , n62626 );
and ( n62769 , n62766 , n62768 );
xor ( n590093 , n62766 , n62768 );
xor ( n62771 , n62643 , n62760 );
xor ( n62772 , n62771 , n62763 );
xor ( n590096 , n62532 , n589904 );
xor ( n62774 , n590096 , n62614 );
xor ( n62775 , n62534 , n62543 );
xor ( n62776 , n62775 , n62578 );
xor ( n62777 , n62606 , n589931 );
xor ( n590101 , n62777 , n62611 );
and ( n62779 , n62776 , n590101 );
xor ( n62780 , n62598 , n62600 );
xor ( n62781 , n62780 , n589926 );
xor ( n62782 , n589909 , n62590 );
xor ( n62783 , n62782 , n62595 );
and ( n590107 , n52272 , n52137 );
xor ( n590108 , n589995 , n589997 );
xor ( n590109 , n590108 , n590000 );
and ( n62787 , n590107 , n590109 );
nor ( n590111 , n52707 , n52705 );
xnor ( n590112 , n590111 , n52526 );
nor ( n590113 , n52509 , n52507 );
xnor ( n62791 , n590113 , n52383 );
and ( n590115 , n590112 , n62791 );
nor ( n62793 , n52432 , n52430 );
xnor ( n62794 , n62793 , n52255 );
and ( n590118 , n62791 , n62794 );
and ( n590119 , n590112 , n62794 );
or ( n62797 , n590115 , n590118 , n590119 );
and ( n590121 , n590109 , n62797 );
and ( n62799 , n590107 , n62797 );
or ( n62800 , n62787 , n590121 , n62799 );
and ( n62801 , n62783 , n62800 );
and ( n62802 , n585973 , n52976 );
nor ( n590126 , n52978 , n62802 );
xnor ( n590127 , n590126 , n52680 );
and ( n590128 , n590127 , n52271 );
and ( n62806 , n57058 , n55013 );
and ( n590130 , n56909 , n55010 );
nor ( n590131 , n62806 , n590130 );
xnor ( n590132 , n590131 , n53762 );
and ( n590133 , n57283 , n54532 );
and ( n62811 , n584529 , n54530 );
nor ( n590135 , n590133 , n62811 );
xnor ( n590136 , n590135 , n53769 );
and ( n62814 , n590132 , n590136 );
and ( n590138 , n57482 , n54414 );
and ( n590139 , n57484 , n54412 );
nor ( n62817 , n590138 , n590139 );
xnor ( n590141 , n62817 , n53650 );
and ( n590142 , n590136 , n590141 );
and ( n62820 , n590132 , n590141 );
or ( n62821 , n62814 , n590142 , n62820 );
and ( n62822 , n590128 , n62821 );
and ( n590146 , n57900 , n53996 );
and ( n590147 , n585062 , n53994 );
nor ( n590148 , n590146 , n590147 );
xnor ( n62826 , n590148 , n53376 );
and ( n590150 , n58219 , n53683 );
and ( n590151 , n585221 , n53681 );
nor ( n590152 , n590150 , n590151 );
xnor ( n590153 , n590152 , n53118 );
and ( n62831 , n62826 , n590153 );
and ( n590155 , n585586 , n53468 );
and ( n590156 , n58246 , n53466 );
nor ( n62834 , n590155 , n590156 );
xnor ( n590158 , n62834 , n52945 );
and ( n590159 , n590153 , n590158 );
and ( n62837 , n62826 , n590158 );
or ( n590161 , n62831 , n590159 , n62837 );
and ( n590162 , n62821 , n590161 );
and ( n62840 , n590128 , n590161 );
or ( n62841 , n62822 , n590162 , n62840 );
and ( n62842 , n62800 , n62841 );
and ( n590166 , n62783 , n62841 );
or ( n62844 , n62801 , n62842 , n590166 );
and ( n62845 , n62781 , n62844 );
xor ( n590169 , n62685 , n62689 );
xor ( n590170 , n590169 , n590017 );
xor ( n62848 , n590031 , n62712 );
xor ( n590172 , n62848 , n590040 );
and ( n62850 , n590170 , n590172 );
xor ( n62851 , n62724 , n62728 );
xor ( n62852 , n62851 , n62731 );
and ( n62853 , n590172 , n62852 );
and ( n62854 , n590170 , n62852 );
or ( n590178 , n62850 , n62853 , n62854 );
xor ( n62856 , n589981 , n62662 );
xor ( n590180 , n62856 , n589988 );
and ( n590181 , n590178 , n590180 );
xor ( n62859 , n589993 , n590003 );
xor ( n590183 , n62859 , n590020 );
and ( n590184 , n590180 , n590183 );
and ( n62862 , n590178 , n590183 );
or ( n62863 , n590181 , n590184 , n62862 );
and ( n590187 , n62844 , n62863 );
and ( n62865 , n62781 , n62863 );
or ( n62866 , n62845 , n590187 , n62865 );
and ( n590190 , n590101 , n62866 );
and ( n62868 , n62776 , n62866 );
or ( n590192 , n62779 , n590190 , n62868 );
and ( n590193 , n62774 , n590192 );
xor ( n62871 , n62647 , n62649 );
xor ( n62872 , n62871 , n590074 );
and ( n62873 , n590192 , n62872 );
and ( n590197 , n62774 , n62872 );
or ( n590198 , n590193 , n62873 , n590197 );
xor ( n590199 , n589968 , n62754 );
xor ( n590200 , n590199 , n62757 );
and ( n62878 , n590198 , n590200 );
xor ( n590202 , n590198 , n590200 );
xor ( n590203 , n62652 , n590026 );
xor ( n62881 , n590203 , n590071 );
xor ( n590205 , n62654 , n589991 );
xor ( n590206 , n590205 , n590023 );
xor ( n62884 , n590063 , n62742 );
xor ( n590208 , n62884 , n62745 );
and ( n590209 , n590206 , n590208 );
xor ( n62887 , n62720 , n62734 );
xor ( n62888 , n62887 , n590060 );
xor ( n590212 , n590112 , n62791 );
xor ( n590213 , n590212 , n62794 );
xor ( n62891 , n590127 , n52271 );
and ( n590215 , n590213 , n62891 );
nor ( n590216 , n52707 , n52705 );
xnor ( n62894 , n590216 , n52526 );
nor ( n590218 , n52509 , n52507 );
xnor ( n590219 , n590218 , n52383 );
and ( n62897 , n62894 , n590219 );
nor ( n590221 , n52432 , n52430 );
xnor ( n590222 , n590221 , n52255 );
and ( n62900 , n590219 , n590222 );
and ( n590224 , n62894 , n590222 );
or ( n62902 , n62897 , n62900 , n590224 );
and ( n62903 , n62891 , n62902 );
and ( n62904 , n590213 , n62902 );
or ( n590228 , n590215 , n62903 , n62904 );
nor ( n62906 , n52978 , n52976 );
xnor ( n590230 , n62906 , n52680 );
and ( n62908 , n52431 , n52255 );
and ( n62909 , n590230 , n62908 );
and ( n590233 , n584529 , n55013 );
and ( n590234 , n57058 , n55010 );
nor ( n62912 , n590233 , n590234 );
xnor ( n62913 , n62912 , n53762 );
and ( n590237 , n57484 , n54532 );
and ( n590238 , n57283 , n54530 );
nor ( n62916 , n590237 , n590238 );
xnor ( n590240 , n62916 , n53769 );
and ( n62918 , n62913 , n590240 );
and ( n62919 , n585062 , n54414 );
and ( n590243 , n57482 , n54412 );
nor ( n590244 , n62919 , n590243 );
xnor ( n62922 , n590244 , n53650 );
and ( n62923 , n590240 , n62922 );
and ( n590247 , n62913 , n62922 );
or ( n62925 , n62918 , n62923 , n590247 );
and ( n62926 , n62909 , n62925 );
and ( n62927 , n585221 , n53996 );
and ( n62928 , n57900 , n53994 );
nor ( n62929 , n62927 , n62928 );
xnor ( n62930 , n62929 , n53376 );
and ( n590254 , n58246 , n53683 );
and ( n62932 , n58219 , n53681 );
nor ( n62933 , n590254 , n62932 );
xnor ( n62934 , n62933 , n53118 );
and ( n62935 , n62930 , n62934 );
and ( n590259 , n585909 , n53468 );
and ( n590260 , n585586 , n53466 );
nor ( n62938 , n590259 , n590260 );
xnor ( n62939 , n62938 , n52945 );
and ( n62940 , n62934 , n62939 );
and ( n590264 , n62930 , n62939 );
or ( n590265 , n62935 , n62940 , n590264 );
and ( n62943 , n62925 , n590265 );
and ( n590267 , n62909 , n590265 );
or ( n590268 , n62926 , n62943 , n590267 );
and ( n62946 , n590228 , n590268 );
xor ( n62947 , n590107 , n590109 );
xor ( n590271 , n62947 , n62797 );
and ( n62949 , n590268 , n590271 );
and ( n62950 , n590228 , n590271 );
or ( n62951 , n62946 , n62949 , n62950 );
and ( n62952 , n62888 , n62951 );
xor ( n590276 , n62783 , n62800 );
xor ( n62954 , n590276 , n62841 );
and ( n62955 , n62951 , n62954 );
and ( n590279 , n62888 , n62954 );
or ( n590280 , n62952 , n62955 , n590279 );
and ( n62958 , n590208 , n590280 );
and ( n62959 , n590206 , n590280 );
or ( n590283 , n590209 , n62958 , n62959 );
and ( n590284 , n62881 , n590283 );
xor ( n62962 , n62776 , n590101 );
xor ( n590286 , n62962 , n62866 );
and ( n62964 , n590283 , n590286 );
and ( n62965 , n62881 , n590286 );
or ( n590289 , n590284 , n62964 , n62965 );
xor ( n590290 , n62774 , n590192 );
xor ( n62968 , n590290 , n62872 );
and ( n62969 , n590289 , n62968 );
xor ( n590293 , n590289 , n62968 );
xor ( n590294 , n62781 , n62844 );
xor ( n62972 , n590294 , n62863 );
xor ( n62973 , n590178 , n590180 );
xor ( n590297 , n62973 , n590183 );
xor ( n590298 , n590128 , n62821 );
xor ( n62976 , n590298 , n590161 );
xor ( n590300 , n590170 , n590172 );
xor ( n590301 , n590300 , n62852 );
and ( n62979 , n62976 , n590301 );
xor ( n590303 , n590230 , n62908 );
and ( n590304 , n585973 , n53175 );
nor ( n62982 , n53177 , n590304 );
xnor ( n590306 , n62982 , n52827 );
nor ( n62984 , n52978 , n52976 );
xnor ( n62985 , n62984 , n52680 );
and ( n62986 , n590306 , n62985 );
and ( n590310 , n62985 , n52430 );
and ( n590311 , n590306 , n52430 );
or ( n62989 , n62986 , n590310 , n590311 );
and ( n590313 , n590303 , n62989 );
and ( n62991 , n585973 , n53177 );
and ( n590315 , n58623 , n53175 );
nor ( n62993 , n62991 , n590315 );
xnor ( n62994 , n62993 , n52827 );
and ( n590318 , n62989 , n62994 );
and ( n62996 , n590303 , n62994 );
or ( n590320 , n590313 , n590318 , n62996 );
and ( n62998 , n58623 , n53177 );
and ( n590322 , n585909 , n53175 );
nor ( n590323 , n62998 , n590322 );
xnor ( n63001 , n590323 , n52827 );
and ( n590325 , n590320 , n63001 );
and ( n590326 , n590301 , n590325 );
and ( n63004 , n62976 , n590325 );
or ( n63005 , n62979 , n590326 , n63004 );
and ( n63006 , n590297 , n63005 );
xor ( n63007 , n62888 , n62951 );
xor ( n63008 , n63007 , n62954 );
and ( n590332 , n63005 , n63008 );
and ( n63010 , n590297 , n63008 );
or ( n63011 , n63006 , n590332 , n63010 );
and ( n590335 , n62972 , n63011 );
xor ( n63013 , n590206 , n590208 );
xor ( n63014 , n63013 , n590280 );
and ( n63015 , n63011 , n63014 );
and ( n63016 , n62972 , n63014 );
or ( n590340 , n590335 , n63015 , n63016 );
xor ( n63018 , n62881 , n590283 );
xor ( n63019 , n63018 , n590286 );
and ( n63020 , n590340 , n63019 );
xor ( n63021 , n590340 , n63019 );
xor ( n63022 , n62972 , n63011 );
xor ( n590346 , n63022 , n63014 );
xor ( n63024 , n590132 , n590136 );
xor ( n63025 , n63024 , n590141 );
xor ( n63026 , n62826 , n590153 );
xor ( n63027 , n63026 , n590158 );
and ( n63028 , n63025 , n63027 );
xor ( n63029 , n62894 , n590219 );
xor ( n63030 , n63029 , n590222 );
and ( n590354 , n57283 , n55013 );
and ( n63032 , n584529 , n55010 );
nor ( n590356 , n590354 , n63032 );
xnor ( n590357 , n590356 , n53762 );
and ( n63035 , n57482 , n54532 );
and ( n590359 , n57484 , n54530 );
nor ( n590360 , n63035 , n590359 );
xnor ( n63038 , n590360 , n53769 );
and ( n63039 , n590357 , n63038 );
and ( n590363 , n57900 , n54414 );
and ( n590364 , n585062 , n54412 );
nor ( n63042 , n590363 , n590364 );
xnor ( n63043 , n63042 , n53650 );
and ( n590367 , n63038 , n63043 );
and ( n63045 , n590357 , n63043 );
or ( n63046 , n63039 , n590367 , n63045 );
and ( n590370 , n63030 , n63046 );
and ( n590371 , n58219 , n53996 );
and ( n63049 , n585221 , n53994 );
nor ( n590373 , n590371 , n63049 );
xnor ( n590374 , n590373 , n53376 );
and ( n590375 , n585586 , n53683 );
and ( n590376 , n58246 , n53681 );
nor ( n63054 , n590375 , n590376 );
xnor ( n590378 , n63054 , n53118 );
and ( n590379 , n590374 , n590378 );
and ( n63057 , n58623 , n53468 );
and ( n590381 , n585909 , n53466 );
nor ( n590382 , n63057 , n590381 );
xnor ( n63060 , n590382 , n52945 );
and ( n590384 , n590378 , n63060 );
and ( n590385 , n590374 , n63060 );
or ( n63063 , n590379 , n590384 , n590385 );
and ( n63064 , n63046 , n63063 );
and ( n63065 , n63030 , n63063 );
or ( n590389 , n590370 , n63064 , n63065 );
and ( n63067 , n63027 , n590389 );
and ( n590391 , n63025 , n590389 );
or ( n590392 , n63028 , n63067 , n590391 );
xor ( n63070 , n590228 , n590268 );
xor ( n590394 , n63070 , n590271 );
and ( n590395 , n590392 , n590394 );
xor ( n590396 , n590213 , n62891 );
xor ( n63074 , n590396 , n62902 );
xor ( n590398 , n62909 , n62925 );
xor ( n63076 , n590398 , n590265 );
and ( n63077 , n63074 , n63076 );
xor ( n63078 , n590320 , n63001 );
and ( n63079 , n63076 , n63078 );
and ( n63080 , n63074 , n63078 );
or ( n63081 , n63077 , n63079 , n63080 );
and ( n63082 , n590394 , n63081 );
and ( n63083 , n590392 , n63081 );
or ( n63084 , n590395 , n63082 , n63083 );
xor ( n63085 , n590297 , n63005 );
xor ( n63086 , n63085 , n63008 );
and ( n63087 , n63084 , n63086 );
xor ( n63088 , n62913 , n590240 );
xor ( n63089 , n63088 , n62922 );
xor ( n63090 , n62930 , n62934 );
xor ( n590414 , n63090 , n62939 );
and ( n63092 , n63089 , n590414 );
xor ( n63093 , n590303 , n62989 );
xor ( n590417 , n63093 , n62994 );
and ( n590418 , n590414 , n590417 );
and ( n63096 , n63089 , n590417 );
or ( n63097 , n63092 , n590418 , n63096 );
nor ( n590421 , n52707 , n52705 );
xnor ( n63099 , n590421 , n52526 );
nor ( n63100 , n52509 , n52507 );
xnor ( n63101 , n63100 , n52383 );
and ( n63102 , n63099 , n63101 );
xor ( n590426 , n590306 , n62985 );
xor ( n590427 , n590426 , n52430 );
and ( n590428 , n63101 , n590427 );
and ( n63106 , n63099 , n590427 );
or ( n590430 , n63102 , n590428 , n63106 );
nor ( n590431 , n53177 , n53175 );
xnor ( n590432 , n590431 , n52827 );
nor ( n590433 , n52978 , n52976 );
xnor ( n63111 , n590433 , n52680 );
and ( n590435 , n590432 , n63111 );
nor ( n590436 , n52707 , n52705 );
xnor ( n63114 , n590436 , n52526 );
and ( n590438 , n63111 , n63114 );
and ( n590439 , n590432 , n63114 );
or ( n63117 , n590435 , n590438 , n590439 );
and ( n590441 , n57484 , n55013 );
and ( n590442 , n57283 , n55010 );
nor ( n63120 , n590441 , n590442 );
xnor ( n63121 , n63120 , n53762 );
and ( n63122 , n585062 , n54532 );
and ( n590446 , n57482 , n54530 );
nor ( n590447 , n63122 , n590446 );
xnor ( n63125 , n590447 , n53769 );
and ( n63126 , n63121 , n63125 );
and ( n63127 , n585221 , n54414 );
and ( n590451 , n57900 , n54412 );
nor ( n63129 , n63127 , n590451 );
xnor ( n590453 , n63129 , n53650 );
and ( n590454 , n63125 , n590453 );
and ( n63132 , n63121 , n590453 );
or ( n590456 , n63126 , n590454 , n63132 );
and ( n590457 , n63117 , n590456 );
and ( n590458 , n58246 , n53996 );
and ( n63136 , n58219 , n53994 );
nor ( n590460 , n590458 , n63136 );
xnor ( n63138 , n590460 , n53376 );
and ( n63139 , n585909 , n53683 );
and ( n63140 , n585586 , n53681 );
nor ( n63141 , n63139 , n63140 );
xnor ( n63142 , n63141 , n53118 );
and ( n63143 , n63138 , n63142 );
and ( n590467 , n585973 , n53468 );
and ( n63145 , n58623 , n53466 );
nor ( n63146 , n590467 , n63145 );
xnor ( n63147 , n63146 , n52945 );
and ( n590471 , n63142 , n63147 );
and ( n590472 , n63138 , n63147 );
or ( n590473 , n63143 , n590471 , n590472 );
and ( n590474 , n590456 , n590473 );
and ( n63152 , n63117 , n590473 );
or ( n590476 , n590457 , n590474 , n63152 );
and ( n590477 , n590430 , n590476 );
xor ( n590478 , n63030 , n63046 );
xor ( n590479 , n590478 , n63063 );
and ( n63157 , n590476 , n590479 );
and ( n590481 , n590430 , n590479 );
or ( n590482 , n590477 , n63157 , n590481 );
and ( n63160 , n63097 , n590482 );
xor ( n590484 , n63025 , n63027 );
xor ( n590485 , n590484 , n590389 );
and ( n63163 , n590482 , n590485 );
and ( n590487 , n63097 , n590485 );
or ( n590488 , n63160 , n63163 , n590487 );
xor ( n63166 , n62976 , n590301 );
xor ( n590490 , n63166 , n590325 );
and ( n590491 , n590488 , n590490 );
xor ( n63169 , n590357 , n63038 );
xor ( n63170 , n63169 , n63043 );
xor ( n590494 , n590374 , n590378 );
xor ( n590495 , n590494 , n63060 );
and ( n63173 , n63170 , n590495 );
nor ( n590497 , n52509 , n52507 );
xnor ( n63175 , n590497 , n52383 );
and ( n63176 , n52508 , n52383 );
and ( n63177 , n63175 , n63176 );
xor ( n63178 , n590432 , n63111 );
xor ( n63179 , n63178 , n63114 );
and ( n590503 , n63176 , n63179 );
and ( n590504 , n63175 , n63179 );
or ( n63182 , n63177 , n590503 , n590504 );
and ( n590506 , n590495 , n63182 );
and ( n63184 , n63170 , n63182 );
or ( n590508 , n63173 , n590506 , n63184 );
nor ( n590509 , n53177 , n53175 );
xnor ( n63187 , n590509 , n52827 );
nor ( n590511 , n52978 , n52976 );
xnor ( n63189 , n590511 , n52680 );
and ( n63190 , n63187 , n63189 );
nor ( n590514 , n52707 , n52705 );
xnor ( n590515 , n590514 , n52526 );
and ( n63193 , n63189 , n590515 );
and ( n590517 , n63187 , n590515 );
or ( n590518 , n63190 , n63193 , n590517 );
and ( n63196 , n57482 , n55013 );
and ( n590520 , n57484 , n55010 );
nor ( n590521 , n63196 , n590520 );
xnor ( n63199 , n590521 , n53762 );
and ( n590523 , n57900 , n54532 );
and ( n63201 , n585062 , n54530 );
nor ( n63202 , n590523 , n63201 );
xnor ( n63203 , n63202 , n53769 );
and ( n63204 , n63199 , n63203 );
and ( n590528 , n58219 , n54414 );
and ( n63206 , n585221 , n54412 );
nor ( n63207 , n590528 , n63206 );
xnor ( n63208 , n63207 , n53650 );
and ( n63209 , n63203 , n63208 );
and ( n63210 , n63199 , n63208 );
or ( n63211 , n63204 , n63209 , n63210 );
and ( n63212 , n590518 , n63211 );
and ( n63213 , n585586 , n53996 );
and ( n63214 , n58246 , n53994 );
nor ( n63215 , n63213 , n63214 );
xnor ( n590539 , n63215 , n53376 );
and ( n63217 , n58623 , n53683 );
and ( n63218 , n585909 , n53681 );
nor ( n63219 , n63217 , n63218 );
xnor ( n63220 , n63219 , n53118 );
and ( n63221 , n590539 , n63220 );
and ( n63222 , n585973 , n53466 );
nor ( n590546 , n53468 , n63222 );
xnor ( n590547 , n590546 , n52945 );
and ( n63225 , n63220 , n590547 );
and ( n590549 , n590539 , n590547 );
or ( n63227 , n63221 , n63225 , n590549 );
and ( n63228 , n63211 , n63227 );
and ( n63229 , n590518 , n63227 );
or ( n63230 , n63212 , n63228 , n63229 );
xor ( n63231 , n63099 , n63101 );
xor ( n63232 , n63231 , n590427 );
and ( n63233 , n63230 , n63232 );
xor ( n63234 , n63117 , n590456 );
xor ( n63235 , n63234 , n590473 );
and ( n63236 , n63232 , n63235 );
and ( n63237 , n63230 , n63235 );
or ( n63238 , n63233 , n63236 , n63237 );
and ( n590562 , n590508 , n63238 );
xor ( n63240 , n63089 , n590414 );
xor ( n63241 , n63240 , n590417 );
and ( n63242 , n63238 , n63241 );
and ( n590566 , n590508 , n63241 );
or ( n590567 , n590562 , n63242 , n590566 );
xor ( n590568 , n63074 , n63076 );
xor ( n590569 , n590568 , n63078 );
and ( n63247 , n590567 , n590569 );
xor ( n590571 , n63097 , n590482 );
xor ( n590572 , n590571 , n590485 );
and ( n590573 , n590569 , n590572 );
and ( n63251 , n590567 , n590572 );
or ( n590575 , n63247 , n590573 , n63251 );
and ( n63253 , n590490 , n590575 );
and ( n590577 , n590488 , n590575 );
or ( n590578 , n590491 , n63253 , n590577 );
and ( n63256 , n63086 , n590578 );
and ( n590580 , n63084 , n590578 );
or ( n63258 , n63087 , n63256 , n590580 );
and ( n63259 , n590346 , n63258 );
xor ( n63260 , n590346 , n63258 );
xor ( n63261 , n63084 , n63086 );
xor ( n63262 , n63261 , n590578 );
xor ( n63263 , n590392 , n590394 );
xor ( n63264 , n63263 , n63081 );
xor ( n63265 , n590488 , n590490 );
xor ( n63266 , n63265 , n590575 );
and ( n63267 , n63264 , n63266 );
xor ( n590591 , n63264 , n63266 );
xor ( n590592 , n590430 , n590476 );
xor ( n63270 , n590592 , n590479 );
xor ( n590594 , n63121 , n63125 );
xor ( n63272 , n590594 , n590453 );
xor ( n63273 , n63138 , n63142 );
xor ( n63274 , n63273 , n63147 );
and ( n63275 , n63272 , n63274 );
xor ( n63276 , n63187 , n63189 );
xor ( n590600 , n63276 , n590515 );
and ( n63278 , n52507 , n590600 );
nor ( n63279 , n53468 , n53466 );
xnor ( n63280 , n63279 , n52945 );
nor ( n63281 , n53177 , n53175 );
xnor ( n63282 , n63281 , n52827 );
and ( n63283 , n63280 , n63282 );
nor ( n63284 , n52978 , n52976 );
xnor ( n63285 , n63284 , n52680 );
and ( n590609 , n63282 , n63285 );
and ( n63287 , n63280 , n63285 );
or ( n63288 , n63283 , n590609 , n63287 );
and ( n590612 , n590600 , n63288 );
and ( n63290 , n52507 , n63288 );
or ( n63291 , n63278 , n590612 , n63290 );
and ( n63292 , n63274 , n63291 );
and ( n63293 , n63272 , n63291 );
or ( n590617 , n63275 , n63292 , n63293 );
and ( n590618 , n585062 , n55013 );
and ( n63296 , n57482 , n55010 );
nor ( n590620 , n590618 , n63296 );
xnor ( n63298 , n590620 , n53762 );
and ( n63299 , n585221 , n54532 );
and ( n590623 , n57900 , n54530 );
nor ( n590624 , n63299 , n590623 );
xnor ( n63302 , n590624 , n53769 );
and ( n590626 , n63298 , n63302 );
and ( n63304 , n58246 , n54414 );
and ( n590628 , n58219 , n54412 );
nor ( n590629 , n63304 , n590628 );
xnor ( n63307 , n590629 , n53650 );
and ( n590631 , n63302 , n63307 );
and ( n590632 , n63298 , n63307 );
or ( n63310 , n590626 , n590631 , n590632 );
and ( n590634 , n585909 , n53996 );
and ( n590635 , n585586 , n53994 );
nor ( n590636 , n590634 , n590635 );
xnor ( n590637 , n590636 , n53376 );
and ( n63315 , n585973 , n53683 );
and ( n590639 , n58623 , n53681 );
nor ( n63317 , n63315 , n590639 );
xnor ( n63318 , n63317 , n53118 );
and ( n63319 , n590637 , n63318 );
nor ( n63320 , n52707 , n52705 );
xnor ( n63321 , n63320 , n52526 );
and ( n63322 , n63318 , n63321 );
and ( n63323 , n590637 , n63321 );
or ( n63324 , n63319 , n63322 , n63323 );
and ( n63325 , n63310 , n63324 );
xor ( n63326 , n63199 , n63203 );
xor ( n63327 , n63326 , n63208 );
and ( n63328 , n63324 , n63327 );
and ( n590652 , n63310 , n63327 );
or ( n63330 , n63325 , n63328 , n590652 );
xor ( n590654 , n63175 , n63176 );
xor ( n63332 , n590654 , n63179 );
and ( n590656 , n63330 , n63332 );
xor ( n590657 , n590518 , n63211 );
xor ( n63335 , n590657 , n63227 );
and ( n590659 , n63332 , n63335 );
and ( n590660 , n63330 , n63335 );
or ( n63338 , n590656 , n590659 , n590660 );
and ( n63339 , n590617 , n63338 );
xor ( n590663 , n63170 , n590495 );
xor ( n590664 , n590663 , n63182 );
and ( n63342 , n63338 , n590664 );
and ( n63343 , n590617 , n590664 );
or ( n590667 , n63339 , n63342 , n63343 );
and ( n590668 , n63270 , n590667 );
xor ( n590669 , n590508 , n63238 );
xor ( n63347 , n590669 , n63241 );
and ( n590671 , n590667 , n63347 );
and ( n590672 , n63270 , n63347 );
or ( n63350 , n590668 , n590671 , n590672 );
xor ( n590674 , n590567 , n590569 );
xor ( n590675 , n590674 , n590572 );
and ( n63353 , n63350 , n590675 );
xor ( n63354 , n63350 , n590675 );
xor ( n590678 , n63230 , n63232 );
xor ( n590679 , n590678 , n63235 );
xor ( n63357 , n590539 , n63220 );
xor ( n63358 , n63357 , n590547 );
and ( n590682 , n52706 , n52526 );
xor ( n590683 , n63280 , n63282 );
xor ( n63361 , n590683 , n63285 );
and ( n63362 , n590682 , n63361 );
nor ( n63363 , n53468 , n53466 );
xnor ( n63364 , n63363 , n52945 );
nor ( n63365 , n53177 , n53175 );
xnor ( n63366 , n63365 , n52827 );
and ( n63367 , n63364 , n63366 );
nor ( n590691 , n52978 , n52976 );
xnor ( n63369 , n590691 , n52680 );
and ( n63370 , n63366 , n63369 );
and ( n63371 , n63364 , n63369 );
or ( n590695 , n63367 , n63370 , n63371 );
and ( n590696 , n63361 , n590695 );
and ( n63374 , n590682 , n590695 );
or ( n590698 , n63362 , n590696 , n63374 );
and ( n590699 , n63358 , n590698 );
and ( n63377 , n585973 , n53681 );
nor ( n63378 , n53683 , n63377 );
xnor ( n63379 , n63378 , n53118 );
and ( n63380 , n63379 , n52705 );
and ( n63381 , n57900 , n55013 );
and ( n63382 , n585062 , n55010 );
nor ( n63383 , n63381 , n63382 );
xnor ( n63384 , n63383 , n53762 );
and ( n63385 , n58219 , n54532 );
and ( n590709 , n585221 , n54530 );
nor ( n63387 , n63385 , n590709 );
xnor ( n590711 , n63387 , n53769 );
and ( n590712 , n63384 , n590711 );
and ( n63390 , n585586 , n54414 );
and ( n590714 , n58246 , n54412 );
nor ( n590715 , n63390 , n590714 );
xnor ( n63393 , n590715 , n53650 );
and ( n63394 , n590711 , n63393 );
and ( n590718 , n63384 , n63393 );
or ( n590719 , n590712 , n63394 , n590718 );
and ( n63397 , n63380 , n590719 );
xor ( n63398 , n63298 , n63302 );
xor ( n590722 , n63398 , n63307 );
and ( n63400 , n590719 , n590722 );
and ( n63401 , n63380 , n590722 );
or ( n63402 , n63397 , n63400 , n63401 );
and ( n63403 , n590698 , n63402 );
and ( n63404 , n63358 , n63402 );
or ( n63405 , n590699 , n63403 , n63404 );
xor ( n63406 , n63272 , n63274 );
xor ( n63407 , n63406 , n63291 );
and ( n63408 , n63405 , n63407 );
xor ( n63409 , n63330 , n63332 );
xor ( n63410 , n63409 , n63335 );
and ( n63411 , n63407 , n63410 );
and ( n63412 , n63405 , n63410 );
or ( n590736 , n63408 , n63411 , n63412 );
and ( n63414 , n590679 , n590736 );
xor ( n590738 , n590617 , n63338 );
xor ( n590739 , n590738 , n590664 );
and ( n63417 , n590736 , n590739 );
and ( n63418 , n590679 , n590739 );
or ( n590742 , n63414 , n63417 , n63418 );
xor ( n63420 , n63270 , n590667 );
xor ( n590744 , n63420 , n63347 );
and ( n590745 , n590742 , n590744 );
xor ( n590746 , n590742 , n590744 );
xor ( n590747 , n590679 , n590736 );
xor ( n63425 , n590747 , n590739 );
xor ( n590749 , n52507 , n590600 );
xor ( n63427 , n590749 , n63288 );
xor ( n590751 , n63310 , n63324 );
xor ( n590752 , n590751 , n63327 );
and ( n63430 , n63427 , n590752 );
xor ( n63431 , n590637 , n63318 );
xor ( n63432 , n63431 , n63321 );
and ( n63433 , n58623 , n53996 );
and ( n590757 , n585909 , n53994 );
nor ( n63435 , n63433 , n590757 );
xnor ( n63436 , n63435 , n53376 );
xor ( n590760 , n63364 , n63366 );
xor ( n590761 , n590760 , n63369 );
and ( n63439 , n63436 , n590761 );
xor ( n590763 , n63379 , n52705 );
and ( n63441 , n590761 , n590763 );
and ( n590765 , n63436 , n590763 );
or ( n590766 , n63439 , n63441 , n590765 );
and ( n63444 , n63432 , n590766 );
nor ( n590768 , n53683 , n53681 );
xnor ( n590769 , n590768 , n53118 );
nor ( n590770 , n53468 , n53466 );
xnor ( n63448 , n590770 , n52945 );
and ( n590772 , n590769 , n63448 );
nor ( n63450 , n53177 , n53175 );
xnor ( n63451 , n63450 , n52827 );
and ( n63452 , n63448 , n63451 );
and ( n63453 , n590769 , n63451 );
or ( n63454 , n590772 , n63452 , n63453 );
and ( n63455 , n585221 , n55013 );
and ( n590779 , n57900 , n55010 );
nor ( n590780 , n63455 , n590779 );
xnor ( n590781 , n590780 , n53762 );
and ( n63459 , n58246 , n54532 );
and ( n590783 , n58219 , n54530 );
nor ( n590784 , n63459 , n590783 );
xnor ( n590785 , n590784 , n53769 );
and ( n590786 , n590781 , n590785 );
and ( n63464 , n585909 , n54414 );
and ( n590788 , n585586 , n54412 );
nor ( n590789 , n63464 , n590788 );
xnor ( n63467 , n590789 , n53650 );
and ( n590791 , n590785 , n63467 );
and ( n590792 , n590781 , n63467 );
or ( n63470 , n590786 , n590791 , n590792 );
and ( n590794 , n63454 , n63470 );
and ( n590795 , n585973 , n53996 );
and ( n63473 , n58623 , n53994 );
nor ( n590797 , n590795 , n63473 );
xnor ( n590798 , n590797 , n53376 );
nor ( n63476 , n52978 , n52976 );
xnor ( n63477 , n63476 , n52680 );
and ( n63478 , n590798 , n63477 );
and ( n63479 , n52977 , n52680 );
and ( n63480 , n63477 , n63479 );
and ( n63481 , n590798 , n63479 );
or ( n63482 , n63478 , n63480 , n63481 );
and ( n63483 , n63470 , n63482 );
and ( n63484 , n63454 , n63482 );
or ( n63485 , n590794 , n63483 , n63484 );
and ( n63486 , n590766 , n63485 );
and ( n63487 , n63432 , n63485 );
or ( n63488 , n63444 , n63486 , n63487 );
and ( n63489 , n590752 , n63488 );
and ( n63490 , n63427 , n63488 );
or ( n63491 , n63430 , n63489 , n63490 );
xor ( n63492 , n63405 , n63407 );
xor ( n590816 , n63492 , n63410 );
and ( n63494 , n63491 , n590816 );
xor ( n63495 , n63358 , n590698 );
xor ( n63496 , n63495 , n63402 );
xor ( n63497 , n590682 , n63361 );
xor ( n63498 , n63497 , n590695 );
xor ( n63499 , n63380 , n590719 );
xor ( n63500 , n63499 , n590722 );
and ( n63501 , n63498 , n63500 );
xor ( n63502 , n63384 , n590711 );
xor ( n63503 , n63502 , n63393 );
xor ( n590827 , n590769 , n63448 );
xor ( n63505 , n590827 , n63451 );
nor ( n63506 , n53683 , n53681 );
xnor ( n63507 , n63506 , n53118 );
nor ( n590831 , n53468 , n53466 );
xnor ( n590832 , n590831 , n52945 );
and ( n590833 , n63507 , n590832 );
nor ( n590834 , n53177 , n53175 );
xnor ( n63512 , n590834 , n52827 );
and ( n590836 , n590832 , n63512 );
and ( n590837 , n63507 , n63512 );
or ( n63515 , n590833 , n590836 , n590837 );
and ( n63516 , n63505 , n63515 );
xor ( n63517 , n590781 , n590785 );
xor ( n63518 , n63517 , n63467 );
and ( n590842 , n63515 , n63518 );
and ( n590843 , n63505 , n63518 );
or ( n63521 , n63516 , n590842 , n590843 );
and ( n63522 , n63503 , n63521 );
xor ( n63523 , n63436 , n590761 );
xor ( n63524 , n63523 , n590763 );
and ( n63525 , n63521 , n63524 );
and ( n590849 , n63503 , n63524 );
or ( n63527 , n63522 , n63525 , n590849 );
and ( n590851 , n63500 , n63527 );
and ( n590852 , n63498 , n63527 );
or ( n63530 , n63501 , n590851 , n590852 );
and ( n63531 , n63496 , n63530 );
xor ( n590855 , n63427 , n590752 );
xor ( n63533 , n590855 , n63488 );
and ( n63534 , n63530 , n63533 );
and ( n63535 , n63496 , n63533 );
or ( n63536 , n63531 , n63534 , n63535 );
and ( n590860 , n590816 , n63536 );
and ( n63538 , n63491 , n63536 );
or ( n63539 , n63494 , n590860 , n63538 );
and ( n590863 , n63425 , n63539 );
xor ( n63541 , n63425 , n63539 );
xor ( n63542 , n63491 , n590816 );
xor ( n590866 , n63542 , n63536 );
xor ( n63544 , n63432 , n590766 );
xor ( n63545 , n63544 , n63485 );
xor ( n590869 , n63454 , n63470 );
xor ( n63547 , n590869 , n63482 );
xor ( n63548 , n590798 , n63477 );
xor ( n63549 , n63548 , n63479 );
nor ( n63550 , n53996 , n53994 );
xnor ( n590874 , n63550 , n53376 );
and ( n63552 , n53176 , n52827 );
and ( n63553 , n590874 , n63552 );
and ( n590877 , n585973 , n53994 );
nor ( n63555 , n53996 , n590877 );
xnor ( n63556 , n63555 , n53376 );
and ( n63557 , n63553 , n63556 );
and ( n63558 , n63556 , n52976 );
and ( n590882 , n63553 , n52976 );
or ( n63560 , n63557 , n63558 , n590882 );
and ( n63561 , n63549 , n63560 );
xor ( n63562 , n63505 , n63515 );
xor ( n63563 , n63562 , n63518 );
and ( n63564 , n63560 , n63563 );
and ( n63565 , n63549 , n63563 );
or ( n63566 , n63561 , n63564 , n63565 );
and ( n63567 , n63547 , n63566 );
xor ( n590891 , n63503 , n63521 );
xor ( n63569 , n590891 , n63524 );
and ( n63570 , n63566 , n63569 );
and ( n590894 , n63547 , n63569 );
or ( n590895 , n63567 , n63570 , n590894 );
and ( n63573 , n63545 , n590895 );
xor ( n590897 , n63498 , n63500 );
xor ( n590898 , n590897 , n63527 );
and ( n63576 , n590895 , n590898 );
and ( n63577 , n63545 , n590898 );
or ( n590901 , n63573 , n63576 , n63577 );
xor ( n590902 , n63496 , n63530 );
xor ( n590903 , n590902 , n63533 );
and ( n590904 , n590901 , n590903 );
xor ( n63582 , n590901 , n590903 );
xor ( n590906 , n63545 , n590895 );
xor ( n590907 , n590906 , n590898 );
xor ( n63585 , n63547 , n63566 );
xor ( n63586 , n63585 , n63569 );
nor ( n63587 , n53683 , n53681 );
xnor ( n63588 , n63587 , n53118 );
nor ( n590912 , n53468 , n53466 );
xnor ( n590913 , n590912 , n52945 );
and ( n590914 , n63588 , n590913 );
nor ( n63592 , n53177 , n53175 );
xnor ( n590916 , n63592 , n52827 );
and ( n590917 , n590913 , n590916 );
and ( n63595 , n63588 , n590916 );
or ( n63596 , n590914 , n590917 , n63595 );
xor ( n63597 , n63507 , n590832 );
xor ( n63598 , n63597 , n63512 );
and ( n63599 , n63596 , n63598 );
xor ( n590923 , n63553 , n63556 );
xor ( n590924 , n590923 , n52976 );
and ( n590925 , n63598 , n590924 );
and ( n63603 , n63596 , n590924 );
or ( n590927 , n63599 , n590925 , n63603 );
xor ( n590928 , n63549 , n63560 );
xor ( n63606 , n590928 , n63563 );
and ( n63607 , n590927 , n63606 );
xor ( n63608 , n590874 , n63552 );
and ( n63609 , n585973 , n54412 );
nor ( n590933 , n54414 , n63609 );
xnor ( n590934 , n590933 , n53650 );
nor ( n63612 , n53996 , n53994 );
xnor ( n590936 , n63612 , n53376 );
and ( n63614 , n590934 , n590936 );
and ( n63615 , n590936 , n53175 );
and ( n63616 , n590934 , n53175 );
or ( n63617 , n63614 , n63615 , n63616 );
and ( n63618 , n63608 , n63617 );
nor ( n63619 , n54414 , n54412 );
xnor ( n590943 , n63619 , n53650 );
nor ( n63621 , n53996 , n53994 );
xnor ( n63622 , n63621 , n53376 );
and ( n63623 , n590943 , n63622 );
nor ( n63624 , n53683 , n53681 );
xnor ( n590948 , n63624 , n53118 );
and ( n590949 , n63623 , n590948 );
nor ( n590950 , n53468 , n53466 );
xnor ( n590951 , n590950 , n52945 );
and ( n63629 , n590948 , n590951 );
and ( n590953 , n63623 , n590951 );
or ( n590954 , n590949 , n63629 , n590953 );
and ( n590955 , n63617 , n590954 );
and ( n63633 , n63608 , n590954 );
or ( n590957 , n63618 , n590955 , n63633 );
and ( n590958 , n58623 , n54414 );
and ( n590959 , n585909 , n54412 );
nor ( n63637 , n590958 , n590959 );
xnor ( n590961 , n63637 , n53650 );
and ( n63639 , n590957 , n590961 );
xor ( n63640 , n63596 , n63598 );
xor ( n63641 , n63640 , n590924 );
and ( n590965 , n590961 , n63641 );
and ( n63643 , n590957 , n63641 );
or ( n63644 , n63639 , n590965 , n63643 );
and ( n590968 , n63606 , n63644 );
and ( n63646 , n590927 , n63644 );
or ( n63647 , n63607 , n590968 , n63646 );
and ( n63648 , n63586 , n63647 );
and ( n63649 , n585973 , n54414 );
and ( n590973 , n58623 , n54412 );
nor ( n63651 , n63649 , n590973 );
xnor ( n63652 , n63651 , n53650 );
xor ( n590976 , n63588 , n590913 );
xor ( n63654 , n590976 , n590916 );
and ( n63655 , n63652 , n63654 );
xor ( n63656 , n63608 , n63617 );
xor ( n63657 , n63656 , n590954 );
and ( n590981 , n63654 , n63657 );
and ( n590982 , n63652 , n63657 );
or ( n590983 , n63655 , n590981 , n590982 );
and ( n63661 , n585586 , n54532 );
and ( n590985 , n58246 , n54530 );
nor ( n590986 , n63661 , n590985 );
xnor ( n63664 , n590986 , n53769 );
and ( n590988 , n590983 , n63664 );
xor ( n590989 , n590957 , n590961 );
xor ( n63667 , n590989 , n63641 );
and ( n590991 , n63664 , n63667 );
and ( n590992 , n590983 , n63667 );
or ( n63670 , n590988 , n590991 , n590992 );
xor ( n63671 , n590927 , n63606 );
xor ( n590995 , n63671 , n63644 );
and ( n590996 , n63670 , n590995 );
and ( n63674 , n58219 , n55013 );
and ( n63675 , n585221 , n55010 );
nor ( n590999 , n63674 , n63675 );
xnor ( n591000 , n590999 , n53762 );
and ( n63678 , n58246 , n55013 );
and ( n591002 , n58219 , n55010 );
nor ( n591003 , n63678 , n591002 );
xnor ( n63681 , n591003 , n53762 );
and ( n591005 , n585909 , n54532 );
and ( n591006 , n585586 , n54530 );
nor ( n63684 , n591005 , n591006 );
xnor ( n63685 , n63684 , n53769 );
and ( n591009 , n63681 , n63685 );
and ( n591010 , n585586 , n55013 );
and ( n63688 , n58246 , n55010 );
nor ( n63689 , n591010 , n63688 );
xnor ( n591013 , n63689 , n53762 );
and ( n591014 , n58623 , n54532 );
and ( n63692 , n585909 , n54530 );
nor ( n591016 , n591014 , n63692 );
xnor ( n591017 , n591016 , n53769 );
and ( n63695 , n591013 , n591017 );
and ( n591019 , n585973 , n54530 );
nor ( n591020 , n54532 , n591019 );
xnor ( n63698 , n591020 , n53769 );
nor ( n591022 , n53996 , n53994 );
xnor ( n63700 , n591022 , n53376 );
and ( n591024 , n63698 , n63700 );
and ( n591025 , n63700 , n53466 );
and ( n63703 , n63698 , n53466 );
or ( n591027 , n591024 , n591025 , n63703 );
nor ( n591028 , n53468 , n53466 );
xnor ( n63706 , n591028 , n52945 );
and ( n591030 , n591027 , n63706 );
and ( n591031 , n591017 , n591030 );
and ( n63709 , n591013 , n591030 );
or ( n591033 , n63695 , n591031 , n63709 );
and ( n591034 , n63685 , n591033 );
and ( n591035 , n63681 , n591033 );
or ( n591036 , n591009 , n591034 , n591035 );
and ( n63714 , n591000 , n591036 );
xor ( n591038 , n590983 , n63664 );
xor ( n591039 , n591038 , n63667 );
and ( n63717 , n591036 , n591039 );
and ( n591041 , n591000 , n591039 );
or ( n591042 , n63714 , n63717 , n591041 );
and ( n63720 , n590995 , n591042 );
and ( n591044 , n63670 , n591042 );
or ( n591045 , n590996 , n63720 , n591044 );
and ( n63723 , n63647 , n591045 );
and ( n63724 , n63586 , n591045 );
or ( n63725 , n63648 , n63723 , n63724 );
and ( n591049 , n590907 , n63725 );
xor ( n591050 , n590907 , n63725 );
xor ( n63728 , n63586 , n63647 );
xor ( n63729 , n63728 , n591045 );
xor ( n591053 , n590943 , n63622 );
nor ( n591054 , n53683 , n53681 );
xnor ( n63732 , n591054 , n53118 );
and ( n63733 , n591053 , n63732 );
and ( n591057 , n53467 , n52945 );
and ( n591058 , n63732 , n591057 );
and ( n63736 , n591053 , n591057 );
or ( n591060 , n63733 , n591058 , n63736 );
xor ( n591061 , n590934 , n590936 );
xor ( n63739 , n591061 , n53175 );
and ( n591063 , n591060 , n63739 );
xor ( n591064 , n63623 , n590948 );
xor ( n591065 , n591064 , n590951 );
and ( n591066 , n63739 , n591065 );
and ( n63744 , n591060 , n591065 );
or ( n591068 , n591063 , n591066 , n63744 );
xor ( n591069 , n63652 , n63654 );
xor ( n63747 , n591069 , n63657 );
and ( n591071 , n591068 , n63747 );
xor ( n63749 , n591060 , n63739 );
xor ( n63750 , n63749 , n591065 );
and ( n591074 , n585973 , n54532 );
and ( n63752 , n58623 , n54530 );
nor ( n63753 , n591074 , n63752 );
xnor ( n591077 , n63753 , n53769 );
xor ( n591078 , n591053 , n63732 );
xor ( n63756 , n591078 , n591057 );
and ( n591080 , n591077 , n63756 );
and ( n591081 , n63750 , n591080 );
and ( n63759 , n585909 , n55013 );
and ( n591083 , n585586 , n55010 );
nor ( n591084 , n63759 , n591083 );
xnor ( n63762 , n591084 , n53762 );
and ( n591086 , n58623 , n55013 );
and ( n591087 , n585909 , n55010 );
nor ( n63765 , n591086 , n591087 );
xnor ( n63766 , n63765 , n53762 );
nor ( n591090 , n54414 , n54412 );
xnor ( n63768 , n591090 , n53650 );
and ( n591092 , n63766 , n63768 );
nor ( n591093 , n53683 , n53681 );
xnor ( n591094 , n591093 , n53118 );
and ( n63772 , n63768 , n591094 );
and ( n591096 , n63766 , n591094 );
or ( n591097 , n591092 , n63772 , n591096 );
and ( n63775 , n63762 , n591097 );
xor ( n591099 , n591027 , n63706 );
and ( n591100 , n591097 , n591099 );
and ( n63778 , n63762 , n591099 );
or ( n591102 , n63775 , n591100 , n63778 );
and ( n591103 , n591080 , n591102 );
and ( n63781 , n63750 , n591102 );
or ( n591105 , n591081 , n591103 , n63781 );
xor ( n591106 , n63681 , n63685 );
xor ( n63784 , n591106 , n591033 );
and ( n63785 , n591105 , n63784 );
xor ( n591109 , n591068 , n63747 );
and ( n591110 , n63784 , n591109 );
and ( n63788 , n591105 , n591109 );
or ( n591112 , n63785 , n591110 , n63788 );
and ( n591113 , n591071 , n591112 );
xor ( n591114 , n591000 , n591036 );
xor ( n591115 , n591114 , n591039 );
and ( n63793 , n591112 , n591115 );
and ( n591117 , n591071 , n591115 );
or ( n591118 , n591113 , n63793 , n591117 );
xor ( n63796 , n63670 , n590995 );
xor ( n591120 , n63796 , n591042 );
and ( n63798 , n591118 , n591120 );
xor ( n591122 , n591118 , n591120 );
xor ( n63800 , n591071 , n591112 );
xor ( n63801 , n63800 , n591115 );
xor ( n591125 , n591013 , n591017 );
xor ( n591126 , n591125 , n591030 );
xor ( n63804 , n63698 , n63700 );
xor ( n591128 , n63804 , n53466 );
nor ( n591129 , n54532 , n54530 );
xnor ( n63807 , n591129 , n53769 );
nor ( n591131 , n54414 , n54412 );
xnor ( n591132 , n591131 , n53650 );
and ( n63810 , n63807 , n591132 );
nor ( n591134 , n53996 , n53994 );
xnor ( n591135 , n591134 , n53376 );
and ( n591136 , n591132 , n591135 );
and ( n591137 , n63807 , n591135 );
or ( n63815 , n63810 , n591136 , n591137 );
and ( n591139 , n591128 , n63815 );
and ( n591140 , n585973 , n55013 );
and ( n63818 , n58623 , n55010 );
nor ( n591142 , n591140 , n63818 );
xnor ( n63820 , n591142 , n53762 );
nor ( n591144 , n53683 , n53681 );
xnor ( n63822 , n591144 , n53118 );
and ( n63823 , n63820 , n63822 );
and ( n591147 , n53682 , n53118 );
and ( n591148 , n63822 , n591147 );
and ( n63826 , n63820 , n591147 );
or ( n63827 , n63823 , n591148 , n63826 );
and ( n591151 , n63815 , n63827 );
and ( n591152 , n591128 , n63827 );
or ( n63830 , n591139 , n591151 , n591152 );
xor ( n63831 , n591077 , n63756 );
and ( n63832 , n63830 , n63831 );
xor ( n591156 , n63766 , n63768 );
xor ( n591157 , n591156 , n591094 );
xor ( n63835 , n63807 , n591132 );
xor ( n591159 , n63835 , n591135 );
nor ( n591160 , n54532 , n54530 );
xnor ( n591161 , n591160 , n53769 );
nor ( n63839 , n54414 , n54412 );
xnor ( n591163 , n63839 , n53650 );
and ( n63841 , n591161 , n591163 );
nor ( n591165 , n53996 , n53994 );
xnor ( n591166 , n591165 , n53376 );
and ( n63844 , n591163 , n591166 );
and ( n591168 , n591161 , n591166 );
or ( n591169 , n63841 , n63844 , n591168 );
and ( n63847 , n591159 , n591169 );
and ( n591171 , n585973 , n55010 );
nor ( n591172 , n55013 , n591171 );
xnor ( n63850 , n591172 , n53762 );
and ( n591174 , n63850 , n53681 );
and ( n63852 , n591169 , n591174 );
and ( n591176 , n591159 , n591174 );
or ( n591177 , n63847 , n63852 , n591176 );
and ( n591178 , n591157 , n591177 );
xor ( n591179 , n591128 , n63815 );
xor ( n63857 , n591179 , n63827 );
and ( n591181 , n591177 , n63857 );
and ( n63859 , n591157 , n63857 );
or ( n591183 , n591178 , n591181 , n63859 );
and ( n591184 , n63831 , n591183 );
and ( n63862 , n63830 , n591183 );
or ( n63863 , n63832 , n591184 , n63862 );
and ( n63864 , n591126 , n63863 );
xor ( n63865 , n63750 , n591080 );
xor ( n591189 , n63865 , n591102 );
and ( n63867 , n63863 , n591189 );
and ( n63868 , n591126 , n591189 );
or ( n591192 , n63864 , n63867 , n63868 );
xor ( n591193 , n591105 , n63784 );
xor ( n63871 , n591193 , n591109 );
and ( n591195 , n591192 , n63871 );
xor ( n63873 , n591192 , n63871 );
xor ( n591197 , n591126 , n63863 );
xor ( n63875 , n591197 , n591189 );
xor ( n63876 , n63762 , n591097 );
xor ( n591200 , n63876 , n591099 );
xor ( n591201 , n63830 , n63831 );
xor ( n63879 , n591201 , n591183 );
and ( n63880 , n591200 , n63879 );
xor ( n591204 , n591200 , n63879 );
xor ( n63882 , n63820 , n63822 );
xor ( n63883 , n63882 , n591147 );
xor ( n63884 , n591161 , n591163 );
xor ( n63885 , n63884 , n591166 );
xor ( n63886 , n63850 , n53681 );
and ( n63887 , n63885 , n63886 );
nor ( n591211 , n54532 , n54530 );
xnor ( n63889 , n591211 , n53769 );
nor ( n591213 , n54414 , n54412 );
xnor ( n63891 , n591213 , n53650 );
and ( n591215 , n63889 , n63891 );
nor ( n591216 , n53996 , n53994 );
xnor ( n63894 , n591216 , n53376 );
and ( n591218 , n63891 , n63894 );
and ( n63896 , n63889 , n63894 );
or ( n63897 , n591215 , n591218 , n63896 );
and ( n63898 , n63886 , n63897 );
and ( n63899 , n63885 , n63897 );
or ( n63900 , n63887 , n63898 , n63899 );
and ( n63901 , n63883 , n63900 );
xor ( n63902 , n591159 , n591169 );
xor ( n63903 , n63902 , n591174 );
and ( n591227 , n63900 , n63903 );
and ( n63905 , n63883 , n63903 );
or ( n591229 , n63901 , n591227 , n63905 );
xor ( n591230 , n591157 , n591177 );
xor ( n63908 , n591230 , n63857 );
and ( n63909 , n591229 , n63908 );
xor ( n591233 , n591229 , n63908 );
nor ( n591234 , n55013 , n55010 );
xnor ( n591235 , n591234 , n53762 );
and ( n63913 , n53995 , n53376 );
and ( n591237 , n591235 , n63913 );
xor ( n63915 , n591235 , n63913 );
nor ( n591239 , n55013 , n55010 );
xnor ( n591240 , n591239 , n53762 );
nor ( n63918 , n54532 , n54530 );
xnor ( n63919 , n63918 , n53769 );
and ( n63920 , n591240 , n63919 );
and ( n63921 , n63919 , n53994 );
and ( n591245 , n591240 , n53994 );
or ( n591246 , n63920 , n63921 , n591245 );
and ( n591247 , n63915 , n591246 );
xor ( n63925 , n63889 , n63891 );
xor ( n591249 , n63925 , n63894 );
and ( n591250 , n591246 , n591249 );
and ( n591251 , n63915 , n591249 );
or ( n63929 , n591247 , n591250 , n591251 );
and ( n591253 , n591237 , n63929 );
xor ( n591254 , n63885 , n63886 );
xor ( n63932 , n591254 , n63897 );
and ( n591256 , n63929 , n63932 );
and ( n63934 , n591237 , n63932 );
or ( n63935 , n591253 , n591256 , n63934 );
xor ( n591259 , n63883 , n63900 );
xor ( n63937 , n591259 , n63903 );
and ( n63938 , n63935 , n63937 );
xor ( n591262 , n63935 , n63937 );
xor ( n591263 , n591237 , n63929 );
xor ( n63941 , n591263 , n63932 );
xor ( n63942 , n63915 , n591246 );
xor ( n63943 , n63942 , n591249 );
nor ( n63944 , n55013 , n55010 );
xnor ( n63945 , n63944 , n53762 );
and ( n591269 , n54413 , n53650 );
and ( n63947 , n63945 , n591269 );
nor ( n591271 , n54414 , n54412 );
xnor ( n591272 , n591271 , n53650 );
and ( n591273 , n63947 , n591272 );
xor ( n63951 , n591240 , n63919 );
xor ( n591275 , n63951 , n53994 );
and ( n591276 , n591272 , n591275 );
and ( n591277 , n63947 , n591275 );
or ( n63955 , n591273 , n591276 , n591277 );
and ( n591279 , n63943 , n63955 );
xor ( n591280 , n63943 , n63955 );
xor ( n63958 , n63947 , n591272 );
xor ( n591282 , n63958 , n591275 );
xor ( n63960 , n63945 , n591269 );
nor ( n63961 , n54532 , n54530 );
xnor ( n591285 , n63961 , n53769 );
and ( n591286 , n63960 , n591285 );
nor ( n591287 , n54414 , n54412 );
xnor ( n63965 , n591287 , n53650 );
and ( n591289 , n591285 , n63965 );
and ( n591290 , n63960 , n63965 );
or ( n591291 , n591286 , n591289 , n591290 );
and ( n591292 , n591282 , n591291 );
xor ( n63970 , n591282 , n591291 );
nor ( n591294 , n55013 , n55010 );
xnor ( n591295 , n591294 , n53762 );
nor ( n63973 , n54532 , n54530 );
xnor ( n63974 , n63973 , n53769 );
and ( n591298 , n591295 , n63974 );
and ( n63976 , n63974 , n54412 );
and ( n63977 , n591295 , n54412 );
or ( n63978 , n591298 , n63976 , n63977 );
xor ( n591302 , n63960 , n591285 );
xor ( n591303 , n591302 , n63965 );
and ( n63981 , n63978 , n591303 );
xor ( n591305 , n63978 , n591303 );
xor ( n63983 , n591295 , n63974 );
xor ( n591307 , n63983 , n54412 );
nor ( n63985 , n55013 , n55010 );
xnor ( n63986 , n63985 , n53762 );
and ( n591310 , n54531 , n53769 );
and ( n591311 , n63986 , n591310 );
and ( n63989 , n591307 , n591311 );
xor ( n63990 , n591307 , n591311 );
nor ( n591314 , n54532 , n54530 );
xnor ( n591315 , n591314 , n53769 );
xor ( n63993 , n63986 , n591310 );
and ( n591317 , n591315 , n63993 );
xor ( n63995 , n591315 , n63993 );
nor ( n63996 , n55013 , n55010 );
xnor ( n591320 , n63996 , n53762 );
and ( n591321 , n591320 , n54530 );
xor ( n63999 , n591320 , n54530 );
nor ( n64000 , n55013 , n55010 );
xnor ( n591324 , n64000 , n53762 );
and ( n591325 , n55012 , n53762 );
and ( n64003 , n591324 , n591325 );
and ( n591327 , n63999 , n64003 );
or ( n591328 , n591321 , n591327 );
and ( n64006 , n63995 , n591328 );
or ( n64007 , n591317 , n64006 );
and ( n64008 , n63990 , n64007 );
or ( n64009 , n63989 , n64008 );
and ( n64010 , n591305 , n64009 );
or ( n64011 , n63981 , n64010 );
and ( n64012 , n63970 , n64011 );
or ( n64013 , n591292 , n64012 );
and ( n64014 , n591280 , n64013 );
or ( n64015 , n591279 , n64014 );
and ( n591339 , n63941 , n64015 );
and ( n591340 , n591262 , n591339 );
or ( n64018 , n63938 , n591340 );
and ( n591342 , n591233 , n64018 );
or ( n64020 , n63909 , n591342 );
and ( n591344 , n591204 , n64020 );
or ( n591345 , n63880 , n591344 );
and ( n64023 , n63875 , n591345 );
and ( n64024 , n63873 , n64023 );
or ( n64025 , n591195 , n64024 );
and ( n64026 , n63801 , n64025 );
and ( n591350 , n591122 , n64026 );
or ( n591351 , n63798 , n591350 );
and ( n591352 , n63729 , n591351 );
and ( n64030 , n591050 , n591352 );
or ( n591354 , n591049 , n64030 );
and ( n591355 , n63582 , n591354 );
or ( n64033 , n590904 , n591355 );
and ( n591357 , n590866 , n64033 );
and ( n591358 , n63541 , n591357 );
or ( n64036 , n590863 , n591358 );
and ( n591360 , n590746 , n64036 );
or ( n64038 , n590745 , n591360 );
and ( n591362 , n63354 , n64038 );
or ( n591363 , n63353 , n591362 );
and ( n591364 , n590591 , n591363 );
or ( n591365 , n63267 , n591364 );
and ( n64043 , n63262 , n591365 );
and ( n591367 , n63260 , n64043 );
or ( n64045 , n63259 , n591367 );
and ( n591369 , n63021 , n64045 );
or ( n591370 , n63020 , n591369 );
and ( n64048 , n590293 , n591370 );
or ( n64049 , n62969 , n64048 );
and ( n64050 , n590202 , n64049 );
or ( n64051 , n62878 , n64050 );
and ( n591375 , n62772 , n64051 );
and ( n591376 , n590093 , n591375 );
or ( n591377 , n62769 , n591376 );
and ( n591378 , n62641 , n591377 );
and ( n591379 , n62639 , n591378 );
or ( n64057 , n62638 , n591379 );
and ( n64058 , n62310 , n64057 );
and ( n64059 , n62308 , n64058 );
or ( n64060 , n62307 , n64059 );
and ( n64061 , n62303 , n64060 );
or ( n591385 , n62302 , n64061 );
and ( n591386 , n589301 , n591385 );
or ( n591387 , n61977 , n591386 );
and ( n64065 , n589296 , n591387 );
and ( n591389 , n589294 , n64065 );
and ( n64067 , n61969 , n591389 );
or ( n591391 , n61968 , n64067 );
and ( n64069 , n589272 , n591391 );
and ( n64070 , n589270 , n64069 );
and ( n591394 , n61945 , n64070 );
and ( n64072 , n589266 , n591394 );
and ( n591396 , n589264 , n64072 );
and ( n591397 , n61939 , n591396 );
and ( n64075 , n589260 , n591397 );
and ( n591399 , n589258 , n64075 );
and ( n591400 , n589256 , n591399 );
and ( n64078 , n61931 , n591400 );
and ( n591402 , n589252 , n64078 );
and ( n64080 , n589250 , n591402 );
and ( n591404 , n589248 , n64080 );
and ( n591405 , n589246 , n591404 );
and ( n64083 , n61921 , n591405 );
and ( n591407 , n61919 , n64083 );
and ( n591408 , n61917 , n591407 );
and ( n64086 , n61915 , n591408 );
and ( n64087 , n589236 , n64086 );
and ( n591411 , n61911 , n64087 );
and ( n591412 , n589232 , n591411 );
and ( n64090 , n61907 , n591412 );
and ( n64091 , n589228 , n64090 );
and ( n591415 , n61903 , n64091 );
and ( n591416 , n589224 , n591415 );
and ( n64094 , n61899 , n591416 );
and ( n64095 , n61897 , n64094 );
and ( n591419 , n589218 , n64095 );
and ( n591420 , n589216 , n591419 );
and ( n64098 , n61891 , n591420 );
and ( n64099 , n589212 , n64098 );
and ( n591423 , n61887 , n64099 );
and ( n591424 , n61885 , n591423 );
and ( n64102 , n589206 , n591424 );
and ( n591426 , n61881 , n64102 );
and ( n591427 , n589202 , n591426 );
and ( n591428 , n589200 , n591427 );
and ( n64106 , n589198 , n591428 );
and ( n591430 , n61873 , n64106 );
and ( n591431 , n589194 , n591430 );
and ( n591432 , n589192 , n591431 );
and ( n591433 , n61867 , n591432 );
and ( n64111 , n589188 , n591433 );
and ( n591435 , n61863 , n64111 );
and ( n591436 , n589184 , n591435 );
and ( n64114 , n61859 , n591436 );
and ( n591438 , n589180 , n64114 );
and ( n591439 , n589178 , n591438 );
and ( n64117 , n589176 , n591439 );
and ( n64118 , n61851 , n64117 );
and ( n591442 , n589172 , n64118 );
and ( n64120 , n61847 , n591442 );
and ( n64121 , n589168 , n64120 );
and ( n64122 , n61843 , n64121 );
and ( n64123 , n589164 , n64122 );
and ( n591447 , n61839 , n64123 );
and ( n64125 , n61837 , n591447 );
and ( n591449 , n61835 , n64125 );
and ( n591450 , n61833 , n591449 );
and ( n591451 , n589154 , n591450 );
and ( n64129 , n61829 , n591451 );
and ( n591453 , n589150 , n64129 );
and ( n591454 , n61825 , n591453 );
and ( n591455 , n589146 , n591454 );
and ( n591456 , n61821 , n591455 );
xor ( n64134 , n589142 , n591456 );
buf ( n591458 , n64134 );
xor ( n591459 , n61821 , n591455 );
buf ( n591460 , n591459 );
xor ( n591461 , n589146 , n591454 );
buf ( n591462 , n591461 );
xor ( n64140 , n61825 , n591453 );
buf ( n591464 , n64140 );
xor ( n591465 , n589150 , n64129 );
buf ( n591466 , n591465 );
xor ( n591467 , n61829 , n591451 );
buf ( n591468 , n591467 );
xor ( n64146 , n589154 , n591450 );
buf ( n591470 , n64146 );
xor ( n591471 , n61833 , n591449 );
buf ( n591472 , n591471 );
xor ( n64150 , n61835 , n64125 );
buf ( n591474 , n64150 );
xor ( n591475 , n61837 , n591447 );
buf ( n591476 , n591475 );
xor ( n591477 , n61839 , n64123 );
buf ( n591478 , n591477 );
xor ( n64156 , n589164 , n64122 );
buf ( n591480 , n64156 );
xor ( n591481 , n61843 , n64121 );
buf ( n591482 , n591481 );
xor ( n64160 , n589168 , n64120 );
buf ( n591484 , n64160 );
xor ( n591485 , n61847 , n591442 );
buf ( n591486 , n591485 );
xor ( n64164 , n589172 , n64118 );
buf ( n591488 , n64164 );
xor ( n591489 , n61851 , n64117 );
buf ( n591490 , n591489 );
xor ( n591491 , n589176 , n591439 );
buf ( n591492 , n591491 );
xor ( n64170 , n589178 , n591438 );
buf ( n591494 , n64170 );
xor ( n64172 , n589180 , n64114 );
buf ( n591496 , n64172 );
xor ( n64174 , n61859 , n591436 );
buf ( n591498 , n64174 );
xor ( n591499 , n589184 , n591435 );
buf ( n591500 , n591499 );
xor ( n64178 , n61863 , n64111 );
buf ( n591502 , n64178 );
xor ( n591503 , n589188 , n591433 );
buf ( n591504 , n591503 );
xor ( n591505 , n61867 , n591432 );
buf ( n591506 , n591505 );
xor ( n64184 , n589192 , n591431 );
buf ( n591508 , n64184 );
xor ( n591509 , n589194 , n591430 );
buf ( n591510 , n591509 );
xor ( n591511 , n61873 , n64106 );
buf ( n591512 , n591511 );
xor ( n591513 , n589198 , n591428 );
buf ( n591514 , n591513 );
xor ( n591515 , n589200 , n591427 );
buf ( n591516 , n591515 );
xor ( n64194 , n589202 , n591426 );
buf ( n591518 , n64194 );
xor ( n591519 , n61881 , n64102 );
buf ( n591520 , n591519 );
xor ( n64198 , n589206 , n591424 );
buf ( n591522 , n64198 );
xor ( n591523 , n61885 , n591423 );
buf ( n591524 , n591523 );
xor ( n64202 , n61887 , n64099 );
buf ( n591526 , n64202 );
xor ( n591527 , n589212 , n64098 );
buf ( n591528 , n591527 );
xor ( n64206 , n61891 , n591420 );
buf ( n591530 , n64206 );
xor ( n64208 , n589216 , n591419 );
buf ( n591532 , n64208 );
xor ( n64210 , n589218 , n64095 );
buf ( n591534 , n64210 );
xor ( n591535 , n61897 , n64094 );
buf ( n591536 , n591535 );
xor ( n64214 , n61899 , n591416 );
buf ( n591538 , n64214 );
xor ( n64216 , n589224 , n591415 );
buf ( n591540 , n64216 );
xor ( n64218 , n61903 , n64091 );
buf ( n591542 , n64218 );
xor ( n64220 , n589228 , n64090 );
buf ( n591544 , n64220 );
xor ( n591545 , n61907 , n591412 );
buf ( n591546 , n591545 );
xor ( n64224 , n589232 , n591411 );
buf ( n591548 , n64224 );
xor ( n64226 , n61911 , n64087 );
buf ( n591550 , n64226 );
xor ( n591551 , n589236 , n64086 );
buf ( n591552 , n591551 );
xor ( n591553 , n61915 , n591408 );
buf ( n591554 , n591553 );
xor ( n591555 , n61917 , n591407 );
buf ( n591556 , n591555 );
xor ( n64234 , n61919 , n64083 );
buf ( n591558 , n64234 );
xor ( n591559 , n61921 , n591405 );
buf ( n591560 , n591559 );
xor ( n64238 , n589246 , n591404 );
buf ( n591562 , n64238 );
xor ( n64240 , n589248 , n64080 );
buf ( n591564 , n64240 );
xor ( n64242 , n589250 , n591402 );
buf ( n591566 , n64242 );
xor ( n591567 , n589252 , n64078 );
buf ( n591568 , n591567 );
xor ( n64246 , n61931 , n591400 );
buf ( n591570 , n64246 );
xor ( n64248 , n589256 , n591399 );
buf ( n591572 , n64248 );
xor ( n591573 , n589258 , n64075 );
buf ( n591574 , n591573 );
xor ( n591575 , n589260 , n591397 );
buf ( n591576 , n591575 );
xor ( n591577 , n61939 , n591396 );
buf ( n591578 , n591577 );
xor ( n591579 , n589264 , n64072 );
buf ( n591580 , n591579 );
xor ( n64258 , n589266 , n591394 );
buf ( n591582 , n64258 );
xor ( n64260 , n61945 , n64070 );
buf ( n591584 , n64260 );
xor ( n591585 , n589270 , n64069 );
buf ( n591586 , n591585 );
xor ( n591587 , n589272 , n591391 );
buf ( n591588 , n591587 );
xor ( n64266 , n61969 , n591389 );
buf ( n591590 , n64266 );
xor ( n591591 , n589294 , n64065 );
buf ( n591592 , n591591 );
xor ( n64270 , n589296 , n591387 );
buf ( n591594 , n64270 );
xor ( n64272 , n589301 , n591385 );
buf ( n591596 , n64272 );
xor ( n591597 , n62303 , n64060 );
buf ( n591598 , n591597 );
xor ( n64276 , n62308 , n64058 );
buf ( n591600 , n64276 );
xor ( n591601 , n62310 , n64057 );
buf ( n591602 , n591601 );
xor ( n64280 , n62639 , n591378 );
buf ( n591604 , n64280 );
xor ( n64282 , n62641 , n591377 );
buf ( n591606 , n64282 );
xor ( n64284 , n590093 , n591375 );
buf ( n591608 , n64284 );
xor ( n591609 , n62772 , n64051 );
buf ( n591610 , n591609 );
xor ( n591611 , n590202 , n64049 );
buf ( n591612 , n591611 );
xor ( n591613 , n590293 , n591370 );
buf ( n591614 , n591613 );
xor ( n591615 , n63021 , n64045 );
buf ( n591616 , n591615 );
xor ( n591617 , n63260 , n64043 );
buf ( n591618 , n591617 );
xor ( n64296 , n63262 , n591365 );
buf ( n591620 , n64296 );
xor ( n591621 , n590591 , n591363 );
buf ( n591622 , n591621 );
xor ( n64300 , n63354 , n64038 );
buf ( n591624 , n64300 );
xor ( n591625 , n590746 , n64036 );
buf ( n591626 , n591625 );
xor ( n591627 , n63541 , n591357 );
buf ( n591628 , n591627 );
xor ( n591629 , n590866 , n64033 );
buf ( n591630 , n591629 );
xor ( n64308 , n63582 , n591354 );
buf ( n591632 , n64308 );
xor ( n64310 , n591050 , n591352 );
buf ( n591634 , n64310 );
xor ( n591635 , n63729 , n591351 );
buf ( n591636 , n591635 );
xor ( n591637 , n591122 , n64026 );
buf ( n591638 , n591637 );
xor ( n591639 , n63801 , n64025 );
buf ( n591640 , n591639 );
xor ( n591641 , n63873 , n64023 );
buf ( n591642 , n591641 );
xor ( n591643 , n63875 , n591345 );
buf ( n591644 , n591643 );
xor ( n591645 , n591204 , n64020 );
buf ( n591646 , n591645 );
xor ( n591647 , n591233 , n64018 );
buf ( n591648 , n591647 );
xor ( n591649 , n591262 , n591339 );
buf ( n591650 , n591649 );
xor ( n591651 , n63941 , n64015 );
buf ( n591652 , n591651 );
xor ( n591653 , n591280 , n64013 );
buf ( n591654 , n591653 );
xor ( n591655 , n63970 , n64011 );
buf ( n591656 , n591655 );
xor ( n591657 , n591305 , n64009 );
buf ( n591658 , n591657 );
xor ( n591659 , n63990 , n64007 );
buf ( n591660 , n591659 );
xor ( n591661 , n63995 , n591328 );
buf ( n591662 , n591661 );
xor ( n591663 , n63999 , n64003 );
buf ( n591664 , n591663 );
xor ( n591665 , n591324 , n591325 );
buf ( n591666 , n591665 );
buf ( n591667 , n55010 );
buf ( n591668 , n591667 );
buf ( n591669 , n557576 );
buf ( n591670 , n557579 );
buf ( n591671 , n557582 );
buf ( n591672 , n557585 );
buf ( n591673 , n557588 );
buf ( n591674 , n557591 );
buf ( n591675 , n557594 );
buf ( n591676 , n557597 );
buf ( n591677 , n557600 );
buf ( n591678 , n557603 );
buf ( n591679 , n557606 );
buf ( n591680 , n557609 );
buf ( n591681 , n557612 );
buf ( n591682 , n557615 );
buf ( n591683 , n557618 );
buf ( n591684 , n557621 );
buf ( n591685 , n557624 );
buf ( n591686 , n557627 );
buf ( n591687 , n557630 );
buf ( n591688 , n557633 );
buf ( n591689 , n557636 );
buf ( n591690 , n557639 );
buf ( n591691 , n557642 );
buf ( n591692 , n557645 );
buf ( n591693 , n557648 );
buf ( n591694 , n557651 );
buf ( n591695 , n557654 );
buf ( n591696 , n557657 );
buf ( n591697 , n557660 );
buf ( n591698 , n557663 );
buf ( n591699 , n557666 );
buf ( n591700 , n557669 );
buf ( n591701 , n557672 );
buf ( n591702 , n557675 );
buf ( n591703 , n557678 );
buf ( n591704 , n557681 );
buf ( n591705 , n557684 );
buf ( n591706 , n557687 );
buf ( n591707 , n557690 );
buf ( n591708 , n557693 );
buf ( n591709 , n557696 );
buf ( n591710 , n557699 );
buf ( n591711 , n557702 );
buf ( n591712 , n557705 );
buf ( n591713 , n557708 );
buf ( n591714 , n557711 );
buf ( n591715 , n557714 );
buf ( n591716 , n557717 );
buf ( n591717 , n557720 );
buf ( n591718 , n557723 );
buf ( n591719 , n557726 );
buf ( n591720 , n557729 );
buf ( n591721 , n557732 );
buf ( n591722 , n557735 );
buf ( n591723 , n557738 );
buf ( n591724 , n557741 );
buf ( n591725 , n557744 );
buf ( n591726 , n557747 );
buf ( n591727 , n557750 );
buf ( n591728 , n557753 );
buf ( n591729 , n557756 );
buf ( n591730 , n557759 );
buf ( n591731 , n557762 );
buf ( n591732 , n557765 );
buf ( n591733 , n557767 );
buf ( n591734 , n1186 );
buf ( n591735 , n1187 );
buf ( n591736 , n1188 );
buf ( n591737 , n1189 );
buf ( n591738 , n1190 );
buf ( n591739 , n1191 );
buf ( n591740 , n1192 );
buf ( n591741 , n1193 );
buf ( n591742 , n1194 );
buf ( n591743 , n1195 );
buf ( n591744 , n1196 );
buf ( n591745 , n1197 );
buf ( n591746 , n1198 );
buf ( n591747 , n1199 );
buf ( n591748 , n1200 );
buf ( n591749 , n1201 );
buf ( n591750 , n1202 );
buf ( n591751 , n1203 );
buf ( n591752 , n1204 );
buf ( n591753 , n1205 );
buf ( n591754 , n1206 );
buf ( n591755 , n1207 );
buf ( n591756 , n1208 );
buf ( n591757 , n1209 );
buf ( n591758 , n1210 );
buf ( n591759 , n1211 );
buf ( n591760 , n1212 );
buf ( n591761 , n1213 );
buf ( n591762 , n1214 );
buf ( n591763 , n1215 );
buf ( n591764 , n1216 );
buf ( n591765 , n1217 );
buf ( n64443 , n591736 );
buf ( n64444 , n591737 );
buf ( n64445 , n591738 );
and ( n64446 , n64444 , n64445 );
not ( n64447 , n64446 );
and ( n64448 , n64443 , n64447 );
not ( n64449 , n64448 );
buf ( n64450 , n591670 );
buf ( n64451 , n591734 );
buf ( n64452 , n591735 );
xor ( n64453 , n64451 , n64452 );
xor ( n64454 , n64452 , n64443 );
not ( n64455 , n64454 );
and ( n64456 , n64453 , n64455 );
and ( n64457 , n64450 , n64456 );
buf ( n64458 , n591669 );
and ( n64459 , n64458 , n64454 );
nor ( n591783 , n64457 , n64459 );
and ( n64461 , n64452 , n64443 );
not ( n591785 , n64461 );
and ( n591786 , n64451 , n591785 );
xnor ( n64464 , n591783 , n591786 );
and ( n64465 , n64449 , n64464 );
buf ( n64466 , n591671 );
and ( n64467 , n64466 , n64451 );
and ( n591791 , n64464 , n64467 );
and ( n64469 , n64449 , n64467 );
or ( n64470 , n64465 , n591791 , n64469 );
and ( n64471 , n64458 , n64456 );
not ( n64472 , n64471 );
xnor ( n591796 , n64472 , n591786 );
not ( n64474 , n591796 );
and ( n64475 , n64470 , n64474 );
and ( n64476 , n64450 , n64451 );
and ( n64477 , n64474 , n64476 );
and ( n64478 , n64470 , n64476 );
or ( n64479 , n64475 , n64477 , n64478 );
buf ( n591803 , n591796 );
not ( n64481 , n591786 );
xor ( n591805 , n591803 , n64481 );
and ( n64483 , n64458 , n64451 );
xor ( n64484 , n591805 , n64483 );
xor ( n64485 , n64479 , n64484 );
xor ( n64486 , n64470 , n64474 );
xor ( n64487 , n64486 , n64476 );
xor ( n64488 , n64443 , n64444 );
xor ( n64489 , n64444 , n64445 );
not ( n64490 , n64489 );
and ( n64491 , n64488 , n64490 );
and ( n64492 , n64458 , n64491 );
not ( n64493 , n64492 );
xnor ( n64494 , n64493 , n64448 );
not ( n64495 , n64494 );
and ( n591819 , n64466 , n64456 );
and ( n64497 , n64450 , n64454 );
nor ( n64498 , n591819 , n64497 );
xnor ( n64499 , n64498 , n591786 );
and ( n64500 , n64495 , n64499 );
buf ( n64501 , n591672 );
and ( n64502 , n64501 , n64451 );
and ( n591826 , n64499 , n64502 );
and ( n591827 , n64495 , n64502 );
or ( n64505 , n64500 , n591826 , n591827 );
buf ( n591829 , n64494 );
and ( n591830 , n64505 , n591829 );
xor ( n591831 , n64449 , n64464 );
xor ( n591832 , n591831 , n64467 );
and ( n64510 , n591829 , n591832 );
and ( n64511 , n64505 , n591832 );
or ( n64512 , n591830 , n64510 , n64511 );
and ( n64513 , n64487 , n64512 );
xor ( n64514 , n64487 , n64512 );
xor ( n591838 , n64505 , n591829 );
xor ( n64516 , n591838 , n591832 );
buf ( n591840 , n591739 );
buf ( n591841 , n591740 );
and ( n64519 , n591840 , n591841 );
not ( n64520 , n64519 );
and ( n64521 , n64445 , n64520 );
not ( n591845 , n64521 );
and ( n64523 , n64501 , n64456 );
and ( n591847 , n64466 , n64454 );
nor ( n64525 , n64523 , n591847 );
xnor ( n64526 , n64525 , n591786 );
and ( n64527 , n591845 , n64526 );
buf ( n591851 , n591673 );
and ( n64529 , n591851 , n64451 );
and ( n591853 , n64526 , n64529 );
and ( n591854 , n591845 , n64529 );
or ( n64532 , n64527 , n591853 , n591854 );
buf ( n64533 , n591674 );
and ( n64534 , n64533 , n64451 );
buf ( n64535 , n64534 );
and ( n64536 , n64450 , n64491 );
and ( n64537 , n64458 , n64489 );
nor ( n64538 , n64536 , n64537 );
xnor ( n64539 , n64538 , n64448 );
and ( n591863 , n64535 , n64539 );
xor ( n591864 , n591845 , n64526 );
xor ( n64542 , n591864 , n64529 );
and ( n64543 , n64539 , n64542 );
and ( n64544 , n64535 , n64542 );
or ( n64545 , n591863 , n64543 , n64544 );
and ( n64546 , n64532 , n64545 );
xor ( n64547 , n64495 , n64499 );
xor ( n64548 , n64547 , n64502 );
and ( n64549 , n64545 , n64548 );
and ( n64550 , n64532 , n64548 );
or ( n64551 , n64546 , n64549 , n64550 );
and ( n64552 , n64516 , n64551 );
xor ( n64553 , n64516 , n64551 );
xor ( n64554 , n64532 , n64545 );
xor ( n591878 , n64554 , n64548 );
xor ( n64556 , n64445 , n591840 );
xor ( n591880 , n591840 , n591841 );
not ( n591881 , n591880 );
and ( n64559 , n64556 , n591881 );
and ( n591883 , n64458 , n64559 );
not ( n591884 , n591883 );
xnor ( n64562 , n591884 , n64521 );
and ( n591886 , n64466 , n64491 );
and ( n64564 , n64450 , n64489 );
nor ( n64565 , n591886 , n64564 );
xnor ( n64566 , n64565 , n64448 );
and ( n591890 , n64562 , n64566 );
and ( n591891 , n591851 , n64456 );
and ( n64569 , n64501 , n64454 );
nor ( n591893 , n591891 , n64569 );
xnor ( n64571 , n591893 , n591786 );
and ( n64572 , n64566 , n64571 );
and ( n64573 , n64562 , n64571 );
or ( n64574 , n591890 , n64572 , n64573 );
buf ( n64575 , n591741 );
buf ( n64576 , n591742 );
and ( n591900 , n64575 , n64576 );
not ( n64578 , n591900 );
and ( n591902 , n591841 , n64578 );
not ( n591903 , n591902 );
and ( n64581 , n64533 , n64456 );
and ( n64582 , n591851 , n64454 );
nor ( n64583 , n64581 , n64582 );
xnor ( n64584 , n64583 , n591786 );
and ( n64585 , n591903 , n64584 );
buf ( n64586 , n591675 );
and ( n64587 , n64586 , n64451 );
and ( n64588 , n64584 , n64587 );
and ( n64589 , n591903 , n64587 );
or ( n64590 , n64585 , n64588 , n64589 );
buf ( n64591 , n591676 );
and ( n64592 , n64591 , n64451 );
buf ( n591916 , n64592 );
and ( n64594 , n64450 , n64559 );
and ( n591918 , n64458 , n591880 );
nor ( n591919 , n64594 , n591918 );
xnor ( n64597 , n591919 , n64521 );
and ( n591921 , n591916 , n64597 );
and ( n64599 , n64501 , n64491 );
and ( n64600 , n64466 , n64489 );
nor ( n64601 , n64599 , n64600 );
xnor ( n64602 , n64601 , n64448 );
and ( n64603 , n64597 , n64602 );
and ( n64604 , n591916 , n64602 );
or ( n64605 , n591921 , n64603 , n64604 );
and ( n64606 , n64590 , n64605 );
not ( n64607 , n64534 );
and ( n64608 , n64605 , n64607 );
and ( n64609 , n64590 , n64607 );
or ( n64610 , n64606 , n64608 , n64609 );
and ( n64611 , n64574 , n64610 );
xor ( n64612 , n64535 , n64539 );
xor ( n64613 , n64612 , n64542 );
and ( n64614 , n64610 , n64613 );
and ( n64615 , n64574 , n64613 );
or ( n64616 , n64611 , n64614 , n64615 );
and ( n64617 , n591878 , n64616 );
xor ( n64618 , n591878 , n64616 );
buf ( n64619 , n591743 );
buf ( n64620 , n591744 );
and ( n64621 , n64619 , n64620 );
not ( n64622 , n64621 );
and ( n64623 , n64576 , n64622 );
not ( n64624 , n64623 );
and ( n64625 , n64591 , n64456 );
and ( n64626 , n64586 , n64454 );
nor ( n64627 , n64625 , n64626 );
xnor ( n64628 , n64627 , n591786 );
and ( n64629 , n64624 , n64628 );
buf ( n64630 , n591677 );
and ( n64631 , n64630 , n64451 );
and ( n64632 , n64628 , n64631 );
and ( n64633 , n64624 , n64631 );
or ( n64634 , n64629 , n64632 , n64633 );
and ( n64635 , n64466 , n64559 );
and ( n64636 , n64450 , n591880 );
nor ( n64637 , n64635 , n64636 );
xnor ( n591961 , n64637 , n64521 );
and ( n64639 , n64634 , n591961 );
and ( n591963 , n591851 , n64491 );
and ( n591964 , n64501 , n64489 );
nor ( n64642 , n591963 , n591964 );
xnor ( n591966 , n64642 , n64448 );
and ( n591967 , n591961 , n591966 );
and ( n64645 , n64634 , n591966 );
or ( n591969 , n64639 , n591967 , n64645 );
xor ( n591970 , n591841 , n64575 );
xor ( n64648 , n64575 , n64576 );
not ( n64649 , n64648 );
and ( n64650 , n591970 , n64649 );
and ( n64651 , n64458 , n64650 );
not ( n591975 , n64651 );
xnor ( n591976 , n591975 , n591902 );
and ( n64654 , n64586 , n64456 );
and ( n64655 , n64533 , n64454 );
nor ( n64656 , n64654 , n64655 );
xnor ( n64657 , n64656 , n591786 );
and ( n591981 , n591976 , n64657 );
not ( n591982 , n64592 );
and ( n64660 , n64657 , n591982 );
and ( n64661 , n591976 , n591982 );
or ( n64662 , n591981 , n64660 , n64661 );
and ( n64663 , n591969 , n64662 );
xor ( n591987 , n591903 , n64584 );
xor ( n591988 , n591987 , n64587 );
and ( n64666 , n64662 , n591988 );
and ( n591990 , n591969 , n591988 );
or ( n64668 , n64663 , n64666 , n591990 );
xor ( n591992 , n64562 , n64566 );
xor ( n591993 , n591992 , n64571 );
and ( n64671 , n64668 , n591993 );
xor ( n591995 , n64590 , n64605 );
xor ( n591996 , n591995 , n64607 );
and ( n64674 , n591993 , n591996 );
and ( n591998 , n64668 , n591996 );
or ( n591999 , n64671 , n64674 , n591998 );
xor ( n592000 , n64574 , n64610 );
xor ( n592001 , n592000 , n64613 );
and ( n64679 , n591999 , n592001 );
xor ( n592003 , n591999 , n592001 );
xor ( n592004 , n64668 , n591993 );
xor ( n64682 , n592004 , n591996 );
buf ( n64683 , n591678 );
and ( n64684 , n64683 , n64451 );
buf ( n64685 , n64684 );
and ( n64686 , n64501 , n64559 );
and ( n592010 , n64466 , n591880 );
nor ( n64688 , n64686 , n592010 );
xnor ( n592012 , n64688 , n64521 );
and ( n592013 , n64685 , n592012 );
and ( n64691 , n64533 , n64491 );
and ( n592015 , n591851 , n64489 );
nor ( n592016 , n64691 , n592015 );
xnor ( n64694 , n592016 , n64448 );
and ( n592018 , n592012 , n64694 );
and ( n64696 , n64685 , n64694 );
or ( n64697 , n592013 , n592018 , n64696 );
xor ( n64698 , n64634 , n591961 );
xor ( n64699 , n64698 , n591966 );
and ( n592023 , n64697 , n64699 );
xor ( n592024 , n591976 , n64657 );
xor ( n64702 , n592024 , n591982 );
and ( n592026 , n64699 , n64702 );
and ( n64704 , n64697 , n64702 );
or ( n64705 , n592023 , n592026 , n64704 );
xor ( n64706 , n591916 , n64597 );
xor ( n64707 , n64706 , n64602 );
and ( n592031 , n64705 , n64707 );
xor ( n592032 , n591969 , n64662 );
xor ( n64710 , n592032 , n591988 );
and ( n592034 , n64707 , n64710 );
and ( n64712 , n64705 , n64710 );
or ( n64713 , n592031 , n592034 , n64712 );
and ( n592037 , n64682 , n64713 );
xor ( n592038 , n64682 , n64713 );
xor ( n64716 , n64705 , n64707 );
xor ( n592040 , n64716 , n64710 );
and ( n592041 , n64586 , n64491 );
and ( n64719 , n64533 , n64489 );
nor ( n592043 , n592041 , n64719 );
xnor ( n64721 , n592043 , n64448 );
and ( n64722 , n64630 , n64456 );
and ( n592046 , n64591 , n64454 );
nor ( n64724 , n64722 , n592046 );
xnor ( n592048 , n64724 , n591786 );
and ( n592049 , n64721 , n592048 );
not ( n64727 , n64684 );
and ( n592051 , n592048 , n64727 );
and ( n64729 , n64721 , n64727 );
or ( n592053 , n592049 , n592051 , n64729 );
and ( n592054 , n64450 , n64650 );
and ( n64732 , n64458 , n64648 );
nor ( n592056 , n592054 , n64732 );
xnor ( n64734 , n592056 , n591902 );
and ( n64735 , n592053 , n64734 );
xor ( n592059 , n64624 , n64628 );
xor ( n592060 , n592059 , n64631 );
and ( n64738 , n64734 , n592060 );
and ( n592062 , n592053 , n592060 );
or ( n64740 , n64735 , n64738 , n592062 );
xor ( n64741 , n64576 , n64619 );
xor ( n64742 , n64619 , n64620 );
not ( n64743 , n64742 );
and ( n64744 , n64741 , n64743 );
and ( n64745 , n64458 , n64744 );
not ( n64746 , n64745 );
xnor ( n64747 , n64746 , n64623 );
and ( n64748 , n64466 , n64650 );
and ( n64749 , n64450 , n64648 );
nor ( n64750 , n64748 , n64749 );
xnor ( n64751 , n64750 , n591902 );
and ( n64752 , n64747 , n64751 );
and ( n64753 , n591851 , n64559 );
and ( n64754 , n64501 , n591880 );
nor ( n64755 , n64753 , n64754 );
xnor ( n592079 , n64755 , n64521 );
and ( n64757 , n64751 , n592079 );
and ( n592081 , n64747 , n592079 );
or ( n592082 , n64752 , n64757 , n592081 );
buf ( n64760 , n591745 );
buf ( n64761 , n591746 );
and ( n592085 , n64760 , n64761 );
not ( n592086 , n592085 );
and ( n64764 , n64620 , n592086 );
not ( n592088 , n64764 );
and ( n592089 , n64591 , n64491 );
and ( n64767 , n64586 , n64489 );
nor ( n592091 , n592089 , n64767 );
xnor ( n592092 , n592091 , n64448 );
and ( n64770 , n592088 , n592092 );
buf ( n592094 , n591679 );
and ( n64772 , n592094 , n64451 );
and ( n592096 , n592092 , n64772 );
and ( n592097 , n592088 , n64772 );
or ( n64775 , n64770 , n592096 , n592097 );
and ( n64776 , n592094 , n64456 );
and ( n592100 , n64683 , n64454 );
nor ( n64778 , n64776 , n592100 );
xnor ( n592102 , n64778 , n591786 );
buf ( n592103 , n592102 );
and ( n592104 , n64533 , n64559 );
and ( n64782 , n591851 , n591880 );
nor ( n592106 , n592104 , n64782 );
xnor ( n592107 , n592106 , n64521 );
and ( n64785 , n592103 , n592107 );
and ( n592109 , n64683 , n64456 );
and ( n592110 , n64630 , n64454 );
nor ( n64788 , n592109 , n592110 );
xnor ( n592112 , n64788 , n591786 );
and ( n592113 , n592107 , n592112 );
and ( n64791 , n592103 , n592112 );
or ( n592115 , n64785 , n592113 , n64791 );
and ( n64793 , n64775 , n592115 );
xor ( n592117 , n64721 , n592048 );
xor ( n64795 , n592117 , n64727 );
and ( n592119 , n592115 , n64795 );
and ( n592120 , n64775 , n64795 );
or ( n592121 , n64793 , n592119 , n592120 );
and ( n64799 , n592082 , n592121 );
xor ( n592123 , n64685 , n592012 );
xor ( n592124 , n592123 , n64694 );
and ( n64802 , n592121 , n592124 );
and ( n592126 , n592082 , n592124 );
or ( n64804 , n64799 , n64802 , n592126 );
and ( n592128 , n64740 , n64804 );
xor ( n64806 , n64697 , n64699 );
xor ( n592130 , n64806 , n64702 );
and ( n592131 , n64804 , n592130 );
and ( n592132 , n64740 , n592130 );
or ( n64810 , n592128 , n592131 , n592132 );
and ( n592134 , n592040 , n64810 );
xor ( n592135 , n592040 , n64810 );
xor ( n64813 , n64740 , n64804 );
xor ( n592137 , n64813 , n592130 );
and ( n592138 , n64450 , n64744 );
and ( n64816 , n64458 , n64742 );
nor ( n592140 , n592138 , n64816 );
xnor ( n592141 , n592140 , n64623 );
and ( n64819 , n64501 , n64650 );
and ( n592143 , n64466 , n64648 );
nor ( n592144 , n64819 , n592143 );
xnor ( n64822 , n592144 , n591902 );
and ( n592146 , n592141 , n64822 );
xor ( n592147 , n592088 , n592092 );
xor ( n64825 , n592147 , n64772 );
and ( n592149 , n64822 , n64825 );
and ( n64827 , n592141 , n64825 );
or ( n64828 , n592146 , n592149 , n64827 );
and ( n64829 , n64586 , n64559 );
and ( n64830 , n64533 , n591880 );
nor ( n64831 , n64829 , n64830 );
xnor ( n592155 , n64831 , n64521 );
and ( n64833 , n64630 , n64491 );
and ( n64834 , n64591 , n64489 );
nor ( n64835 , n64833 , n64834 );
xnor ( n64836 , n64835 , n64448 );
and ( n64837 , n592155 , n64836 );
buf ( n64838 , n591680 );
and ( n64839 , n64838 , n64451 );
and ( n64840 , n64836 , n64839 );
and ( n64841 , n592155 , n64839 );
or ( n64842 , n64837 , n64840 , n64841 );
buf ( n64843 , n591747 );
buf ( n64844 , n591748 );
and ( n64845 , n64843 , n64844 );
not ( n64846 , n64845 );
and ( n64847 , n64761 , n64846 );
not ( n64848 , n64847 );
and ( n64849 , n64838 , n64456 );
and ( n64850 , n592094 , n64454 );
nor ( n64851 , n64849 , n64850 );
xnor ( n64852 , n64851 , n591786 );
and ( n64853 , n64848 , n64852 );
buf ( n64854 , n591681 );
and ( n64855 , n64854 , n64451 );
and ( n64856 , n64852 , n64855 );
and ( n64857 , n64848 , n64855 );
or ( n64858 , n64853 , n64856 , n64857 );
xor ( n64859 , n64620 , n64760 );
xor ( n64860 , n64760 , n64761 );
not ( n64861 , n64860 );
and ( n64862 , n64859 , n64861 );
and ( n592186 , n64458 , n64862 );
not ( n64864 , n592186 );
xnor ( n592188 , n64864 , n64764 );
and ( n592189 , n64858 , n592188 );
not ( n64867 , n592102 );
and ( n592191 , n592188 , n64867 );
and ( n64869 , n64858 , n64867 );
or ( n592193 , n592189 , n592191 , n64869 );
and ( n592194 , n64842 , n592193 );
xor ( n64872 , n592103 , n592107 );
xor ( n64873 , n64872 , n592112 );
and ( n592197 , n592193 , n64873 );
and ( n592198 , n64842 , n64873 );
or ( n64876 , n592194 , n592197 , n592198 );
and ( n64877 , n64828 , n64876 );
xor ( n592201 , n64747 , n64751 );
xor ( n592202 , n592201 , n592079 );
and ( n64880 , n64876 , n592202 );
and ( n592204 , n64828 , n592202 );
or ( n64882 , n64877 , n64880 , n592204 );
xor ( n64883 , n592053 , n64734 );
xor ( n592207 , n64883 , n592060 );
and ( n592208 , n64882 , n592207 );
xor ( n64886 , n592082 , n592121 );
xor ( n64887 , n64886 , n592124 );
and ( n592211 , n592207 , n64887 );
and ( n64889 , n64882 , n64887 );
or ( n592213 , n592208 , n592211 , n64889 );
and ( n592214 , n592137 , n592213 );
xor ( n64892 , n592137 , n592213 );
xor ( n64893 , n64882 , n592207 );
xor ( n64894 , n64893 , n64887 );
and ( n64895 , n592094 , n64491 );
and ( n64896 , n64683 , n64489 );
nor ( n64897 , n64895 , n64896 );
xnor ( n64898 , n64897 , n64448 );
buf ( n64899 , n64898 );
and ( n592223 , n64591 , n64559 );
and ( n64901 , n64586 , n591880 );
nor ( n64902 , n592223 , n64901 );
xnor ( n64903 , n64902 , n64521 );
and ( n592227 , n64899 , n64903 );
and ( n64905 , n64683 , n64491 );
and ( n64906 , n64630 , n64489 );
nor ( n64907 , n64905 , n64906 );
xnor ( n592231 , n64907 , n64448 );
and ( n592232 , n64903 , n592231 );
and ( n64910 , n64899 , n592231 );
or ( n592234 , n592227 , n592232 , n64910 );
and ( n64912 , n64466 , n64744 );
and ( n64913 , n64450 , n64742 );
nor ( n592237 , n64912 , n64913 );
xnor ( n64915 , n592237 , n64623 );
and ( n592239 , n592234 , n64915 );
and ( n592240 , n591851 , n64650 );
and ( n64918 , n64501 , n64648 );
nor ( n64919 , n592240 , n64918 );
xnor ( n64920 , n64919 , n591902 );
and ( n64921 , n64915 , n64920 );
and ( n592245 , n592234 , n64920 );
or ( n64923 , n592239 , n64921 , n592245 );
and ( n592247 , n64450 , n64862 );
and ( n592248 , n64458 , n64860 );
nor ( n64926 , n592247 , n592248 );
xnor ( n592250 , n64926 , n64764 );
and ( n64928 , n64501 , n64744 );
and ( n64929 , n64466 , n64742 );
nor ( n592253 , n64928 , n64929 );
xnor ( n592254 , n592253 , n64623 );
and ( n64932 , n592250 , n592254 );
and ( n592256 , n64533 , n64650 );
and ( n592257 , n591851 , n64648 );
nor ( n64935 , n592256 , n592257 );
xnor ( n64936 , n64935 , n591902 );
and ( n64937 , n592254 , n64936 );
and ( n64938 , n592250 , n64936 );
or ( n64939 , n64932 , n64937 , n64938 );
xor ( n64940 , n592155 , n64836 );
xor ( n64941 , n64940 , n64839 );
and ( n64942 , n64939 , n64941 );
xor ( n64943 , n64858 , n592188 );
xor ( n64944 , n64943 , n64867 );
and ( n64945 , n64941 , n64944 );
and ( n64946 , n64939 , n64944 );
or ( n64947 , n64942 , n64945 , n64946 );
and ( n64948 , n64923 , n64947 );
xor ( n64949 , n592141 , n64822 );
xor ( n64950 , n64949 , n64825 );
and ( n64951 , n64947 , n64950 );
and ( n592275 , n64923 , n64950 );
or ( n64953 , n64948 , n64951 , n592275 );
xor ( n592277 , n64775 , n592115 );
xor ( n592278 , n592277 , n64795 );
and ( n64956 , n64953 , n592278 );
xor ( n592280 , n64828 , n64876 );
xor ( n592281 , n592280 , n592202 );
and ( n64959 , n592278 , n592281 );
and ( n64960 , n64953 , n592281 );
or ( n64961 , n64956 , n64959 , n64960 );
and ( n592285 , n64894 , n64961 );
xor ( n64963 , n64894 , n64961 );
and ( n64964 , n64630 , n64559 );
and ( n64965 , n64591 , n591880 );
nor ( n64966 , n64964 , n64965 );
xnor ( n592290 , n64966 , n64521 );
and ( n64968 , n64854 , n64456 );
and ( n592292 , n64838 , n64454 );
nor ( n592293 , n64968 , n592292 );
xnor ( n64971 , n592293 , n591786 );
and ( n592295 , n592290 , n64971 );
buf ( n64973 , n591682 );
and ( n64974 , n64973 , n64451 );
and ( n64975 , n64971 , n64974 );
and ( n64976 , n592290 , n64974 );
or ( n64977 , n592295 , n64975 , n64976 );
xor ( n64978 , n64848 , n64852 );
xor ( n64979 , n64978 , n64855 );
and ( n64980 , n64977 , n64979 );
xor ( n64981 , n64899 , n64903 );
xor ( n64982 , n64981 , n592231 );
and ( n64983 , n64979 , n64982 );
and ( n64984 , n64977 , n64982 );
or ( n64985 , n64980 , n64983 , n64984 );
buf ( n64986 , n591749 );
buf ( n64987 , n591750 );
and ( n64988 , n64986 , n64987 );
not ( n64989 , n64988 );
and ( n64990 , n64844 , n64989 );
not ( n64991 , n64990 );
and ( n64992 , n64973 , n64456 );
and ( n64993 , n64854 , n64454 );
nor ( n64994 , n64992 , n64993 );
xnor ( n592318 , n64994 , n591786 );
and ( n592319 , n64991 , n592318 );
buf ( n64997 , n591683 );
and ( n64998 , n64997 , n64451 );
and ( n64999 , n592318 , n64998 );
and ( n592323 , n64991 , n64998 );
or ( n65001 , n592319 , n64999 , n592323 );
and ( n65002 , n64466 , n64862 );
and ( n65003 , n64450 , n64860 );
nor ( n592327 , n65002 , n65003 );
xnor ( n592328 , n592327 , n64764 );
and ( n65006 , n65001 , n592328 );
and ( n592330 , n591851 , n64744 );
and ( n65008 , n64501 , n64742 );
nor ( n65009 , n592330 , n65008 );
xnor ( n65010 , n65009 , n64623 );
and ( n592334 , n592328 , n65010 );
and ( n592335 , n65001 , n65010 );
or ( n65013 , n65006 , n592334 , n592335 );
xor ( n592337 , n64761 , n64843 );
xor ( n65015 , n64843 , n64844 );
not ( n592339 , n65015 );
and ( n592340 , n592337 , n592339 );
and ( n65018 , n64458 , n592340 );
not ( n592342 , n65018 );
xnor ( n65020 , n592342 , n64847 );
and ( n65021 , n64586 , n64650 );
and ( n65022 , n64533 , n64648 );
nor ( n65023 , n65021 , n65022 );
xnor ( n592347 , n65023 , n591902 );
and ( n65025 , n65020 , n592347 );
not ( n592349 , n64898 );
and ( n65027 , n592347 , n592349 );
and ( n592351 , n65020 , n592349 );
or ( n592352 , n65025 , n65027 , n592351 );
and ( n65030 , n65013 , n592352 );
xor ( n592354 , n592250 , n592254 );
xor ( n65032 , n592354 , n64936 );
and ( n65033 , n592352 , n65032 );
and ( n65034 , n65013 , n65032 );
or ( n65035 , n65030 , n65033 , n65034 );
and ( n65036 , n64985 , n65035 );
xor ( n592360 , n592234 , n64915 );
xor ( n65038 , n592360 , n64920 );
and ( n592362 , n65035 , n65038 );
and ( n65040 , n64985 , n65038 );
or ( n65041 , n65036 , n592362 , n65040 );
xor ( n65042 , n64842 , n592193 );
xor ( n592366 , n65042 , n64873 );
and ( n592367 , n65041 , n592366 );
xor ( n65045 , n64923 , n64947 );
xor ( n592369 , n65045 , n64950 );
and ( n592370 , n592366 , n592369 );
and ( n65048 , n65041 , n592369 );
or ( n592372 , n592367 , n592370 , n65048 );
xor ( n65050 , n64953 , n592278 );
xor ( n65051 , n65050 , n592281 );
and ( n65052 , n592372 , n65051 );
xor ( n65053 , n592372 , n65051 );
xor ( n65054 , n65041 , n592366 );
xor ( n65055 , n65054 , n592369 );
and ( n65056 , n64591 , n64650 );
and ( n65057 , n64586 , n64648 );
nor ( n65058 , n65056 , n65057 );
xnor ( n65059 , n65058 , n591902 );
and ( n592383 , n64683 , n64559 );
and ( n592384 , n64630 , n591880 );
nor ( n65062 , n592383 , n592384 );
xnor ( n592386 , n65062 , n64521 );
and ( n65064 , n65059 , n592386 );
and ( n65065 , n64838 , n64491 );
and ( n65066 , n592094 , n64489 );
nor ( n65067 , n65065 , n65066 );
xnor ( n65068 , n65067 , n64448 );
and ( n592392 , n592386 , n65068 );
and ( n592393 , n65059 , n65068 );
or ( n65071 , n65064 , n592392 , n592393 );
and ( n592395 , n64854 , n64491 );
and ( n592396 , n64838 , n64489 );
nor ( n65074 , n592395 , n592396 );
xnor ( n592398 , n65074 , n64448 );
and ( n592399 , n64997 , n64456 );
and ( n65077 , n64973 , n64454 );
nor ( n592401 , n592399 , n65077 );
xnor ( n65079 , n592401 , n591786 );
and ( n65080 , n592398 , n65079 );
buf ( n592404 , n591684 );
and ( n65082 , n592404 , n64451 );
and ( n592406 , n65079 , n65082 );
and ( n65084 , n592398 , n65082 );
or ( n592408 , n65080 , n592406 , n65084 );
and ( n592409 , n592094 , n64559 );
and ( n65087 , n64683 , n591880 );
nor ( n592411 , n592409 , n65087 );
xnor ( n65089 , n592411 , n64521 );
buf ( n65090 , n65089 );
and ( n65091 , n592408 , n65090 );
and ( n65092 , n64533 , n64744 );
and ( n65093 , n591851 , n64742 );
nor ( n592417 , n65092 , n65093 );
xnor ( n592418 , n592417 , n64623 );
and ( n65096 , n65090 , n592418 );
and ( n592420 , n592408 , n592418 );
or ( n592421 , n65091 , n65096 , n592420 );
and ( n65099 , n65071 , n592421 );
xor ( n592423 , n592290 , n64971 );
xor ( n65101 , n592423 , n64974 );
and ( n65102 , n592421 , n65101 );
and ( n65103 , n65071 , n65101 );
or ( n65104 , n65099 , n65102 , n65103 );
and ( n592428 , n64450 , n592340 );
and ( n65106 , n64458 , n65015 );
nor ( n592430 , n592428 , n65106 );
xnor ( n592431 , n592430 , n64847 );
and ( n592432 , n64501 , n64862 );
and ( n65110 , n64466 , n64860 );
nor ( n592434 , n592432 , n65110 );
xnor ( n592435 , n592434 , n64764 );
and ( n65113 , n592431 , n592435 );
xor ( n592437 , n64991 , n592318 );
xor ( n65115 , n592437 , n64998 );
and ( n65116 , n592435 , n65115 );
and ( n592440 , n592431 , n65115 );
or ( n65118 , n65113 , n65116 , n592440 );
xor ( n592442 , n65001 , n592328 );
xor ( n65120 , n592442 , n65010 );
and ( n65121 , n65118 , n65120 );
xor ( n65122 , n65020 , n592347 );
xor ( n592446 , n65122 , n592349 );
and ( n65124 , n65120 , n592446 );
and ( n592448 , n65118 , n592446 );
or ( n65126 , n65121 , n65124 , n592448 );
and ( n592450 , n65104 , n65126 );
xor ( n592451 , n64977 , n64979 );
xor ( n592452 , n592451 , n64982 );
and ( n65130 , n65126 , n592452 );
and ( n592454 , n65104 , n592452 );
or ( n592455 , n592450 , n65130 , n592454 );
xor ( n65133 , n64939 , n64941 );
xor ( n592457 , n65133 , n64944 );
and ( n592458 , n592455 , n592457 );
xor ( n592459 , n64985 , n65035 );
xor ( n592460 , n592459 , n65038 );
and ( n592461 , n592457 , n592460 );
and ( n592462 , n592455 , n592460 );
or ( n65140 , n592458 , n592461 , n592462 );
and ( n592464 , n65055 , n65140 );
xor ( n592465 , n65055 , n65140 );
xor ( n65143 , n592455 , n592457 );
xor ( n592467 , n65143 , n592460 );
buf ( n592468 , n591686 );
and ( n65146 , n592468 , n64451 );
buf ( n592470 , n65146 );
buf ( n592471 , n591751 );
buf ( n65149 , n591752 );
and ( n592473 , n592471 , n65149 );
not ( n65151 , n592473 );
and ( n592475 , n64987 , n65151 );
not ( n65153 , n592475 );
and ( n592477 , n592470 , n65153 );
buf ( n592478 , n591685 );
and ( n65156 , n592478 , n64451 );
and ( n592480 , n65153 , n65156 );
and ( n592481 , n592470 , n65156 );
or ( n65159 , n592477 , n592480 , n592481 );
xor ( n592483 , n64844 , n64986 );
xor ( n592484 , n64986 , n64987 );
not ( n65162 , n592484 );
and ( n592486 , n592483 , n65162 );
and ( n65164 , n64458 , n592486 );
not ( n65165 , n65164 );
xnor ( n65166 , n65165 , n64990 );
and ( n65167 , n65159 , n65166 );
and ( n65168 , n591851 , n64862 );
and ( n65169 , n64501 , n64860 );
nor ( n65170 , n65168 , n65169 );
xnor ( n65171 , n65170 , n64764 );
and ( n65172 , n65166 , n65171 );
and ( n65173 , n65159 , n65171 );
or ( n65174 , n65167 , n65172 , n65173 );
and ( n65175 , n64586 , n64744 );
and ( n65176 , n64533 , n64742 );
nor ( n65177 , n65175 , n65176 );
xnor ( n65178 , n65177 , n64623 );
and ( n65179 , n64630 , n64650 );
and ( n65180 , n64591 , n64648 );
nor ( n65181 , n65179 , n65180 );
xnor ( n65182 , n65181 , n591902 );
and ( n65183 , n65178 , n65182 );
not ( n65184 , n65089 );
and ( n65185 , n65182 , n65184 );
and ( n65186 , n65178 , n65184 );
or ( n65187 , n65183 , n65185 , n65186 );
and ( n65188 , n65174 , n65187 );
xor ( n65189 , n65059 , n592386 );
xor ( n65190 , n65189 , n65068 );
and ( n65191 , n65187 , n65190 );
and ( n65192 , n65174 , n65190 );
or ( n65193 , n65188 , n65191 , n65192 );
and ( n65194 , n64838 , n64559 );
and ( n65195 , n592094 , n591880 );
nor ( n65196 , n65194 , n65195 );
xnor ( n65197 , n65196 , n64521 );
and ( n65198 , n64973 , n64491 );
and ( n65199 , n64854 , n64489 );
nor ( n65200 , n65198 , n65199 );
xnor ( n65201 , n65200 , n64448 );
and ( n65202 , n65197 , n65201 );
and ( n65203 , n592404 , n64456 );
and ( n65204 , n64997 , n64454 );
nor ( n65205 , n65203 , n65204 );
xnor ( n65206 , n65205 , n591786 );
and ( n65207 , n65201 , n65206 );
and ( n65208 , n65197 , n65206 );
or ( n65209 , n65202 , n65207 , n65208 );
and ( n65210 , n64466 , n592340 );
and ( n65211 , n64450 , n65015 );
nor ( n65212 , n65210 , n65211 );
xnor ( n65213 , n65212 , n64847 );
and ( n65214 , n65209 , n65213 );
xor ( n592538 , n592398 , n65079 );
xor ( n65216 , n592538 , n65082 );
and ( n65217 , n65213 , n65216 );
and ( n65218 , n65209 , n65216 );
or ( n65219 , n65214 , n65217 , n65218 );
xor ( n65220 , n592408 , n65090 );
xor ( n65221 , n65220 , n592418 );
and ( n65222 , n65219 , n65221 );
xor ( n65223 , n592431 , n592435 );
xor ( n592547 , n65223 , n65115 );
and ( n65225 , n65221 , n592547 );
and ( n592549 , n65219 , n592547 );
or ( n65227 , n65222 , n65225 , n592549 );
and ( n65228 , n65193 , n65227 );
xor ( n65229 , n65071 , n592421 );
xor ( n65230 , n65229 , n65101 );
and ( n65231 , n65227 , n65230 );
and ( n65232 , n65193 , n65230 );
or ( n65233 , n65228 , n65231 , n65232 );
xor ( n65234 , n65013 , n592352 );
xor ( n65235 , n65234 , n65032 );
and ( n65236 , n65233 , n65235 );
xor ( n65237 , n65104 , n65126 );
xor ( n592561 , n65237 , n592452 );
and ( n65239 , n65235 , n592561 );
and ( n592563 , n65233 , n592561 );
or ( n592564 , n65236 , n65239 , n592563 );
and ( n65242 , n592467 , n592564 );
xor ( n65243 , n592467 , n592564 );
xor ( n592567 , n65233 , n65235 );
xor ( n65245 , n592567 , n592561 );
and ( n592569 , n592094 , n64650 );
and ( n65247 , n64683 , n64648 );
nor ( n592571 , n592569 , n65247 );
xnor ( n592572 , n592571 , n591902 );
and ( n65250 , n592478 , n64456 );
and ( n592574 , n592404 , n64454 );
nor ( n592575 , n65250 , n592574 );
xnor ( n65253 , n592575 , n591786 );
and ( n65254 , n592572 , n65253 );
not ( n592578 , n65146 );
and ( n65256 , n65253 , n592578 );
and ( n65257 , n592572 , n592578 );
or ( n592581 , n65254 , n65256 , n65257 );
and ( n65259 , n64501 , n592340 );
and ( n592583 , n64466 , n65015 );
nor ( n65261 , n65259 , n592583 );
xnor ( n592585 , n65261 , n64847 );
and ( n65263 , n592581 , n592585 );
and ( n592587 , n64533 , n64862 );
and ( n592588 , n591851 , n64860 );
nor ( n65266 , n592587 , n592588 );
xnor ( n592590 , n65266 , n64764 );
and ( n592591 , n592585 , n592590 );
and ( n65269 , n592581 , n592590 );
or ( n592593 , n65263 , n592591 , n65269 );
and ( n592594 , n64591 , n64744 );
and ( n65272 , n64586 , n64742 );
nor ( n592596 , n592594 , n65272 );
xnor ( n592597 , n592596 , n64623 );
and ( n65275 , n64683 , n64650 );
and ( n65276 , n64630 , n64648 );
nor ( n65277 , n65275 , n65276 );
xnor ( n65278 , n65277 , n591902 );
and ( n65279 , n592597 , n65278 );
xor ( n65280 , n592470 , n65153 );
xor ( n65281 , n65280 , n65156 );
and ( n65282 , n65278 , n65281 );
and ( n65283 , n592597 , n65281 );
or ( n65284 , n65279 , n65282 , n65283 );
and ( n592608 , n592593 , n65284 );
xor ( n65286 , n65178 , n65182 );
xor ( n592610 , n65286 , n65184 );
and ( n592611 , n65284 , n592610 );
and ( n65289 , n592593 , n592610 );
or ( n592613 , n592608 , n592611 , n65289 );
xor ( n65291 , n65174 , n65187 );
xor ( n592615 , n65291 , n65190 );
and ( n65293 , n592613 , n592615 );
xor ( n592617 , n65219 , n65221 );
xor ( n592618 , n592617 , n592547 );
and ( n65296 , n592615 , n592618 );
and ( n592620 , n592613 , n592618 );
or ( n65298 , n65293 , n65296 , n592620 );
xor ( n65299 , n65118 , n65120 );
xor ( n592623 , n65299 , n592446 );
and ( n65301 , n65298 , n592623 );
xor ( n592625 , n65193 , n65227 );
xor ( n592626 , n592625 , n65230 );
and ( n592627 , n592623 , n592626 );
and ( n592628 , n65298 , n592626 );
or ( n65306 , n65301 , n592627 , n592628 );
and ( n592630 , n65245 , n65306 );
xor ( n592631 , n65245 , n65306 );
xor ( n592632 , n65298 , n592623 );
xor ( n65310 , n592632 , n592626 );
buf ( n592634 , n591753 );
buf ( n592635 , n591754 );
and ( n65313 , n592634 , n592635 );
not ( n592637 , n65313 );
and ( n592638 , n65149 , n592637 );
not ( n592639 , n592638 );
and ( n65317 , n592468 , n64456 );
and ( n592641 , n592478 , n64454 );
nor ( n592642 , n65317 , n592641 );
xnor ( n65320 , n592642 , n591786 );
and ( n592644 , n592639 , n65320 );
buf ( n592645 , n591687 );
and ( n65323 , n592645 , n64451 );
and ( n592647 , n65320 , n65323 );
and ( n592648 , n592639 , n65323 );
or ( n65326 , n592644 , n592647 , n592648 );
and ( n592650 , n64854 , n64559 );
and ( n592651 , n64838 , n591880 );
nor ( n65329 , n592650 , n592651 );
xnor ( n592653 , n65329 , n64521 );
and ( n65331 , n65326 , n592653 );
and ( n65332 , n64997 , n64491 );
and ( n65333 , n64973 , n64489 );
nor ( n65334 , n65332 , n65333 );
xnor ( n65335 , n65334 , n64448 );
and ( n592659 , n592653 , n65335 );
and ( n65337 , n65326 , n65335 );
or ( n592661 , n65331 , n592659 , n65337 );
and ( n65339 , n64450 , n592486 );
and ( n65340 , n64458 , n592484 );
nor ( n592664 , n65339 , n65340 );
xnor ( n65342 , n592664 , n64990 );
and ( n65343 , n592661 , n65342 );
xor ( n592667 , n65197 , n65201 );
xor ( n592668 , n592667 , n65206 );
and ( n592669 , n65342 , n592668 );
and ( n65347 , n592661 , n592668 );
or ( n592671 , n65343 , n592669 , n65347 );
xor ( n592672 , n65159 , n65166 );
xor ( n65350 , n592672 , n65171 );
and ( n592674 , n592671 , n65350 );
xor ( n592675 , n65209 , n65213 );
xor ( n65353 , n592675 , n65216 );
and ( n592677 , n65350 , n65353 );
and ( n592678 , n592671 , n65353 );
or ( n65356 , n592674 , n592677 , n592678 );
xor ( n592680 , n64987 , n592471 );
xor ( n592681 , n592471 , n65149 );
not ( n65359 , n592681 );
and ( n592683 , n592680 , n65359 );
and ( n592684 , n64458 , n592683 );
not ( n65362 , n592684 );
xnor ( n592686 , n65362 , n592475 );
and ( n592687 , n64586 , n64862 );
and ( n65365 , n64533 , n64860 );
nor ( n592689 , n592687 , n65365 );
xnor ( n65367 , n592689 , n64764 );
and ( n65368 , n592686 , n65367 );
and ( n65369 , n64630 , n64744 );
and ( n65370 , n64591 , n64742 );
nor ( n65371 , n65369 , n65370 );
xnor ( n65372 , n65371 , n64623 );
and ( n65373 , n65367 , n65372 );
and ( n65374 , n592686 , n65372 );
or ( n65375 , n65368 , n65373 , n65374 );
xor ( n65376 , n592581 , n592585 );
xor ( n65377 , n65376 , n592590 );
and ( n65378 , n65375 , n65377 );
xor ( n65379 , n592597 , n65278 );
xor ( n65380 , n65379 , n65281 );
and ( n65381 , n65377 , n65380 );
and ( n65382 , n65375 , n65380 );
or ( n65383 , n65378 , n65381 , n65382 );
buf ( n65384 , n591688 );
and ( n65385 , n65384 , n64451 );
buf ( n65386 , n65385 );
and ( n65387 , n64973 , n64559 );
and ( n65388 , n64854 , n591880 );
nor ( n65389 , n65387 , n65388 );
xnor ( n65390 , n65389 , n64521 );
and ( n592714 , n65386 , n65390 );
and ( n65392 , n592404 , n64491 );
and ( n592716 , n64997 , n64489 );
nor ( n592717 , n65392 , n592716 );
xnor ( n65395 , n592717 , n64448 );
and ( n65396 , n65390 , n65395 );
and ( n65397 , n65386 , n65395 );
or ( n592721 , n592714 , n65396 , n65397 );
and ( n65399 , n64466 , n592486 );
and ( n592723 , n64450 , n592484 );
nor ( n65401 , n65399 , n592723 );
xnor ( n65402 , n65401 , n64990 );
and ( n65403 , n592721 , n65402 );
and ( n65404 , n591851 , n592340 );
and ( n592728 , n64501 , n65015 );
nor ( n65406 , n65404 , n592728 );
xnor ( n65407 , n65406 , n64847 );
and ( n65408 , n65402 , n65407 );
and ( n65409 , n592721 , n65407 );
or ( n592733 , n65403 , n65408 , n65409 );
and ( n65411 , n64591 , n64862 );
and ( n592735 , n64586 , n64860 );
nor ( n65413 , n65411 , n592735 );
xnor ( n65414 , n65413 , n64764 );
and ( n65415 , n64838 , n64650 );
and ( n65416 , n592094 , n64648 );
nor ( n592740 , n65415 , n65416 );
xnor ( n65418 , n592740 , n591902 );
and ( n592742 , n65414 , n65418 );
xor ( n65420 , n592639 , n65320 );
xor ( n592744 , n65420 , n65323 );
and ( n65422 , n65418 , n592744 );
and ( n592746 , n65414 , n592744 );
or ( n65424 , n592742 , n65422 , n592746 );
xor ( n592748 , n65326 , n592653 );
xor ( n592749 , n592748 , n65335 );
and ( n592750 , n65424 , n592749 );
xor ( n65428 , n592572 , n65253 );
xor ( n592752 , n65428 , n592578 );
and ( n592753 , n592749 , n592752 );
and ( n65431 , n65424 , n592752 );
or ( n65432 , n592750 , n592753 , n65431 );
and ( n592756 , n592733 , n65432 );
xor ( n65434 , n592661 , n65342 );
xor ( n65435 , n65434 , n592668 );
and ( n592759 , n65432 , n65435 );
and ( n592760 , n592733 , n65435 );
or ( n65438 , n592756 , n592759 , n592760 );
and ( n592762 , n65383 , n65438 );
xor ( n592763 , n592593 , n65284 );
xor ( n65441 , n592763 , n592610 );
and ( n65442 , n65438 , n65441 );
and ( n592766 , n65383 , n65441 );
or ( n592767 , n592762 , n65442 , n592766 );
and ( n65445 , n65356 , n592767 );
xor ( n65446 , n592613 , n592615 );
xor ( n592770 , n65446 , n592618 );
and ( n65448 , n592767 , n592770 );
and ( n65449 , n65356 , n592770 );
or ( n592773 , n65445 , n65448 , n65449 );
and ( n592774 , n65310 , n592773 );
xor ( n65452 , n65310 , n592773 );
xor ( n65453 , n65356 , n592767 );
xor ( n592777 , n65453 , n592770 );
and ( n592778 , n592094 , n64744 );
and ( n65456 , n64683 , n64742 );
nor ( n592780 , n592778 , n65456 );
xnor ( n65458 , n592780 , n64623 );
and ( n65459 , n64997 , n64559 );
and ( n592783 , n64973 , n591880 );
nor ( n65461 , n65459 , n592783 );
xnor ( n592785 , n65461 , n64521 );
and ( n65463 , n65458 , n592785 );
and ( n592787 , n592478 , n64491 );
and ( n592788 , n592404 , n64489 );
nor ( n65466 , n592787 , n592788 );
xnor ( n592790 , n65466 , n64448 );
and ( n65468 , n592785 , n592790 );
and ( n65469 , n65458 , n592790 );
or ( n592793 , n65463 , n65468 , n65469 );
and ( n65471 , n64450 , n592683 );
and ( n65472 , n64458 , n592681 );
nor ( n592796 , n65471 , n65472 );
xnor ( n65474 , n592796 , n592475 );
and ( n592798 , n592793 , n65474 );
and ( n592799 , n64501 , n592486 );
and ( n65477 , n64466 , n592484 );
nor ( n65478 , n592799 , n65477 );
xnor ( n592802 , n65478 , n64990 );
and ( n592803 , n65474 , n592802 );
and ( n65481 , n592793 , n592802 );
or ( n592805 , n592798 , n592803 , n65481 );
buf ( n592806 , n591690 );
and ( n65484 , n592806 , n64451 );
buf ( n592808 , n65484 );
buf ( n65486 , n591755 );
buf ( n65487 , n591756 );
and ( n592811 , n65486 , n65487 );
not ( n592812 , n592811 );
and ( n65490 , n592635 , n592812 );
not ( n592814 , n65490 );
and ( n65492 , n592808 , n592814 );
buf ( n65493 , n591689 );
and ( n65494 , n65493 , n64451 );
and ( n65495 , n592814 , n65494 );
and ( n65496 , n592808 , n65494 );
or ( n65497 , n65492 , n65495 , n65496 );
and ( n65498 , n592645 , n64456 );
and ( n65499 , n592468 , n64454 );
nor ( n592823 , n65498 , n65499 );
xnor ( n65501 , n592823 , n591786 );
and ( n592825 , n65497 , n65501 );
not ( n65503 , n65385 );
and ( n65504 , n65501 , n65503 );
and ( n65505 , n65497 , n65503 );
or ( n65506 , n592825 , n65504 , n65505 );
and ( n65507 , n64533 , n592340 );
and ( n592831 , n591851 , n65015 );
nor ( n65509 , n65507 , n592831 );
xnor ( n592833 , n65509 , n64847 );
and ( n592834 , n65506 , n592833 );
and ( n592835 , n64683 , n64744 );
and ( n65513 , n64630 , n64742 );
nor ( n592837 , n592835 , n65513 );
xnor ( n592838 , n592837 , n64623 );
and ( n65516 , n592833 , n592838 );
and ( n592840 , n65506 , n592838 );
or ( n592841 , n592834 , n65516 , n592840 );
and ( n65519 , n592805 , n592841 );
xor ( n65520 , n592686 , n65367 );
xor ( n65521 , n65520 , n65372 );
and ( n65522 , n592841 , n65521 );
and ( n65523 , n592805 , n65521 );
or ( n65524 , n65519 , n65522 , n65523 );
and ( n65525 , n64586 , n592340 );
and ( n65526 , n64533 , n65015 );
nor ( n65527 , n65525 , n65526 );
xnor ( n65528 , n65527 , n64847 );
and ( n65529 , n64630 , n64862 );
and ( n65530 , n64591 , n64860 );
nor ( n65531 , n65529 , n65530 );
xnor ( n65532 , n65531 , n64764 );
and ( n65533 , n65528 , n65532 );
and ( n592857 , n64854 , n64650 );
and ( n65535 , n64838 , n64648 );
nor ( n592859 , n592857 , n65535 );
xnor ( n65537 , n592859 , n591902 );
and ( n592861 , n65532 , n65537 );
and ( n592862 , n65528 , n65537 );
or ( n592863 , n65533 , n592861 , n592862 );
xor ( n65541 , n65386 , n65390 );
xor ( n65542 , n65541 , n65395 );
and ( n65543 , n592863 , n65542 );
xor ( n592867 , n65414 , n65418 );
xor ( n65545 , n592867 , n592744 );
and ( n592869 , n65542 , n65545 );
and ( n65547 , n592863 , n65545 );
or ( n65548 , n65543 , n592869 , n65547 );
xor ( n65549 , n592721 , n65402 );
xor ( n65550 , n65549 , n65407 );
and ( n65551 , n65548 , n65550 );
xor ( n65552 , n65424 , n592749 );
xor ( n65553 , n65552 , n592752 );
and ( n65554 , n65550 , n65553 );
and ( n65555 , n65548 , n65553 );
or ( n65556 , n65551 , n65554 , n65555 );
and ( n65557 , n65524 , n65556 );
xor ( n65558 , n65375 , n65377 );
xor ( n65559 , n65558 , n65380 );
and ( n592883 , n65556 , n65559 );
and ( n65561 , n65524 , n65559 );
or ( n592885 , n65557 , n592883 , n65561 );
xor ( n65563 , n592671 , n65350 );
xor ( n592887 , n65563 , n65353 );
and ( n65565 , n592885 , n592887 );
xor ( n65566 , n65383 , n65438 );
xor ( n65567 , n65566 , n65441 );
and ( n65568 , n592887 , n65567 );
and ( n65569 , n592885 , n65567 );
or ( n65570 , n65565 , n65568 , n65569 );
and ( n65571 , n592777 , n65570 );
xor ( n65572 , n592777 , n65570 );
xor ( n592896 , n592885 , n592887 );
xor ( n592897 , n592896 , n65567 );
and ( n65575 , n592468 , n64491 );
and ( n592899 , n592478 , n64489 );
nor ( n592900 , n65575 , n592899 );
xnor ( n65578 , n592900 , n64448 );
and ( n592902 , n65384 , n64456 );
and ( n65580 , n592645 , n64454 );
nor ( n65581 , n592902 , n65580 );
xnor ( n592905 , n65581 , n591786 );
and ( n592906 , n65578 , n592905 );
xor ( n65584 , n592808 , n592814 );
xor ( n592908 , n65584 , n65494 );
and ( n65586 , n592905 , n592908 );
and ( n592910 , n65578 , n592908 );
or ( n592911 , n592906 , n65586 , n592910 );
xor ( n65589 , n65149 , n592634 );
xor ( n592913 , n592634 , n592635 );
not ( n592914 , n592913 );
and ( n65592 , n65589 , n592914 );
and ( n592916 , n64458 , n65592 );
not ( n65594 , n592916 );
xnor ( n592918 , n65594 , n592638 );
and ( n592919 , n592911 , n592918 );
xor ( n65597 , n65497 , n65501 );
xor ( n592921 , n65597 , n65503 );
and ( n592922 , n592918 , n592921 );
and ( n592923 , n592911 , n592921 );
or ( n65601 , n592919 , n592922 , n592923 );
xor ( n592925 , n592793 , n65474 );
xor ( n592926 , n592925 , n592802 );
and ( n592927 , n65601 , n592926 );
xor ( n65605 , n65506 , n592833 );
xor ( n592929 , n65605 , n592838 );
and ( n592930 , n592926 , n592929 );
and ( n65608 , n65601 , n592929 );
or ( n592932 , n592927 , n592930 , n65608 );
xor ( n592933 , n592805 , n592841 );
xor ( n65611 , n592933 , n65521 );
and ( n592935 , n592932 , n65611 );
xor ( n65613 , n65548 , n65550 );
xor ( n65614 , n65613 , n65553 );
and ( n65615 , n65611 , n65614 );
and ( n592939 , n592932 , n65614 );
or ( n592940 , n592935 , n65615 , n592939 );
xor ( n65618 , n592733 , n65432 );
xor ( n592942 , n65618 , n65435 );
and ( n592943 , n592940 , n592942 );
xor ( n592944 , n65524 , n65556 );
xor ( n65622 , n592944 , n65559 );
and ( n592946 , n592942 , n65622 );
and ( n592947 , n592940 , n65622 );
or ( n65625 , n592943 , n592946 , n592947 );
and ( n592949 , n592897 , n65625 );
xor ( n592950 , n592897 , n65625 );
xor ( n65628 , n592940 , n592942 );
xor ( n592952 , n65628 , n65622 );
buf ( n65630 , n591692 );
and ( n592954 , n65630 , n64451 );
buf ( n592955 , n592954 );
buf ( n65633 , n591757 );
buf ( n592957 , n591758 );
and ( n65635 , n65633 , n592957 );
not ( n65636 , n65635 );
and ( n592960 , n65487 , n65636 );
not ( n65638 , n592960 );
and ( n592962 , n592955 , n65638 );
buf ( n65640 , n591691 );
and ( n65641 , n65640 , n64451 );
and ( n592965 , n65638 , n65641 );
and ( n592966 , n592955 , n65641 );
or ( n592967 , n592962 , n592965 , n592966 );
and ( n65645 , n592478 , n64559 );
and ( n592969 , n592404 , n591880 );
nor ( n592970 , n65645 , n592969 );
xnor ( n65648 , n592970 , n64521 );
and ( n65649 , n592967 , n65648 );
and ( n65650 , n592645 , n64491 );
and ( n592974 , n592468 , n64489 );
nor ( n65652 , n65650 , n592974 );
xnor ( n592976 , n65652 , n64448 );
and ( n65654 , n65493 , n64456 );
and ( n65655 , n65384 , n64454 );
nor ( n65656 , n65654 , n65655 );
xnor ( n65657 , n65656 , n591786 );
xor ( n65658 , n592976 , n65657 );
not ( n65659 , n65484 );
xor ( n592983 , n65658 , n65659 );
and ( n592984 , n65648 , n592983 );
and ( n65662 , n592967 , n592983 );
or ( n592986 , n65649 , n592984 , n65662 );
and ( n65664 , n64450 , n65592 );
and ( n65665 , n64458 , n592913 );
nor ( n592989 , n65664 , n65665 );
xnor ( n65667 , n592989 , n592638 );
and ( n592991 , n592986 , n65667 );
and ( n592992 , n64501 , n592683 );
and ( n65670 , n64466 , n592681 );
nor ( n592994 , n592992 , n65670 );
xnor ( n592995 , n592994 , n592475 );
and ( n65673 , n65667 , n592995 );
and ( n65674 , n592986 , n592995 );
or ( n65675 , n592991 , n65673 , n65674 );
and ( n65676 , n592094 , n64862 );
and ( n593000 , n64683 , n64860 );
nor ( n593001 , n65676 , n593000 );
xnor ( n65679 , n593001 , n64764 );
and ( n593003 , n64854 , n64744 );
and ( n593004 , n64838 , n64742 );
nor ( n65682 , n593003 , n593004 );
xnor ( n593006 , n65682 , n64623 );
and ( n593007 , n65679 , n593006 );
and ( n65685 , n64997 , n64650 );
and ( n593009 , n64973 , n64648 );
nor ( n593010 , n65685 , n593009 );
xnor ( n65688 , n593010 , n591902 );
and ( n593012 , n593006 , n65688 );
and ( n65690 , n65679 , n65688 );
or ( n65691 , n593007 , n593012 , n65690 );
and ( n65692 , n64533 , n592486 );
and ( n65693 , n591851 , n592484 );
nor ( n65694 , n65692 , n65693 );
xnor ( n65695 , n65694 , n64990 );
and ( n593019 , n65691 , n65695 );
xor ( n65697 , n65578 , n592905 );
xor ( n593021 , n65697 , n592908 );
and ( n593022 , n65695 , n593021 );
and ( n65700 , n65691 , n593021 );
or ( n593024 , n593019 , n593022 , n65700 );
and ( n593025 , n65675 , n593024 );
xor ( n65703 , n592911 , n592918 );
xor ( n593027 , n65703 , n592921 );
and ( n65705 , n593024 , n593027 );
and ( n65706 , n65675 , n593027 );
or ( n593030 , n593025 , n65705 , n65706 );
and ( n65708 , n65384 , n64491 );
and ( n593032 , n592645 , n64489 );
nor ( n65710 , n65708 , n593032 );
xnor ( n65711 , n65710 , n64448 );
and ( n65712 , n592806 , n64456 );
and ( n593036 , n65493 , n64454 );
nor ( n593037 , n65712 , n593036 );
xnor ( n65715 , n593037 , n591786 );
and ( n593039 , n65711 , n65715 );
xor ( n65717 , n592955 , n65638 );
xor ( n65718 , n65717 , n65641 );
and ( n593042 , n65715 , n65718 );
and ( n593043 , n65711 , n65718 );
or ( n65721 , n593039 , n593042 , n593043 );
and ( n593045 , n64586 , n592486 );
and ( n593046 , n64533 , n592484 );
nor ( n65724 , n593045 , n593046 );
xnor ( n593048 , n65724 , n64990 );
and ( n65726 , n65721 , n593048 );
and ( n65727 , n64630 , n592340 );
and ( n65728 , n64591 , n65015 );
nor ( n65729 , n65727 , n65728 );
xnor ( n593053 , n65729 , n64847 );
and ( n65731 , n593048 , n593053 );
and ( n593055 , n65721 , n593053 );
or ( n65733 , n65726 , n65731 , n593055 );
and ( n65734 , n64838 , n64744 );
and ( n65735 , n592094 , n64742 );
nor ( n65736 , n65734 , n65735 );
xnor ( n65737 , n65736 , n64623 );
and ( n65738 , n64973 , n64650 );
and ( n65739 , n64854 , n64648 );
nor ( n65740 , n65738 , n65739 );
xnor ( n65741 , n65740 , n591902 );
xor ( n65742 , n65737 , n65741 );
and ( n65743 , n592404 , n64559 );
and ( n65744 , n64997 , n591880 );
nor ( n65745 , n65743 , n65744 );
xnor ( n65746 , n65745 , n64521 );
xor ( n65747 , n65742 , n65746 );
and ( n65748 , n65733 , n65747 );
and ( n65749 , n592976 , n65657 );
and ( n65750 , n65657 , n65659 );
and ( n65751 , n592976 , n65659 );
or ( n65752 , n65749 , n65750 , n65751 );
and ( n65753 , n64591 , n592340 );
and ( n65754 , n64586 , n65015 );
nor ( n65755 , n65753 , n65754 );
xnor ( n65756 , n65755 , n64847 );
xor ( n65757 , n65752 , n65756 );
and ( n65758 , n64683 , n64862 );
and ( n65759 , n64630 , n64860 );
nor ( n65760 , n65758 , n65759 );
xnor ( n65761 , n65760 , n64764 );
xor ( n65762 , n65757 , n65761 );
and ( n65763 , n65747 , n65762 );
and ( n65764 , n65733 , n65762 );
or ( n65765 , n65748 , n65763 , n65764 );
and ( n65766 , n65737 , n65741 );
and ( n65767 , n65741 , n65746 );
and ( n65768 , n65737 , n65746 );
or ( n65769 , n65766 , n65767 , n65768 );
and ( n65770 , n64466 , n592683 );
and ( n65771 , n64450 , n592681 );
nor ( n65772 , n65770 , n65771 );
xnor ( n65773 , n65772 , n592475 );
xor ( n65774 , n65769 , n65773 );
and ( n65775 , n591851 , n592486 );
and ( n65776 , n64501 , n592484 );
nor ( n65777 , n65775 , n65776 );
xnor ( n65778 , n65777 , n64990 );
xor ( n65779 , n65774 , n65778 );
and ( n65780 , n65765 , n65779 );
and ( n65781 , n65752 , n65756 );
and ( n65782 , n65756 , n65761 );
and ( n593106 , n65752 , n65761 );
or ( n65784 , n65781 , n65782 , n593106 );
xor ( n65785 , n65458 , n592785 );
xor ( n65786 , n65785 , n592790 );
xor ( n65787 , n65784 , n65786 );
xor ( n65788 , n65528 , n65532 );
xor ( n65789 , n65788 , n65537 );
xor ( n65790 , n65787 , n65789 );
and ( n65791 , n65779 , n65790 );
and ( n65792 , n65765 , n65790 );
or ( n65793 , n65780 , n65791 , n65792 );
and ( n65794 , n593030 , n65793 );
xor ( n593118 , n65601 , n592926 );
xor ( n65796 , n593118 , n592929 );
and ( n593120 , n65793 , n65796 );
and ( n593121 , n593030 , n65796 );
or ( n65799 , n65794 , n593120 , n593121 );
and ( n65800 , n65769 , n65773 );
and ( n65801 , n65773 , n65778 );
and ( n65802 , n65769 , n65778 );
or ( n593126 , n65800 , n65801 , n65802 );
and ( n65804 , n65784 , n65786 );
and ( n593128 , n65786 , n65789 );
and ( n593129 , n65784 , n65789 );
or ( n65807 , n65804 , n593128 , n593129 );
and ( n593131 , n593126 , n65807 );
xor ( n593132 , n592863 , n65542 );
xor ( n65810 , n593132 , n65545 );
and ( n593134 , n65807 , n65810 );
and ( n593135 , n593126 , n65810 );
or ( n65813 , n593131 , n593134 , n593135 );
and ( n593137 , n65799 , n65813 );
xor ( n65815 , n592932 , n65611 );
xor ( n593139 , n65815 , n65614 );
and ( n593140 , n65813 , n593139 );
and ( n65818 , n65799 , n593139 );
or ( n593142 , n593137 , n593140 , n65818 );
and ( n593143 , n592952 , n593142 );
xor ( n65821 , n592952 , n593142 );
xor ( n65822 , n65799 , n65813 );
xor ( n65823 , n65822 , n593139 );
and ( n65824 , n592645 , n64559 );
and ( n65825 , n592468 , n591880 );
nor ( n65826 , n65824 , n65825 );
xnor ( n65827 , n65826 , n64521 );
and ( n65828 , n65493 , n64491 );
and ( n65829 , n65384 , n64489 );
nor ( n65830 , n65828 , n65829 );
xnor ( n593154 , n65830 , n64448 );
and ( n65832 , n65827 , n593154 );
buf ( n593156 , n591759 );
buf ( n65834 , n591760 );
and ( n65835 , n593156 , n65834 );
not ( n593159 , n65835 );
and ( n593160 , n592957 , n593159 );
not ( n65838 , n593160 );
and ( n593162 , n65630 , n64456 );
and ( n65840 , n65640 , n64454 );
nor ( n65841 , n593162 , n65840 );
xnor ( n65842 , n65841 , n591786 );
and ( n65843 , n65838 , n65842 );
buf ( n65844 , n591693 );
and ( n65845 , n65844 , n64451 );
and ( n65846 , n65842 , n65845 );
and ( n65847 , n65838 , n65845 );
or ( n65848 , n65843 , n65846 , n65847 );
and ( n593172 , n65640 , n64456 );
and ( n593173 , n592806 , n64454 );
nor ( n65851 , n593172 , n593173 );
xnor ( n593175 , n65851 , n591786 );
xor ( n593176 , n65848 , n593175 );
not ( n593177 , n592954 );
xor ( n593178 , n593176 , n593177 );
and ( n65856 , n593154 , n593178 );
and ( n593180 , n65827 , n593178 );
or ( n593181 , n65832 , n65856 , n593180 );
and ( n65859 , n64591 , n592486 );
and ( n593183 , n64586 , n592484 );
nor ( n593184 , n65859 , n593183 );
xnor ( n65862 , n593184 , n64990 );
and ( n593186 , n593181 , n65862 );
and ( n593187 , n64683 , n592340 );
and ( n65865 , n64630 , n65015 );
nor ( n593189 , n593187 , n65865 );
xnor ( n65867 , n593189 , n64847 );
and ( n65868 , n65862 , n65867 );
and ( n65869 , n593181 , n65867 );
or ( n593193 , n593186 , n65868 , n65869 );
and ( n65871 , n64466 , n65592 );
and ( n593195 , n64450 , n592913 );
nor ( n593196 , n65871 , n593195 );
xnor ( n65874 , n593196 , n592638 );
and ( n593198 , n593193 , n65874 );
and ( n65876 , n591851 , n592683 );
and ( n65877 , n64501 , n592681 );
nor ( n65878 , n65876 , n65877 );
xnor ( n65879 , n65878 , n592475 );
and ( n65880 , n65874 , n65879 );
and ( n65881 , n593193 , n65879 );
or ( n65882 , n593198 , n65880 , n65881 );
xor ( n65883 , n65679 , n593006 );
xor ( n593207 , n65883 , n65688 );
xor ( n65885 , n65721 , n593048 );
xor ( n593209 , n65885 , n593053 );
and ( n65887 , n593207 , n593209 );
xor ( n65888 , n592967 , n65648 );
xor ( n593212 , n65888 , n592983 );
and ( n65890 , n593209 , n593212 );
and ( n593214 , n593207 , n593212 );
or ( n593215 , n65887 , n65890 , n593214 );
and ( n65893 , n65882 , n593215 );
xor ( n593217 , n65733 , n65747 );
xor ( n65895 , n593217 , n65762 );
and ( n593219 , n593215 , n65895 );
and ( n593220 , n65882 , n65895 );
or ( n65898 , n65893 , n593219 , n593220 );
and ( n593222 , n65848 , n593175 );
and ( n593223 , n593175 , n593177 );
and ( n65901 , n65848 , n593177 );
or ( n593225 , n593222 , n593223 , n65901 );
and ( n593226 , n592404 , n64650 );
and ( n65904 , n64997 , n64648 );
nor ( n593228 , n593226 , n65904 );
xnor ( n593229 , n593228 , n591902 );
and ( n65907 , n593225 , n593229 );
and ( n593231 , n592468 , n64559 );
and ( n593232 , n592478 , n591880 );
nor ( n65910 , n593231 , n593232 );
xnor ( n593234 , n65910 , n64521 );
and ( n593235 , n593229 , n593234 );
and ( n65913 , n593225 , n593234 );
or ( n593237 , n65907 , n593235 , n65913 );
and ( n65915 , n64838 , n64862 );
and ( n65916 , n592094 , n64860 );
nor ( n65917 , n65915 , n65916 );
xnor ( n65918 , n65917 , n64764 );
and ( n65919 , n64973 , n64744 );
and ( n593243 , n64854 , n64742 );
nor ( n593244 , n65919 , n593243 );
xnor ( n65922 , n593244 , n64623 );
and ( n593246 , n65918 , n65922 );
xor ( n65924 , n65711 , n65715 );
xor ( n65925 , n65924 , n65718 );
and ( n65926 , n65922 , n65925 );
and ( n65927 , n65918 , n65925 );
or ( n65928 , n593246 , n65926 , n65927 );
and ( n65929 , n593237 , n65928 );
xor ( n65930 , n592635 , n65486 );
xor ( n593254 , n65486 , n65487 );
not ( n65932 , n593254 );
and ( n593256 , n65930 , n65932 );
and ( n65934 , n64458 , n593256 );
not ( n593258 , n65934 );
xnor ( n593259 , n593258 , n65490 );
and ( n65937 , n65928 , n593259 );
and ( n593261 , n593237 , n593259 );
or ( n65939 , n65929 , n65937 , n593261 );
xor ( n65940 , n592986 , n65667 );
xor ( n593264 , n65940 , n592995 );
and ( n65942 , n65939 , n593264 );
xor ( n593266 , n65691 , n65695 );
xor ( n593267 , n593266 , n593021 );
and ( n65945 , n593264 , n593267 );
and ( n65946 , n65939 , n593267 );
or ( n593270 , n65942 , n65945 , n65946 );
and ( n65948 , n65898 , n593270 );
xor ( n65949 , n65675 , n593024 );
xor ( n593273 , n65949 , n593027 );
and ( n593274 , n593270 , n593273 );
and ( n65952 , n65898 , n593273 );
or ( n593276 , n65948 , n593274 , n65952 );
xor ( n593277 , n593030 , n65793 );
xor ( n65955 , n593277 , n65796 );
and ( n593279 , n593276 , n65955 );
xor ( n65957 , n593126 , n65807 );
xor ( n65958 , n65957 , n65810 );
and ( n65959 , n65955 , n65958 );
and ( n65960 , n593276 , n65958 );
or ( n593284 , n593279 , n65959 , n65960 );
and ( n65962 , n65823 , n593284 );
xor ( n593286 , n65823 , n593284 );
xor ( n593287 , n593276 , n65955 );
xor ( n593288 , n593287 , n65958 );
and ( n593289 , n65640 , n64491 );
and ( n65967 , n592806 , n64489 );
nor ( n593291 , n593289 , n65967 );
xnor ( n593292 , n593291 , n64448 );
and ( n65970 , n65844 , n64456 );
and ( n593294 , n65630 , n64454 );
nor ( n593295 , n65970 , n593294 );
xnor ( n65973 , n593295 , n591786 );
and ( n593297 , n593292 , n65973 );
buf ( n593298 , n591694 );
and ( n65976 , n593298 , n64451 );
not ( n593300 , n65976 );
and ( n65978 , n65973 , n593300 );
and ( n593302 , n593292 , n593300 );
or ( n65980 , n593297 , n65978 , n593302 );
and ( n593304 , n592468 , n64650 );
and ( n65982 , n592478 , n64648 );
nor ( n65983 , n593304 , n65982 );
xnor ( n65984 , n65983 , n591902 );
and ( n65985 , n65980 , n65984 );
xor ( n65986 , n65838 , n65842 );
xor ( n65987 , n65986 , n65845 );
and ( n65988 , n65984 , n65987 );
and ( n593312 , n65980 , n65987 );
or ( n65990 , n65985 , n65988 , n593312 );
and ( n65991 , n64854 , n64862 );
and ( n593315 , n64838 , n64860 );
nor ( n593316 , n65991 , n593315 );
xnor ( n593317 , n593316 , n64764 );
and ( n65995 , n65990 , n593317 );
and ( n593319 , n64997 , n64744 );
and ( n593320 , n64973 , n64742 );
nor ( n65998 , n593319 , n593320 );
xnor ( n593322 , n65998 , n64623 );
and ( n593323 , n593317 , n593322 );
and ( n66001 , n65990 , n593322 );
or ( n593325 , n65995 , n593323 , n66001 );
and ( n593326 , n64450 , n593256 );
and ( n66004 , n64458 , n593254 );
nor ( n593328 , n593326 , n66004 );
xnor ( n593329 , n593328 , n65490 );
and ( n66007 , n593325 , n593329 );
and ( n593331 , n64501 , n65592 );
and ( n66009 , n64466 , n592913 );
nor ( n66010 , n593331 , n66009 );
xnor ( n593334 , n66010 , n592638 );
and ( n66012 , n593329 , n593334 );
and ( n593336 , n593325 , n593334 );
or ( n593337 , n66007 , n66012 , n593336 );
buf ( n66015 , n65976 );
and ( n593339 , n65384 , n64559 );
and ( n593340 , n592645 , n591880 );
nor ( n66018 , n593339 , n593340 );
xnor ( n593342 , n66018 , n64521 );
and ( n593343 , n66015 , n593342 );
and ( n66021 , n592806 , n64491 );
and ( n593345 , n65493 , n64489 );
nor ( n66023 , n66021 , n593345 );
xnor ( n66024 , n66023 , n64448 );
and ( n593348 , n593342 , n66024 );
and ( n66026 , n66015 , n66024 );
or ( n593350 , n593343 , n593348 , n66026 );
and ( n66028 , n592094 , n592340 );
and ( n66029 , n64683 , n65015 );
nor ( n66030 , n66028 , n66029 );
xnor ( n66031 , n66030 , n64847 );
and ( n66032 , n593350 , n66031 );
and ( n66033 , n592478 , n64650 );
and ( n593357 , n592404 , n64648 );
nor ( n66035 , n66033 , n593357 );
xnor ( n593359 , n66035 , n591902 );
and ( n66037 , n66031 , n593359 );
and ( n593361 , n593350 , n593359 );
or ( n593362 , n66032 , n66037 , n593361 );
and ( n66040 , n64533 , n592683 );
and ( n593364 , n591851 , n592681 );
nor ( n593365 , n66040 , n593364 );
xnor ( n66043 , n593365 , n592475 );
and ( n593367 , n593362 , n66043 );
xor ( n593368 , n593225 , n593229 );
xor ( n66046 , n593368 , n593234 );
and ( n593370 , n66043 , n66046 );
and ( n593371 , n593362 , n66046 );
or ( n66049 , n593367 , n593370 , n593371 );
and ( n593373 , n593337 , n66049 );
xor ( n66051 , n593237 , n65928 );
xor ( n66052 , n66051 , n593259 );
and ( n66053 , n66049 , n66052 );
and ( n66054 , n593337 , n66052 );
or ( n593378 , n593373 , n66053 , n66054 );
and ( n66056 , n64586 , n592683 );
and ( n593380 , n64533 , n592681 );
nor ( n66058 , n66056 , n593380 );
xnor ( n66059 , n66058 , n592475 );
and ( n593383 , n64630 , n592486 );
and ( n66061 , n64591 , n592484 );
nor ( n593385 , n593383 , n66061 );
xnor ( n66063 , n593385 , n64990 );
and ( n66064 , n66059 , n66063 );
xor ( n66065 , n65827 , n593154 );
xor ( n66066 , n66065 , n593178 );
and ( n66067 , n66063 , n66066 );
and ( n593391 , n66059 , n66066 );
or ( n593392 , n66064 , n66067 , n593391 );
xor ( n66070 , n593181 , n65862 );
xor ( n593394 , n66070 , n65867 );
and ( n593395 , n593392 , n593394 );
xor ( n66073 , n65918 , n65922 );
xor ( n593397 , n66073 , n65925 );
and ( n593398 , n593394 , n593397 );
and ( n593399 , n593392 , n593397 );
or ( n66077 , n593395 , n593398 , n593399 );
xor ( n593401 , n593193 , n65874 );
xor ( n66079 , n593401 , n65879 );
and ( n593403 , n66077 , n66079 );
xor ( n66081 , n593207 , n593209 );
xor ( n593405 , n66081 , n593212 );
and ( n593406 , n66079 , n593405 );
and ( n66084 , n66077 , n593405 );
or ( n593408 , n593403 , n593406 , n66084 );
and ( n66086 , n593378 , n593408 );
xor ( n66087 , n65939 , n593264 );
xor ( n66088 , n66087 , n593267 );
and ( n593412 , n593408 , n66088 );
and ( n66090 , n593378 , n66088 );
or ( n593414 , n66086 , n593412 , n66090 );
xor ( n593415 , n65765 , n65779 );
xor ( n593416 , n593415 , n65790 );
and ( n593417 , n593414 , n593416 );
xor ( n66095 , n65898 , n593270 );
xor ( n593419 , n66095 , n593273 );
and ( n593420 , n593416 , n593419 );
and ( n66098 , n593414 , n593419 );
or ( n593422 , n593417 , n593420 , n66098 );
and ( n66100 , n593288 , n593422 );
xor ( n593424 , n593288 , n593422 );
xor ( n593425 , n593414 , n593416 );
xor ( n593426 , n593425 , n593419 );
buf ( n66104 , n591696 );
and ( n593428 , n66104 , n64451 );
buf ( n593429 , n593428 );
buf ( n66107 , n591761 );
buf ( n593431 , n591762 );
and ( n593432 , n66107 , n593431 );
not ( n66110 , n593432 );
and ( n593434 , n65834 , n66110 );
not ( n66112 , n593434 );
and ( n66113 , n593429 , n66112 );
buf ( n593437 , n591695 );
and ( n66115 , n593437 , n64451 );
and ( n593439 , n66112 , n66115 );
and ( n593440 , n593429 , n66115 );
or ( n593441 , n66113 , n593439 , n593440 );
and ( n66119 , n65493 , n64559 );
and ( n593443 , n65384 , n591880 );
nor ( n66121 , n66119 , n593443 );
xnor ( n593445 , n66121 , n64521 );
and ( n66123 , n593441 , n593445 );
xor ( n593447 , n593292 , n65973 );
xor ( n66125 , n593447 , n593300 );
and ( n66126 , n593445 , n66125 );
and ( n66127 , n593441 , n66125 );
or ( n66128 , n66123 , n66126 , n66127 );
and ( n593452 , n592404 , n64744 );
and ( n593453 , n64997 , n64742 );
nor ( n66131 , n593452 , n593453 );
xnor ( n593455 , n66131 , n64623 );
and ( n593456 , n66128 , n593455 );
xor ( n66134 , n66015 , n593342 );
xor ( n593458 , n66134 , n66024 );
and ( n593459 , n593455 , n593458 );
and ( n593460 , n66128 , n593458 );
or ( n66138 , n593456 , n593459 , n593460 );
xor ( n593462 , n65487 , n65633 );
xor ( n66140 , n65633 , n592957 );
not ( n66141 , n66140 );
and ( n66142 , n593462 , n66141 );
and ( n66143 , n64458 , n66142 );
not ( n66144 , n66143 );
xnor ( n66145 , n66144 , n592960 );
and ( n66146 , n66138 , n66145 );
and ( n66147 , n591851 , n65592 );
and ( n593471 , n64501 , n592913 );
nor ( n66149 , n66147 , n593471 );
xnor ( n593473 , n66149 , n592638 );
and ( n66151 , n66145 , n593473 );
and ( n593475 , n66138 , n593473 );
or ( n66153 , n66146 , n66151 , n593475 );
and ( n593477 , n64591 , n592683 );
and ( n593478 , n64586 , n592681 );
nor ( n593479 , n593477 , n593478 );
xnor ( n66157 , n593479 , n592475 );
and ( n593481 , n64838 , n592340 );
and ( n66159 , n592094 , n65015 );
nor ( n593483 , n593481 , n66159 );
xnor ( n66161 , n593483 , n64847 );
and ( n593485 , n66157 , n66161 );
and ( n66163 , n64973 , n64862 );
and ( n593487 , n64854 , n64860 );
nor ( n66165 , n66163 , n593487 );
xnor ( n593489 , n66165 , n64764 );
and ( n593490 , n66161 , n593489 );
and ( n66168 , n66157 , n593489 );
or ( n593492 , n593485 , n593490 , n66168 );
and ( n66170 , n64466 , n593256 );
and ( n593494 , n64450 , n593254 );
nor ( n66172 , n66170 , n593494 );
xnor ( n593496 , n66172 , n65490 );
and ( n593497 , n593492 , n593496 );
xor ( n593498 , n65990 , n593317 );
xor ( n66176 , n593498 , n593322 );
and ( n593500 , n593496 , n66176 );
and ( n66178 , n593492 , n66176 );
or ( n593502 , n593497 , n593500 , n66178 );
and ( n593503 , n66153 , n593502 );
xor ( n66181 , n593362 , n66043 );
xor ( n593505 , n66181 , n66046 );
and ( n66183 , n593502 , n593505 );
and ( n66184 , n66153 , n593505 );
or ( n66185 , n593503 , n66183 , n66184 );
buf ( n66186 , n591763 );
buf ( n66187 , n591764 );
and ( n66188 , n66186 , n66187 );
not ( n593512 , n66188 );
and ( n66190 , n593431 , n593512 );
not ( n593514 , n66190 );
and ( n593515 , n66104 , n64456 );
and ( n66193 , n593437 , n64454 );
nor ( n593517 , n593515 , n66193 );
xnor ( n66195 , n593517 , n591786 );
and ( n593519 , n593514 , n66195 );
buf ( n593520 , n591697 );
and ( n66198 , n593520 , n64451 );
and ( n593522 , n66195 , n66198 );
and ( n593523 , n593514 , n66198 );
or ( n593524 , n593519 , n593522 , n593523 );
and ( n593525 , n593437 , n64456 );
and ( n66203 , n593298 , n64454 );
nor ( n593527 , n593525 , n66203 );
xnor ( n593528 , n593527 , n591786 );
and ( n66206 , n593524 , n593528 );
not ( n593530 , n593428 );
and ( n66208 , n593528 , n593530 );
and ( n593532 , n593524 , n593530 );
or ( n593533 , n66206 , n66208 , n593532 );
and ( n66211 , n65384 , n64650 );
and ( n593535 , n592645 , n64648 );
nor ( n593536 , n66211 , n593535 );
xnor ( n66214 , n593536 , n591902 );
and ( n593538 , n593533 , n66214 );
and ( n593539 , n592806 , n64559 );
and ( n66217 , n65493 , n591880 );
nor ( n593541 , n593539 , n66217 );
xnor ( n66219 , n593541 , n64521 );
and ( n66220 , n66214 , n66219 );
and ( n66221 , n593533 , n66219 );
or ( n593545 , n593538 , n66220 , n66221 );
and ( n593546 , n65630 , n64491 );
and ( n66224 , n65640 , n64489 );
nor ( n593548 , n593546 , n66224 );
xnor ( n66226 , n593548 , n64448 );
and ( n593550 , n593298 , n64456 );
and ( n593551 , n65844 , n64454 );
nor ( n66229 , n593550 , n593551 );
xnor ( n593553 , n66229 , n591786 );
and ( n593554 , n66226 , n593553 );
xor ( n66232 , n593429 , n66112 );
xor ( n593556 , n66232 , n66115 );
and ( n593557 , n593553 , n593556 );
and ( n66235 , n66226 , n593556 );
or ( n593559 , n593554 , n593557 , n66235 );
and ( n66237 , n593545 , n593559 );
and ( n593561 , n592645 , n64650 );
and ( n593562 , n592468 , n64648 );
nor ( n66240 , n593561 , n593562 );
xnor ( n593564 , n66240 , n591902 );
and ( n66242 , n593559 , n593564 );
and ( n593566 , n593545 , n593564 );
or ( n66244 , n66237 , n66242 , n593566 );
and ( n593568 , n64683 , n592486 );
and ( n593569 , n64630 , n592484 );
nor ( n66247 , n593568 , n593569 );
xnor ( n66248 , n66247 , n64990 );
and ( n66249 , n66244 , n66248 );
xor ( n66250 , n65980 , n65984 );
xor ( n593574 , n66250 , n65987 );
and ( n593575 , n66248 , n593574 );
and ( n66253 , n66244 , n593574 );
or ( n593577 , n66249 , n593575 , n66253 );
xor ( n66255 , n593350 , n66031 );
xor ( n593579 , n66255 , n593359 );
and ( n593580 , n593577 , n593579 );
xor ( n66258 , n66059 , n66063 );
xor ( n593582 , n66258 , n66066 );
and ( n66260 , n593579 , n593582 );
and ( n66261 , n593577 , n593582 );
or ( n66262 , n593580 , n66260 , n66261 );
xor ( n66263 , n593325 , n593329 );
xor ( n66264 , n66263 , n593334 );
and ( n593588 , n66262 , n66264 );
xor ( n66266 , n593392 , n593394 );
xor ( n593590 , n66266 , n593397 );
and ( n593591 , n66264 , n593590 );
and ( n593592 , n66262 , n593590 );
or ( n593593 , n593588 , n593591 , n593592 );
and ( n593594 , n66185 , n593593 );
xor ( n66272 , n593337 , n66049 );
xor ( n593596 , n66272 , n66052 );
and ( n593597 , n593593 , n593596 );
and ( n66275 , n66185 , n593596 );
or ( n66276 , n593594 , n593597 , n66275 );
xor ( n593600 , n65882 , n593215 );
xor ( n66278 , n593600 , n65895 );
and ( n593602 , n66276 , n66278 );
xor ( n593603 , n593378 , n593408 );
xor ( n66281 , n593603 , n66088 );
and ( n593605 , n66278 , n66281 );
and ( n593606 , n66276 , n66281 );
or ( n66284 , n593602 , n593605 , n593606 );
and ( n593608 , n593426 , n66284 );
xor ( n66286 , n593426 , n66284 );
xor ( n593610 , n66276 , n66278 );
xor ( n66288 , n593610 , n66281 );
and ( n593612 , n592094 , n592486 );
and ( n593613 , n64683 , n592484 );
nor ( n66291 , n593612 , n593613 );
xnor ( n593615 , n66291 , n64990 );
and ( n593616 , n64997 , n64862 );
and ( n66294 , n64973 , n64860 );
nor ( n66295 , n593616 , n66294 );
xnor ( n593619 , n66295 , n64764 );
and ( n593620 , n593615 , n593619 );
and ( n66298 , n592478 , n64744 );
and ( n593622 , n592404 , n64742 );
nor ( n66300 , n66298 , n593622 );
xnor ( n593624 , n66300 , n64623 );
and ( n66302 , n593619 , n593624 );
and ( n593626 , n593615 , n593624 );
or ( n593627 , n593620 , n66302 , n593626 );
and ( n66305 , n64501 , n593256 );
and ( n66306 , n64466 , n593254 );
nor ( n593630 , n66305 , n66306 );
xnor ( n66308 , n593630 , n65490 );
and ( n593632 , n593627 , n66308 );
and ( n593633 , n64533 , n65592 );
and ( n66311 , n591851 , n592913 );
nor ( n593635 , n593633 , n66311 );
xnor ( n593636 , n593635 , n592638 );
and ( n66314 , n66308 , n593636 );
and ( n593638 , n593627 , n593636 );
or ( n593639 , n593632 , n66314 , n593638 );
and ( n593640 , n64450 , n66142 );
and ( n66318 , n64458 , n66140 );
nor ( n593642 , n593640 , n66318 );
xnor ( n593643 , n593642 , n592960 );
xor ( n593644 , n66157 , n66161 );
xor ( n66322 , n593644 , n593489 );
and ( n593646 , n593643 , n66322 );
xor ( n593647 , n66128 , n593455 );
xor ( n66325 , n593647 , n593458 );
and ( n593649 , n66322 , n66325 );
and ( n593650 , n593643 , n66325 );
or ( n66328 , n593646 , n593649 , n593650 );
and ( n593652 , n593639 , n66328 );
xor ( n593653 , n66138 , n66145 );
xor ( n593654 , n593653 , n593473 );
and ( n593655 , n66328 , n593654 );
and ( n593656 , n593639 , n593654 );
or ( n66334 , n593652 , n593655 , n593656 );
and ( n66335 , n64586 , n65592 );
and ( n593659 , n64533 , n592913 );
nor ( n593660 , n66335 , n593659 );
xnor ( n66338 , n593660 , n592638 );
and ( n593662 , n64630 , n592683 );
and ( n593663 , n64591 , n592681 );
nor ( n66341 , n593662 , n593663 );
xnor ( n593665 , n66341 , n592475 );
and ( n66343 , n66338 , n593665 );
xor ( n593667 , n593545 , n593559 );
xor ( n593668 , n593667 , n593564 );
and ( n593669 , n593665 , n593668 );
and ( n593670 , n66338 , n593668 );
or ( n593671 , n66343 , n593669 , n593670 );
and ( n66349 , n593520 , n64456 );
and ( n66350 , n66104 , n64454 );
nor ( n66351 , n66349 , n66350 );
xnor ( n66352 , n66351 , n591786 );
buf ( n66353 , n66352 );
and ( n593677 , n65630 , n64559 );
and ( n593678 , n65640 , n591880 );
nor ( n593679 , n593677 , n593678 );
xnor ( n593680 , n593679 , n64521 );
and ( n66358 , n66353 , n593680 );
and ( n593682 , n593298 , n64491 );
and ( n593683 , n65844 , n64489 );
nor ( n66361 , n593682 , n593683 );
xnor ( n593685 , n66361 , n64448 );
and ( n593686 , n593680 , n593685 );
and ( n593687 , n66353 , n593685 );
or ( n66365 , n66358 , n593686 , n593687 );
and ( n593689 , n65640 , n64559 );
and ( n593690 , n592806 , n591880 );
nor ( n66368 , n593689 , n593690 );
xnor ( n593692 , n66368 , n64521 );
and ( n593693 , n66365 , n593692 );
and ( n593694 , n65844 , n64491 );
and ( n593695 , n65630 , n64489 );
nor ( n66373 , n593694 , n593695 );
xnor ( n593697 , n66373 , n64448 );
and ( n593698 , n593692 , n593697 );
and ( n593699 , n66365 , n593697 );
or ( n66377 , n593693 , n593698 , n593699 );
and ( n593701 , n592468 , n64744 );
and ( n593702 , n592478 , n64742 );
nor ( n593703 , n593701 , n593702 );
xnor ( n66381 , n593703 , n64623 );
and ( n593705 , n66377 , n66381 );
xor ( n66383 , n66226 , n593553 );
xor ( n66384 , n66383 , n593556 );
and ( n593708 , n66381 , n66384 );
and ( n593709 , n66377 , n66384 );
or ( n593710 , n593705 , n593708 , n593709 );
and ( n66388 , n64854 , n592340 );
and ( n593712 , n64838 , n65015 );
nor ( n66390 , n66388 , n593712 );
xnor ( n593714 , n66390 , n64847 );
and ( n593715 , n593710 , n593714 );
xor ( n593716 , n593441 , n593445 );
xor ( n66394 , n593716 , n66125 );
and ( n593718 , n593714 , n66394 );
and ( n66396 , n593710 , n66394 );
or ( n593720 , n593715 , n593718 , n66396 );
and ( n66398 , n593671 , n593720 );
xor ( n593722 , n66244 , n66248 );
xor ( n593723 , n593722 , n593574 );
and ( n593724 , n593720 , n593723 );
and ( n66402 , n593671 , n593723 );
or ( n593726 , n66398 , n593724 , n66402 );
xor ( n66404 , n593492 , n593496 );
xor ( n66405 , n66404 , n66176 );
and ( n66406 , n593726 , n66405 );
xor ( n66407 , n593577 , n593579 );
xor ( n66408 , n66407 , n593582 );
and ( n593732 , n66405 , n66408 );
and ( n66410 , n593726 , n66408 );
or ( n593734 , n66406 , n593732 , n66410 );
and ( n593735 , n66334 , n593734 );
xor ( n593736 , n66153 , n593502 );
xor ( n66414 , n593736 , n593505 );
and ( n593738 , n593734 , n66414 );
and ( n593739 , n66334 , n66414 );
or ( n593740 , n593735 , n593738 , n593739 );
xor ( n593741 , n66185 , n593593 );
xor ( n66419 , n593741 , n593596 );
and ( n593743 , n593740 , n66419 );
xor ( n593744 , n66077 , n66079 );
xor ( n593745 , n593744 , n593405 );
and ( n593746 , n66419 , n593745 );
and ( n66424 , n593740 , n593745 );
or ( n593748 , n593743 , n593746 , n66424 );
and ( n593749 , n66288 , n593748 );
xor ( n593750 , n66288 , n593748 );
xor ( n593751 , n593740 , n66419 );
xor ( n66429 , n593751 , n593745 );
and ( n593753 , n592645 , n64744 );
and ( n593754 , n592468 , n64742 );
nor ( n593755 , n593753 , n593754 );
xnor ( n66433 , n593755 , n64623 );
and ( n593757 , n65493 , n64650 );
and ( n66435 , n65384 , n64648 );
nor ( n593759 , n593757 , n66435 );
xnor ( n66437 , n593759 , n591902 );
and ( n593761 , n66433 , n66437 );
xor ( n593762 , n593524 , n593528 );
xor ( n593763 , n593762 , n593530 );
and ( n593764 , n66437 , n593763 );
and ( n66442 , n66433 , n593763 );
or ( n593766 , n593761 , n593764 , n66442 );
and ( n593767 , n592404 , n64862 );
and ( n593768 , n64997 , n64860 );
nor ( n66446 , n593767 , n593768 );
xnor ( n593770 , n66446 , n64764 );
and ( n66448 , n593766 , n593770 );
xor ( n66449 , n593533 , n66214 );
xor ( n593773 , n66449 , n66219 );
and ( n66451 , n593770 , n593773 );
and ( n593775 , n593766 , n593773 );
or ( n593776 , n66448 , n66451 , n593775 );
xor ( n66454 , n592957 , n593156 );
xor ( n593778 , n593156 , n65834 );
not ( n593779 , n593778 );
and ( n66457 , n66454 , n593779 );
and ( n593781 , n64458 , n66457 );
not ( n593782 , n593781 );
xnor ( n593783 , n593782 , n593160 );
and ( n66461 , n593776 , n593783 );
and ( n593785 , n591851 , n593256 );
and ( n593786 , n64501 , n593254 );
nor ( n593787 , n593785 , n593786 );
xnor ( n66465 , n593787 , n65490 );
and ( n593789 , n593783 , n66465 );
and ( n593790 , n593776 , n66465 );
or ( n66468 , n66461 , n593789 , n593790 );
and ( n593792 , n64591 , n65592 );
and ( n593793 , n64586 , n592913 );
nor ( n66471 , n593792 , n593793 );
xnor ( n593795 , n66471 , n592638 );
and ( n66473 , n64838 , n592486 );
and ( n593797 , n592094 , n592484 );
nor ( n593798 , n66473 , n593797 );
xnor ( n66476 , n593798 , n64990 );
and ( n593800 , n593795 , n66476 );
and ( n593801 , n64973 , n592340 );
and ( n66479 , n64854 , n65015 );
nor ( n593803 , n593801 , n66479 );
xnor ( n66481 , n593803 , n64847 );
and ( n593805 , n66476 , n66481 );
and ( n593806 , n593795 , n66481 );
or ( n593807 , n593800 , n593805 , n593806 );
and ( n66485 , n64466 , n66142 );
and ( n593809 , n64450 , n66140 );
nor ( n593810 , n66485 , n593809 );
xnor ( n66488 , n593810 , n592960 );
and ( n66489 , n593807 , n66488 );
xor ( n593813 , n593710 , n593714 );
xor ( n593814 , n593813 , n66394 );
and ( n593815 , n66488 , n593814 );
and ( n66493 , n593807 , n593814 );
or ( n593817 , n66489 , n593815 , n66493 );
and ( n66495 , n66468 , n593817 );
xor ( n593819 , n593627 , n66308 );
xor ( n593820 , n593819 , n593636 );
and ( n593821 , n593817 , n593820 );
and ( n66499 , n66468 , n593820 );
or ( n593823 , n66495 , n593821 , n66499 );
and ( n593824 , n593437 , n64491 );
and ( n66502 , n593298 , n64489 );
nor ( n66503 , n593824 , n66502 );
xnor ( n593827 , n66503 , n64448 );
not ( n593828 , n66352 );
and ( n593829 , n593827 , n593828 );
buf ( n66507 , n591698 );
and ( n593831 , n66507 , n64451 );
and ( n593832 , n593828 , n593831 );
and ( n66510 , n593827 , n593831 );
or ( n593834 , n593829 , n593832 , n66510 );
and ( n593835 , n592806 , n64650 );
and ( n66513 , n65493 , n64648 );
nor ( n66514 , n593835 , n66513 );
xnor ( n66515 , n66514 , n591902 );
and ( n66516 , n593834 , n66515 );
xor ( n66517 , n593514 , n66195 );
xor ( n66518 , n66517 , n66198 );
and ( n593842 , n66515 , n66518 );
and ( n593843 , n593834 , n66518 );
or ( n66521 , n66516 , n593842 , n593843 );
not ( n593845 , n66187 );
and ( n593846 , n66507 , n64456 );
and ( n593847 , n593520 , n64454 );
nor ( n66525 , n593846 , n593847 );
xnor ( n593849 , n66525 , n591786 );
or ( n593850 , n593845 , n593849 );
and ( n66528 , n65640 , n64650 );
and ( n66529 , n592806 , n64648 );
nor ( n66530 , n66528 , n66529 );
xnor ( n66531 , n66530 , n591902 );
and ( n593855 , n593850 , n66531 );
and ( n593856 , n65844 , n64559 );
and ( n66534 , n65630 , n591880 );
nor ( n593858 , n593856 , n66534 );
xnor ( n66536 , n593858 , n64521 );
and ( n593860 , n66531 , n66536 );
and ( n593861 , n593850 , n66536 );
or ( n593862 , n593855 , n593860 , n593861 );
and ( n66540 , n65384 , n64744 );
and ( n593864 , n592645 , n64742 );
nor ( n593865 , n66540 , n593864 );
xnor ( n66543 , n593865 , n64623 );
and ( n593867 , n593862 , n66543 );
xor ( n593868 , n66353 , n593680 );
xor ( n66546 , n593868 , n593685 );
and ( n593870 , n66543 , n66546 );
and ( n593871 , n593862 , n66546 );
or ( n593872 , n593867 , n593870 , n593871 );
and ( n66550 , n66521 , n593872 );
xor ( n593874 , n66365 , n593692 );
xor ( n66552 , n593874 , n593697 );
and ( n593876 , n593872 , n66552 );
and ( n66554 , n66521 , n66552 );
or ( n593878 , n66550 , n593876 , n66554 );
and ( n593879 , n64533 , n593256 );
and ( n593880 , n591851 , n593254 );
nor ( n66558 , n593879 , n593880 );
xnor ( n593882 , n66558 , n65490 );
and ( n66560 , n593878 , n593882 );
and ( n593884 , n64683 , n592683 );
and ( n593885 , n64630 , n592681 );
nor ( n66563 , n593884 , n593885 );
xnor ( n593887 , n66563 , n592475 );
and ( n66565 , n593882 , n593887 );
and ( n593889 , n593878 , n593887 );
or ( n66567 , n66560 , n66565 , n593889 );
xor ( n66568 , n593615 , n593619 );
xor ( n66569 , n66568 , n593624 );
and ( n66570 , n66567 , n66569 );
xor ( n593894 , n66338 , n593665 );
xor ( n593895 , n593894 , n593668 );
and ( n66573 , n66569 , n593895 );
and ( n593897 , n66567 , n593895 );
or ( n66575 , n66570 , n66573 , n593897 );
xor ( n593899 , n593643 , n66322 );
xor ( n593900 , n593899 , n66325 );
and ( n593901 , n66575 , n593900 );
xor ( n66579 , n593671 , n593720 );
xor ( n593903 , n66579 , n593723 );
and ( n593904 , n593900 , n593903 );
and ( n593905 , n66575 , n593903 );
or ( n66583 , n593901 , n593904 , n593905 );
and ( n593907 , n593823 , n66583 );
xor ( n66585 , n593639 , n66328 );
xor ( n593909 , n66585 , n593654 );
and ( n593910 , n66583 , n593909 );
and ( n593911 , n593823 , n593909 );
or ( n593912 , n593907 , n593910 , n593911 );
xor ( n593913 , n66334 , n593734 );
xor ( n66591 , n593913 , n66414 );
and ( n593915 , n593912 , n66591 );
xor ( n593916 , n66262 , n66264 );
xor ( n66594 , n593916 , n593590 );
and ( n593918 , n66591 , n66594 );
and ( n593919 , n593912 , n66594 );
or ( n593920 , n593915 , n593918 , n593919 );
and ( n66598 , n66429 , n593920 );
xor ( n593922 , n66429 , n593920 );
xor ( n593923 , n593912 , n66591 );
xor ( n593924 , n593923 , n66594 );
and ( n593925 , n593520 , n64491 );
and ( n66603 , n66104 , n64489 );
nor ( n593927 , n593925 , n66603 );
xnor ( n593928 , n593927 , n64448 );
buf ( n66606 , n591699 );
and ( n66607 , n66606 , n64456 );
and ( n66608 , n66507 , n64454 );
nor ( n66609 , n66607 , n66608 );
xnor ( n593933 , n66609 , n591786 );
and ( n593934 , n593928 , n593933 );
and ( n593935 , n66104 , n64491 );
and ( n593936 , n593437 , n64489 );
nor ( n66614 , n593935 , n593936 );
xnor ( n66615 , n66614 , n64448 );
and ( n593939 , n593934 , n66615 );
and ( n593940 , n66606 , n64451 );
and ( n593941 , n66615 , n593940 );
and ( n66619 , n593934 , n593940 );
or ( n593943 , n593939 , n593941 , n66619 );
xnor ( n593944 , n593845 , n593849 );
and ( n593945 , n65630 , n64650 );
and ( n66623 , n65640 , n64648 );
nor ( n593947 , n593945 , n66623 );
xnor ( n593948 , n593947 , n591902 );
and ( n66626 , n593944 , n593948 );
and ( n593950 , n593298 , n64559 );
and ( n593951 , n65844 , n591880 );
nor ( n593952 , n593950 , n593951 );
xnor ( n66630 , n593952 , n64521 );
and ( n593954 , n593948 , n66630 );
and ( n593955 , n593944 , n66630 );
or ( n66633 , n66626 , n593954 , n593955 );
and ( n593957 , n593943 , n66633 );
xor ( n593958 , n593827 , n593828 );
xor ( n593959 , n593958 , n593831 );
and ( n66637 , n66633 , n593959 );
and ( n593961 , n593943 , n593959 );
or ( n593962 , n593957 , n66637 , n593961 );
and ( n66640 , n592468 , n64862 );
and ( n593964 , n592478 , n64860 );
nor ( n66642 , n66640 , n593964 );
xnor ( n66643 , n66642 , n64764 );
and ( n593967 , n593962 , n66643 );
xor ( n66645 , n593834 , n66515 );
xor ( n593969 , n66645 , n66518 );
and ( n593970 , n66643 , n593969 );
and ( n66648 , n593962 , n593969 );
or ( n593972 , n593967 , n593970 , n66648 );
and ( n66650 , n64854 , n592486 );
and ( n593974 , n64838 , n592484 );
nor ( n593975 , n66650 , n593974 );
xnor ( n66653 , n593975 , n64990 );
and ( n593977 , n593972 , n66653 );
xor ( n593978 , n66433 , n66437 );
xor ( n66656 , n593978 , n593763 );
and ( n66657 , n66653 , n66656 );
and ( n66658 , n593972 , n66656 );
or ( n66659 , n593977 , n66657 , n66658 );
and ( n66660 , n64450 , n66457 );
and ( n593984 , n64458 , n593778 );
nor ( n66662 , n66660 , n593984 );
xnor ( n593986 , n66662 , n593160 );
and ( n593987 , n66659 , n593986 );
xor ( n593988 , n593795 , n66476 );
xor ( n593989 , n593988 , n66481 );
and ( n66667 , n593986 , n593989 );
and ( n593991 , n66659 , n593989 );
or ( n66669 , n593987 , n66667 , n593991 );
and ( n66670 , n592094 , n592683 );
and ( n593994 , n64683 , n592681 );
nor ( n66672 , n66670 , n593994 );
xnor ( n593996 , n66672 , n592475 );
and ( n593997 , n64997 , n592340 );
and ( n66675 , n64973 , n65015 );
nor ( n593999 , n593997 , n66675 );
xnor ( n594000 , n593999 , n64847 );
and ( n594001 , n593996 , n594000 );
and ( n66679 , n592478 , n64862 );
and ( n594003 , n592404 , n64860 );
nor ( n594004 , n66679 , n594003 );
xnor ( n594005 , n594004 , n64764 );
and ( n66683 , n594000 , n594005 );
and ( n594007 , n593996 , n594005 );
or ( n594008 , n594001 , n66683 , n594007 );
and ( n594009 , n64501 , n66142 );
and ( n66687 , n64466 , n66140 );
nor ( n594011 , n594009 , n66687 );
xnor ( n594012 , n594011 , n592960 );
and ( n594013 , n594008 , n594012 );
xor ( n66691 , n66377 , n66381 );
xor ( n594015 , n66691 , n66384 );
and ( n66693 , n594012 , n594015 );
and ( n594017 , n594008 , n594015 );
or ( n594018 , n594013 , n66693 , n594017 );
and ( n66696 , n66669 , n594018 );
xor ( n594020 , n593776 , n593783 );
xor ( n66698 , n594020 , n66465 );
and ( n66699 , n594018 , n66698 );
and ( n594023 , n66669 , n66698 );
or ( n594024 , n66696 , n66699 , n594023 );
and ( n66702 , n64586 , n593256 );
and ( n594026 , n64533 , n593254 );
nor ( n594027 , n66702 , n594026 );
xnor ( n594028 , n594027 , n65490 );
and ( n66706 , n64630 , n65592 );
and ( n594030 , n64591 , n592913 );
nor ( n594031 , n66706 , n594030 );
xnor ( n594032 , n594031 , n592638 );
and ( n66710 , n594028 , n594032 );
xor ( n594034 , n66521 , n593872 );
xor ( n594035 , n594034 , n66552 );
and ( n594036 , n594032 , n594035 );
and ( n66714 , n594028 , n594035 );
or ( n594038 , n66710 , n594036 , n66714 );
xor ( n594039 , n593878 , n593882 );
xor ( n66717 , n594039 , n593887 );
and ( n66718 , n594038 , n66717 );
xor ( n594042 , n593766 , n593770 );
xor ( n66720 , n594042 , n593773 );
and ( n594044 , n66717 , n66720 );
and ( n594045 , n594038 , n66720 );
or ( n594046 , n66718 , n594044 , n594045 );
xor ( n66724 , n66567 , n66569 );
xor ( n594048 , n66724 , n593895 );
and ( n594049 , n594046 , n594048 );
xor ( n66727 , n593807 , n66488 );
xor ( n594051 , n66727 , n593814 );
and ( n594052 , n594048 , n594051 );
and ( n66730 , n594046 , n594051 );
or ( n66731 , n594049 , n594052 , n66730 );
and ( n594055 , n594024 , n66731 );
xor ( n66733 , n66468 , n593817 );
xor ( n66734 , n66733 , n593820 );
and ( n66735 , n66731 , n66734 );
and ( n66736 , n594024 , n66734 );
or ( n66737 , n594055 , n66735 , n66736 );
xor ( n66738 , n593823 , n66583 );
xor ( n66739 , n66738 , n593909 );
and ( n66740 , n66737 , n66739 );
xor ( n66741 , n593726 , n66405 );
xor ( n66742 , n66741 , n66408 );
and ( n66743 , n66739 , n66742 );
and ( n594067 , n66737 , n66742 );
or ( n66745 , n66740 , n66743 , n594067 );
and ( n66746 , n593924 , n66745 );
xor ( n66747 , n593924 , n66745 );
xor ( n66748 , n66737 , n66739 );
xor ( n66749 , n66748 , n66742 );
and ( n66750 , n592094 , n65592 );
and ( n66751 , n64683 , n592913 );
nor ( n66752 , n66750 , n66751 );
xnor ( n66753 , n66752 , n592638 );
and ( n66754 , n64997 , n592486 );
and ( n66755 , n64973 , n592484 );
nor ( n66756 , n66754 , n66755 );
xnor ( n66757 , n66756 , n64990 );
and ( n66758 , n66753 , n66757 );
and ( n66759 , n592478 , n592340 );
and ( n66760 , n592404 , n65015 );
nor ( n66761 , n66759 , n66760 );
xnor ( n66762 , n66761 , n64847 );
and ( n66763 , n66757 , n66762 );
and ( n66764 , n66753 , n66762 );
or ( n66765 , n66758 , n66763 , n66764 );
xor ( n66766 , n593928 , n593933 );
and ( n66767 , n65640 , n64744 );
and ( n66768 , n592806 , n64742 );
nor ( n66769 , n66767 , n66768 );
xnor ( n66770 , n66769 , n64623 );
and ( n66771 , n66766 , n66770 );
and ( n66772 , n65844 , n64650 );
and ( n66773 , n65630 , n64648 );
nor ( n66774 , n66772 , n66773 );
xnor ( n66775 , n66774 , n591902 );
and ( n66776 , n66770 , n66775 );
and ( n594100 , n66766 , n66775 );
or ( n66778 , n66771 , n66776 , n594100 );
and ( n594102 , n65384 , n64862 );
and ( n594103 , n592645 , n64860 );
nor ( n66781 , n594102 , n594103 );
xnor ( n594105 , n66781 , n64764 );
and ( n594106 , n66778 , n594105 );
xor ( n66784 , n593944 , n593948 );
xor ( n66785 , n66784 , n66630 );
and ( n66786 , n594105 , n66785 );
and ( n66787 , n66778 , n66785 );
or ( n594111 , n594106 , n66786 , n66787 );
and ( n66789 , n66104 , n64559 );
and ( n594113 , n593437 , n591880 );
nor ( n594114 , n66789 , n594113 );
xnor ( n594115 , n594114 , n64521 );
buf ( n66793 , n591701 );
and ( n594117 , n66793 , n64451 );
and ( n594118 , n594115 , n594117 );
and ( n66796 , n593437 , n64559 );
and ( n594120 , n593298 , n591880 );
nor ( n594121 , n66796 , n594120 );
xnor ( n66799 , n594121 , n64521 );
and ( n594123 , n594118 , n66799 );
buf ( n594124 , n591700 );
and ( n66802 , n594124 , n64451 );
and ( n66803 , n66799 , n66802 );
and ( n594127 , n594118 , n66802 );
or ( n594128 , n594123 , n66803 , n594127 );
and ( n66806 , n592806 , n64744 );
and ( n594130 , n65493 , n64742 );
nor ( n66808 , n66806 , n594130 );
xnor ( n66809 , n66808 , n64623 );
and ( n594133 , n594128 , n66809 );
xor ( n594134 , n593934 , n66615 );
xor ( n66812 , n594134 , n593940 );
and ( n594136 , n66809 , n66812 );
and ( n66814 , n594128 , n66812 );
or ( n594138 , n594133 , n594136 , n66814 );
and ( n66816 , n594111 , n594138 );
xor ( n66817 , n593943 , n66633 );
xor ( n594141 , n66817 , n593959 );
and ( n594142 , n594138 , n594141 );
and ( n66820 , n594111 , n594141 );
or ( n594144 , n66816 , n594142 , n66820 );
and ( n594145 , n66765 , n594144 );
and ( n66823 , n64501 , n66457 );
and ( n594147 , n64466 , n593778 );
nor ( n594148 , n66823 , n594147 );
xnor ( n594149 , n594148 , n593160 );
and ( n66827 , n594144 , n594149 );
and ( n594151 , n66765 , n594149 );
or ( n594152 , n594145 , n66827 , n594151 );
and ( n66830 , n64533 , n66142 );
and ( n594154 , n591851 , n66140 );
nor ( n594155 , n66830 , n594154 );
xnor ( n66833 , n594155 , n592960 );
and ( n594157 , n64683 , n65592 );
and ( n594158 , n64630 , n592913 );
nor ( n66836 , n594157 , n594158 );
xnor ( n594160 , n66836 , n592638 );
and ( n66838 , n66833 , n594160 );
xor ( n594162 , n593962 , n66643 );
xor ( n594163 , n594162 , n593969 );
and ( n66841 , n594160 , n594163 );
and ( n594165 , n66833 , n594163 );
or ( n66843 , n66838 , n66841 , n594165 );
and ( n66844 , n594152 , n66843 );
xor ( n66845 , n593996 , n594000 );
xor ( n66846 , n66845 , n594005 );
and ( n66847 , n66843 , n66846 );
and ( n66848 , n594152 , n66846 );
or ( n66849 , n66844 , n66847 , n66848 );
xor ( n594173 , n66659 , n593986 );
xor ( n66851 , n594173 , n593989 );
and ( n594175 , n66849 , n66851 );
xor ( n66853 , n594038 , n66717 );
xor ( n594177 , n66853 , n66720 );
and ( n594178 , n66851 , n594177 );
and ( n594179 , n66849 , n594177 );
or ( n66857 , n594175 , n594178 , n594179 );
and ( n594181 , n592645 , n64862 );
and ( n594182 , n592468 , n64860 );
nor ( n66860 , n594181 , n594182 );
xnor ( n66861 , n66860 , n64764 );
and ( n594185 , n65493 , n64744 );
and ( n66863 , n65384 , n64742 );
nor ( n594187 , n594185 , n66863 );
xnor ( n66865 , n594187 , n64623 );
and ( n66866 , n66861 , n66865 );
xor ( n594190 , n593850 , n66531 );
xor ( n66868 , n594190 , n66536 );
and ( n66869 , n66865 , n66868 );
and ( n66870 , n66861 , n66868 );
or ( n66871 , n66866 , n66869 , n66870 );
and ( n594195 , n64973 , n592486 );
and ( n594196 , n64854 , n592484 );
nor ( n594197 , n594195 , n594196 );
xnor ( n66875 , n594197 , n64990 );
and ( n66876 , n66871 , n66875 );
and ( n66877 , n592404 , n592340 );
and ( n594201 , n64997 , n65015 );
nor ( n594202 , n66877 , n594201 );
xnor ( n66880 , n594202 , n64847 );
and ( n594204 , n66875 , n66880 );
and ( n594205 , n66871 , n66880 );
or ( n66883 , n66876 , n594204 , n594205 );
xor ( n66884 , n65834 , n66107 );
xor ( n66885 , n66107 , n593431 );
not ( n66886 , n66885 );
and ( n594210 , n66884 , n66886 );
and ( n594211 , n64458 , n594210 );
not ( n66889 , n594211 );
xnor ( n594213 , n66889 , n593434 );
and ( n594214 , n66883 , n594213 );
and ( n66892 , n591851 , n66142 );
and ( n594216 , n64501 , n66140 );
nor ( n594217 , n66892 , n594216 );
xnor ( n66895 , n594217 , n592960 );
and ( n594219 , n594213 , n66895 );
and ( n594220 , n66883 , n66895 );
or ( n66898 , n594214 , n594219 , n594220 );
and ( n594222 , n64591 , n593256 );
and ( n594223 , n64586 , n593254 );
nor ( n594224 , n594222 , n594223 );
xnor ( n66902 , n594224 , n65490 );
and ( n594226 , n64838 , n592683 );
and ( n66904 , n592094 , n592681 );
nor ( n66905 , n594226 , n66904 );
xnor ( n66906 , n66905 , n592475 );
and ( n66907 , n66902 , n66906 );
xor ( n66908 , n593862 , n66543 );
xor ( n66909 , n66908 , n66546 );
and ( n594233 , n66906 , n66909 );
and ( n66911 , n66902 , n66909 );
or ( n594235 , n66907 , n594233 , n66911 );
and ( n66913 , n64466 , n66457 );
and ( n66914 , n64450 , n593778 );
nor ( n594238 , n66913 , n66914 );
xnor ( n594239 , n594238 , n593160 );
and ( n66917 , n594235 , n594239 );
xor ( n594241 , n593972 , n66653 );
xor ( n594242 , n594241 , n66656 );
and ( n66920 , n594239 , n594242 );
and ( n594244 , n594235 , n594242 );
or ( n594245 , n66917 , n66920 , n594244 );
and ( n66923 , n66898 , n594245 );
xor ( n594247 , n594008 , n594012 );
xor ( n594248 , n594247 , n594015 );
and ( n66926 , n594245 , n594248 );
and ( n594250 , n66898 , n594248 );
or ( n594251 , n66923 , n66926 , n594250 );
and ( n66929 , n66857 , n594251 );
xor ( n66930 , n66669 , n594018 );
xor ( n594254 , n66930 , n66698 );
and ( n594255 , n594251 , n594254 );
and ( n66933 , n66857 , n594254 );
or ( n594257 , n66929 , n594255 , n66933 );
xor ( n594258 , n594024 , n66731 );
xor ( n594259 , n594258 , n66734 );
and ( n594260 , n594257 , n594259 );
xor ( n66938 , n66575 , n593900 );
xor ( n594262 , n66938 , n593903 );
and ( n66940 , n594259 , n594262 );
and ( n66941 , n594257 , n594262 );
or ( n594265 , n594260 , n66940 , n66941 );
and ( n66943 , n66749 , n594265 );
xor ( n594267 , n66749 , n594265 );
xor ( n594268 , n594257 , n594259 );
xor ( n66946 , n594268 , n594262 );
and ( n66947 , n593520 , n64559 );
and ( n594271 , n66104 , n591880 );
nor ( n594272 , n66947 , n594271 );
xnor ( n594273 , n594272 , n64521 );
buf ( n66951 , n591702 );
and ( n594275 , n66951 , n64451 );
and ( n594276 , n594273 , n594275 );
and ( n66954 , n66507 , n64491 );
and ( n594278 , n593520 , n64489 );
nor ( n594279 , n66954 , n594278 );
xnor ( n594280 , n594279 , n64448 );
and ( n66958 , n594276 , n594280 );
and ( n594282 , n594124 , n64456 );
and ( n594283 , n66606 , n64454 );
nor ( n594284 , n594282 , n594283 );
xnor ( n66962 , n594284 , n591786 );
and ( n594286 , n594280 , n66962 );
and ( n66964 , n594276 , n66962 );
or ( n594288 , n66958 , n594286 , n66964 );
xor ( n594289 , n594115 , n594117 );
buf ( n66967 , n591703 );
and ( n594291 , n66967 , n64456 );
and ( n594292 , n66951 , n64454 );
nor ( n66970 , n594291 , n594292 );
xnor ( n594294 , n66970 , n591786 );
buf ( n594295 , n591704 );
and ( n66973 , n594295 , n64451 );
and ( n594297 , n594294 , n66973 );
and ( n594298 , n66967 , n64451 );
and ( n66976 , n594297 , n594298 );
and ( n594300 , n66606 , n64491 );
and ( n594301 , n66507 , n64489 );
nor ( n594302 , n594300 , n594301 );
xnor ( n66980 , n594302 , n64448 );
and ( n594304 , n66976 , n66980 );
and ( n594305 , n66793 , n64456 );
and ( n594306 , n594124 , n64454 );
nor ( n66984 , n594305 , n594306 );
xnor ( n594308 , n66984 , n591786 );
and ( n594309 , n66980 , n594308 );
and ( n66987 , n66976 , n594308 );
or ( n66988 , n594304 , n594309 , n66987 );
and ( n594312 , n594289 , n66988 );
and ( n594313 , n65630 , n64744 );
and ( n66991 , n65640 , n64742 );
nor ( n594315 , n594313 , n66991 );
xnor ( n594316 , n594315 , n64623 );
and ( n594317 , n66988 , n594316 );
and ( n594318 , n594289 , n594316 );
or ( n66996 , n594312 , n594317 , n594318 );
and ( n66997 , n594288 , n66996 );
xor ( n594321 , n594118 , n66799 );
xor ( n594322 , n594321 , n66802 );
and ( n594323 , n66996 , n594322 );
and ( n594324 , n594288 , n594322 );
or ( n67002 , n66997 , n594323 , n594324 );
and ( n594326 , n592468 , n592340 );
and ( n594327 , n592478 , n65015 );
nor ( n67005 , n594326 , n594327 );
xnor ( n67006 , n67005 , n64847 );
and ( n594330 , n67002 , n67006 );
xor ( n67008 , n594128 , n66809 );
xor ( n67009 , n67008 , n66812 );
and ( n594333 , n67006 , n67009 );
and ( n67011 , n67002 , n67009 );
or ( n594335 , n594330 , n594333 , n67011 );
and ( n594336 , n64854 , n592683 );
and ( n594337 , n64838 , n592681 );
nor ( n67015 , n594336 , n594337 );
xnor ( n594339 , n67015 , n592475 );
and ( n594340 , n594335 , n594339 );
xor ( n67018 , n66861 , n66865 );
xor ( n67019 , n67018 , n66868 );
and ( n67020 , n594339 , n67019 );
and ( n67021 , n594335 , n67019 );
or ( n67022 , n594340 , n67020 , n67021 );
and ( n594346 , n64450 , n594210 );
and ( n67024 , n64458 , n66885 );
nor ( n594348 , n594346 , n67024 );
xnor ( n594349 , n594348 , n593434 );
and ( n67027 , n67022 , n594349 );
xor ( n594351 , n66902 , n66906 );
xor ( n594352 , n594351 , n66909 );
and ( n594353 , n594349 , n594352 );
and ( n67031 , n67022 , n594352 );
or ( n594355 , n67027 , n594353 , n67031 );
xor ( n594356 , n66883 , n594213 );
xor ( n594357 , n594356 , n66895 );
and ( n67035 , n594355 , n594357 );
xor ( n594359 , n594028 , n594032 );
xor ( n594360 , n594359 , n594035 );
and ( n67038 , n594357 , n594360 );
and ( n594362 , n594355 , n594360 );
or ( n67040 , n67035 , n67038 , n594362 );
and ( n67041 , n64586 , n66142 );
and ( n67042 , n64533 , n66140 );
nor ( n594366 , n67041 , n67042 );
xnor ( n67044 , n594366 , n592960 );
and ( n594368 , n64630 , n593256 );
and ( n594369 , n64591 , n593254 );
nor ( n67047 , n594368 , n594369 );
xnor ( n594371 , n67047 , n65490 );
and ( n594372 , n67044 , n594371 );
xor ( n67050 , n594111 , n594138 );
xor ( n594374 , n67050 , n594141 );
and ( n594375 , n594371 , n594374 );
and ( n67053 , n67044 , n594374 );
or ( n594377 , n594372 , n594375 , n67053 );
xor ( n67055 , n66871 , n66875 );
xor ( n594379 , n67055 , n66880 );
and ( n594380 , n594377 , n594379 );
xor ( n67058 , n66833 , n594160 );
xor ( n594382 , n67058 , n594163 );
and ( n594383 , n594379 , n594382 );
and ( n67061 , n594377 , n594382 );
or ( n594385 , n594380 , n594383 , n67061 );
xor ( n594386 , n594152 , n66843 );
xor ( n594387 , n594386 , n66846 );
and ( n67065 , n594385 , n594387 );
xor ( n594389 , n594235 , n594239 );
xor ( n594390 , n594389 , n594242 );
and ( n594391 , n594387 , n594390 );
and ( n67069 , n594385 , n594390 );
or ( n594393 , n67065 , n594391 , n67069 );
and ( n594394 , n67040 , n594393 );
xor ( n594395 , n66898 , n594245 );
xor ( n67073 , n594395 , n594248 );
and ( n594397 , n594393 , n67073 );
and ( n594398 , n67040 , n67073 );
or ( n67076 , n594394 , n594397 , n594398 );
xor ( n594400 , n66857 , n594251 );
xor ( n594401 , n594400 , n594254 );
and ( n594402 , n67076 , n594401 );
xor ( n67080 , n594046 , n594048 );
xor ( n594404 , n67080 , n594051 );
and ( n594405 , n594401 , n594404 );
and ( n67083 , n67076 , n594404 );
or ( n594407 , n594402 , n594405 , n67083 );
and ( n594408 , n66946 , n594407 );
xor ( n594409 , n66946 , n594407 );
xor ( n67087 , n67076 , n594401 );
xor ( n594411 , n67087 , n594404 );
and ( n594412 , n592645 , n592340 );
and ( n594413 , n592468 , n65015 );
nor ( n67091 , n594412 , n594413 );
xnor ( n594415 , n67091 , n64847 );
and ( n594416 , n65493 , n64862 );
and ( n594417 , n65384 , n64860 );
nor ( n67095 , n594416 , n594417 );
xnor ( n594419 , n67095 , n64764 );
and ( n594420 , n594415 , n594419 );
xor ( n67098 , n66766 , n66770 );
xor ( n594422 , n67098 , n66775 );
and ( n594423 , n594419 , n594422 );
and ( n67101 , n594415 , n594422 );
or ( n594425 , n594420 , n594423 , n67101 );
and ( n594426 , n64973 , n592683 );
and ( n67104 , n64854 , n592681 );
nor ( n594428 , n594426 , n67104 );
xnor ( n594429 , n594428 , n592475 );
and ( n67107 , n594425 , n594429 );
and ( n594431 , n592404 , n592486 );
and ( n594432 , n64997 , n592484 );
nor ( n67110 , n594431 , n594432 );
xnor ( n594434 , n67110 , n64990 );
and ( n594435 , n594429 , n594434 );
and ( n67113 , n594425 , n594434 );
or ( n594437 , n67107 , n594435 , n67113 );
xor ( n594438 , n593431 , n66186 );
xor ( n67116 , n66186 , n66187 );
not ( n594440 , n67116 );
and ( n594441 , n594438 , n594440 );
and ( n67119 , n64458 , n594441 );
not ( n594443 , n67119 );
xnor ( n594444 , n594443 , n66190 );
and ( n67122 , n594437 , n594444 );
and ( n594446 , n591851 , n66457 );
and ( n594447 , n64501 , n593778 );
nor ( n67125 , n594446 , n594447 );
xnor ( n67126 , n67125 , n593160 );
and ( n67127 , n594444 , n67126 );
and ( n67128 , n594437 , n67126 );
or ( n594452 , n67122 , n67127 , n67128 );
and ( n594453 , n64591 , n66142 );
and ( n594454 , n64586 , n66140 );
nor ( n594455 , n594453 , n594454 );
xnor ( n67133 , n594455 , n592960 );
and ( n67134 , n64838 , n65592 );
and ( n594458 , n592094 , n592913 );
nor ( n594459 , n67134 , n594458 );
xnor ( n594460 , n594459 , n592638 );
and ( n67138 , n67133 , n594460 );
xor ( n67139 , n66778 , n594105 );
xor ( n594463 , n67139 , n66785 );
and ( n594464 , n594460 , n594463 );
and ( n594465 , n67133 , n594463 );
or ( n67143 , n67138 , n594464 , n594465 );
and ( n67144 , n64466 , n594210 );
and ( n594468 , n64450 , n66885 );
nor ( n594469 , n67144 , n594468 );
xnor ( n594470 , n594469 , n593434 );
and ( n67148 , n67143 , n594470 );
xor ( n67149 , n594335 , n594339 );
xor ( n594473 , n67149 , n67019 );
and ( n594474 , n594470 , n594473 );
and ( n594475 , n67143 , n594473 );
or ( n67153 , n67148 , n594474 , n594475 );
and ( n67154 , n594452 , n67153 );
xor ( n594478 , n66765 , n594144 );
xor ( n594479 , n594478 , n594149 );
and ( n594480 , n67153 , n594479 );
and ( n67158 , n594452 , n594479 );
or ( n67159 , n67154 , n594480 , n67158 );
and ( n594483 , n65640 , n64862 );
and ( n594484 , n592806 , n64860 );
nor ( n594485 , n594483 , n594484 );
xnor ( n67163 , n594485 , n64764 );
and ( n67164 , n65844 , n64744 );
and ( n594488 , n65630 , n64742 );
nor ( n594489 , n67164 , n594488 );
xnor ( n594490 , n594489 , n64623 );
and ( n67168 , n67163 , n594490 );
xor ( n67169 , n66976 , n66980 );
xor ( n594493 , n67169 , n594308 );
and ( n594494 , n594490 , n594493 );
and ( n594495 , n67163 , n594493 );
or ( n67173 , n67168 , n594494 , n594495 );
and ( n67174 , n65384 , n592340 );
and ( n594498 , n592645 , n65015 );
nor ( n594499 , n67174 , n594498 );
xnor ( n594500 , n594499 , n64847 );
and ( n67178 , n67173 , n594500 );
and ( n67179 , n592806 , n64862 );
and ( n594503 , n65493 , n64860 );
nor ( n67181 , n67179 , n594503 );
xnor ( n67182 , n67181 , n64764 );
and ( n67183 , n594500 , n67182 );
and ( n67184 , n67173 , n67182 );
or ( n594508 , n67178 , n67183 , n67184 );
xor ( n67186 , n594273 , n594275 );
xor ( n594510 , n594297 , n594298 );
and ( n594511 , n66104 , n64650 );
and ( n67189 , n593437 , n64648 );
nor ( n594513 , n594511 , n67189 );
xnor ( n594514 , n594513 , n591902 );
and ( n67192 , n594510 , n594514 );
and ( n594516 , n66951 , n64456 );
and ( n67194 , n66793 , n64454 );
nor ( n67195 , n594516 , n67194 );
xnor ( n67196 , n67195 , n591786 );
and ( n67197 , n594514 , n67196 );
and ( n67198 , n594510 , n67196 );
or ( n67199 , n67192 , n67197 , n67198 );
and ( n67200 , n67186 , n67199 );
and ( n67201 , n593437 , n64650 );
and ( n67202 , n593298 , n64648 );
nor ( n594526 , n67201 , n67202 );
xnor ( n67204 , n594526 , n591902 );
and ( n594528 , n67199 , n67204 );
and ( n594529 , n67186 , n67204 );
or ( n67207 , n67200 , n594528 , n594529 );
and ( n67208 , n593298 , n64650 );
and ( n594532 , n65844 , n64648 );
nor ( n67210 , n67208 , n594532 );
xnor ( n594534 , n67210 , n591902 );
and ( n594535 , n67207 , n594534 );
xor ( n67213 , n594276 , n594280 );
xor ( n594537 , n67213 , n66962 );
and ( n67215 , n594534 , n594537 );
and ( n594539 , n67207 , n594537 );
or ( n594540 , n594535 , n67215 , n594539 );
and ( n67218 , n594508 , n594540 );
xor ( n594542 , n594288 , n66996 );
xor ( n594543 , n594542 , n594322 );
and ( n67221 , n594540 , n594543 );
and ( n67222 , n594508 , n594543 );
or ( n594546 , n67218 , n67221 , n67222 );
and ( n67224 , n64533 , n66457 );
and ( n67225 , n591851 , n593778 );
nor ( n67226 , n67224 , n67225 );
xnor ( n67227 , n67226 , n593160 );
and ( n67228 , n594546 , n67227 );
and ( n67229 , n64683 , n593256 );
and ( n67230 , n64630 , n593254 );
nor ( n67231 , n67229 , n67230 );
xnor ( n67232 , n67231 , n65490 );
and ( n67233 , n67227 , n67232 );
and ( n67234 , n594546 , n67232 );
or ( n594558 , n67228 , n67233 , n67234 );
and ( n67236 , n592094 , n593256 );
and ( n594560 , n64683 , n593254 );
nor ( n594561 , n67236 , n594560 );
xnor ( n67239 , n594561 , n65490 );
and ( n67240 , n64997 , n592683 );
and ( n67241 , n64973 , n592681 );
nor ( n67242 , n67240 , n67241 );
xnor ( n67243 , n67242 , n592475 );
and ( n67244 , n67239 , n67243 );
and ( n67245 , n592478 , n592486 );
and ( n594569 , n592404 , n592484 );
nor ( n67247 , n67245 , n594569 );
xnor ( n594571 , n67247 , n64990 );
and ( n594572 , n67243 , n594571 );
and ( n67250 , n67239 , n594571 );
or ( n594574 , n67244 , n594572 , n67250 );
and ( n594575 , n64501 , n594210 );
and ( n67253 , n64466 , n66885 );
nor ( n594577 , n594575 , n67253 );
xnor ( n594578 , n594577 , n593434 );
and ( n67256 , n594574 , n594578 );
xor ( n67257 , n67002 , n67006 );
xor ( n67258 , n67257 , n67009 );
and ( n594582 , n594578 , n67258 );
and ( n67260 , n594574 , n67258 );
or ( n594584 , n67256 , n594582 , n67260 );
and ( n594585 , n594558 , n594584 );
xor ( n67263 , n66753 , n66757 );
xor ( n594587 , n67263 , n66762 );
and ( n67265 , n594584 , n594587 );
and ( n67266 , n594558 , n594587 );
or ( n67267 , n594585 , n67265 , n67266 );
xor ( n67268 , n67022 , n594349 );
xor ( n67269 , n67268 , n594352 );
and ( n67270 , n67267 , n67269 );
xor ( n67271 , n594377 , n594379 );
xor ( n67272 , n67271 , n594382 );
and ( n67273 , n67269 , n67272 );
and ( n67274 , n67267 , n67272 );
or ( n67275 , n67270 , n67273 , n67274 );
and ( n67276 , n67159 , n67275 );
xor ( n67277 , n594355 , n594357 );
xor ( n594601 , n67277 , n594360 );
and ( n67279 , n67275 , n594601 );
and ( n594603 , n67159 , n594601 );
or ( n594604 , n67276 , n67279 , n594603 );
xor ( n67282 , n66849 , n66851 );
xor ( n594606 , n67282 , n594177 );
and ( n594607 , n594604 , n594606 );
xor ( n67285 , n67040 , n594393 );
xor ( n594609 , n67285 , n67073 );
and ( n594610 , n594606 , n594609 );
and ( n67288 , n594604 , n594609 );
or ( n594612 , n594607 , n594610 , n67288 );
and ( n594613 , n594411 , n594612 );
xor ( n67291 , n594411 , n594612 );
xor ( n67292 , n594604 , n594606 );
xor ( n594616 , n67292 , n594609 );
and ( n67294 , n592468 , n592486 );
and ( n594618 , n592478 , n592484 );
nor ( n594619 , n67294 , n594618 );
xnor ( n67297 , n594619 , n64990 );
xor ( n594621 , n594289 , n66988 );
xor ( n594622 , n594621 , n594316 );
and ( n594623 , n67297 , n594622 );
xor ( n67301 , n67207 , n594534 );
xor ( n594625 , n67301 , n594537 );
and ( n594626 , n594622 , n594625 );
and ( n67304 , n67297 , n594625 );
or ( n594628 , n594623 , n594626 , n67304 );
and ( n594629 , n64854 , n65592 );
and ( n67307 , n64838 , n592913 );
nor ( n67308 , n594629 , n67307 );
xnor ( n594632 , n67308 , n592638 );
and ( n67310 , n594628 , n594632 );
xor ( n67311 , n594415 , n594419 );
xor ( n67312 , n67311 , n594422 );
and ( n67313 , n594632 , n67312 );
and ( n67314 , n594628 , n67312 );
or ( n67315 , n67310 , n67313 , n67314 );
and ( n67316 , n64450 , n594441 );
and ( n67317 , n64458 , n67116 );
nor ( n67318 , n67316 , n67317 );
xnor ( n67319 , n67318 , n66190 );
and ( n67320 , n67315 , n67319 );
xor ( n67321 , n67133 , n594460 );
xor ( n594645 , n67321 , n594463 );
and ( n67323 , n67319 , n594645 );
and ( n594647 , n67315 , n594645 );
or ( n594648 , n67320 , n67323 , n594647 );
xor ( n67326 , n594437 , n594444 );
xor ( n67327 , n67326 , n67126 );
and ( n594651 , n594648 , n67327 );
xor ( n594652 , n67044 , n594371 );
xor ( n67330 , n594652 , n594374 );
and ( n594654 , n67327 , n67330 );
and ( n594655 , n594648 , n67330 );
or ( n67333 , n594651 , n594654 , n594655 );
and ( n594657 , n64586 , n66457 );
and ( n594658 , n64533 , n593778 );
nor ( n594659 , n594657 , n594658 );
xnor ( n594660 , n594659 , n593160 );
and ( n67338 , n64630 , n66142 );
and ( n594662 , n64591 , n66140 );
nor ( n594663 , n67338 , n594662 );
xnor ( n594664 , n594663 , n592960 );
and ( n67342 , n594660 , n594664 );
xor ( n594666 , n594508 , n594540 );
xor ( n594667 , n594666 , n594543 );
and ( n67345 , n594664 , n594667 );
and ( n594669 , n594660 , n594667 );
or ( n594670 , n67342 , n67345 , n594669 );
xor ( n67348 , n594425 , n594429 );
xor ( n594672 , n67348 , n594434 );
and ( n594673 , n594670 , n594672 );
xor ( n67351 , n594546 , n67227 );
xor ( n594675 , n67351 , n67232 );
and ( n594676 , n594672 , n594675 );
and ( n67354 , n594670 , n594675 );
or ( n594678 , n594673 , n594676 , n67354 );
xor ( n594679 , n594558 , n594584 );
xor ( n67357 , n594679 , n594587 );
and ( n67358 , n594678 , n67357 );
xor ( n67359 , n67143 , n594470 );
xor ( n67360 , n67359 , n594473 );
and ( n67361 , n67357 , n67360 );
and ( n67362 , n594678 , n67360 );
or ( n67363 , n67358 , n67361 , n67362 );
and ( n67364 , n67333 , n67363 );
xor ( n67365 , n594452 , n67153 );
xor ( n67366 , n67365 , n594479 );
and ( n594690 , n67363 , n67366 );
and ( n67368 , n67333 , n67366 );
or ( n594692 , n67364 , n594690 , n67368 );
xor ( n67370 , n594385 , n594387 );
xor ( n594694 , n67370 , n594390 );
and ( n67372 , n594692 , n594694 );
xor ( n67373 , n67159 , n67275 );
xor ( n67374 , n67373 , n594601 );
and ( n67375 , n594694 , n67374 );
and ( n67376 , n594692 , n67374 );
or ( n67377 , n67372 , n67375 , n67376 );
and ( n67378 , n594616 , n67377 );
xor ( n67379 , n594616 , n67377 );
xor ( n67380 , n594692 , n594694 );
xor ( n67381 , n67380 , n67374 );
xor ( n67382 , n594294 , n66973 );
and ( n67383 , n594295 , n64456 );
and ( n67384 , n66967 , n64454 );
nor ( n67385 , n67383 , n67384 );
xnor ( n67386 , n67385 , n591786 );
buf ( n594710 , n591705 );
and ( n67388 , n594710 , n64451 );
and ( n67389 , n67386 , n67388 );
and ( n67390 , n67382 , n67389 );
and ( n67391 , n593520 , n64650 );
and ( n594715 , n66104 , n64648 );
nor ( n67393 , n67391 , n594715 );
xnor ( n594717 , n67393 , n591902 );
and ( n67395 , n67389 , n594717 );
and ( n594719 , n67382 , n594717 );
or ( n594720 , n67390 , n67395 , n594719 );
and ( n67398 , n66507 , n64559 );
and ( n594722 , n593520 , n591880 );
nor ( n67400 , n67398 , n594722 );
xnor ( n67401 , n67400 , n64521 );
and ( n594725 , n594720 , n67401 );
and ( n67403 , n594124 , n64491 );
and ( n67404 , n66606 , n64489 );
nor ( n67405 , n67403 , n67404 );
xnor ( n67406 , n67405 , n64448 );
and ( n67407 , n67401 , n67406 );
and ( n67408 , n594720 , n67406 );
or ( n67409 , n594725 , n67407 , n67408 );
and ( n67410 , n65493 , n592340 );
and ( n67411 , n65384 , n65015 );
nor ( n67412 , n67410 , n67411 );
xnor ( n67413 , n67412 , n64847 );
and ( n594737 , n67409 , n67413 );
xor ( n67415 , n67186 , n67199 );
xor ( n594739 , n67415 , n67204 );
and ( n594740 , n67413 , n594739 );
and ( n67418 , n67409 , n594739 );
or ( n594742 , n594737 , n594740 , n67418 );
and ( n594743 , n64838 , n593256 );
and ( n67421 , n592094 , n593254 );
nor ( n67422 , n594743 , n67421 );
xnor ( n594746 , n67422 , n65490 );
and ( n67424 , n594742 , n594746 );
and ( n594748 , n592404 , n592683 );
and ( n594749 , n64997 , n592681 );
nor ( n594750 , n594748 , n594749 );
xnor ( n67428 , n594750 , n592475 );
and ( n594752 , n594746 , n67428 );
and ( n594753 , n594742 , n67428 );
or ( n67431 , n67424 , n594752 , n594753 );
and ( n594755 , n593437 , n64744 );
and ( n67433 , n593298 , n64742 );
nor ( n594757 , n594755 , n67433 );
xnor ( n67435 , n594757 , n64623 );
and ( n594759 , n66606 , n64559 );
and ( n67437 , n66507 , n591880 );
nor ( n67438 , n594759 , n67437 );
xnor ( n594762 , n67438 , n64521 );
and ( n67440 , n67435 , n594762 );
and ( n594764 , n66793 , n64491 );
and ( n594765 , n594124 , n64489 );
nor ( n67443 , n594764 , n594765 );
xnor ( n67444 , n67443 , n64448 );
and ( n67445 , n594762 , n67444 );
and ( n67446 , n67435 , n67444 );
or ( n67447 , n67440 , n67445 , n67446 );
and ( n67448 , n65630 , n64862 );
and ( n67449 , n65640 , n64860 );
nor ( n594773 , n67448 , n67449 );
xnor ( n67451 , n594773 , n64764 );
and ( n594775 , n67447 , n67451 );
and ( n594776 , n593298 , n64744 );
and ( n67454 , n65844 , n64742 );
nor ( n594778 , n594776 , n67454 );
xnor ( n67456 , n594778 , n64623 );
and ( n67457 , n67451 , n67456 );
and ( n67458 , n67447 , n67456 );
or ( n67459 , n594775 , n67457 , n67458 );
and ( n67460 , n592645 , n592486 );
and ( n67461 , n592468 , n592484 );
nor ( n67462 , n67460 , n67461 );
xnor ( n67463 , n67462 , n64990 );
and ( n67464 , n67459 , n67463 );
xor ( n67465 , n67163 , n594490 );
xor ( n67466 , n67465 , n594493 );
and ( n67467 , n67463 , n67466 );
and ( n67468 , n67459 , n67466 );
or ( n67469 , n67464 , n67467 , n67468 );
and ( n67470 , n64973 , n65592 );
and ( n594794 , n64854 , n592913 );
nor ( n67472 , n67470 , n594794 );
xnor ( n67473 , n67472 , n592638 );
and ( n67474 , n67469 , n67473 );
xor ( n594798 , n67173 , n594500 );
xor ( n594799 , n594798 , n67182 );
and ( n67477 , n67473 , n594799 );
and ( n594801 , n67469 , n594799 );
or ( n594802 , n67474 , n67477 , n594801 );
and ( n67480 , n67431 , n594802 );
buf ( n594804 , n591765 );
xor ( n594805 , n66187 , n594804 );
not ( n67483 , n594804 );
and ( n594807 , n594805 , n67483 );
and ( n594808 , n64458 , n594807 );
not ( n67486 , n594808 );
xnor ( n67487 , n67486 , n66187 );
and ( n67488 , n594802 , n67487 );
and ( n67489 , n67431 , n67487 );
or ( n594813 , n67480 , n67488 , n67489 );
and ( n67491 , n64466 , n594441 );
and ( n594815 , n64450 , n67116 );
nor ( n594816 , n67491 , n594815 );
xnor ( n67494 , n594816 , n66190 );
and ( n594818 , n591851 , n594210 );
and ( n594819 , n64501 , n66885 );
nor ( n67497 , n594818 , n594819 );
xnor ( n594821 , n67497 , n593434 );
and ( n594822 , n67494 , n594821 );
xor ( n67500 , n594628 , n594632 );
xor ( n594824 , n67500 , n67312 );
and ( n67502 , n594821 , n594824 );
and ( n67503 , n67494 , n594824 );
or ( n67504 , n594822 , n67502 , n67503 );
and ( n67505 , n594813 , n67504 );
xor ( n67506 , n594574 , n594578 );
xor ( n67507 , n67506 , n67258 );
and ( n67508 , n67504 , n67507 );
and ( n67509 , n594813 , n67507 );
or ( n67510 , n67505 , n67508 , n67509 );
and ( n67511 , n64533 , n594210 );
and ( n67512 , n591851 , n66885 );
nor ( n594836 , n67511 , n67512 );
xnor ( n67514 , n594836 , n593434 );
and ( n67515 , n64591 , n66457 );
and ( n67516 , n64586 , n593778 );
nor ( n594840 , n67515 , n67516 );
xnor ( n594841 , n594840 , n593160 );
and ( n67519 , n67514 , n594841 );
and ( n594843 , n64683 , n66142 );
and ( n594844 , n64630 , n66140 );
nor ( n67522 , n594843 , n594844 );
xnor ( n594846 , n67522 , n592960 );
and ( n594847 , n594841 , n594846 );
and ( n67525 , n67514 , n594846 );
or ( n594849 , n67519 , n594847 , n67525 );
xor ( n594850 , n67239 , n67243 );
xor ( n67528 , n594850 , n594571 );
and ( n594852 , n594849 , n67528 );
xor ( n594853 , n594660 , n594664 );
xor ( n67531 , n594853 , n594667 );
and ( n594855 , n67528 , n67531 );
and ( n594856 , n594849 , n67531 );
or ( n67534 , n594852 , n594855 , n594856 );
xor ( n594858 , n594670 , n594672 );
xor ( n594859 , n594858 , n594675 );
and ( n67537 , n67534 , n594859 );
xor ( n594861 , n67315 , n67319 );
xor ( n594862 , n594861 , n594645 );
and ( n67540 , n594859 , n594862 );
and ( n594864 , n67534 , n594862 );
or ( n594865 , n67537 , n67540 , n594864 );
and ( n67543 , n67510 , n594865 );
xor ( n594867 , n594648 , n67327 );
xor ( n594868 , n594867 , n67330 );
and ( n67546 , n594865 , n594868 );
and ( n67547 , n67510 , n594868 );
or ( n594871 , n67543 , n67546 , n67547 );
xor ( n594872 , n67333 , n67363 );
xor ( n67550 , n594872 , n67366 );
and ( n594874 , n594871 , n67550 );
xor ( n594875 , n67267 , n67269 );
xor ( n67553 , n594875 , n67272 );
and ( n594877 , n67550 , n67553 );
and ( n594878 , n594871 , n67553 );
or ( n67556 , n594874 , n594877 , n594878 );
and ( n67557 , n67381 , n67556 );
xor ( n67558 , n67381 , n67556 );
xor ( n594882 , n594871 , n67550 );
xor ( n67560 , n594882 , n67553 );
and ( n67561 , n64630 , n66457 );
and ( n67562 , n64591 , n593778 );
nor ( n67563 , n67561 , n67562 );
xnor ( n67564 , n67563 , n593160 );
and ( n67565 , n64997 , n65592 );
and ( n67566 , n64973 , n592913 );
nor ( n67567 , n67565 , n67566 );
xnor ( n67568 , n67567 , n592638 );
and ( n67569 , n67564 , n67568 );
xor ( n594893 , n67459 , n67463 );
xor ( n67571 , n594893 , n67466 );
and ( n67572 , n67568 , n67571 );
and ( n67573 , n67564 , n67571 );
or ( n594897 , n67569 , n67572 , n67573 );
and ( n67575 , n64450 , n594807 );
and ( n594899 , n64458 , n594804 );
nor ( n594900 , n67575 , n594899 );
xnor ( n67578 , n594900 , n66187 );
and ( n67579 , n594897 , n67578 );
and ( n594903 , n64501 , n594441 );
and ( n594904 , n64466 , n67116 );
nor ( n67582 , n594903 , n594904 );
xnor ( n67583 , n67582 , n66190 );
and ( n594907 , n67578 , n67583 );
and ( n67585 , n594897 , n67583 );
or ( n67586 , n67579 , n594907 , n67585 );
and ( n67587 , n592094 , n66142 );
and ( n67588 , n64683 , n66140 );
nor ( n67589 , n67587 , n67588 );
xnor ( n67590 , n67589 , n592960 );
and ( n594914 , n64854 , n593256 );
and ( n67592 , n64838 , n593254 );
nor ( n594916 , n594914 , n67592 );
xnor ( n67594 , n594916 , n65490 );
and ( n67595 , n67590 , n67594 );
and ( n594919 , n592478 , n592683 );
and ( n67597 , n592404 , n592681 );
nor ( n594921 , n594919 , n67597 );
xnor ( n67599 , n594921 , n592475 );
and ( n67600 , n67594 , n67599 );
and ( n67601 , n67590 , n67599 );
or ( n67602 , n67595 , n67600 , n67601 );
and ( n67603 , n65640 , n592340 );
and ( n67604 , n592806 , n65015 );
nor ( n67605 , n67603 , n67604 );
xnor ( n594929 , n67605 , n64847 );
xor ( n67607 , n67435 , n594762 );
xor ( n594931 , n67607 , n67444 );
and ( n594932 , n594929 , n594931 );
xor ( n67610 , n67382 , n67389 );
xor ( n594934 , n67610 , n594717 );
and ( n594935 , n594931 , n594934 );
and ( n67613 , n594929 , n594934 );
or ( n67614 , n594932 , n594935 , n67613 );
and ( n594938 , n65384 , n592486 );
and ( n67616 , n592645 , n592484 );
nor ( n594940 , n594938 , n67616 );
xnor ( n594941 , n594940 , n64990 );
and ( n594942 , n67614 , n594941 );
xor ( n67620 , n594720 , n67401 );
xor ( n594944 , n67620 , n67406 );
and ( n594945 , n594941 , n594944 );
and ( n67623 , n67614 , n594944 );
or ( n594947 , n594942 , n594945 , n67623 );
and ( n594948 , n594710 , n64456 );
and ( n594949 , n594295 , n64454 );
nor ( n67627 , n594948 , n594949 );
xnor ( n594951 , n67627 , n591786 );
buf ( n594952 , n591706 );
and ( n67630 , n594952 , n64451 );
xor ( n594954 , n594951 , n67630 );
and ( n594955 , n594952 , n64456 );
and ( n67633 , n594710 , n64454 );
nor ( n594957 , n594955 , n67633 );
xnor ( n594958 , n594957 , n591786 );
buf ( n67636 , n591707 );
and ( n594960 , n67636 , n64451 );
and ( n594961 , n594958 , n594960 );
and ( n67639 , n594954 , n594961 );
and ( n67640 , n66967 , n64491 );
and ( n594964 , n66951 , n64489 );
nor ( n594965 , n67640 , n594964 );
xnor ( n67643 , n594965 , n64448 );
and ( n67644 , n594961 , n67643 );
and ( n67645 , n594954 , n67643 );
or ( n594969 , n67639 , n67644 , n67645 );
and ( n594970 , n66104 , n64744 );
and ( n67648 , n593437 , n64742 );
nor ( n67649 , n594970 , n67648 );
xnor ( n594973 , n67649 , n64623 );
and ( n67651 , n594969 , n594973 );
and ( n67652 , n66507 , n64650 );
and ( n594976 , n593520 , n64648 );
nor ( n67654 , n67652 , n594976 );
xnor ( n67655 , n67654 , n591902 );
and ( n594979 , n594973 , n67655 );
and ( n67657 , n594969 , n67655 );
or ( n594981 , n67651 , n594979 , n67657 );
xor ( n594982 , n67386 , n67388 );
and ( n67660 , n594951 , n67630 );
and ( n594984 , n594982 , n67660 );
and ( n67662 , n66951 , n64491 );
and ( n594986 , n66793 , n64489 );
nor ( n67664 , n67662 , n594986 );
xnor ( n594988 , n67664 , n64448 );
and ( n67666 , n67660 , n594988 );
and ( n67667 , n594982 , n594988 );
or ( n594991 , n594984 , n67666 , n67667 );
and ( n67669 , n594981 , n594991 );
and ( n594993 , n65844 , n64862 );
and ( n594994 , n65630 , n64860 );
nor ( n67672 , n594993 , n594994 );
xnor ( n67673 , n67672 , n64764 );
and ( n67674 , n594991 , n67673 );
and ( n594998 , n594981 , n67673 );
or ( n67676 , n67669 , n67674 , n594998 );
and ( n67677 , n592806 , n592340 );
and ( n595001 , n65493 , n65015 );
nor ( n67679 , n67677 , n595001 );
xnor ( n595003 , n67679 , n64847 );
and ( n595004 , n67676 , n595003 );
xor ( n67682 , n594510 , n594514 );
xor ( n595006 , n67682 , n67196 );
and ( n595007 , n595003 , n595006 );
and ( n67685 , n67676 , n595006 );
or ( n595009 , n595004 , n595007 , n67685 );
and ( n595010 , n594947 , n595009 );
xor ( n67688 , n67409 , n67413 );
xor ( n67689 , n67688 , n594739 );
and ( n595013 , n595009 , n67689 );
and ( n67691 , n594947 , n67689 );
or ( n595015 , n595010 , n595013 , n67691 );
and ( n595016 , n67602 , n595015 );
xor ( n67694 , n67297 , n594622 );
xor ( n67695 , n67694 , n594625 );
and ( n595019 , n595015 , n67695 );
and ( n67697 , n67602 , n67695 );
or ( n595021 , n595016 , n595019 , n67697 );
and ( n595022 , n67586 , n595021 );
xor ( n67700 , n67431 , n594802 );
xor ( n595024 , n67700 , n67487 );
and ( n595025 , n595021 , n595024 );
and ( n67703 , n67586 , n595024 );
or ( n67704 , n595022 , n595025 , n67703 );
xor ( n67705 , n67514 , n594841 );
xor ( n595029 , n67705 , n594846 );
xor ( n67707 , n594742 , n594746 );
xor ( n595031 , n67707 , n67428 );
and ( n595032 , n595029 , n595031 );
xor ( n595033 , n67469 , n67473 );
xor ( n67711 , n595033 , n594799 );
and ( n595035 , n595031 , n67711 );
and ( n595036 , n595029 , n67711 );
or ( n67714 , n595032 , n595035 , n595036 );
and ( n595038 , n64838 , n66142 );
and ( n595039 , n592094 , n66140 );
nor ( n67717 , n595038 , n595039 );
xnor ( n595041 , n67717 , n592960 );
and ( n595042 , n64973 , n593256 );
and ( n67720 , n64854 , n593254 );
nor ( n595044 , n595042 , n67720 );
xnor ( n595045 , n595044 , n65490 );
and ( n67723 , n595041 , n595045 );
xor ( n595047 , n67676 , n595003 );
xor ( n67725 , n595047 , n595006 );
and ( n595049 , n595045 , n67725 );
and ( n67727 , n595041 , n67725 );
or ( n67728 , n67723 , n595049 , n67727 );
and ( n595052 , n592645 , n592683 );
and ( n67730 , n592468 , n592681 );
nor ( n595054 , n595052 , n67730 );
xnor ( n67732 , n595054 , n592475 );
xor ( n67733 , n594981 , n594991 );
xor ( n595057 , n67733 , n67673 );
and ( n67735 , n67732 , n595057 );
xor ( n595059 , n594929 , n594931 );
xor ( n67737 , n595059 , n594934 );
and ( n595061 , n595057 , n67737 );
and ( n595062 , n67732 , n67737 );
or ( n67740 , n67735 , n595061 , n595062 );
and ( n595064 , n592404 , n65592 );
and ( n595065 , n64997 , n592913 );
nor ( n595066 , n595064 , n595065 );
xnor ( n67744 , n595066 , n592638 );
and ( n595068 , n67740 , n67744 );
xor ( n595069 , n67614 , n594941 );
xor ( n67747 , n595069 , n594944 );
and ( n595071 , n67744 , n67747 );
and ( n595072 , n67740 , n67747 );
or ( n67750 , n595068 , n595071 , n595072 );
and ( n595074 , n67728 , n67750 );
and ( n595075 , n591851 , n594441 );
and ( n67753 , n64501 , n67116 );
nor ( n67754 , n595075 , n67753 );
xnor ( n595078 , n67754 , n66190 );
and ( n67756 , n67750 , n595078 );
and ( n67757 , n67728 , n595078 );
or ( n595081 , n595074 , n67756 , n67757 );
and ( n595082 , n593437 , n64862 );
and ( n67760 , n593298 , n64860 );
nor ( n595084 , n595082 , n67760 );
xnor ( n595085 , n595084 , n64764 );
and ( n67763 , n66606 , n64650 );
and ( n595087 , n66507 , n64648 );
nor ( n595088 , n67763 , n595087 );
xnor ( n67766 , n595088 , n591902 );
and ( n595090 , n595085 , n67766 );
and ( n67768 , n66793 , n64559 );
and ( n595092 , n594124 , n591880 );
nor ( n67770 , n67768 , n595092 );
xnor ( n595094 , n67770 , n64521 );
and ( n595095 , n67766 , n595094 );
and ( n67773 , n595085 , n595094 );
or ( n595097 , n595090 , n595095 , n67773 );
xor ( n595098 , n594958 , n594960 );
and ( n67776 , n67636 , n64456 );
and ( n67777 , n594952 , n64454 );
nor ( n595101 , n67776 , n67777 );
xnor ( n67779 , n595101 , n591786 );
buf ( n595103 , n591708 );
and ( n595104 , n595103 , n64451 );
and ( n67782 , n67779 , n595104 );
and ( n595106 , n595098 , n67782 );
and ( n67784 , n594295 , n64491 );
and ( n595108 , n66967 , n64489 );
nor ( n595109 , n67784 , n595108 );
xnor ( n67787 , n595109 , n64448 );
and ( n595111 , n67782 , n67787 );
and ( n595112 , n595098 , n67787 );
or ( n67790 , n595106 , n595111 , n595112 );
and ( n67791 , n593520 , n64744 );
and ( n595115 , n66104 , n64742 );
nor ( n67793 , n67791 , n595115 );
xnor ( n595117 , n67793 , n64623 );
and ( n67795 , n67790 , n595117 );
xor ( n67796 , n594954 , n594961 );
xor ( n595120 , n67796 , n67643 );
and ( n595121 , n595117 , n595120 );
and ( n67799 , n67790 , n595120 );
or ( n595123 , n67795 , n595121 , n67799 );
and ( n595124 , n595097 , n595123 );
and ( n67802 , n65630 , n592340 );
and ( n595126 , n65640 , n65015 );
nor ( n595127 , n67802 , n595126 );
xnor ( n595128 , n595127 , n64847 );
and ( n595129 , n595123 , n595128 );
and ( n67807 , n595097 , n595128 );
or ( n595131 , n595124 , n595129 , n67807 );
and ( n595132 , n593298 , n64862 );
and ( n595133 , n65844 , n64860 );
nor ( n67811 , n595132 , n595133 );
xnor ( n595135 , n67811 , n64764 );
and ( n595136 , n594124 , n64559 );
and ( n67814 , n66606 , n591880 );
nor ( n595138 , n595136 , n67814 );
xnor ( n595139 , n595138 , n64521 );
and ( n67817 , n595135 , n595139 );
xor ( n595141 , n594982 , n67660 );
xor ( n595142 , n595141 , n594988 );
and ( n67820 , n595139 , n595142 );
and ( n595144 , n595135 , n595142 );
or ( n595145 , n67817 , n67820 , n595144 );
and ( n67823 , n595131 , n595145 );
and ( n595147 , n65493 , n592486 );
and ( n595148 , n65384 , n592484 );
nor ( n67826 , n595147 , n595148 );
xnor ( n595150 , n67826 , n64990 );
and ( n595151 , n595145 , n595150 );
and ( n67829 , n595131 , n595150 );
or ( n67830 , n67823 , n595151 , n67829 );
and ( n67831 , n592468 , n592683 );
and ( n595155 , n592478 , n592681 );
nor ( n595156 , n67831 , n595155 );
xnor ( n67834 , n595156 , n592475 );
and ( n595158 , n67830 , n67834 );
xor ( n595159 , n67447 , n67451 );
xor ( n67837 , n595159 , n67456 );
and ( n67838 , n67834 , n67837 );
and ( n595162 , n67830 , n67837 );
or ( n67840 , n595158 , n67838 , n595162 );
and ( n67841 , n64586 , n594210 );
and ( n595165 , n64533 , n66885 );
nor ( n595166 , n67841 , n595165 );
xnor ( n595167 , n595166 , n593434 );
and ( n595168 , n67840 , n595167 );
xor ( n67846 , n594947 , n595009 );
xor ( n595170 , n67846 , n67689 );
and ( n595171 , n595167 , n595170 );
and ( n67849 , n67840 , n595170 );
or ( n595173 , n595168 , n595171 , n67849 );
and ( n595174 , n595081 , n595173 );
xor ( n67852 , n67602 , n595015 );
xor ( n595176 , n67852 , n67695 );
and ( n595177 , n595173 , n595176 );
and ( n67855 , n595081 , n595176 );
or ( n595179 , n595174 , n595177 , n67855 );
and ( n67857 , n67714 , n595179 );
xor ( n595181 , n67494 , n594821 );
xor ( n67859 , n595181 , n594824 );
and ( n595183 , n595179 , n67859 );
and ( n595184 , n67714 , n67859 );
or ( n595185 , n67857 , n595183 , n595184 );
and ( n595186 , n67704 , n595185 );
xor ( n67864 , n594813 , n67504 );
xor ( n595188 , n67864 , n67507 );
and ( n595189 , n595185 , n595188 );
and ( n67867 , n67704 , n595188 );
or ( n595191 , n595186 , n595189 , n67867 );
xor ( n595192 , n594678 , n67357 );
xor ( n67870 , n595192 , n67360 );
and ( n595194 , n595191 , n67870 );
xor ( n595195 , n67510 , n594865 );
xor ( n67873 , n595195 , n594868 );
and ( n595197 , n67870 , n67873 );
and ( n67875 , n595191 , n67873 );
or ( n595199 , n595194 , n595197 , n67875 );
and ( n67877 , n67560 , n595199 );
xor ( n67878 , n67560 , n595199 );
xor ( n67879 , n595191 , n67870 );
xor ( n67880 , n67879 , n67873 );
and ( n67881 , n64466 , n594807 );
and ( n67882 , n64450 , n594804 );
nor ( n67883 , n67881 , n67882 );
xnor ( n67884 , n67883 , n66187 );
xor ( n67885 , n67590 , n67594 );
xor ( n67886 , n67885 , n67599 );
and ( n67887 , n67884 , n67886 );
xor ( n67888 , n67564 , n67568 );
xor ( n595212 , n67888 , n67571 );
and ( n67890 , n67886 , n595212 );
and ( n595214 , n67884 , n595212 );
or ( n595215 , n67887 , n67890 , n595214 );
xor ( n67893 , n594897 , n67578 );
xor ( n67894 , n67893 , n67583 );
and ( n67895 , n595215 , n67894 );
xor ( n67896 , n595029 , n595031 );
xor ( n67897 , n67896 , n67711 );
and ( n595221 , n67894 , n67897 );
and ( n67899 , n595215 , n67897 );
or ( n595223 , n67895 , n595221 , n67899 );
xor ( n67901 , n67586 , n595021 );
xor ( n595225 , n67901 , n595024 );
and ( n595226 , n595223 , n595225 );
xor ( n67904 , n594849 , n67528 );
xor ( n595228 , n67904 , n67531 );
and ( n595229 , n595225 , n595228 );
and ( n67907 , n595223 , n595228 );
or ( n67908 , n595226 , n595229 , n67907 );
xor ( n595232 , n67534 , n594859 );
xor ( n67910 , n595232 , n594862 );
and ( n595234 , n67908 , n67910 );
xor ( n595235 , n67704 , n595185 );
xor ( n595236 , n595235 , n595188 );
and ( n67914 , n67910 , n595236 );
and ( n595238 , n67908 , n595236 );
or ( n595239 , n595234 , n67914 , n595238 );
and ( n67917 , n67880 , n595239 );
xor ( n67918 , n67880 , n595239 );
and ( n595242 , n66104 , n64862 );
and ( n595243 , n593437 , n64860 );
nor ( n67921 , n595242 , n595243 );
xnor ( n67922 , n67921 , n64764 );
and ( n67923 , n66507 , n64744 );
and ( n595247 , n593520 , n64742 );
nor ( n67925 , n67923 , n595247 );
xnor ( n595249 , n67925 , n64623 );
and ( n67927 , n67922 , n595249 );
and ( n595251 , n594124 , n64650 );
and ( n595252 , n66606 , n64648 );
nor ( n67930 , n595251 , n595252 );
xnor ( n67931 , n67930 , n591902 );
and ( n67932 , n595249 , n67931 );
and ( n595256 , n67922 , n67931 );
or ( n595257 , n67927 , n67932 , n595256 );
xor ( n595258 , n67779 , n595104 );
and ( n595259 , n595103 , n64456 );
and ( n67937 , n67636 , n64454 );
nor ( n595261 , n595259 , n67937 );
xnor ( n595262 , n595261 , n591786 );
buf ( n67940 , n591709 );
and ( n67941 , n67940 , n64451 );
and ( n595265 , n595262 , n67941 );
and ( n67943 , n595258 , n595265 );
and ( n67944 , n594710 , n64491 );
and ( n595268 , n594295 , n64489 );
nor ( n595269 , n67944 , n595268 );
xnor ( n595270 , n595269 , n64448 );
and ( n595271 , n595265 , n595270 );
and ( n67949 , n595258 , n595270 );
or ( n595273 , n67943 , n595271 , n67949 );
and ( n595274 , n66951 , n64559 );
and ( n67952 , n66793 , n591880 );
nor ( n595276 , n595274 , n67952 );
xnor ( n595277 , n595276 , n64521 );
and ( n67955 , n595273 , n595277 );
xor ( n595279 , n595098 , n67782 );
xor ( n67957 , n595279 , n67787 );
and ( n67958 , n595277 , n67957 );
and ( n595282 , n595273 , n67957 );
or ( n67960 , n67955 , n67958 , n595282 );
and ( n595284 , n595257 , n67960 );
and ( n595285 , n65844 , n592340 );
and ( n67963 , n65630 , n65015 );
nor ( n595287 , n595285 , n67963 );
xnor ( n67965 , n595287 , n64847 );
and ( n67966 , n67960 , n67965 );
and ( n595290 , n595257 , n67965 );
or ( n67968 , n595284 , n67966 , n595290 );
and ( n595292 , n592806 , n592486 );
and ( n67970 , n65493 , n592484 );
nor ( n595294 , n595292 , n67970 );
xnor ( n67972 , n595294 , n64990 );
and ( n67973 , n67968 , n67972 );
xor ( n67974 , n594969 , n594973 );
xor ( n67975 , n67974 , n67655 );
and ( n595299 , n67972 , n67975 );
and ( n67977 , n67968 , n67975 );
or ( n595301 , n67973 , n595299 , n67977 );
and ( n595302 , n65640 , n592486 );
and ( n595303 , n592806 , n592484 );
nor ( n67981 , n595302 , n595303 );
xnor ( n595305 , n67981 , n64990 );
xor ( n67983 , n595085 , n67766 );
xor ( n595307 , n67983 , n595094 );
and ( n595308 , n595305 , n595307 );
xor ( n67986 , n67790 , n595117 );
xor ( n595310 , n67986 , n595120 );
and ( n67988 , n595307 , n595310 );
and ( n595312 , n595305 , n595310 );
or ( n67990 , n595308 , n67988 , n595312 );
and ( n67991 , n65384 , n592683 );
and ( n595315 , n592645 , n592681 );
nor ( n67993 , n67991 , n595315 );
xnor ( n595317 , n67993 , n592475 );
and ( n595318 , n67990 , n595317 );
xor ( n67996 , n595135 , n595139 );
xor ( n595320 , n67996 , n595142 );
and ( n595321 , n595317 , n595320 );
and ( n595322 , n67990 , n595320 );
or ( n68000 , n595318 , n595321 , n595322 );
and ( n595324 , n595301 , n68000 );
and ( n595325 , n592478 , n65592 );
and ( n68003 , n592404 , n592913 );
nor ( n595327 , n595325 , n68003 );
xnor ( n595328 , n595327 , n592638 );
and ( n68006 , n68000 , n595328 );
and ( n68007 , n595301 , n595328 );
or ( n595331 , n595324 , n68006 , n68007 );
and ( n68009 , n64501 , n594807 );
and ( n595333 , n64466 , n594804 );
nor ( n68011 , n68009 , n595333 );
xnor ( n595335 , n68011 , n66187 );
and ( n595336 , n595331 , n595335 );
and ( n68014 , n64533 , n594441 );
and ( n595338 , n591851 , n67116 );
nor ( n595339 , n68014 , n595338 );
xnor ( n68017 , n595339 , n66190 );
and ( n68018 , n595335 , n68017 );
and ( n595342 , n595331 , n68017 );
or ( n595343 , n595336 , n68018 , n595342 );
and ( n68021 , n64591 , n594210 );
and ( n595345 , n64586 , n66885 );
nor ( n595346 , n68021 , n595345 );
xnor ( n68024 , n595346 , n593434 );
and ( n595348 , n64683 , n66457 );
and ( n595349 , n64630 , n593778 );
nor ( n595350 , n595348 , n595349 );
xnor ( n68028 , n595350 , n593160 );
and ( n595352 , n68024 , n68028 );
xor ( n595353 , n67830 , n67834 );
xor ( n68031 , n595353 , n67837 );
and ( n595355 , n68028 , n68031 );
and ( n595356 , n68024 , n68031 );
or ( n68034 , n595352 , n595355 , n595356 );
and ( n595358 , n595343 , n68034 );
xor ( n68036 , n67840 , n595167 );
xor ( n595360 , n68036 , n595170 );
and ( n68038 , n68034 , n595360 );
and ( n68039 , n595343 , n595360 );
or ( n595363 , n595358 , n68038 , n68039 );
and ( n595364 , n592094 , n66457 );
and ( n68042 , n64683 , n593778 );
nor ( n595366 , n595364 , n68042 );
xnor ( n595367 , n595366 , n593160 );
and ( n68045 , n64854 , n66142 );
and ( n595369 , n64838 , n66140 );
nor ( n595370 , n68045 , n595369 );
xnor ( n595371 , n595370 , n592960 );
and ( n68049 , n595367 , n595371 );
and ( n595373 , n64997 , n593256 );
and ( n68051 , n64973 , n593254 );
nor ( n595375 , n595373 , n68051 );
xnor ( n68053 , n595375 , n65490 );
and ( n595377 , n595371 , n68053 );
and ( n595378 , n595367 , n68053 );
or ( n68056 , n68049 , n595377 , n595378 );
and ( n595380 , n64630 , n594210 );
and ( n595381 , n64591 , n66885 );
nor ( n68059 , n595380 , n595381 );
xnor ( n595383 , n68059 , n593434 );
xor ( n595384 , n595131 , n595145 );
xor ( n68062 , n595384 , n595150 );
and ( n595386 , n595383 , n68062 );
xor ( n595387 , n67732 , n595057 );
xor ( n595388 , n595387 , n67737 );
and ( n68066 , n68062 , n595388 );
and ( n595390 , n595383 , n595388 );
or ( n68068 , n595386 , n68066 , n595390 );
and ( n68069 , n68056 , n68068 );
xor ( n595393 , n595041 , n595045 );
xor ( n595394 , n595393 , n67725 );
and ( n68072 , n68068 , n595394 );
and ( n595396 , n68056 , n595394 );
or ( n595397 , n68069 , n68072 , n595396 );
xor ( n68075 , n67728 , n67750 );
xor ( n595399 , n68075 , n595078 );
and ( n595400 , n595397 , n595399 );
xor ( n595401 , n67884 , n67886 );
xor ( n68079 , n595401 , n595212 );
and ( n595403 , n595399 , n68079 );
and ( n68081 , n595397 , n68079 );
or ( n68082 , n595400 , n595403 , n68081 );
and ( n68083 , n595363 , n68082 );
xor ( n68084 , n595081 , n595173 );
xor ( n68085 , n68084 , n595176 );
and ( n68086 , n68082 , n68085 );
and ( n68087 , n595363 , n68085 );
or ( n68088 , n68083 , n68086 , n68087 );
xor ( n68089 , n67714 , n595179 );
xor ( n68090 , n68089 , n67859 );
and ( n68091 , n68088 , n68090 );
xor ( n68092 , n595223 , n595225 );
xor ( n68093 , n68092 , n595228 );
and ( n68094 , n68090 , n68093 );
and ( n68095 , n68088 , n68093 );
or ( n68096 , n68091 , n68094 , n68095 );
xor ( n68097 , n67908 , n67910 );
xor ( n68098 , n68097 , n595236 );
and ( n68099 , n68096 , n68098 );
xor ( n68100 , n68096 , n68098 );
xor ( n68101 , n68088 , n68090 );
xor ( n595425 , n68101 , n68093 );
and ( n68103 , n592645 , n65592 );
and ( n595427 , n592468 , n592913 );
nor ( n595428 , n68103 , n595427 );
xnor ( n68106 , n595428 , n592638 );
xor ( n595430 , n595257 , n67960 );
xor ( n595431 , n595430 , n67965 );
and ( n68109 , n68106 , n595431 );
xor ( n595433 , n595305 , n595307 );
xor ( n595434 , n595433 , n595310 );
and ( n68112 , n595431 , n595434 );
and ( n68113 , n68106 , n595434 );
or ( n595437 , n68109 , n68112 , n68113 );
and ( n68115 , n64838 , n66457 );
and ( n595439 , n592094 , n593778 );
nor ( n595440 , n68115 , n595439 );
xnor ( n68118 , n595440 , n593160 );
and ( n595442 , n595437 , n68118 );
and ( n595443 , n592404 , n593256 );
and ( n595444 , n64997 , n593254 );
nor ( n68122 , n595443 , n595444 );
xnor ( n595446 , n68122 , n65490 );
and ( n595447 , n68118 , n595446 );
and ( n68125 , n595437 , n595446 );
or ( n595449 , n595442 , n595447 , n68125 );
and ( n595450 , n592468 , n65592 );
and ( n68128 , n592478 , n592913 );
nor ( n68129 , n595450 , n68128 );
xnor ( n595453 , n68129 , n592638 );
xor ( n595454 , n595097 , n595123 );
xor ( n68132 , n595454 , n595128 );
and ( n595456 , n595453 , n68132 );
xor ( n595457 , n67968 , n67972 );
xor ( n68135 , n595457 , n67975 );
and ( n595459 , n68132 , n68135 );
and ( n595460 , n595453 , n68135 );
or ( n68138 , n595456 , n595459 , n595460 );
and ( n68139 , n595449 , n68138 );
and ( n68140 , n64586 , n594441 );
and ( n68141 , n64533 , n67116 );
nor ( n68142 , n68140 , n68141 );
xnor ( n68143 , n68142 , n66190 );
and ( n595467 , n68138 , n68143 );
and ( n68145 , n595449 , n68143 );
or ( n595469 , n68139 , n595467 , n68145 );
xor ( n595470 , n67740 , n67744 );
xor ( n68148 , n595470 , n67747 );
and ( n595472 , n595469 , n68148 );
xor ( n68150 , n68024 , n68028 );
xor ( n595474 , n68150 , n68031 );
and ( n68152 , n68148 , n595474 );
and ( n595476 , n595469 , n595474 );
or ( n68154 , n595472 , n68152 , n595476 );
xor ( n68155 , n595262 , n67941 );
and ( n68156 , n67940 , n64456 );
and ( n68157 , n595103 , n64454 );
nor ( n68158 , n68156 , n68157 );
xnor ( n68159 , n68158 , n591786 );
buf ( n68160 , n591710 );
and ( n68161 , n68160 , n64451 );
and ( n68162 , n68159 , n68161 );
and ( n595486 , n68155 , n68162 );
and ( n595487 , n594952 , n64491 );
and ( n595488 , n594710 , n64489 );
nor ( n68166 , n595487 , n595488 );
xnor ( n595490 , n68166 , n64448 );
and ( n595491 , n68162 , n595490 );
and ( n68169 , n68155 , n595490 );
or ( n595493 , n595486 , n595491 , n68169 );
and ( n595494 , n66967 , n64559 );
and ( n68172 , n66951 , n591880 );
nor ( n68173 , n595494 , n68172 );
xnor ( n595497 , n68173 , n64521 );
and ( n68175 , n595493 , n595497 );
xor ( n68176 , n595258 , n595265 );
xor ( n595500 , n68176 , n595270 );
and ( n595501 , n595497 , n595500 );
and ( n68179 , n595493 , n595500 );
or ( n595503 , n68175 , n595501 , n68179 );
and ( n595504 , n65630 , n592486 );
and ( n68182 , n65640 , n592484 );
nor ( n68183 , n595504 , n68182 );
xnor ( n68184 , n68183 , n64990 );
and ( n68185 , n595503 , n68184 );
and ( n68186 , n593298 , n592340 );
and ( n68187 , n65844 , n65015 );
nor ( n68188 , n68186 , n68187 );
xnor ( n68189 , n68188 , n64847 );
and ( n68190 , n68184 , n68189 );
and ( n595514 , n595503 , n68189 );
or ( n68192 , n68185 , n68190 , n595514 );
xor ( n595516 , n68159 , n68161 );
and ( n595517 , n595103 , n64491 );
and ( n68195 , n67636 , n64489 );
nor ( n595519 , n595517 , n68195 );
xnor ( n595520 , n595519 , n64448 );
buf ( n595521 , n591711 );
and ( n68199 , n595521 , n64451 );
and ( n595523 , n595520 , n68199 );
and ( n595524 , n595516 , n595523 );
and ( n68202 , n67636 , n64491 );
and ( n595526 , n594952 , n64489 );
nor ( n595527 , n68202 , n595526 );
xnor ( n68205 , n595527 , n64448 );
and ( n68206 , n595523 , n68205 );
and ( n68207 , n595516 , n68205 );
or ( n68208 , n595524 , n68206 , n68207 );
and ( n68209 , n594295 , n64559 );
and ( n68210 , n66967 , n591880 );
nor ( n595534 , n68209 , n68210 );
xnor ( n68212 , n595534 , n64521 );
and ( n595536 , n68208 , n68212 );
xor ( n595537 , n68155 , n68162 );
xor ( n68215 , n595537 , n595490 );
and ( n595539 , n68212 , n68215 );
and ( n595540 , n68208 , n68215 );
or ( n595541 , n595536 , n595539 , n595540 );
and ( n68219 , n66606 , n64744 );
and ( n68220 , n66507 , n64742 );
nor ( n68221 , n68219 , n68220 );
xnor ( n68222 , n68221 , n64623 );
and ( n68223 , n595541 , n68222 );
and ( n68224 , n66793 , n64650 );
and ( n68225 , n594124 , n64648 );
nor ( n68226 , n68224 , n68225 );
xnor ( n68227 , n68226 , n591902 );
and ( n68228 , n68222 , n68227 );
and ( n595552 , n595541 , n68227 );
or ( n68230 , n68223 , n68228 , n595552 );
and ( n595554 , n593437 , n592340 );
and ( n595555 , n593298 , n65015 );
nor ( n68233 , n595554 , n595555 );
xnor ( n595557 , n68233 , n64847 );
and ( n595558 , n593520 , n64862 );
and ( n68236 , n66104 , n64860 );
nor ( n595560 , n595558 , n68236 );
xnor ( n595561 , n595560 , n64764 );
and ( n68239 , n595557 , n595561 );
xor ( n68240 , n595493 , n595497 );
xor ( n595564 , n68240 , n595500 );
and ( n595565 , n595561 , n595564 );
and ( n68243 , n595557 , n595564 );
or ( n595567 , n68239 , n595565 , n68243 );
and ( n595568 , n68230 , n595567 );
xor ( n68246 , n595273 , n595277 );
xor ( n595570 , n68246 , n67957 );
and ( n595571 , n595567 , n595570 );
and ( n68249 , n68230 , n595570 );
or ( n595573 , n595568 , n595571 , n68249 );
and ( n595574 , n68192 , n595573 );
and ( n68252 , n65493 , n592683 );
and ( n595576 , n65384 , n592681 );
nor ( n595577 , n68252 , n595576 );
xnor ( n68255 , n595577 , n592475 );
and ( n68256 , n595573 , n68255 );
and ( n68257 , n68192 , n68255 );
or ( n595581 , n595574 , n68256 , n68257 );
and ( n595582 , n64973 , n66142 );
and ( n68260 , n64854 , n66140 );
nor ( n68261 , n595582 , n68260 );
xnor ( n595585 , n68261 , n592960 );
and ( n595586 , n595581 , n595585 );
xor ( n68264 , n67990 , n595317 );
xor ( n595588 , n68264 , n595320 );
and ( n595589 , n595585 , n595588 );
and ( n68267 , n595581 , n595588 );
or ( n595591 , n595586 , n595589 , n68267 );
and ( n68269 , n591851 , n594807 );
and ( n595593 , n64501 , n594804 );
nor ( n68271 , n68269 , n595593 );
xnor ( n595595 , n68271 , n66187 );
and ( n68273 , n595591 , n595595 );
xor ( n68274 , n595301 , n68000 );
xor ( n595598 , n68274 , n595328 );
and ( n68276 , n595595 , n595598 );
and ( n68277 , n595591 , n595598 );
or ( n595601 , n68273 , n68276 , n68277 );
xor ( n595602 , n595331 , n595335 );
xor ( n68280 , n595602 , n68017 );
and ( n595604 , n595601 , n68280 );
xor ( n595605 , n68056 , n68068 );
xor ( n68283 , n595605 , n595394 );
and ( n595607 , n68280 , n68283 );
and ( n595608 , n595601 , n68283 );
or ( n68286 , n595604 , n595607 , n595608 );
and ( n68287 , n68154 , n68286 );
xor ( n595611 , n595343 , n68034 );
xor ( n68289 , n595611 , n595360 );
and ( n595613 , n68286 , n68289 );
and ( n595614 , n68154 , n68289 );
or ( n595615 , n68287 , n595613 , n595614 );
xor ( n68293 , n595215 , n67894 );
xor ( n595617 , n68293 , n67897 );
and ( n595618 , n595615 , n595617 );
xor ( n68296 , n595363 , n68082 );
xor ( n595620 , n68296 , n68085 );
and ( n595621 , n595617 , n595620 );
and ( n595622 , n595615 , n595620 );
or ( n68300 , n595618 , n595621 , n595622 );
and ( n595624 , n595425 , n68300 );
xor ( n595625 , n595425 , n68300 );
xor ( n68303 , n595615 , n595617 );
xor ( n595627 , n68303 , n595620 );
xor ( n68305 , n595520 , n68199 );
and ( n68306 , n595521 , n64456 );
and ( n68307 , n68160 , n64454 );
nor ( n595631 , n68306 , n68307 );
xnor ( n68309 , n595631 , n591786 );
buf ( n595633 , n591712 );
and ( n595634 , n595633 , n64451 );
and ( n68312 , n68309 , n595634 );
and ( n68313 , n68305 , n68312 );
and ( n595637 , n68160 , n64456 );
and ( n68315 , n67940 , n64454 );
nor ( n68316 , n595637 , n68315 );
xnor ( n595640 , n68316 , n591786 );
and ( n68318 , n68312 , n595640 );
and ( n595642 , n68305 , n595640 );
or ( n68320 , n68313 , n68318 , n595642 );
and ( n595644 , n66967 , n64650 );
and ( n68322 , n66951 , n64648 );
nor ( n68323 , n595644 , n68322 );
xnor ( n68324 , n68323 , n591902 );
and ( n68325 , n68320 , n68324 );
and ( n68326 , n594710 , n64559 );
and ( n68327 , n594295 , n591880 );
nor ( n68328 , n68326 , n68327 );
xnor ( n68329 , n68328 , n64521 );
and ( n68330 , n68324 , n68329 );
and ( n68331 , n68320 , n68329 );
or ( n68332 , n68325 , n68330 , n68331 );
and ( n68333 , n66507 , n64862 );
and ( n68334 , n593520 , n64860 );
nor ( n68335 , n68333 , n68334 );
xnor ( n68336 , n68335 , n64764 );
and ( n68337 , n68332 , n68336 );
and ( n68338 , n66951 , n64650 );
and ( n68339 , n66793 , n64648 );
nor ( n68340 , n68338 , n68339 );
xnor ( n68341 , n68340 , n591902 );
and ( n68342 , n68336 , n68341 );
and ( n68343 , n68332 , n68341 );
or ( n68344 , n68337 , n68342 , n68343 );
and ( n68345 , n66104 , n592340 );
and ( n68346 , n593437 , n65015 );
nor ( n68347 , n68345 , n68346 );
xnor ( n68348 , n68347 , n64847 );
and ( n68349 , n594124 , n64744 );
and ( n595673 , n66606 , n64742 );
nor ( n68351 , n68349 , n595673 );
xnor ( n595675 , n68351 , n64623 );
and ( n595676 , n68348 , n595675 );
xor ( n68354 , n68208 , n68212 );
xor ( n595678 , n68354 , n68215 );
and ( n68356 , n595675 , n595678 );
and ( n68357 , n68348 , n595678 );
or ( n68358 , n595676 , n68356 , n68357 );
and ( n68359 , n68344 , n68358 );
and ( n68360 , n65844 , n592486 );
and ( n68361 , n65630 , n592484 );
nor ( n68362 , n68360 , n68361 );
xnor ( n68363 , n68362 , n64990 );
and ( n68364 , n68358 , n68363 );
and ( n595688 , n68344 , n68363 );
or ( n68366 , n68359 , n68364 , n595688 );
and ( n595690 , n592806 , n592683 );
and ( n595691 , n65493 , n592681 );
nor ( n68369 , n595690 , n595691 );
xnor ( n595693 , n68369 , n592475 );
and ( n68371 , n68366 , n595693 );
xor ( n68372 , n67922 , n595249 );
xor ( n68373 , n68372 , n67931 );
and ( n68374 , n595693 , n68373 );
and ( n68375 , n68366 , n68373 );
or ( n68376 , n68371 , n68374 , n68375 );
and ( n68377 , n65384 , n65592 );
and ( n68378 , n592645 , n592913 );
nor ( n68379 , n68377 , n68378 );
xnor ( n68380 , n68379 , n592638 );
xor ( n68381 , n595503 , n68184 );
xor ( n68382 , n68381 , n68189 );
and ( n68383 , n68380 , n68382 );
xor ( n68384 , n68230 , n595567 );
xor ( n68385 , n68384 , n595570 );
and ( n68386 , n68382 , n68385 );
and ( n68387 , n68380 , n68385 );
or ( n595711 , n68383 , n68386 , n68387 );
and ( n68389 , n68376 , n595711 );
and ( n595713 , n64854 , n66457 );
and ( n68391 , n64838 , n593778 );
nor ( n68392 , n595713 , n68391 );
xnor ( n68393 , n68392 , n593160 );
and ( n68394 , n595711 , n68393 );
and ( n68395 , n68376 , n68393 );
or ( n595719 , n68389 , n68394 , n68395 );
and ( n68397 , n592094 , n594210 );
and ( n595721 , n64683 , n66885 );
nor ( n68399 , n68397 , n595721 );
xnor ( n595723 , n68399 , n593434 );
and ( n595724 , n64997 , n66142 );
and ( n68402 , n64973 , n66140 );
nor ( n595726 , n595724 , n68402 );
xnor ( n68404 , n595726 , n592960 );
and ( n595728 , n595723 , n68404 );
xor ( n68406 , n68192 , n595573 );
xor ( n595730 , n68406 , n68255 );
and ( n595731 , n68404 , n595730 );
and ( n68409 , n595723 , n595730 );
or ( n595733 , n595728 , n595731 , n68409 );
and ( n595734 , n595719 , n595733 );
xor ( n68412 , n595453 , n68132 );
xor ( n595736 , n68412 , n68135 );
and ( n595737 , n595733 , n595736 );
and ( n595738 , n595719 , n595736 );
or ( n595739 , n595734 , n595737 , n595738 );
xor ( n68417 , n595449 , n68138 );
xor ( n68418 , n68417 , n68143 );
and ( n595742 , n595739 , n68418 );
xor ( n68420 , n595591 , n595595 );
xor ( n68421 , n68420 , n595598 );
and ( n595745 , n68418 , n68421 );
and ( n595746 , n595739 , n68421 );
or ( n68424 , n595742 , n595745 , n595746 );
and ( n595748 , n64533 , n594807 );
and ( n595749 , n591851 , n594804 );
nor ( n68427 , n595748 , n595749 );
xnor ( n595751 , n68427 , n66187 );
and ( n595752 , n64591 , n594441 );
and ( n68430 , n64586 , n67116 );
nor ( n68431 , n595752 , n68430 );
xnor ( n68432 , n68431 , n66190 );
and ( n68433 , n595751 , n68432 );
and ( n68434 , n64683 , n594210 );
and ( n68435 , n64630 , n66885 );
nor ( n595759 , n68434 , n68435 );
xnor ( n68437 , n595759 , n593434 );
and ( n595761 , n68432 , n68437 );
and ( n68439 , n595751 , n68437 );
or ( n595763 , n68433 , n595761 , n68439 );
xor ( n595764 , n595367 , n595371 );
xor ( n68442 , n595764 , n68053 );
and ( n595766 , n595763 , n68442 );
xor ( n595767 , n595383 , n68062 );
xor ( n68445 , n595767 , n595388 );
and ( n68446 , n68442 , n68445 );
and ( n595770 , n595763 , n68445 );
or ( n68448 , n595766 , n68446 , n595770 );
and ( n595772 , n68424 , n68448 );
xor ( n595773 , n595469 , n68148 );
xor ( n68451 , n595773 , n595474 );
and ( n595775 , n68448 , n68451 );
and ( n595776 , n68424 , n68451 );
or ( n68454 , n595772 , n595775 , n595776 );
xor ( n595778 , n595397 , n595399 );
xor ( n68456 , n595778 , n68079 );
and ( n595780 , n68454 , n68456 );
xor ( n595781 , n68154 , n68286 );
xor ( n68459 , n595781 , n68289 );
and ( n595783 , n68456 , n68459 );
and ( n595784 , n68454 , n68459 );
or ( n68462 , n595780 , n595783 , n595784 );
and ( n68463 , n595627 , n68462 );
xor ( n595787 , n595627 , n68462 );
xor ( n68465 , n68454 , n68456 );
xor ( n68466 , n68465 , n68459 );
and ( n68467 , n65640 , n592683 );
and ( n68468 , n592806 , n592681 );
nor ( n68469 , n68467 , n68468 );
xnor ( n595793 , n68469 , n592475 );
xor ( n595794 , n595541 , n68222 );
xor ( n68472 , n595794 , n68227 );
and ( n595796 , n595793 , n68472 );
xor ( n595797 , n595557 , n595561 );
xor ( n595798 , n595797 , n595564 );
and ( n68476 , n68472 , n595798 );
and ( n595800 , n595793 , n595798 );
or ( n68478 , n595796 , n68476 , n595800 );
and ( n68479 , n592468 , n593256 );
and ( n68480 , n592478 , n593254 );
nor ( n68481 , n68479 , n68480 );
xnor ( n68482 , n68481 , n65490 );
and ( n68483 , n68478 , n68482 );
xor ( n68484 , n68366 , n595693 );
xor ( n68485 , n68484 , n68373 );
and ( n68486 , n68482 , n68485 );
and ( n595810 , n68478 , n68485 );
or ( n68488 , n68483 , n68486 , n595810 );
and ( n595812 , n64586 , n594807 );
and ( n595813 , n64533 , n594804 );
nor ( n68491 , n595812 , n595813 );
xnor ( n68492 , n68491 , n66187 );
and ( n595816 , n68488 , n68492 );
xor ( n68494 , n68376 , n595711 );
xor ( n595818 , n68494 , n68393 );
and ( n595819 , n68492 , n595818 );
and ( n595820 , n68488 , n595818 );
or ( n68498 , n595816 , n595819 , n595820 );
xor ( n595822 , n68309 , n595634 );
and ( n595823 , n595633 , n64456 );
and ( n68501 , n595521 , n64454 );
nor ( n595825 , n595823 , n68501 );
xnor ( n595826 , n595825 , n591786 );
buf ( n595827 , n591713 );
and ( n68505 , n595827 , n64451 );
and ( n595829 , n595826 , n68505 );
and ( n595830 , n595822 , n595829 );
and ( n68508 , n67940 , n64491 );
and ( n595832 , n595103 , n64489 );
nor ( n595833 , n68508 , n595832 );
xnor ( n68511 , n595833 , n64448 );
and ( n595835 , n595829 , n68511 );
and ( n595836 , n595822 , n68511 );
or ( n68514 , n595830 , n595835 , n595836 );
and ( n595838 , n594295 , n64650 );
and ( n595839 , n66967 , n64648 );
nor ( n68517 , n595838 , n595839 );
xnor ( n68518 , n68517 , n591902 );
and ( n68519 , n68514 , n68518 );
and ( n595843 , n594952 , n64559 );
and ( n595844 , n594710 , n591880 );
nor ( n68522 , n595843 , n595844 );
xnor ( n595846 , n68522 , n64521 );
and ( n595847 , n68518 , n595846 );
and ( n68525 , n68514 , n595846 );
or ( n595849 , n68519 , n595847 , n68525 );
and ( n68527 , n66606 , n64862 );
and ( n595851 , n66507 , n64860 );
nor ( n68529 , n68527 , n595851 );
xnor ( n595853 , n68529 , n64764 );
and ( n68531 , n595849 , n595853 );
xor ( n595855 , n595516 , n595523 );
xor ( n595856 , n595855 , n68205 );
and ( n68534 , n595853 , n595856 );
and ( n68535 , n595849 , n595856 );
or ( n595859 , n68531 , n68534 , n68535 );
and ( n595860 , n65630 , n592683 );
and ( n68538 , n65640 , n592681 );
nor ( n595862 , n595860 , n68538 );
xnor ( n595863 , n595862 , n592475 );
and ( n68541 , n595859 , n595863 );
and ( n595865 , n593298 , n592486 );
and ( n595866 , n65844 , n592484 );
nor ( n68544 , n595865 , n595866 );
xnor ( n68545 , n68544 , n64990 );
and ( n595869 , n595863 , n68545 );
and ( n595870 , n595859 , n68545 );
or ( n68548 , n68541 , n595869 , n595870 );
and ( n595872 , n65493 , n65592 );
and ( n595873 , n65384 , n592913 );
nor ( n68551 , n595872 , n595873 );
xnor ( n595875 , n68551 , n592638 );
and ( n68553 , n68548 , n595875 );
xor ( n68554 , n68344 , n68358 );
xor ( n595878 , n68554 , n68363 );
and ( n68556 , n595875 , n595878 );
and ( n68557 , n68548 , n595878 );
or ( n68558 , n68553 , n68556 , n68557 );
and ( n68559 , n593520 , n592340 );
and ( n68560 , n66104 , n65015 );
nor ( n595884 , n68559 , n68560 );
xnor ( n68562 , n595884 , n64847 );
and ( n68563 , n66793 , n64744 );
and ( n595887 , n594124 , n64742 );
nor ( n595888 , n68563 , n595887 );
xnor ( n68566 , n595888 , n64623 );
and ( n595890 , n68562 , n68566 );
xor ( n595891 , n68320 , n68324 );
xor ( n68569 , n595891 , n68329 );
and ( n595893 , n68566 , n68569 );
and ( n68571 , n68562 , n68569 );
or ( n68572 , n595890 , n595893 , n68571 );
xor ( n68573 , n68332 , n68336 );
xor ( n68574 , n68573 , n68341 );
and ( n68575 , n68572 , n68574 );
xor ( n68576 , n68348 , n595675 );
xor ( n68577 , n68576 , n595678 );
and ( n68578 , n68574 , n68577 );
and ( n68579 , n68572 , n68577 );
or ( n68580 , n68575 , n68578 , n68579 );
and ( n68581 , n592645 , n593256 );
and ( n68582 , n592468 , n593254 );
nor ( n68583 , n68581 , n68582 );
xnor ( n68584 , n68583 , n65490 );
and ( n68585 , n68580 , n68584 );
xor ( n68586 , n595793 , n68472 );
xor ( n595910 , n68586 , n595798 );
and ( n68588 , n68584 , n595910 );
and ( n595912 , n68580 , n595910 );
or ( n68590 , n68585 , n68588 , n595912 );
and ( n68591 , n68558 , n68590 );
and ( n68592 , n64973 , n66457 );
and ( n68593 , n64854 , n593778 );
nor ( n68594 , n68592 , n68593 );
xnor ( n595918 , n68594 , n593160 );
and ( n68596 , n68590 , n595918 );
and ( n595920 , n68558 , n595918 );
or ( n68598 , n68591 , n68596 , n595920 );
and ( n595922 , n64838 , n594210 );
and ( n595923 , n592094 , n66885 );
nor ( n68601 , n595922 , n595923 );
xnor ( n595925 , n68601 , n593434 );
and ( n68603 , n592404 , n66142 );
and ( n68604 , n64997 , n66140 );
nor ( n68605 , n68603 , n68604 );
xnor ( n68606 , n68605 , n592960 );
and ( n68607 , n595925 , n68606 );
xor ( n68608 , n68380 , n68382 );
xor ( n595932 , n68608 , n68385 );
and ( n68610 , n68606 , n595932 );
and ( n68611 , n595925 , n595932 );
or ( n595935 , n68607 , n68610 , n68611 );
and ( n595936 , n68598 , n595935 );
xor ( n68614 , n595723 , n68404 );
xor ( n595938 , n68614 , n595730 );
and ( n595939 , n595935 , n595938 );
and ( n68617 , n68598 , n595938 );
or ( n595941 , n595936 , n595939 , n68617 );
and ( n68619 , n68498 , n595941 );
xor ( n595943 , n595751 , n68432 );
xor ( n595944 , n595943 , n68437 );
and ( n68622 , n595941 , n595944 );
and ( n595946 , n68498 , n595944 );
or ( n595947 , n68619 , n68622 , n595946 );
and ( n68625 , n64630 , n594441 );
and ( n595949 , n64591 , n67116 );
nor ( n68627 , n68625 , n595949 );
xnor ( n595951 , n68627 , n66190 );
and ( n595952 , n592478 , n593256 );
and ( n68630 , n592404 , n593254 );
nor ( n595954 , n595952 , n68630 );
xnor ( n595955 , n595954 , n65490 );
and ( n68633 , n595951 , n595955 );
xor ( n68634 , n68106 , n595431 );
xor ( n595958 , n68634 , n595434 );
and ( n595959 , n595955 , n595958 );
and ( n68637 , n595951 , n595958 );
or ( n595961 , n68633 , n595959 , n68637 );
xor ( n595962 , n595437 , n68118 );
xor ( n68640 , n595962 , n595446 );
and ( n595964 , n595961 , n68640 );
xor ( n595965 , n595581 , n595585 );
xor ( n68643 , n595965 , n595588 );
and ( n595967 , n68640 , n68643 );
and ( n595968 , n595961 , n68643 );
or ( n68646 , n595964 , n595967 , n595968 );
and ( n595970 , n595947 , n68646 );
xor ( n68648 , n595763 , n68442 );
xor ( n595972 , n68648 , n68445 );
and ( n595973 , n68646 , n595972 );
and ( n68651 , n595947 , n595972 );
or ( n595975 , n595970 , n595973 , n68651 );
xor ( n68653 , n595601 , n68280 );
xor ( n595977 , n68653 , n68283 );
and ( n595978 , n595975 , n595977 );
xor ( n68656 , n68424 , n68448 );
xor ( n68657 , n68656 , n68451 );
and ( n595981 , n595977 , n68657 );
and ( n595982 , n595975 , n68657 );
or ( n68660 , n595978 , n595981 , n595982 );
and ( n68661 , n68466 , n68660 );
xor ( n595985 , n68466 , n68660 );
xor ( n68663 , n595975 , n595977 );
xor ( n595987 , n68663 , n68657 );
and ( n68665 , n64591 , n594807 );
and ( n595989 , n64586 , n594804 );
nor ( n595990 , n68665 , n595989 );
xnor ( n68668 , n595990 , n66187 );
and ( n595992 , n64683 , n594441 );
and ( n595993 , n64630 , n67116 );
nor ( n68671 , n595992 , n595993 );
xnor ( n595995 , n68671 , n66190 );
and ( n595996 , n68668 , n595995 );
xor ( n68674 , n68478 , n68482 );
xor ( n68675 , n68674 , n68485 );
and ( n595999 , n595995 , n68675 );
and ( n68677 , n68668 , n68675 );
or ( n68678 , n595996 , n595999 , n68677 );
xor ( n596002 , n68488 , n68492 );
xor ( n596003 , n596002 , n595818 );
and ( n68681 , n68678 , n596003 );
xor ( n596005 , n595951 , n595955 );
xor ( n596006 , n596005 , n595958 );
and ( n68684 , n596003 , n596006 );
and ( n68685 , n68678 , n596006 );
or ( n596009 , n68681 , n68684 , n68685 );
xor ( n596010 , n595719 , n595733 );
xor ( n68688 , n596010 , n595736 );
and ( n596012 , n596009 , n68688 );
xor ( n596013 , n595961 , n68640 );
xor ( n68691 , n596013 , n68643 );
and ( n596015 , n68688 , n68691 );
and ( n68693 , n596009 , n68691 );
or ( n596017 , n596012 , n596015 , n68693 );
xor ( n68695 , n595739 , n68418 );
xor ( n68696 , n68695 , n68421 );
and ( n68697 , n596017 , n68696 );
xor ( n596021 , n595947 , n68646 );
xor ( n596022 , n596021 , n595972 );
and ( n68700 , n68696 , n596022 );
and ( n596024 , n596017 , n596022 );
or ( n596025 , n68697 , n68700 , n596024 );
and ( n596026 , n595987 , n596025 );
xor ( n68704 , n595987 , n596025 );
xor ( n596028 , n596017 , n68696 );
xor ( n68706 , n596028 , n596022 );
and ( n68707 , n64630 , n594807 );
and ( n596031 , n64591 , n594804 );
nor ( n68709 , n68707 , n596031 );
xnor ( n596033 , n68709 , n66187 );
and ( n596034 , n64854 , n594210 );
and ( n68712 , n64838 , n66885 );
nor ( n596036 , n596034 , n68712 );
xnor ( n596037 , n596036 , n593434 );
and ( n596038 , n596033 , n596037 );
xor ( n68716 , n68580 , n68584 );
xor ( n596040 , n68716 , n595910 );
and ( n596041 , n596037 , n596040 );
and ( n68719 , n596033 , n596040 );
or ( n596043 , n596038 , n596041 , n68719 );
xor ( n596044 , n68558 , n68590 );
xor ( n68722 , n596044 , n595918 );
and ( n596046 , n596043 , n68722 );
xor ( n596047 , n68668 , n595995 );
xor ( n68725 , n596047 , n68675 );
and ( n596049 , n68722 , n68725 );
and ( n68727 , n596043 , n68725 );
or ( n68728 , n596046 , n596049 , n68727 );
xor ( n596052 , n595826 , n68505 );
and ( n68730 , n595827 , n64456 );
and ( n596054 , n595633 , n64454 );
nor ( n68732 , n68730 , n596054 );
xnor ( n596056 , n68732 , n591786 );
buf ( n596057 , n591714 );
and ( n68735 , n596057 , n64451 );
and ( n68736 , n596056 , n68735 );
and ( n596060 , n596052 , n68736 );
and ( n68738 , n595103 , n64559 );
and ( n596062 , n67636 , n591880 );
nor ( n68740 , n68738 , n596062 );
xnor ( n596064 , n68740 , n64521 );
and ( n596065 , n68736 , n596064 );
and ( n68743 , n596052 , n596064 );
or ( n596067 , n596060 , n596065 , n68743 );
and ( n596068 , n594710 , n64650 );
and ( n596069 , n594295 , n64648 );
nor ( n68747 , n596068 , n596069 );
xnor ( n68748 , n68747 , n591902 );
and ( n596072 , n596067 , n68748 );
and ( n68750 , n67636 , n64559 );
and ( n596074 , n594952 , n591880 );
nor ( n68752 , n68750 , n596074 );
xnor ( n68753 , n68752 , n64521 );
and ( n596077 , n68748 , n68753 );
and ( n68755 , n596067 , n68753 );
or ( n68756 , n596072 , n596077 , n68755 );
xor ( n596080 , n68514 , n68518 );
xor ( n68758 , n596080 , n595846 );
and ( n68759 , n68756 , n68758 );
xor ( n68760 , n68305 , n68312 );
xor ( n596084 , n68760 , n595640 );
and ( n68762 , n68758 , n596084 );
and ( n68763 , n68756 , n596084 );
or ( n596087 , n68759 , n68762 , n68763 );
and ( n596088 , n65844 , n592683 );
and ( n68766 , n65630 , n592681 );
nor ( n596090 , n596088 , n68766 );
xnor ( n596091 , n596090 , n592475 );
and ( n68769 , n596087 , n596091 );
and ( n596093 , n593437 , n592486 );
and ( n68771 , n593298 , n592484 );
nor ( n596095 , n596093 , n68771 );
xnor ( n68773 , n596095 , n64990 );
and ( n596097 , n596091 , n68773 );
and ( n596098 , n596087 , n68773 );
or ( n68776 , n68769 , n596097 , n596098 );
and ( n596100 , n592806 , n65592 );
and ( n68778 , n65493 , n592913 );
nor ( n596102 , n596100 , n68778 );
xnor ( n68780 , n596102 , n592638 );
and ( n68781 , n68776 , n68780 );
xor ( n68782 , n595859 , n595863 );
xor ( n596106 , n68782 , n68545 );
and ( n68784 , n68780 , n596106 );
and ( n596108 , n68776 , n596106 );
or ( n68786 , n68781 , n68784 , n596108 );
and ( n68787 , n66507 , n592340 );
and ( n596111 , n593520 , n65015 );
nor ( n68789 , n68787 , n596111 );
xnor ( n68790 , n68789 , n64847 );
and ( n596114 , n594124 , n64862 );
and ( n596115 , n66606 , n64860 );
nor ( n68793 , n596114 , n596115 );
xnor ( n596117 , n68793 , n64764 );
and ( n596118 , n68790 , n596117 );
and ( n68796 , n66951 , n64744 );
and ( n596120 , n66793 , n64742 );
nor ( n596121 , n68796 , n596120 );
xnor ( n68799 , n596121 , n64623 );
and ( n68800 , n596117 , n68799 );
and ( n596124 , n68790 , n68799 );
or ( n68802 , n596118 , n68800 , n596124 );
and ( n68803 , n65640 , n65592 );
and ( n596127 , n592806 , n592913 );
nor ( n68805 , n68803 , n596127 );
xnor ( n596129 , n68805 , n592638 );
and ( n596130 , n68802 , n596129 );
xor ( n68808 , n595849 , n595853 );
xor ( n68809 , n68808 , n595856 );
and ( n596133 , n596129 , n68809 );
and ( n596134 , n68802 , n68809 );
or ( n68812 , n596130 , n596133 , n596134 );
and ( n596136 , n65384 , n593256 );
and ( n596137 , n592645 , n593254 );
nor ( n68815 , n596136 , n596137 );
xnor ( n596139 , n68815 , n65490 );
and ( n596140 , n68812 , n596139 );
xor ( n596141 , n68572 , n68574 );
xor ( n68819 , n596141 , n68577 );
and ( n596143 , n596139 , n68819 );
and ( n596144 , n68812 , n68819 );
or ( n68822 , n596140 , n596143 , n596144 );
and ( n596146 , n68786 , n68822 );
and ( n596147 , n592478 , n66142 );
and ( n68825 , n592404 , n66140 );
nor ( n68826 , n596147 , n68825 );
xnor ( n68827 , n68826 , n592960 );
and ( n596151 , n68822 , n68827 );
and ( n68829 , n68786 , n68827 );
or ( n596153 , n596146 , n596151 , n68829 );
and ( n68831 , n592094 , n594441 );
and ( n68832 , n64683 , n67116 );
nor ( n596156 , n68831 , n68832 );
xnor ( n68834 , n596156 , n66190 );
and ( n596158 , n64997 , n66457 );
and ( n68836 , n64973 , n593778 );
nor ( n68837 , n596158 , n68836 );
xnor ( n68838 , n68837 , n593160 );
and ( n68839 , n68834 , n68838 );
xor ( n68840 , n68548 , n595875 );
xor ( n68841 , n68840 , n595878 );
and ( n68842 , n68838 , n68841 );
and ( n68843 , n68834 , n68841 );
or ( n68844 , n68839 , n68842 , n68843 );
and ( n68845 , n596153 , n68844 );
xor ( n596169 , n595925 , n68606 );
xor ( n68847 , n596169 , n595932 );
and ( n596171 , n68844 , n68847 );
and ( n596172 , n596153 , n68847 );
or ( n596173 , n68845 , n596171 , n596172 );
and ( n68851 , n68728 , n596173 );
xor ( n596175 , n68598 , n595935 );
xor ( n596176 , n596175 , n595938 );
and ( n68854 , n596173 , n596176 );
and ( n596178 , n68728 , n596176 );
or ( n596179 , n68851 , n68854 , n596178 );
xor ( n68857 , n68498 , n595941 );
xor ( n596181 , n68857 , n595944 );
and ( n68859 , n596179 , n596181 );
xor ( n596183 , n596009 , n68688 );
xor ( n68861 , n596183 , n68691 );
and ( n596185 , n596181 , n68861 );
and ( n68863 , n596179 , n68861 );
or ( n596187 , n68859 , n596185 , n68863 );
and ( n596188 , n68706 , n596187 );
xor ( n68866 , n68706 , n596187 );
xor ( n596190 , n596179 , n596181 );
xor ( n596191 , n596190 , n68861 );
xor ( n68869 , n596056 , n68735 );
buf ( n596193 , n591715 );
and ( n596194 , n596193 , n64456 );
and ( n68872 , n596057 , n64454 );
nor ( n68873 , n596194 , n68872 );
xnor ( n596197 , n68873 , n591786 );
buf ( n596198 , n591716 );
and ( n68876 , n596198 , n64451 );
and ( n596200 , n596197 , n68876 );
and ( n596201 , n596193 , n64451 );
and ( n68879 , n596200 , n596201 );
and ( n596203 , n68869 , n68879 );
and ( n596204 , n595521 , n64491 );
and ( n68882 , n68160 , n64489 );
nor ( n68883 , n596204 , n68882 );
xnor ( n596207 , n68883 , n64448 );
and ( n596208 , n68879 , n596207 );
and ( n68886 , n68869 , n596207 );
or ( n596210 , n596203 , n596208 , n68886 );
and ( n68888 , n594952 , n64650 );
and ( n596212 , n594710 , n64648 );
nor ( n596213 , n68888 , n596212 );
xnor ( n68891 , n596213 , n591902 );
and ( n68892 , n596210 , n68891 );
and ( n596216 , n68160 , n64491 );
and ( n596217 , n67940 , n64489 );
nor ( n68895 , n596216 , n596217 );
xnor ( n596219 , n68895 , n64448 );
and ( n596220 , n68891 , n596219 );
and ( n68898 , n596210 , n596219 );
or ( n596222 , n68892 , n596220 , n68898 );
and ( n596223 , n66967 , n64744 );
and ( n68901 , n66951 , n64742 );
nor ( n596225 , n596223 , n68901 );
xnor ( n596226 , n596225 , n64623 );
and ( n68904 , n596222 , n596226 );
xor ( n596228 , n595822 , n595829 );
xor ( n596229 , n596228 , n68511 );
and ( n68907 , n596226 , n596229 );
and ( n596231 , n596222 , n596229 );
or ( n596232 , n68904 , n68907 , n596231 );
and ( n68910 , n66104 , n592486 );
and ( n596234 , n593437 , n592484 );
nor ( n596235 , n68910 , n596234 );
xnor ( n68913 , n596235 , n64990 );
and ( n68914 , n596232 , n68913 );
xor ( n596238 , n68756 , n68758 );
xor ( n68916 , n596238 , n596084 );
and ( n596240 , n68913 , n68916 );
and ( n68918 , n596232 , n68916 );
or ( n596242 , n68914 , n596240 , n68918 );
xor ( n596243 , n596087 , n596091 );
xor ( n68921 , n596243 , n68773 );
and ( n596245 , n596242 , n68921 );
xor ( n68923 , n68562 , n68566 );
xor ( n596247 , n68923 , n68569 );
and ( n596248 , n68921 , n596247 );
and ( n68926 , n596242 , n596247 );
or ( n68927 , n596245 , n596248 , n68926 );
and ( n596251 , n592468 , n66142 );
and ( n68929 , n592478 , n66140 );
nor ( n596253 , n596251 , n68929 );
xnor ( n596254 , n596253 , n592960 );
and ( n68932 , n68927 , n596254 );
xor ( n596256 , n68776 , n68780 );
xor ( n596257 , n596256 , n596106 );
and ( n596258 , n596254 , n596257 );
and ( n68936 , n68927 , n596257 );
or ( n596260 , n68932 , n596258 , n68936 );
xor ( n68938 , n596200 , n596201 );
and ( n596262 , n595633 , n64491 );
and ( n68940 , n595521 , n64489 );
nor ( n596264 , n596262 , n68940 );
xnor ( n596265 , n596264 , n64448 );
and ( n68943 , n68938 , n596265 );
and ( n596267 , n596057 , n64456 );
and ( n596268 , n595827 , n64454 );
nor ( n68946 , n596267 , n596268 );
xnor ( n68947 , n68946 , n591786 );
and ( n596271 , n596265 , n68947 );
and ( n596272 , n68938 , n68947 );
or ( n68950 , n68943 , n596271 , n596272 );
and ( n596274 , n67636 , n64650 );
and ( n596275 , n594952 , n64648 );
nor ( n68953 , n596274 , n596275 );
xnor ( n596277 , n68953 , n591902 );
and ( n596278 , n68950 , n596277 );
and ( n68956 , n67940 , n64559 );
and ( n68957 , n595103 , n591880 );
nor ( n596281 , n68956 , n68957 );
xnor ( n68959 , n596281 , n64521 );
and ( n596283 , n596277 , n68959 );
and ( n68961 , n68950 , n68959 );
or ( n68962 , n596278 , n596283 , n68961 );
and ( n596286 , n594295 , n64744 );
and ( n596287 , n66967 , n64742 );
nor ( n68965 , n596286 , n596287 );
xnor ( n596289 , n68965 , n64623 );
and ( n596290 , n68962 , n596289 );
xor ( n68968 , n596052 , n68736 );
xor ( n596292 , n68968 , n596064 );
and ( n596293 , n596289 , n596292 );
and ( n596294 , n68962 , n596292 );
or ( n68972 , n596290 , n596293 , n596294 );
and ( n596296 , n66606 , n592340 );
and ( n596297 , n66507 , n65015 );
nor ( n68975 , n596296 , n596297 );
xnor ( n596299 , n68975 , n64847 );
and ( n596300 , n68972 , n596299 );
xor ( n68978 , n596067 , n68748 );
xor ( n596302 , n68978 , n68753 );
and ( n68980 , n596299 , n596302 );
and ( n596304 , n68972 , n596302 );
or ( n68982 , n596300 , n68980 , n596304 );
and ( n596306 , n65630 , n65592 );
and ( n68984 , n65640 , n592913 );
nor ( n596308 , n596306 , n68984 );
xnor ( n596309 , n596308 , n592638 );
and ( n68987 , n68982 , n596309 );
and ( n596311 , n593298 , n592683 );
and ( n596312 , n65844 , n592681 );
nor ( n68990 , n596311 , n596312 );
xnor ( n68991 , n68990 , n592475 );
and ( n596315 , n596309 , n68991 );
and ( n596316 , n68982 , n68991 );
or ( n68994 , n68987 , n596315 , n596316 );
and ( n596318 , n65493 , n593256 );
and ( n596319 , n65384 , n593254 );
nor ( n68997 , n596318 , n596319 );
xnor ( n596321 , n68997 , n65490 );
and ( n596322 , n68994 , n596321 );
xor ( n69000 , n68802 , n596129 );
xor ( n69001 , n69000 , n68809 );
and ( n596325 , n596321 , n69001 );
and ( n69003 , n68994 , n69001 );
or ( n596327 , n596322 , n596325 , n69003 );
and ( n69005 , n64973 , n594210 );
and ( n69006 , n64854 , n66885 );
nor ( n596330 , n69005 , n69006 );
xnor ( n596331 , n596330 , n593434 );
and ( n69009 , n596327 , n596331 );
xor ( n596333 , n68812 , n596139 );
xor ( n596334 , n596333 , n68819 );
and ( n69012 , n596331 , n596334 );
and ( n596336 , n596327 , n596334 );
or ( n596337 , n69009 , n69012 , n596336 );
and ( n596338 , n596260 , n596337 );
xor ( n69016 , n68786 , n68822 );
xor ( n596340 , n69016 , n68827 );
and ( n596341 , n596337 , n596340 );
and ( n69019 , n596260 , n596340 );
or ( n596343 , n596338 , n596341 , n69019 );
xor ( n596344 , n596043 , n68722 );
xor ( n69022 , n596344 , n68725 );
and ( n69023 , n596343 , n69022 );
xor ( n596347 , n596153 , n68844 );
xor ( n69025 , n596347 , n68847 );
and ( n596349 , n69022 , n69025 );
and ( n596350 , n596343 , n69025 );
or ( n69028 , n69023 , n596349 , n596350 );
xor ( n596352 , n68728 , n596173 );
xor ( n69030 , n596352 , n596176 );
and ( n596354 , n69028 , n69030 );
xor ( n596355 , n68678 , n596003 );
xor ( n69033 , n596355 , n596006 );
and ( n69034 , n69030 , n69033 );
and ( n69035 , n69028 , n69033 );
or ( n69036 , n596354 , n69034 , n69035 );
and ( n69037 , n596191 , n69036 );
xor ( n69038 , n596191 , n69036 );
xor ( n69039 , n69028 , n69030 );
xor ( n69040 , n69039 , n69033 );
and ( n69041 , n66104 , n592683 );
and ( n69042 , n593437 , n592681 );
nor ( n69043 , n69041 , n69042 );
xnor ( n69044 , n69043 , n592475 );
and ( n596368 , n66507 , n592486 );
and ( n69046 , n593520 , n592484 );
nor ( n596370 , n596368 , n69046 );
xnor ( n596371 , n596370 , n64990 );
and ( n69049 , n69044 , n596371 );
xor ( n596373 , n68962 , n596289 );
xor ( n596374 , n596373 , n596292 );
and ( n69052 , n596371 , n596374 );
and ( n596376 , n69044 , n596374 );
or ( n596377 , n69049 , n69052 , n596376 );
xor ( n69055 , n68972 , n596299 );
xor ( n596379 , n69055 , n596302 );
and ( n596380 , n596377 , n596379 );
and ( n596381 , n593520 , n592486 );
and ( n69059 , n66104 , n592484 );
nor ( n596383 , n596381 , n69059 );
xnor ( n596384 , n596383 , n64990 );
and ( n596385 , n66793 , n64862 );
and ( n69063 , n594124 , n64860 );
nor ( n596387 , n596385 , n69063 );
xnor ( n69065 , n596387 , n64764 );
xor ( n69066 , n596384 , n69065 );
xor ( n69067 , n596222 , n596226 );
xor ( n596391 , n69067 , n596229 );
xor ( n596392 , n69066 , n596391 );
and ( n596393 , n596379 , n596392 );
and ( n69071 , n596377 , n596392 );
or ( n596395 , n596380 , n596393 , n69071 );
and ( n596396 , n65384 , n66142 );
and ( n69074 , n592645 , n66140 );
nor ( n596398 , n596396 , n69074 );
xnor ( n596399 , n596398 , n592960 );
and ( n69077 , n596395 , n596399 );
and ( n596401 , n596384 , n69065 );
and ( n69079 , n69065 , n596391 );
and ( n596403 , n596384 , n596391 );
or ( n69081 , n596401 , n69079 , n596403 );
xor ( n596405 , n68790 , n596117 );
xor ( n69083 , n596405 , n68799 );
xor ( n596407 , n69081 , n69083 );
xor ( n596408 , n596232 , n68913 );
xor ( n69086 , n596408 , n68916 );
xor ( n69087 , n596407 , n69086 );
and ( n596411 , n596399 , n69087 );
and ( n596412 , n596395 , n69087 );
or ( n69090 , n69077 , n596411 , n596412 );
and ( n596414 , n592094 , n594807 );
and ( n596415 , n64683 , n594804 );
nor ( n69093 , n596414 , n596415 );
xnor ( n596417 , n69093 , n66187 );
and ( n596418 , n69090 , n596417 );
and ( n69096 , n64854 , n594441 );
and ( n69097 , n64838 , n67116 );
nor ( n596421 , n69096 , n69097 );
xnor ( n596422 , n596421 , n66190 );
and ( n69100 , n596417 , n596422 );
and ( n596424 , n69090 , n596422 );
or ( n596425 , n596418 , n69100 , n596424 );
and ( n69103 , n64683 , n594807 );
and ( n596427 , n64630 , n594804 );
nor ( n596428 , n69103 , n596427 );
xnor ( n69106 , n596428 , n66187 );
and ( n596430 , n596425 , n69106 );
xor ( n596431 , n68927 , n596254 );
xor ( n69109 , n596431 , n596257 );
and ( n596433 , n69106 , n69109 );
and ( n596434 , n596425 , n69109 );
or ( n69112 , n596430 , n596433 , n596434 );
and ( n596436 , n595827 , n64491 );
and ( n596437 , n595633 , n64489 );
nor ( n69115 , n596436 , n596437 );
xnor ( n69116 , n69115 , n64448 );
xor ( n69117 , n596197 , n68876 );
and ( n596441 , n69116 , n69117 );
and ( n69119 , n595103 , n64650 );
and ( n596443 , n67636 , n64648 );
nor ( n69121 , n69119 , n596443 );
xnor ( n596445 , n69121 , n591902 );
and ( n596446 , n596441 , n596445 );
and ( n69124 , n68160 , n64559 );
and ( n69125 , n67940 , n591880 );
nor ( n596449 , n69124 , n69125 );
xnor ( n596450 , n596449 , n64521 );
and ( n69128 , n596445 , n596450 );
and ( n596452 , n596441 , n596450 );
or ( n596453 , n596446 , n69128 , n596452 );
and ( n69131 , n594710 , n64744 );
and ( n596455 , n594295 , n64742 );
nor ( n69133 , n69131 , n596455 );
xnor ( n69134 , n69133 , n64623 );
and ( n596458 , n596453 , n69134 );
xor ( n69136 , n68869 , n68879 );
xor ( n596460 , n69136 , n596207 );
and ( n69138 , n69134 , n596460 );
and ( n69139 , n596453 , n596460 );
or ( n596463 , n596458 , n69138 , n69139 );
and ( n596464 , n66951 , n64862 );
and ( n69142 , n66793 , n64860 );
nor ( n596466 , n596464 , n69142 );
xnor ( n596467 , n596466 , n64764 );
and ( n69145 , n596463 , n596467 );
xor ( n596469 , n596210 , n68891 );
xor ( n596470 , n596469 , n596219 );
and ( n596471 , n596467 , n596470 );
and ( n69149 , n596463 , n596470 );
or ( n596473 , n69145 , n596471 , n69149 );
and ( n69151 , n65844 , n65592 );
and ( n69152 , n65630 , n592913 );
nor ( n596476 , n69151 , n69152 );
xnor ( n69154 , n596476 , n592638 );
and ( n69155 , n596473 , n69154 );
and ( n596479 , n593437 , n592683 );
and ( n69157 , n593298 , n592681 );
nor ( n69158 , n596479 , n69157 );
xnor ( n596482 , n69158 , n592475 );
and ( n596483 , n69154 , n596482 );
and ( n69161 , n596473 , n596482 );
or ( n596485 , n69155 , n596483 , n69161 );
and ( n596486 , n592806 , n593256 );
and ( n69164 , n65493 , n593254 );
nor ( n596488 , n596486 , n69164 );
xnor ( n69166 , n596488 , n65490 );
and ( n69167 , n596485 , n69166 );
xor ( n596491 , n68982 , n596309 );
xor ( n69169 , n596491 , n68991 );
and ( n596493 , n69166 , n69169 );
and ( n69171 , n596485 , n69169 );
or ( n69172 , n69167 , n596493 , n69171 );
and ( n69173 , n64997 , n594210 );
and ( n69174 , n64973 , n66885 );
nor ( n596498 , n69173 , n69174 );
xnor ( n596499 , n596498 , n593434 );
and ( n69177 , n69172 , n596499 );
and ( n596501 , n592478 , n66457 );
and ( n69179 , n592404 , n593778 );
nor ( n69180 , n596501 , n69179 );
xnor ( n69181 , n69180 , n593160 );
and ( n596505 , n596499 , n69181 );
and ( n69183 , n69172 , n69181 );
or ( n596507 , n69177 , n596505 , n69183 );
and ( n69185 , n69081 , n69083 );
and ( n69186 , n69083 , n69086 );
and ( n596510 , n69081 , n69086 );
or ( n596511 , n69185 , n69186 , n596510 );
and ( n69189 , n592645 , n66142 );
and ( n596513 , n592468 , n66140 );
nor ( n596514 , n69189 , n596513 );
xnor ( n69192 , n596514 , n592960 );
and ( n596516 , n596511 , n69192 );
xor ( n69194 , n596242 , n68921 );
xor ( n69195 , n69194 , n596247 );
and ( n596519 , n69192 , n69195 );
and ( n69197 , n596511 , n69195 );
or ( n596521 , n596516 , n596519 , n69197 );
and ( n69199 , n64838 , n594441 );
and ( n596523 , n592094 , n67116 );
nor ( n596524 , n69199 , n596523 );
xnor ( n69202 , n596524 , n66190 );
xor ( n69203 , n596521 , n69202 );
and ( n596527 , n592404 , n66457 );
and ( n596528 , n64997 , n593778 );
nor ( n69206 , n596527 , n596528 );
xnor ( n596530 , n69206 , n593160 );
xor ( n596531 , n69203 , n596530 );
and ( n69209 , n596507 , n596531 );
xor ( n596533 , n596327 , n596331 );
xor ( n596534 , n596533 , n596334 );
and ( n596535 , n596531 , n596534 );
and ( n69213 , n596507 , n596534 );
or ( n596537 , n69209 , n596535 , n69213 );
and ( n69215 , n69112 , n596537 );
xor ( n69216 , n596260 , n596337 );
xor ( n596540 , n69216 , n596340 );
and ( n69218 , n596537 , n596540 );
and ( n596542 , n69112 , n596540 );
or ( n69220 , n69215 , n69218 , n596542 );
and ( n596544 , n596521 , n69202 );
and ( n596545 , n69202 , n596530 );
and ( n69223 , n596521 , n596530 );
or ( n69224 , n596544 , n596545 , n69223 );
xor ( n69225 , n68834 , n68838 );
xor ( n596549 , n69225 , n68841 );
and ( n69227 , n69224 , n596549 );
xor ( n69228 , n596033 , n596037 );
xor ( n69229 , n69228 , n596040 );
and ( n69230 , n596549 , n69229 );
and ( n69231 , n69224 , n69229 );
or ( n596555 , n69227 , n69230 , n69231 );
and ( n596556 , n69220 , n596555 );
xor ( n596557 , n596343 , n69022 );
xor ( n69235 , n596557 , n69025 );
and ( n596559 , n596555 , n69235 );
and ( n69237 , n69220 , n69235 );
or ( n596561 , n596556 , n596559 , n69237 );
and ( n69239 , n69040 , n596561 );
xor ( n69240 , n69040 , n596561 );
xor ( n596564 , n69220 , n596555 );
xor ( n69242 , n596564 , n69235 );
and ( n596566 , n65493 , n66142 );
and ( n596567 , n65384 , n66140 );
nor ( n69245 , n596566 , n596567 );
xnor ( n596569 , n69245 , n592960 );
xor ( n596570 , n596473 , n69154 );
xor ( n596571 , n596570 , n596482 );
and ( n69249 , n596569 , n596571 );
xor ( n596573 , n596377 , n596379 );
xor ( n596574 , n596573 , n596392 );
and ( n69252 , n596571 , n596574 );
and ( n596576 , n596569 , n596574 );
or ( n596577 , n69249 , n69252 , n596576 );
and ( n69255 , n64838 , n594807 );
and ( n69256 , n592094 , n594804 );
nor ( n596580 , n69255 , n69256 );
xnor ( n596581 , n596580 , n66187 );
and ( n69259 , n596577 , n596581 );
xor ( n596583 , n596395 , n596399 );
xor ( n596584 , n596583 , n69087 );
and ( n69262 , n596581 , n596584 );
and ( n596586 , n596577 , n596584 );
or ( n596587 , n69259 , n69262 , n596586 );
xor ( n596588 , n69090 , n596417 );
xor ( n69266 , n596588 , n596422 );
and ( n596590 , n596587 , n69266 );
xor ( n69268 , n69172 , n596499 );
xor ( n69269 , n69268 , n69181 );
and ( n596593 , n69266 , n69269 );
and ( n596594 , n596587 , n69269 );
or ( n69272 , n596590 , n596593 , n596594 );
and ( n596596 , n596193 , n64491 );
and ( n596597 , n596057 , n64489 );
nor ( n69275 , n596596 , n596597 );
xnor ( n596599 , n69275 , n64448 );
buf ( n596600 , n591717 );
and ( n69278 , n596600 , n64456 );
and ( n596602 , n596198 , n64454 );
nor ( n69280 , n69278 , n596602 );
xnor ( n596604 , n69280 , n591786 );
and ( n69282 , n596599 , n596604 );
buf ( n69283 , n591718 );
and ( n596607 , n69283 , n64451 );
and ( n596608 , n596604 , n596607 );
and ( n69286 , n596599 , n596607 );
or ( n596610 , n69282 , n596608 , n69286 );
and ( n596611 , n595633 , n64559 );
and ( n69289 , n595521 , n591880 );
nor ( n596613 , n596611 , n69289 );
xnor ( n596614 , n596613 , n64521 );
and ( n69292 , n596610 , n596614 );
and ( n596616 , n596057 , n64491 );
and ( n596617 , n595827 , n64489 );
nor ( n69295 , n596616 , n596617 );
xnor ( n596619 , n69295 , n64448 );
and ( n69297 , n596198 , n64456 );
and ( n596621 , n596193 , n64454 );
nor ( n596622 , n69297 , n596621 );
xnor ( n596623 , n596622 , n591786 );
xor ( n596624 , n596619 , n596623 );
and ( n69302 , n596600 , n64451 );
xor ( n69303 , n596624 , n69302 );
and ( n596627 , n596614 , n69303 );
and ( n69305 , n596610 , n69303 );
or ( n69306 , n69292 , n596627 , n69305 );
and ( n596630 , n67636 , n64744 );
and ( n69308 , n594952 , n64742 );
nor ( n596632 , n596630 , n69308 );
xnor ( n596633 , n596632 , n64623 );
and ( n69311 , n69306 , n596633 );
and ( n596635 , n67940 , n64650 );
and ( n596636 , n595103 , n64648 );
nor ( n69314 , n596635 , n596636 );
xnor ( n596638 , n69314 , n591902 );
and ( n596639 , n596633 , n596638 );
and ( n69317 , n69306 , n596638 );
or ( n69318 , n69311 , n596639 , n69317 );
and ( n596642 , n594295 , n64862 );
and ( n69320 , n66967 , n64860 );
nor ( n596644 , n596642 , n69320 );
xnor ( n69322 , n596644 , n64764 );
and ( n69323 , n69318 , n69322 );
xor ( n69324 , n596441 , n596445 );
xor ( n69325 , n69324 , n596450 );
and ( n69326 , n69322 , n69325 );
and ( n69327 , n69318 , n69325 );
or ( n69328 , n69323 , n69326 , n69327 );
and ( n69329 , n593520 , n592683 );
and ( n69330 , n66104 , n592681 );
nor ( n69331 , n69329 , n69330 );
xnor ( n69332 , n69331 , n592475 );
and ( n596656 , n69328 , n69332 );
xor ( n69334 , n596453 , n69134 );
xor ( n596658 , n69334 , n596460 );
and ( n69336 , n69332 , n596658 );
and ( n69337 , n69328 , n596658 );
or ( n596661 , n596656 , n69336 , n69337 );
and ( n69339 , n65630 , n593256 );
and ( n596663 , n65640 , n593254 );
nor ( n69341 , n69339 , n596663 );
xnor ( n596665 , n69341 , n65490 );
and ( n69343 , n596661 , n596665 );
and ( n69344 , n593298 , n65592 );
and ( n596668 , n65844 , n592913 );
nor ( n69346 , n69344 , n596668 );
xnor ( n596670 , n69346 , n592638 );
and ( n69348 , n596665 , n596670 );
and ( n596672 , n596661 , n596670 );
or ( n596673 , n69343 , n69348 , n596672 );
xor ( n69351 , n69116 , n69117 );
and ( n596675 , n596619 , n596623 );
and ( n596676 , n596623 , n69302 );
and ( n69354 , n596619 , n69302 );
or ( n596678 , n596675 , n596676 , n69354 );
and ( n596679 , n69351 , n596678 );
and ( n69357 , n595521 , n64559 );
and ( n69358 , n68160 , n591880 );
nor ( n596682 , n69357 , n69358 );
xnor ( n596683 , n596682 , n64521 );
and ( n69361 , n596678 , n596683 );
and ( n596685 , n69351 , n596683 );
or ( n596686 , n596679 , n69361 , n596685 );
and ( n69364 , n594952 , n64744 );
and ( n596688 , n594710 , n64742 );
nor ( n596689 , n69364 , n596688 );
xnor ( n596690 , n596689 , n64623 );
and ( n69368 , n596686 , n596690 );
xor ( n596692 , n68938 , n596265 );
xor ( n596693 , n596692 , n68947 );
and ( n69371 , n596690 , n596693 );
and ( n596695 , n596686 , n596693 );
or ( n596696 , n69368 , n69371 , n596695 );
and ( n69374 , n66967 , n64862 );
and ( n69375 , n66951 , n64860 );
nor ( n69376 , n69374 , n69375 );
xnor ( n69377 , n69376 , n64764 );
and ( n596701 , n596696 , n69377 );
xor ( n69379 , n68950 , n596277 );
xor ( n596703 , n69379 , n68959 );
and ( n596704 , n69377 , n596703 );
and ( n69382 , n596696 , n596703 );
or ( n596706 , n596701 , n596704 , n69382 );
and ( n69384 , n594124 , n592340 );
and ( n596708 , n66606 , n65015 );
nor ( n69386 , n69384 , n596708 );
xnor ( n596710 , n69386 , n64847 );
and ( n69388 , n596706 , n596710 );
xor ( n69389 , n596463 , n596467 );
xor ( n69390 , n69389 , n596470 );
and ( n69391 , n596710 , n69390 );
and ( n596715 , n596706 , n69390 );
or ( n69393 , n69388 , n69391 , n596715 );
and ( n596717 , n596673 , n69393 );
and ( n69395 , n65640 , n593256 );
and ( n596719 , n592806 , n593254 );
nor ( n596720 , n69395 , n596719 );
xnor ( n69398 , n596720 , n65490 );
and ( n596722 , n69393 , n69398 );
and ( n596723 , n596673 , n69398 );
or ( n69401 , n596717 , n596722 , n596723 );
and ( n69402 , n592468 , n66457 );
and ( n69403 , n592478 , n593778 );
nor ( n69404 , n69402 , n69403 );
xnor ( n69405 , n69404 , n593160 );
and ( n596729 , n69401 , n69405 );
xor ( n69407 , n596485 , n69166 );
xor ( n596731 , n69407 , n69169 );
and ( n69409 , n69405 , n596731 );
and ( n69410 , n69401 , n596731 );
or ( n596734 , n596729 , n69409 , n69410 );
xor ( n596735 , n68994 , n596321 );
xor ( n69413 , n596735 , n69001 );
and ( n596737 , n596734 , n69413 );
xor ( n596738 , n596511 , n69192 );
xor ( n69416 , n596738 , n69195 );
and ( n596740 , n69413 , n69416 );
and ( n596741 , n596734 , n69416 );
or ( n69419 , n596737 , n596740 , n596741 );
and ( n69420 , n69272 , n69419 );
xor ( n69421 , n596425 , n69106 );
xor ( n596745 , n69421 , n69109 );
and ( n596746 , n69419 , n596745 );
and ( n69424 , n69272 , n596745 );
or ( n69425 , n69420 , n596746 , n69424 );
xor ( n69426 , n69112 , n596537 );
xor ( n596750 , n69426 , n596540 );
and ( n596751 , n69425 , n596750 );
xor ( n69429 , n69224 , n596549 );
xor ( n69430 , n69429 , n69229 );
and ( n69431 , n596750 , n69430 );
and ( n69432 , n69425 , n69430 );
or ( n69433 , n596751 , n69431 , n69432 );
and ( n69434 , n69242 , n69433 );
xor ( n69435 , n69242 , n69433 );
xor ( n596759 , n69425 , n596750 );
xor ( n69437 , n596759 , n69430 );
and ( n596761 , n66606 , n592486 );
and ( n69439 , n66507 , n592484 );
nor ( n596763 , n596761 , n69439 );
xnor ( n69441 , n596763 , n64990 );
and ( n596765 , n66793 , n592340 );
and ( n69443 , n594124 , n65015 );
nor ( n596767 , n596765 , n69443 );
xnor ( n596768 , n596767 , n64847 );
and ( n69446 , n69441 , n596768 );
xor ( n596770 , n596696 , n69377 );
xor ( n596771 , n596770 , n596703 );
and ( n69449 , n596768 , n596771 );
and ( n69450 , n69441 , n596771 );
or ( n596774 , n69446 , n69449 , n69450 );
xor ( n69452 , n69044 , n596371 );
xor ( n596776 , n69452 , n596374 );
and ( n596777 , n596774 , n596776 );
xor ( n596778 , n596706 , n596710 );
xor ( n69456 , n596778 , n69390 );
and ( n596780 , n596776 , n69456 );
and ( n596781 , n596774 , n69456 );
or ( n69459 , n596777 , n596780 , n596781 );
and ( n596783 , n592645 , n66457 );
and ( n596784 , n592468 , n593778 );
nor ( n69462 , n596783 , n596784 );
xnor ( n69463 , n69462 , n593160 );
and ( n69464 , n69459 , n69463 );
xor ( n596788 , n596673 , n69393 );
xor ( n69466 , n596788 , n69398 );
and ( n596790 , n69463 , n69466 );
and ( n69468 , n69459 , n69466 );
or ( n69469 , n69464 , n596790 , n69468 );
and ( n596793 , n64973 , n594441 );
and ( n69471 , n64854 , n67116 );
nor ( n596795 , n596793 , n69471 );
xnor ( n69473 , n596795 , n66190 );
and ( n69474 , n69469 , n69473 );
and ( n596798 , n592404 , n594210 );
and ( n69476 , n64997 , n66885 );
nor ( n596800 , n596798 , n69476 );
xnor ( n69478 , n596800 , n593434 );
and ( n596802 , n69473 , n69478 );
and ( n69480 , n69469 , n69478 );
or ( n596804 , n69474 , n596802 , n69480 );
and ( n69482 , n596198 , n64491 );
and ( n596806 , n596193 , n64489 );
nor ( n69484 , n69482 , n596806 );
xnor ( n596808 , n69484 , n64448 );
and ( n69486 , n69283 , n64456 );
and ( n596810 , n596600 , n64454 );
nor ( n69488 , n69486 , n596810 );
xnor ( n596812 , n69488 , n591786 );
and ( n69490 , n596808 , n596812 );
buf ( n69491 , n591719 );
and ( n596815 , n69491 , n64451 );
and ( n596816 , n596812 , n596815 );
and ( n69494 , n596808 , n596815 );
or ( n596818 , n69490 , n596816 , n69494 );
and ( n69496 , n595827 , n64559 );
and ( n69497 , n595633 , n591880 );
nor ( n69498 , n69496 , n69497 );
xnor ( n69499 , n69498 , n64521 );
and ( n69500 , n596818 , n69499 );
xor ( n69501 , n596599 , n596604 );
xor ( n596825 , n69501 , n596607 );
and ( n69503 , n69499 , n596825 );
and ( n69504 , n596818 , n596825 );
or ( n69505 , n69500 , n69503 , n69504 );
and ( n69506 , n595103 , n64744 );
and ( n69507 , n67636 , n64742 );
nor ( n596831 , n69506 , n69507 );
xnor ( n69509 , n596831 , n64623 );
and ( n596833 , n69505 , n69509 );
and ( n596834 , n68160 , n64650 );
and ( n69512 , n67940 , n64648 );
nor ( n596836 , n596834 , n69512 );
xnor ( n69514 , n596836 , n591902 );
and ( n69515 , n69509 , n69514 );
and ( n596839 , n69505 , n69514 );
or ( n596840 , n596833 , n69515 , n596839 );
and ( n69518 , n594710 , n64862 );
and ( n69519 , n594295 , n64860 );
nor ( n596843 , n69518 , n69519 );
xnor ( n596844 , n596843 , n64764 );
and ( n69522 , n596840 , n596844 );
xor ( n596846 , n69351 , n596678 );
xor ( n596847 , n596846 , n596683 );
and ( n69525 , n596844 , n596847 );
and ( n596849 , n596840 , n596847 );
or ( n69527 , n69522 , n69525 , n596849 );
and ( n596851 , n66951 , n592340 );
and ( n69529 , n66793 , n65015 );
nor ( n69530 , n596851 , n69529 );
xnor ( n596854 , n69530 , n64847 );
and ( n596855 , n69527 , n596854 );
xor ( n69533 , n596686 , n596690 );
xor ( n596857 , n69533 , n596693 );
and ( n596858 , n596854 , n596857 );
and ( n69536 , n69527 , n596857 );
or ( n596860 , n596855 , n596858 , n69536 );
and ( n596861 , n593437 , n65592 );
and ( n69539 , n593298 , n592913 );
nor ( n69540 , n596861 , n69539 );
xnor ( n596864 , n69540 , n592638 );
and ( n69542 , n596860 , n596864 );
xor ( n596866 , n69328 , n69332 );
xor ( n69544 , n596866 , n596658 );
and ( n596868 , n596864 , n69544 );
and ( n596869 , n596860 , n69544 );
or ( n69547 , n69542 , n596868 , n596869 );
and ( n69548 , n65384 , n66457 );
and ( n596872 , n592645 , n593778 );
nor ( n69550 , n69548 , n596872 );
xnor ( n596874 , n69550 , n593160 );
and ( n69552 , n69547 , n596874 );
and ( n69553 , n592806 , n66142 );
and ( n596877 , n65493 , n66140 );
nor ( n596878 , n69553 , n596877 );
xnor ( n69556 , n596878 , n592960 );
and ( n596880 , n596874 , n69556 );
and ( n596881 , n69547 , n69556 );
or ( n69559 , n69552 , n596880 , n596881 );
and ( n596883 , n64997 , n594441 );
and ( n69561 , n64973 , n67116 );
nor ( n596885 , n596883 , n69561 );
xnor ( n69563 , n596885 , n66190 );
and ( n596887 , n69559 , n69563 );
and ( n596888 , n592478 , n594210 );
and ( n69566 , n592404 , n66885 );
nor ( n596890 , n596888 , n69566 );
xnor ( n596891 , n596890 , n593434 );
and ( n69569 , n69563 , n596891 );
and ( n596893 , n69559 , n596891 );
or ( n69571 , n596887 , n69569 , n596893 );
and ( n69572 , n596193 , n64559 );
and ( n596896 , n596057 , n591880 );
nor ( n596897 , n69572 , n596896 );
xnor ( n69575 , n596897 , n64521 );
and ( n596899 , n69491 , n64456 );
and ( n69577 , n69283 , n64454 );
nor ( n596901 , n596899 , n69577 );
xnor ( n69579 , n596901 , n591786 );
and ( n69580 , n69575 , n69579 );
buf ( n69581 , n591720 );
and ( n69582 , n69581 , n64451 );
and ( n69583 , n69579 , n69582 );
and ( n69584 , n69575 , n69582 );
or ( n69585 , n69580 , n69583 , n69584 );
and ( n69586 , n596057 , n64559 );
and ( n596910 , n595827 , n591880 );
nor ( n596911 , n69586 , n596910 );
xnor ( n596912 , n596911 , n64521 );
and ( n69590 , n69585 , n596912 );
xor ( n596914 , n596808 , n596812 );
xor ( n69592 , n596914 , n596815 );
and ( n69593 , n596912 , n69592 );
and ( n596917 , n69585 , n69592 );
or ( n596918 , n69590 , n69593 , n596917 );
and ( n69596 , n67940 , n64744 );
and ( n596920 , n595103 , n64742 );
nor ( n596921 , n69596 , n596920 );
xnor ( n69599 , n596921 , n64623 );
and ( n596923 , n596918 , n69599 );
and ( n596924 , n595521 , n64650 );
and ( n69602 , n68160 , n64648 );
nor ( n596926 , n596924 , n69602 );
xnor ( n69604 , n596926 , n591902 );
and ( n596928 , n69599 , n69604 );
and ( n69606 , n596918 , n69604 );
or ( n69607 , n596923 , n596928 , n69606 );
and ( n596931 , n594952 , n64862 );
and ( n596932 , n594710 , n64860 );
nor ( n69610 , n596931 , n596932 );
xnor ( n596934 , n69610 , n64764 );
and ( n596935 , n69607 , n596934 );
xor ( n69613 , n596610 , n596614 );
xor ( n596937 , n69613 , n69303 );
and ( n596938 , n596934 , n596937 );
and ( n69616 , n69607 , n596937 );
or ( n69617 , n596935 , n596938 , n69616 );
and ( n69618 , n66967 , n592340 );
and ( n596942 , n66951 , n65015 );
nor ( n69620 , n69618 , n596942 );
xnor ( n69621 , n69620 , n64847 );
and ( n69622 , n69617 , n69621 );
xor ( n69623 , n69306 , n596633 );
xor ( n69624 , n69623 , n596638 );
and ( n69625 , n69621 , n69624 );
and ( n69626 , n69617 , n69624 );
or ( n596950 , n69622 , n69625 , n69626 );
and ( n69628 , n594124 , n592486 );
and ( n596952 , n66606 , n592484 );
nor ( n596953 , n69628 , n596952 );
xnor ( n69631 , n596953 , n64990 );
and ( n69632 , n596950 , n69631 );
xor ( n69633 , n69318 , n69322 );
xor ( n596957 , n69633 , n69325 );
and ( n69635 , n69631 , n596957 );
and ( n596959 , n596950 , n596957 );
or ( n69637 , n69632 , n69635 , n596959 );
and ( n596961 , n65844 , n593256 );
and ( n69639 , n65630 , n593254 );
nor ( n69640 , n596961 , n69639 );
xnor ( n596964 , n69640 , n65490 );
and ( n596965 , n69637 , n596964 );
xor ( n69643 , n69441 , n596768 );
xor ( n596967 , n69643 , n596771 );
and ( n596968 , n596964 , n596967 );
and ( n69646 , n69637 , n596967 );
or ( n596970 , n596965 , n596968 , n69646 );
xor ( n69648 , n596661 , n596665 );
xor ( n596972 , n69648 , n596670 );
and ( n69650 , n596970 , n596972 );
xor ( n596974 , n596774 , n596776 );
xor ( n596975 , n596974 , n69456 );
and ( n69653 , n596972 , n596975 );
and ( n596977 , n596970 , n596975 );
or ( n69655 , n69650 , n69653 , n596977 );
and ( n596979 , n64854 , n594807 );
and ( n596980 , n64838 , n594804 );
nor ( n69658 , n596979 , n596980 );
xnor ( n69659 , n69658 , n66187 );
and ( n596983 , n69655 , n69659 );
xor ( n69661 , n596569 , n596571 );
xor ( n596985 , n69661 , n596574 );
and ( n69663 , n69659 , n596985 );
and ( n69664 , n69655 , n596985 );
or ( n596988 , n596983 , n69663 , n69664 );
and ( n596989 , n69571 , n596988 );
xor ( n69667 , n69401 , n69405 );
xor ( n596991 , n69667 , n596731 );
and ( n596992 , n596988 , n596991 );
and ( n69670 , n69571 , n596991 );
or ( n596994 , n596989 , n596992 , n69670 );
and ( n596995 , n596804 , n596994 );
xor ( n596996 , n596734 , n69413 );
xor ( n69674 , n596996 , n69416 );
and ( n69675 , n596994 , n69674 );
and ( n596999 , n596804 , n69674 );
or ( n69677 , n596995 , n69675 , n596999 );
xor ( n69678 , n69272 , n69419 );
xor ( n597002 , n69678 , n596745 );
and ( n69680 , n69677 , n597002 );
xor ( n597004 , n596507 , n596531 );
xor ( n69682 , n597004 , n596534 );
and ( n69683 , n597002 , n69682 );
and ( n597007 , n69677 , n69682 );
or ( n597008 , n69680 , n69683 , n597007 );
and ( n69686 , n69437 , n597008 );
xor ( n597010 , n69437 , n597008 );
xor ( n597011 , n69677 , n597002 );
xor ( n69689 , n597011 , n69682 );
and ( n597013 , n66104 , n65592 );
and ( n69691 , n593437 , n592913 );
nor ( n69692 , n597013 , n69691 );
xnor ( n597016 , n69692 , n592638 );
and ( n69694 , n66507 , n592683 );
and ( n597018 , n593520 , n592681 );
nor ( n597019 , n69694 , n597018 );
xnor ( n597020 , n597019 , n592475 );
and ( n69698 , n597016 , n597020 );
xor ( n597022 , n69527 , n596854 );
xor ( n69700 , n597022 , n596857 );
and ( n69701 , n597020 , n69700 );
and ( n69702 , n597016 , n69700 );
or ( n69703 , n69698 , n69701 , n69702 );
and ( n69704 , n65640 , n66142 );
and ( n69705 , n592806 , n66140 );
nor ( n69706 , n69704 , n69705 );
xnor ( n69707 , n69706 , n592960 );
and ( n69708 , n69703 , n69707 );
xor ( n69709 , n596860 , n596864 );
xor ( n69710 , n69709 , n69544 );
and ( n69711 , n69707 , n69710 );
and ( n69712 , n69703 , n69710 );
or ( n69713 , n69708 , n69711 , n69712 );
and ( n69714 , n593520 , n65592 );
and ( n597038 , n66104 , n592913 );
nor ( n69716 , n69714 , n597038 );
xnor ( n597040 , n69716 , n592638 );
and ( n69718 , n66606 , n592683 );
and ( n69719 , n66507 , n592681 );
nor ( n597043 , n69718 , n69719 );
xnor ( n69721 , n597043 , n592475 );
and ( n597045 , n597040 , n69721 );
and ( n69723 , n66793 , n592486 );
and ( n69724 , n594124 , n592484 );
nor ( n597048 , n69723 , n69724 );
xnor ( n69726 , n597048 , n64990 );
and ( n597050 , n69721 , n69726 );
and ( n69728 , n597040 , n69726 );
or ( n597052 , n597045 , n597050 , n69728 );
and ( n69730 , n69283 , n64491 );
and ( n69731 , n596600 , n64489 );
nor ( n597055 , n69730 , n69731 );
xnor ( n597056 , n597055 , n64448 );
and ( n69734 , n69581 , n64456 );
and ( n597058 , n69491 , n64454 );
nor ( n69736 , n69734 , n597058 );
xnor ( n597060 , n69736 , n591786 );
and ( n597061 , n597056 , n597060 );
buf ( n69739 , n591721 );
and ( n597063 , n69739 , n64451 );
and ( n597064 , n597060 , n597063 );
and ( n69742 , n597056 , n597063 );
or ( n597066 , n597061 , n597064 , n69742 );
and ( n597067 , n595827 , n64650 );
and ( n69745 , n595633 , n64648 );
nor ( n597069 , n597067 , n69745 );
xnor ( n69747 , n597069 , n591902 );
and ( n597071 , n597066 , n69747 );
and ( n597072 , n596600 , n64491 );
and ( n69750 , n596198 , n64489 );
nor ( n597074 , n597072 , n69750 );
xnor ( n597075 , n597074 , n64448 );
and ( n69753 , n69747 , n597075 );
and ( n69754 , n597066 , n597075 );
or ( n597078 , n597071 , n69753 , n69754 );
and ( n69756 , n68160 , n64744 );
and ( n597080 , n67940 , n64742 );
nor ( n69758 , n69756 , n597080 );
xnor ( n69759 , n69758 , n64623 );
and ( n69760 , n597078 , n69759 );
and ( n69761 , n595633 , n64650 );
and ( n597085 , n595521 , n64648 );
nor ( n597086 , n69761 , n597085 );
xnor ( n69764 , n597086 , n591902 );
and ( n597088 , n69759 , n69764 );
and ( n597089 , n597078 , n69764 );
or ( n69767 , n69760 , n597088 , n597089 );
and ( n597091 , n67636 , n64862 );
and ( n597092 , n594952 , n64860 );
nor ( n69770 , n597091 , n597092 );
xnor ( n597094 , n69770 , n64764 );
and ( n597095 , n69767 , n597094 );
xor ( n597096 , n596818 , n69499 );
xor ( n69774 , n597096 , n596825 );
and ( n597098 , n597094 , n69774 );
and ( n69776 , n69767 , n69774 );
or ( n597100 , n597095 , n597098 , n69776 );
and ( n597101 , n594295 , n592340 );
and ( n69779 , n66967 , n65015 );
nor ( n597103 , n597101 , n69779 );
xnor ( n597104 , n597103 , n64847 );
and ( n69782 , n597100 , n597104 );
xor ( n597106 , n69505 , n69509 );
xor ( n597107 , n597106 , n69514 );
and ( n69785 , n597104 , n597107 );
and ( n69786 , n597100 , n597107 );
or ( n597110 , n69782 , n69785 , n69786 );
xor ( n69788 , n69617 , n69621 );
xor ( n597112 , n69788 , n69624 );
and ( n69790 , n597110 , n597112 );
xor ( n597114 , n596840 , n596844 );
xor ( n597115 , n597114 , n596847 );
and ( n69793 , n597112 , n597115 );
and ( n597117 , n597110 , n597115 );
or ( n597118 , n69790 , n69793 , n597117 );
and ( n69796 , n597052 , n597118 );
and ( n69797 , n65630 , n66142 );
and ( n597121 , n65640 , n66140 );
nor ( n69799 , n69797 , n597121 );
xnor ( n597123 , n69799 , n592960 );
and ( n69801 , n597118 , n597123 );
and ( n597125 , n597052 , n597123 );
or ( n69803 , n69796 , n69801 , n597125 );
and ( n69804 , n65493 , n66457 );
and ( n597128 , n65384 , n593778 );
nor ( n69806 , n69804 , n597128 );
xnor ( n597130 , n69806 , n593160 );
and ( n69808 , n69803 , n597130 );
xor ( n597132 , n69637 , n596964 );
xor ( n69810 , n597132 , n596967 );
and ( n597134 , n597130 , n69810 );
and ( n597135 , n69803 , n69810 );
or ( n69813 , n69808 , n597134 , n597135 );
and ( n597137 , n69713 , n69813 );
and ( n69815 , n592468 , n594210 );
and ( n69816 , n592478 , n66885 );
nor ( n597140 , n69815 , n69816 );
xnor ( n69818 , n597140 , n593434 );
and ( n597142 , n69813 , n69818 );
and ( n69820 , n69713 , n69818 );
or ( n69821 , n597137 , n597142 , n69820 );
and ( n597145 , n64973 , n594807 );
and ( n597146 , n64854 , n594804 );
nor ( n69824 , n597145 , n597146 );
xnor ( n597148 , n69824 , n66187 );
and ( n597149 , n592404 , n594441 );
and ( n69827 , n64997 , n67116 );
nor ( n597151 , n597149 , n69827 );
xnor ( n597152 , n597151 , n66190 );
and ( n597153 , n597148 , n597152 );
xor ( n69831 , n69547 , n596874 );
xor ( n597155 , n69831 , n69556 );
and ( n597156 , n597152 , n597155 );
and ( n69834 , n597148 , n597155 );
or ( n597158 , n597153 , n597156 , n69834 );
and ( n597159 , n69821 , n597158 );
xor ( n69837 , n69459 , n69463 );
xor ( n597161 , n69837 , n69466 );
and ( n597162 , n597158 , n597161 );
and ( n69840 , n69821 , n597161 );
or ( n69841 , n597159 , n597162 , n69840 );
xor ( n69842 , n69469 , n69473 );
xor ( n69843 , n69842 , n69478 );
and ( n69844 , n69841 , n69843 );
xor ( n597168 , n596577 , n596581 );
xor ( n597169 , n597168 , n596584 );
and ( n69847 , n69843 , n597169 );
and ( n597171 , n69841 , n597169 );
or ( n597172 , n69844 , n69847 , n597171 );
xor ( n69850 , n596587 , n69266 );
xor ( n597174 , n69850 , n69269 );
and ( n597175 , n597172 , n597174 );
xor ( n69853 , n596804 , n596994 );
xor ( n597177 , n69853 , n69674 );
and ( n597178 , n597174 , n597177 );
and ( n69856 , n597172 , n597177 );
or ( n69857 , n597175 , n597178 , n69856 );
and ( n597181 , n69689 , n69857 );
xor ( n69859 , n69689 , n69857 );
xor ( n69860 , n597172 , n597174 );
xor ( n597184 , n69860 , n597177 );
and ( n597185 , n593298 , n593256 );
and ( n69863 , n65844 , n593254 );
nor ( n69864 , n597185 , n69863 );
xnor ( n597188 , n69864 , n65490 );
xor ( n69866 , n596950 , n69631 );
xor ( n597190 , n69866 , n596957 );
and ( n69868 , n597188 , n597190 );
xor ( n597192 , n597016 , n597020 );
xor ( n597193 , n597192 , n69700 );
and ( n69871 , n597190 , n597193 );
and ( n597195 , n597188 , n597193 );
or ( n597196 , n69868 , n69871 , n597195 );
and ( n69874 , n592645 , n594210 );
and ( n597198 , n592468 , n66885 );
nor ( n69876 , n69874 , n597198 );
xnor ( n69877 , n69876 , n593434 );
and ( n69878 , n597196 , n69877 );
xor ( n69879 , n69703 , n69707 );
xor ( n597203 , n69879 , n69710 );
and ( n69881 , n69877 , n597203 );
and ( n69882 , n597196 , n597203 );
or ( n597206 , n69878 , n69881 , n69882 );
xor ( n597207 , n69713 , n69813 );
xor ( n69885 , n597207 , n69818 );
and ( n69886 , n597206 , n69885 );
xor ( n597210 , n596970 , n596972 );
xor ( n597211 , n597210 , n596975 );
and ( n69889 , n69885 , n597211 );
and ( n69890 , n597206 , n597211 );
or ( n597214 , n69886 , n69889 , n69890 );
xor ( n69892 , n69559 , n69563 );
xor ( n597216 , n69892 , n596891 );
and ( n69894 , n597214 , n597216 );
xor ( n69895 , n69655 , n69659 );
xor ( n597219 , n69895 , n596985 );
and ( n597220 , n597216 , n597219 );
and ( n69898 , n597214 , n597219 );
or ( n597222 , n69894 , n597220 , n69898 );
xor ( n69900 , n69571 , n596988 );
xor ( n69901 , n69900 , n596991 );
and ( n69902 , n597222 , n69901 );
xor ( n69903 , n69841 , n69843 );
xor ( n69904 , n69903 , n597169 );
and ( n69905 , n69901 , n69904 );
and ( n597229 , n597222 , n69904 );
or ( n69907 , n69902 , n69905 , n597229 );
and ( n597231 , n597184 , n69907 );
xor ( n597232 , n597184 , n69907 );
xor ( n69910 , n597222 , n69901 );
xor ( n597234 , n69910 , n69904 );
and ( n597235 , n66104 , n593256 );
and ( n69913 , n593437 , n593254 );
nor ( n597237 , n597235 , n69913 );
xnor ( n597238 , n597237 , n65490 );
and ( n69916 , n66507 , n65592 );
and ( n69917 , n593520 , n592913 );
nor ( n597241 , n69916 , n69917 );
xnor ( n69919 , n597241 , n592638 );
and ( n69920 , n597238 , n69919 );
and ( n597244 , n594124 , n592683 );
and ( n597245 , n66606 , n592681 );
nor ( n69923 , n597244 , n597245 );
xnor ( n69924 , n69923 , n592475 );
and ( n597248 , n69919 , n69924 );
and ( n597249 , n597238 , n69924 );
or ( n69927 , n69920 , n597248 , n597249 );
and ( n597251 , n69491 , n64491 );
and ( n597252 , n69283 , n64489 );
nor ( n69930 , n597251 , n597252 );
xnor ( n597254 , n69930 , n64448 );
and ( n69932 , n69739 , n64456 );
and ( n597256 , n69581 , n64454 );
nor ( n69934 , n69932 , n597256 );
xnor ( n597258 , n69934 , n591786 );
and ( n69936 , n597254 , n597258 );
buf ( n597260 , n591722 );
and ( n597261 , n597260 , n64451 );
and ( n69939 , n597258 , n597261 );
and ( n69940 , n597254 , n597261 );
or ( n597264 , n69936 , n69939 , n69940 );
and ( n597265 , n596198 , n64559 );
and ( n69943 , n596193 , n591880 );
nor ( n597267 , n597265 , n69943 );
xnor ( n597268 , n597267 , n64521 );
and ( n69946 , n597264 , n597268 );
xor ( n597270 , n597056 , n597060 );
xor ( n597271 , n597270 , n597063 );
and ( n597272 , n597268 , n597271 );
and ( n69950 , n597264 , n597271 );
or ( n597274 , n69946 , n597272 , n69950 );
and ( n597275 , n595521 , n64744 );
and ( n69953 , n68160 , n64742 );
nor ( n597277 , n597275 , n69953 );
xnor ( n597278 , n597277 , n64623 );
and ( n69956 , n597274 , n597278 );
xor ( n597280 , n69575 , n69579 );
xor ( n597281 , n597280 , n69582 );
and ( n69959 , n597278 , n597281 );
and ( n597283 , n597274 , n597281 );
or ( n69961 , n69956 , n69959 , n597283 );
and ( n69962 , n595103 , n64862 );
and ( n597286 , n67636 , n64860 );
nor ( n69964 , n69962 , n597286 );
xnor ( n69965 , n69964 , n64764 );
and ( n69966 , n69961 , n69965 );
xor ( n69967 , n69585 , n596912 );
xor ( n69968 , n69967 , n69592 );
and ( n597292 , n69965 , n69968 );
and ( n597293 , n69961 , n69968 );
or ( n597294 , n69966 , n597292 , n597293 );
and ( n597295 , n594710 , n592340 );
and ( n69973 , n594295 , n65015 );
nor ( n597297 , n597295 , n69973 );
xnor ( n597298 , n597297 , n64847 );
and ( n597299 , n597294 , n597298 );
xor ( n69977 , n596918 , n69599 );
xor ( n597301 , n69977 , n69604 );
and ( n69979 , n597298 , n597301 );
and ( n597303 , n597294 , n597301 );
or ( n69981 , n597299 , n69979 , n597303 );
and ( n597305 , n66951 , n592486 );
and ( n597306 , n66793 , n592484 );
nor ( n69984 , n597305 , n597306 );
xnor ( n69985 , n69984 , n64990 );
and ( n597309 , n69981 , n69985 );
xor ( n597310 , n69607 , n596934 );
xor ( n69988 , n597310 , n596937 );
and ( n597312 , n69985 , n69988 );
and ( n597313 , n69981 , n69988 );
or ( n69991 , n597309 , n597312 , n597313 );
and ( n597315 , n69927 , n69991 );
and ( n597316 , n593437 , n593256 );
and ( n69994 , n593298 , n593254 );
nor ( n69995 , n597316 , n69994 );
xnor ( n597319 , n69995 , n65490 );
and ( n597320 , n69991 , n597319 );
and ( n69998 , n69927 , n597319 );
or ( n597322 , n597315 , n597320 , n69998 );
and ( n597323 , n592806 , n66457 );
and ( n70001 , n65493 , n593778 );
nor ( n597325 , n597323 , n70001 );
xnor ( n597326 , n597325 , n593160 );
and ( n70004 , n597322 , n597326 );
xor ( n597328 , n597052 , n597118 );
xor ( n70006 , n597328 , n597123 );
and ( n597330 , n597326 , n70006 );
and ( n70008 , n597322 , n70006 );
or ( n597332 , n70004 , n597330 , n70008 );
and ( n70010 , n65640 , n66457 );
and ( n70011 , n592806 , n593778 );
nor ( n597335 , n70010 , n70011 );
xnor ( n597336 , n597335 , n593160 );
and ( n70014 , n65844 , n66142 );
and ( n597338 , n65630 , n66140 );
nor ( n597339 , n70014 , n597338 );
xnor ( n70017 , n597339 , n592960 );
and ( n597341 , n597336 , n70017 );
xor ( n597342 , n597040 , n69721 );
xor ( n70020 , n597342 , n69726 );
and ( n70021 , n70017 , n70020 );
and ( n597345 , n597336 , n70020 );
or ( n597346 , n597341 , n70021 , n597345 );
and ( n70024 , n65384 , n594210 );
and ( n597348 , n592645 , n66885 );
nor ( n597349 , n70024 , n597348 );
xnor ( n70027 , n597349 , n593434 );
and ( n597351 , n597346 , n70027 );
xor ( n597352 , n597188 , n597190 );
xor ( n70030 , n597352 , n597193 );
and ( n597354 , n70027 , n70030 );
and ( n597355 , n597346 , n70030 );
or ( n70033 , n597351 , n597354 , n597355 );
and ( n597357 , n597332 , n70033 );
and ( n70035 , n592478 , n594441 );
and ( n597359 , n592404 , n67116 );
nor ( n597360 , n70035 , n597359 );
xnor ( n597361 , n597360 , n66190 );
and ( n70039 , n70033 , n597361 );
and ( n597363 , n597332 , n597361 );
or ( n70041 , n597357 , n70039 , n597363 );
and ( n597365 , n64997 , n594807 );
and ( n597366 , n64973 , n594804 );
nor ( n597367 , n597365 , n597366 );
xnor ( n597368 , n597367 , n66187 );
xor ( n70046 , n69803 , n597130 );
xor ( n597370 , n70046 , n69810 );
and ( n597371 , n597368 , n597370 );
xor ( n70049 , n597196 , n69877 );
xor ( n597373 , n70049 , n597203 );
and ( n597374 , n597370 , n597373 );
and ( n70052 , n597368 , n597373 );
or ( n597376 , n597371 , n597374 , n70052 );
and ( n597377 , n70041 , n597376 );
xor ( n70055 , n597148 , n597152 );
xor ( n597379 , n70055 , n597155 );
and ( n597380 , n597376 , n597379 );
and ( n70058 , n70041 , n597379 );
or ( n70059 , n597377 , n597380 , n70058 );
xor ( n70060 , n69821 , n597158 );
xor ( n597384 , n70060 , n597161 );
and ( n597385 , n70059 , n597384 );
xor ( n70063 , n597214 , n597216 );
xor ( n70064 , n70063 , n597219 );
and ( n597388 , n597384 , n70064 );
and ( n70066 , n70059 , n70064 );
or ( n597390 , n597385 , n597388 , n70066 );
and ( n70068 , n597234 , n597390 );
xor ( n70069 , n597234 , n597390 );
and ( n70070 , n69581 , n64491 );
and ( n597394 , n69491 , n64489 );
nor ( n70072 , n70070 , n597394 );
xnor ( n597396 , n70072 , n64448 );
and ( n70074 , n597260 , n64456 );
and ( n597398 , n69739 , n64454 );
nor ( n70076 , n70074 , n597398 );
xnor ( n70077 , n70076 , n591786 );
and ( n70078 , n597396 , n70077 );
buf ( n597402 , n591723 );
and ( n597403 , n597402 , n64451 );
and ( n70081 , n70077 , n597403 );
and ( n70082 , n597396 , n597403 );
or ( n70083 , n70078 , n70081 , n70082 );
and ( n597407 , n596193 , n64650 );
and ( n597408 , n596057 , n64648 );
nor ( n70086 , n597407 , n597408 );
xnor ( n597410 , n70086 , n591902 );
and ( n597411 , n70083 , n597410 );
xor ( n70089 , n597254 , n597258 );
xor ( n597413 , n70089 , n597261 );
and ( n597414 , n597410 , n597413 );
and ( n70092 , n70083 , n597413 );
or ( n597416 , n597411 , n597414 , n70092 );
and ( n597417 , n595633 , n64744 );
and ( n70095 , n595521 , n64742 );
nor ( n70096 , n597417 , n70095 );
xnor ( n597420 , n70096 , n64623 );
and ( n597421 , n597416 , n597420 );
and ( n597422 , n596057 , n64650 );
and ( n70100 , n595827 , n64648 );
nor ( n597424 , n597422 , n70100 );
xnor ( n70102 , n597424 , n591902 );
and ( n597426 , n597420 , n70102 );
and ( n70104 , n597416 , n70102 );
or ( n70105 , n597421 , n597426 , n70104 );
and ( n597429 , n67940 , n64862 );
and ( n597430 , n595103 , n64860 );
nor ( n70108 , n597429 , n597430 );
xnor ( n597432 , n70108 , n64764 );
and ( n597433 , n70105 , n597432 );
xor ( n70111 , n597066 , n69747 );
xor ( n597435 , n70111 , n597075 );
and ( n597436 , n597432 , n597435 );
and ( n70114 , n70105 , n597435 );
or ( n70115 , n597433 , n597436 , n70114 );
and ( n597439 , n594952 , n592340 );
and ( n597440 , n594710 , n65015 );
nor ( n70118 , n597439 , n597440 );
xnor ( n597442 , n70118 , n64847 );
and ( n597443 , n70115 , n597442 );
xor ( n70121 , n597078 , n69759 );
xor ( n597445 , n70121 , n69764 );
and ( n597446 , n597442 , n597445 );
and ( n70124 , n70115 , n597445 );
or ( n70125 , n597443 , n597446 , n70124 );
and ( n70126 , n66967 , n592486 );
and ( n597450 , n66951 , n592484 );
nor ( n70128 , n70126 , n597450 );
xnor ( n597452 , n70128 , n64990 );
and ( n70130 , n70125 , n597452 );
xor ( n70131 , n69767 , n597094 );
xor ( n70132 , n70131 , n69774 );
and ( n597456 , n597452 , n70132 );
and ( n70134 , n70125 , n70132 );
or ( n597458 , n70130 , n597456 , n70134 );
xor ( n597459 , n597100 , n597104 );
xor ( n597460 , n597459 , n597107 );
and ( n70138 , n597458 , n597460 );
xor ( n597462 , n69981 , n69985 );
xor ( n597463 , n597462 , n69988 );
and ( n70141 , n597460 , n597463 );
and ( n597465 , n597458 , n597463 );
or ( n597466 , n70138 , n70141 , n597465 );
xor ( n597467 , n69927 , n69991 );
xor ( n70145 , n597467 , n597319 );
and ( n597469 , n597466 , n70145 );
xor ( n70147 , n597110 , n597112 );
xor ( n70148 , n70147 , n597115 );
and ( n70149 , n70145 , n70148 );
and ( n70150 , n597466 , n70148 );
or ( n70151 , n597469 , n70149 , n70150 );
and ( n70152 , n592468 , n594441 );
and ( n70153 , n592478 , n67116 );
nor ( n70154 , n70152 , n70153 );
xnor ( n70155 , n70154 , n66190 );
and ( n597479 , n70151 , n70155 );
xor ( n597480 , n597322 , n597326 );
xor ( n70158 , n597480 , n70006 );
and ( n597482 , n70155 , n70158 );
and ( n70160 , n70151 , n70158 );
or ( n70161 , n597479 , n597482 , n70160 );
and ( n597485 , n593520 , n593256 );
and ( n70163 , n66104 , n593254 );
nor ( n597487 , n597485 , n70163 );
xnor ( n70165 , n597487 , n65490 );
and ( n597489 , n66793 , n592683 );
and ( n70167 , n594124 , n592681 );
nor ( n597491 , n597489 , n70167 );
xnor ( n597492 , n597491 , n592475 );
and ( n70170 , n70165 , n597492 );
xor ( n70171 , n597294 , n597298 );
xor ( n597495 , n70171 , n597301 );
and ( n597496 , n597492 , n597495 );
and ( n70174 , n70165 , n597495 );
or ( n597498 , n70170 , n597496 , n70174 );
and ( n597499 , n65630 , n66457 );
and ( n70177 , n65640 , n593778 );
nor ( n597501 , n597499 , n70177 );
xnor ( n597502 , n597501 , n593160 );
and ( n70180 , n597498 , n597502 );
and ( n70181 , n593298 , n66142 );
and ( n597505 , n65844 , n66140 );
nor ( n597506 , n70181 , n597505 );
xnor ( n70184 , n597506 , n592960 );
and ( n597508 , n597502 , n70184 );
and ( n597509 , n597498 , n70184 );
or ( n70187 , n70180 , n597508 , n597509 );
and ( n597511 , n65493 , n594210 );
and ( n597512 , n65384 , n66885 );
nor ( n70190 , n597511 , n597512 );
xnor ( n597514 , n70190 , n593434 );
and ( n70192 , n70187 , n597514 );
xor ( n597516 , n597336 , n70017 );
xor ( n597517 , n597516 , n70020 );
and ( n70195 , n597514 , n597517 );
and ( n70196 , n70187 , n597517 );
or ( n597520 , n70192 , n70195 , n70196 );
and ( n70198 , n592404 , n594807 );
and ( n70199 , n64997 , n594804 );
nor ( n597523 , n70198 , n70199 );
xnor ( n597524 , n597523 , n66187 );
and ( n70202 , n597520 , n597524 );
xor ( n597526 , n597346 , n70027 );
xor ( n597527 , n597526 , n70030 );
and ( n70205 , n597524 , n597527 );
and ( n70206 , n597520 , n597527 );
or ( n70207 , n70202 , n70205 , n70206 );
and ( n597531 , n70161 , n70207 );
xor ( n597532 , n597368 , n597370 );
xor ( n70210 , n597532 , n597373 );
and ( n597534 , n70207 , n70210 );
and ( n597535 , n70161 , n70210 );
or ( n70213 , n597531 , n597534 , n597535 );
xor ( n597537 , n70041 , n597376 );
xor ( n597538 , n597537 , n597379 );
and ( n70216 , n70213 , n597538 );
xor ( n70217 , n597206 , n69885 );
xor ( n597541 , n70217 , n597211 );
and ( n597542 , n597538 , n597541 );
and ( n70220 , n70213 , n597541 );
or ( n597544 , n70216 , n597542 , n70220 );
xor ( n597545 , n70059 , n597384 );
xor ( n70223 , n597545 , n70064 );
and ( n597547 , n597544 , n70223 );
xor ( n70225 , n597544 , n70223 );
xor ( n597549 , n70213 , n597538 );
xor ( n70227 , n597549 , n597541 );
and ( n597551 , n596198 , n64650 );
and ( n70229 , n596193 , n64648 );
nor ( n597553 , n597551 , n70229 );
xnor ( n70231 , n597553 , n591902 );
and ( n70232 , n69283 , n64559 );
and ( n597556 , n596600 , n591880 );
nor ( n597557 , n70232 , n597556 );
xnor ( n70235 , n597557 , n64521 );
and ( n597559 , n70231 , n70235 );
and ( n597560 , n69739 , n64491 );
and ( n70238 , n69581 , n64489 );
nor ( n597562 , n597560 , n70238 );
xnor ( n597563 , n597562 , n64448 );
and ( n70241 , n597402 , n64456 );
and ( n70242 , n597260 , n64454 );
nor ( n597566 , n70241 , n70242 );
xnor ( n597567 , n597566 , n591786 );
and ( n70245 , n597563 , n597567 );
buf ( n597569 , n591724 );
and ( n597570 , n597569 , n64451 );
and ( n70248 , n597567 , n597570 );
and ( n597572 , n597563 , n597570 );
or ( n70250 , n70245 , n70248 , n597572 );
and ( n70251 , n597402 , n64491 );
and ( n70252 , n597260 , n64489 );
nor ( n70253 , n70251 , n70252 );
xnor ( n70254 , n70253 , n64448 );
buf ( n70255 , n591725 );
and ( n597579 , n70255 , n64456 );
and ( n70257 , n597569 , n64454 );
nor ( n70258 , n597579 , n70257 );
xnor ( n70259 , n70258 , n591786 );
and ( n70260 , n70254 , n70259 );
buf ( n70261 , n591726 );
and ( n70262 , n70261 , n64451 );
and ( n70263 , n70259 , n70262 );
and ( n597587 , n70254 , n70262 );
or ( n597588 , n70260 , n70263 , n597587 );
and ( n70266 , n597569 , n64456 );
and ( n597590 , n597402 , n64454 );
nor ( n70268 , n70266 , n597590 );
xnor ( n70269 , n70268 , n591786 );
and ( n597593 , n597588 , n70269 );
and ( n70271 , n70255 , n64451 );
and ( n597595 , n70269 , n70271 );
and ( n70273 , n597588 , n70271 );
or ( n597597 , n597593 , n597595 , n70273 );
and ( n597598 , n69491 , n64559 );
and ( n70276 , n69283 , n591880 );
nor ( n70277 , n597598 , n70276 );
xnor ( n597601 , n70277 , n64521 );
and ( n597602 , n597597 , n597601 );
xor ( n70280 , n597563 , n597567 );
xor ( n597604 , n70280 , n597570 );
and ( n597605 , n597601 , n597604 );
and ( n70283 , n597597 , n597604 );
or ( n597607 , n597602 , n597605 , n70283 );
xor ( n597608 , n70250 , n597607 );
xor ( n597609 , n597396 , n70077 );
xor ( n70287 , n597609 , n597403 );
xor ( n597611 , n597608 , n70287 );
and ( n597612 , n70235 , n597611 );
and ( n70290 , n70231 , n597611 );
or ( n597614 , n597559 , n597612 , n70290 );
and ( n597615 , n595521 , n64862 );
and ( n70293 , n68160 , n64860 );
nor ( n597617 , n597615 , n70293 );
xnor ( n70295 , n597617 , n64764 );
and ( n597619 , n597614 , n70295 );
xor ( n70297 , n70083 , n597410 );
xor ( n70298 , n70297 , n597413 );
and ( n597622 , n70295 , n70298 );
and ( n70300 , n597614 , n70298 );
or ( n597624 , n597619 , n597622 , n70300 );
and ( n70302 , n595103 , n592340 );
and ( n70303 , n67636 , n65015 );
nor ( n597627 , n70302 , n70303 );
xnor ( n70305 , n597627 , n64847 );
and ( n597629 , n597624 , n70305 );
xor ( n70307 , n597416 , n597420 );
xor ( n597631 , n70307 , n70102 );
and ( n597632 , n70305 , n597631 );
and ( n70310 , n597624 , n597631 );
or ( n597634 , n597629 , n597632 , n70310 );
and ( n597635 , n594710 , n592486 );
and ( n597636 , n594295 , n592484 );
nor ( n70314 , n597635 , n597636 );
xnor ( n597638 , n70314 , n64990 );
and ( n597639 , n597634 , n597638 );
xor ( n70317 , n70105 , n597432 );
xor ( n597641 , n70317 , n597435 );
and ( n597642 , n597638 , n597641 );
and ( n70320 , n597634 , n597641 );
or ( n70321 , n597639 , n597642 , n70320 );
and ( n70322 , n66951 , n592683 );
and ( n597646 , n66793 , n592681 );
nor ( n597647 , n70322 , n597646 );
xnor ( n70325 , n597647 , n592475 );
and ( n70326 , n70321 , n70325 );
xor ( n70327 , n70115 , n597442 );
xor ( n597651 , n70327 , n597445 );
and ( n597652 , n70325 , n597651 );
and ( n70330 , n70321 , n597651 );
or ( n70331 , n70326 , n597652 , n70330 );
and ( n597655 , n69581 , n64559 );
and ( n597656 , n69491 , n591880 );
nor ( n70334 , n597655 , n597656 );
xnor ( n70335 , n70334 , n64521 );
and ( n70336 , n597260 , n64491 );
and ( n597660 , n69739 , n64489 );
nor ( n70338 , n70336 , n597660 );
xnor ( n597662 , n70338 , n64448 );
and ( n70340 , n70335 , n597662 );
xor ( n597664 , n597588 , n70269 );
xor ( n70342 , n597664 , n70271 );
and ( n70343 , n597662 , n70342 );
and ( n70344 , n70335 , n70342 );
or ( n597668 , n70340 , n70343 , n70344 );
and ( n70346 , n596600 , n64650 );
and ( n597670 , n596198 , n64648 );
nor ( n70348 , n70346 , n597670 );
xnor ( n70349 , n70348 , n591902 );
and ( n597673 , n597668 , n70349 );
xor ( n70351 , n597597 , n597601 );
xor ( n597675 , n70351 , n597604 );
and ( n597676 , n70349 , n597675 );
and ( n70354 , n597668 , n597675 );
or ( n597678 , n597673 , n597676 , n70354 );
and ( n70356 , n595633 , n64862 );
and ( n597680 , n595521 , n64860 );
nor ( n597681 , n70356 , n597680 );
xnor ( n70359 , n597681 , n64764 );
and ( n597683 , n597678 , n70359 );
and ( n70361 , n596057 , n64744 );
and ( n70362 , n595827 , n64742 );
nor ( n70363 , n70361 , n70362 );
xnor ( n70364 , n70363 , n64623 );
and ( n70365 , n70359 , n70364 );
and ( n597689 , n597678 , n70364 );
or ( n597690 , n597683 , n70365 , n597689 );
and ( n70368 , n67940 , n592340 );
and ( n70369 , n595103 , n65015 );
nor ( n597693 , n70368 , n70369 );
xnor ( n70371 , n597693 , n64847 );
and ( n70372 , n597690 , n70371 );
and ( n597696 , n70250 , n597607 );
and ( n70374 , n597607 , n70287 );
and ( n70375 , n70250 , n70287 );
or ( n597699 , n597696 , n70374 , n70375 );
and ( n597700 , n595827 , n64744 );
and ( n70378 , n595633 , n64742 );
nor ( n597702 , n597700 , n70378 );
xnor ( n70380 , n597702 , n64623 );
xor ( n70381 , n597699 , n70380 );
and ( n70382 , n596600 , n64559 );
and ( n70383 , n596198 , n591880 );
nor ( n597707 , n70382 , n70383 );
xnor ( n597708 , n597707 , n64521 );
xor ( n70386 , n70381 , n597708 );
and ( n597710 , n70371 , n70386 );
and ( n597711 , n597690 , n70386 );
or ( n70389 , n70372 , n597710 , n597711 );
and ( n597713 , n594952 , n592486 );
and ( n597714 , n594710 , n592484 );
nor ( n70392 , n597713 , n597714 );
xnor ( n70393 , n70392 , n64990 );
and ( n597717 , n70389 , n70393 );
and ( n597718 , n597699 , n70380 );
and ( n597719 , n70380 , n597708 );
and ( n597720 , n597699 , n597708 );
or ( n70398 , n597718 , n597719 , n597720 );
and ( n597722 , n68160 , n64862 );
and ( n597723 , n67940 , n64860 );
nor ( n70401 , n597722 , n597723 );
xnor ( n597725 , n70401 , n64764 );
xor ( n597726 , n70398 , n597725 );
xor ( n597727 , n597264 , n597268 );
xor ( n70405 , n597727 , n597271 );
xor ( n597729 , n597726 , n70405 );
and ( n597730 , n70393 , n597729 );
and ( n70408 , n70389 , n597729 );
or ( n597732 , n597717 , n597730 , n70408 );
and ( n70410 , n66967 , n592683 );
and ( n597734 , n66951 , n592681 );
nor ( n597735 , n70410 , n597734 );
xnor ( n597736 , n597735 , n592475 );
and ( n597737 , n597732 , n597736 );
and ( n597738 , n70398 , n597725 );
and ( n70416 , n597725 , n70405 );
and ( n597740 , n70398 , n70405 );
or ( n70418 , n597738 , n70416 , n597740 );
and ( n70419 , n67636 , n592340 );
and ( n70420 , n594952 , n65015 );
nor ( n70421 , n70419 , n70420 );
xnor ( n70422 , n70421 , n64847 );
xor ( n70423 , n70418 , n70422 );
xor ( n70424 , n597274 , n597278 );
xor ( n597748 , n70424 , n597281 );
xor ( n70426 , n70423 , n597748 );
and ( n597750 , n597736 , n70426 );
and ( n597751 , n597732 , n70426 );
or ( n70429 , n597737 , n597750 , n597751 );
and ( n597753 , n66104 , n66142 );
and ( n597754 , n593437 , n66140 );
nor ( n70432 , n597753 , n597754 );
xnor ( n597756 , n70432 , n592960 );
and ( n597757 , n70429 , n597756 );
and ( n597758 , n70418 , n70422 );
and ( n70436 , n70422 , n597748 );
and ( n597760 , n70418 , n597748 );
or ( n597761 , n597758 , n70436 , n597760 );
and ( n70439 , n594295 , n592486 );
and ( n597763 , n66967 , n592484 );
nor ( n597764 , n70439 , n597763 );
xnor ( n70442 , n597764 , n64990 );
xor ( n597766 , n597761 , n70442 );
xor ( n70444 , n69961 , n69965 );
xor ( n70445 , n70444 , n69968 );
xor ( n70446 , n597766 , n70445 );
and ( n70447 , n597756 , n70446 );
and ( n70448 , n70429 , n70446 );
or ( n70449 , n597757 , n70447 , n70448 );
and ( n70450 , n70331 , n70449 );
and ( n70451 , n593437 , n66142 );
and ( n70452 , n593298 , n66140 );
nor ( n70453 , n70451 , n70452 );
xnor ( n597777 , n70453 , n592960 );
and ( n70455 , n70449 , n597777 );
and ( n597779 , n70331 , n597777 );
or ( n597780 , n70450 , n70455 , n597779 );
and ( n70458 , n65640 , n594210 );
and ( n597782 , n592806 , n66885 );
nor ( n597783 , n70458 , n597782 );
xnor ( n70461 , n597783 , n593434 );
and ( n597785 , n65844 , n66457 );
and ( n597786 , n65630 , n593778 );
nor ( n70464 , n597785 , n597786 );
xnor ( n70465 , n70464 , n593160 );
and ( n70466 , n70461 , n70465 );
and ( n597790 , n597761 , n70442 );
and ( n70468 , n70442 , n70445 );
and ( n597792 , n597761 , n70445 );
or ( n70470 , n597790 , n70468 , n597792 );
and ( n597794 , n66606 , n65592 );
and ( n70472 , n66507 , n592913 );
nor ( n70473 , n597794 , n70472 );
xnor ( n597797 , n70473 , n592638 );
xor ( n70475 , n70470 , n597797 );
xor ( n597799 , n70125 , n597452 );
xor ( n70477 , n597799 , n70132 );
xor ( n597801 , n70475 , n70477 );
and ( n597802 , n70465 , n597801 );
and ( n70480 , n70461 , n597801 );
or ( n70481 , n70466 , n597802 , n70480 );
and ( n597805 , n597780 , n70481 );
and ( n597806 , n592806 , n594210 );
and ( n70484 , n65493 , n66885 );
nor ( n597808 , n597806 , n70484 );
xnor ( n597809 , n597808 , n593434 );
and ( n70487 , n70481 , n597809 );
and ( n597811 , n597780 , n597809 );
or ( n597812 , n597805 , n70487 , n597811 );
and ( n597813 , n65384 , n594441 );
and ( n70491 , n592645 , n67116 );
nor ( n597815 , n597813 , n70491 );
xnor ( n597816 , n597815 , n66190 );
xor ( n70494 , n597498 , n597502 );
xor ( n597818 , n70494 , n70184 );
and ( n70496 , n597816 , n597818 );
and ( n70497 , n70470 , n597797 );
and ( n70498 , n597797 , n70477 );
and ( n70499 , n70470 , n70477 );
or ( n70500 , n70497 , n70498 , n70499 );
xor ( n70501 , n597238 , n69919 );
xor ( n597825 , n70501 , n69924 );
xor ( n70503 , n70500 , n597825 );
xor ( n597827 , n597458 , n597460 );
xor ( n70505 , n597827 , n597463 );
xor ( n597829 , n70503 , n70505 );
and ( n70507 , n597818 , n597829 );
and ( n70508 , n597816 , n597829 );
or ( n597832 , n70496 , n70507 , n70508 );
and ( n70510 , n597812 , n597832 );
xor ( n597834 , n70187 , n597514 );
xor ( n70512 , n597834 , n597517 );
and ( n597836 , n597832 , n70512 );
and ( n597837 , n597812 , n70512 );
or ( n70515 , n70510 , n597836 , n597837 );
and ( n597839 , n70500 , n597825 );
and ( n597840 , n597825 , n70505 );
and ( n70518 , n70500 , n70505 );
or ( n70519 , n597839 , n597840 , n70518 );
and ( n597843 , n592645 , n594441 );
and ( n597844 , n592468 , n67116 );
nor ( n70522 , n597843 , n597844 );
xnor ( n597846 , n70522 , n66190 );
and ( n597847 , n70519 , n597846 );
xor ( n70525 , n597466 , n70145 );
xor ( n597849 , n70525 , n70148 );
and ( n597850 , n597846 , n597849 );
and ( n70528 , n70519 , n597849 );
or ( n70529 , n597847 , n597850 , n70528 );
and ( n597853 , n70515 , n70529 );
xor ( n70531 , n70151 , n70155 );
xor ( n597855 , n70531 , n70158 );
and ( n70533 , n70529 , n597855 );
and ( n597857 , n70515 , n597855 );
or ( n70535 , n597853 , n70533 , n597857 );
xor ( n70536 , n597332 , n70033 );
xor ( n597860 , n70536 , n597361 );
and ( n70538 , n70535 , n597860 );
xor ( n597862 , n70161 , n70207 );
xor ( n70540 , n597862 , n70210 );
and ( n597864 , n597860 , n70540 );
and ( n597865 , n70535 , n70540 );
or ( n70543 , n70538 , n597864 , n597865 );
and ( n70544 , n70227 , n70543 );
xor ( n597868 , n70227 , n70543 );
xor ( n70546 , n70535 , n597860 );
xor ( n597870 , n70546 , n70540 );
and ( n70548 , n66507 , n593256 );
and ( n597872 , n593520 , n593254 );
nor ( n597873 , n70548 , n597872 );
xnor ( n70551 , n597873 , n65490 );
and ( n597875 , n594124 , n65592 );
and ( n597876 , n66606 , n592913 );
nor ( n597877 , n597875 , n597876 );
xnor ( n70555 , n597877 , n592638 );
and ( n597879 , n70551 , n70555 );
xor ( n597880 , n70321 , n70325 );
xor ( n70558 , n597880 , n597651 );
and ( n597882 , n70555 , n70558 );
and ( n597883 , n70551 , n70558 );
or ( n70561 , n597879 , n597882 , n597883 );
xor ( n70562 , n70331 , n70449 );
xor ( n70563 , n70562 , n597777 );
and ( n597887 , n70561 , n70563 );
xor ( n70565 , n70165 , n597492 );
xor ( n70566 , n70565 , n597495 );
and ( n70567 , n70563 , n70566 );
and ( n597891 , n70561 , n70566 );
or ( n70569 , n597887 , n70567 , n597891 );
and ( n70570 , n592468 , n594807 );
and ( n70571 , n592478 , n594804 );
nor ( n597895 , n70570 , n70571 );
xnor ( n597896 , n597895 , n66187 );
and ( n597897 , n70569 , n597896 );
xor ( n70575 , n597780 , n70481 );
xor ( n597899 , n70575 , n597809 );
and ( n597900 , n597896 , n597899 );
and ( n70578 , n70569 , n597899 );
or ( n70579 , n597897 , n597900 , n70578 );
and ( n70580 , n592478 , n594807 );
and ( n70581 , n592404 , n594804 );
nor ( n70582 , n70580 , n70581 );
xnor ( n70583 , n70582 , n66187 );
and ( n597907 , n70579 , n70583 );
xor ( n70585 , n70519 , n597846 );
xor ( n70586 , n70585 , n597849 );
and ( n597910 , n70583 , n70586 );
and ( n597911 , n70579 , n70586 );
or ( n70589 , n597907 , n597910 , n597911 );
xor ( n70590 , n70515 , n70529 );
xor ( n597914 , n70590 , n597855 );
and ( n597915 , n70589 , n597914 );
xor ( n70593 , n597520 , n597524 );
xor ( n70594 , n70593 , n597527 );
and ( n70595 , n597914 , n70594 );
and ( n597919 , n70589 , n70594 );
or ( n70597 , n597915 , n70595 , n597919 );
and ( n70598 , n597870 , n70597 );
xor ( n70599 , n597870 , n70597 );
xor ( n70600 , n70589 , n597914 );
xor ( n597924 , n70600 , n70594 );
and ( n70602 , n593520 , n66142 );
and ( n597926 , n66104 , n66140 );
nor ( n70604 , n70602 , n597926 );
xnor ( n70605 , n70604 , n592960 );
and ( n597929 , n66606 , n593256 );
and ( n597930 , n66507 , n593254 );
nor ( n70608 , n597929 , n597930 );
xnor ( n597932 , n70608 , n65490 );
and ( n597933 , n70605 , n597932 );
xor ( n70611 , n597634 , n597638 );
xor ( n597935 , n70611 , n597641 );
and ( n70613 , n597932 , n597935 );
and ( n70614 , n70605 , n597935 );
or ( n70615 , n597933 , n70613 , n70614 );
and ( n70616 , n65630 , n594210 );
and ( n70617 , n65640 , n66885 );
nor ( n70618 , n70616 , n70617 );
xnor ( n70619 , n70618 , n593434 );
and ( n70620 , n70615 , n70619 );
and ( n597944 , n593298 , n66457 );
and ( n70622 , n65844 , n593778 );
nor ( n597946 , n597944 , n70622 );
xnor ( n70624 , n597946 , n593160 );
and ( n70625 , n70619 , n70624 );
and ( n597949 , n70615 , n70624 );
or ( n597950 , n70620 , n70625 , n597949 );
and ( n70628 , n597569 , n64491 );
and ( n70629 , n597402 , n64489 );
nor ( n597953 , n70628 , n70629 );
xnor ( n70631 , n597953 , n64448 );
and ( n597955 , n70261 , n64456 );
and ( n70633 , n70255 , n64454 );
nor ( n597957 , n597955 , n70633 );
xnor ( n70635 , n597957 , n591786 );
and ( n70636 , n70631 , n70635 );
buf ( n70637 , n591727 );
and ( n70638 , n70637 , n64451 );
and ( n70639 , n70635 , n70638 );
and ( n70640 , n70631 , n70638 );
or ( n597964 , n70636 , n70639 , n70640 );
and ( n70642 , n69739 , n64559 );
and ( n597966 , n69581 , n591880 );
nor ( n70644 , n70642 , n597966 );
xnor ( n70645 , n70644 , n64521 );
and ( n70646 , n597964 , n70645 );
xor ( n70647 , n70254 , n70259 );
xor ( n70648 , n70647 , n70262 );
and ( n70649 , n70645 , n70648 );
and ( n597973 , n597964 , n70648 );
or ( n70651 , n70646 , n70649 , n597973 );
buf ( n70652 , n591733 );
and ( n70653 , n70652 , n64454 );
not ( n597977 , n70653 );
and ( n597978 , n597977 , n591786 );
and ( n70656 , n70652 , n64456 );
buf ( n597980 , n591732 );
and ( n70658 , n597980 , n64454 );
nor ( n597982 , n70656 , n70658 );
xnor ( n70660 , n597982 , n591786 );
and ( n597984 , n597978 , n70660 );
and ( n70662 , n597980 , n64456 );
buf ( n70663 , n591731 );
and ( n597987 , n70663 , n64454 );
nor ( n597988 , n70662 , n597987 );
xnor ( n70666 , n597988 , n591786 );
and ( n70667 , n597984 , n70666 );
and ( n597991 , n70652 , n64451 );
and ( n597992 , n70666 , n597991 );
and ( n70670 , n597984 , n597991 );
or ( n70671 , n70667 , n597992 , n70670 );
and ( n597995 , n70663 , n64456 );
buf ( n597996 , n591730 );
and ( n70674 , n597996 , n64454 );
nor ( n70675 , n597995 , n70674 );
xnor ( n597999 , n70675 , n591786 );
and ( n598000 , n70671 , n597999 );
and ( n70678 , n597980 , n64451 );
and ( n70679 , n597999 , n70678 );
and ( n70680 , n70671 , n70678 );
or ( n598004 , n598000 , n70679 , n70680 );
and ( n598005 , n597996 , n64456 );
buf ( n70683 , n591729 );
and ( n598007 , n70683 , n64454 );
nor ( n598008 , n598005 , n598007 );
xnor ( n70686 , n598008 , n591786 );
and ( n598010 , n598004 , n70686 );
and ( n70688 , n70663 , n64451 );
and ( n70689 , n70686 , n70688 );
and ( n70690 , n598004 , n70688 );
or ( n598014 , n598010 , n70689 , n70690 );
and ( n598015 , n70683 , n64456 );
buf ( n70693 , n591728 );
and ( n598017 , n70693 , n64454 );
nor ( n598018 , n598015 , n598017 );
xnor ( n598019 , n598018 , n591786 );
and ( n70697 , n598014 , n598019 );
and ( n598021 , n597996 , n64451 );
and ( n70699 , n598019 , n598021 );
and ( n598023 , n598014 , n598021 );
or ( n70701 , n70697 , n70699 , n598023 );
and ( n70702 , n70693 , n64456 );
and ( n598026 , n70637 , n64454 );
nor ( n598027 , n70702 , n598026 );
xnor ( n70705 , n598027 , n591786 );
and ( n70706 , n70701 , n70705 );
and ( n598030 , n70683 , n64451 );
and ( n598031 , n70705 , n598030 );
and ( n70709 , n70701 , n598030 );
or ( n70710 , n70706 , n598031 , n70709 );
and ( n598034 , n70637 , n64456 );
and ( n598035 , n70261 , n64454 );
nor ( n70713 , n598034 , n598035 );
xnor ( n70714 , n70713 , n591786 );
and ( n598038 , n70710 , n70714 );
and ( n598039 , n70693 , n64451 );
and ( n598040 , n70714 , n598039 );
and ( n70718 , n70710 , n598039 );
or ( n598042 , n598038 , n598040 , n70718 );
and ( n70720 , n597402 , n64559 );
and ( n70721 , n597260 , n591880 );
nor ( n598045 , n70720 , n70721 );
xnor ( n70723 , n598045 , n64521 );
and ( n598047 , n70255 , n64491 );
and ( n70725 , n597569 , n64489 );
nor ( n70726 , n598047 , n70725 );
xnor ( n598050 , n70726 , n64448 );
and ( n70728 , n70723 , n598050 );
xor ( n598052 , n70710 , n70714 );
xor ( n598053 , n598052 , n598039 );
and ( n70731 , n598050 , n598053 );
and ( n598055 , n70723 , n598053 );
or ( n70733 , n70728 , n70731 , n598055 );
and ( n598057 , n598042 , n70733 );
xor ( n598058 , n70631 , n70635 );
xor ( n70736 , n598058 , n70638 );
and ( n598060 , n70733 , n70736 );
and ( n598061 , n598042 , n70736 );
or ( n598062 , n598057 , n598060 , n598061 );
and ( n70740 , n69491 , n64650 );
and ( n598064 , n69283 , n64648 );
nor ( n598065 , n70740 , n598064 );
xnor ( n70743 , n598065 , n591902 );
and ( n598067 , n598062 , n70743 );
xor ( n598068 , n597964 , n70645 );
xor ( n70746 , n598068 , n70648 );
and ( n598070 , n70743 , n70746 );
and ( n70748 , n598062 , n70746 );
or ( n598072 , n598067 , n598070 , n70748 );
and ( n70750 , n70651 , n598072 );
xor ( n70751 , n70335 , n597662 );
xor ( n598075 , n70751 , n70342 );
and ( n70753 , n598072 , n598075 );
and ( n598077 , n70651 , n598075 );
or ( n70755 , n70750 , n70753 , n598077 );
and ( n70756 , n595827 , n64862 );
and ( n598080 , n595633 , n64860 );
nor ( n598081 , n70756 , n598080 );
xnor ( n70759 , n598081 , n64764 );
and ( n598083 , n70755 , n70759 );
and ( n598084 , n596193 , n64744 );
and ( n70762 , n596057 , n64742 );
nor ( n598086 , n598084 , n70762 );
xnor ( n598087 , n598086 , n64623 );
and ( n598088 , n70759 , n598087 );
and ( n70766 , n70755 , n598087 );
or ( n598090 , n598083 , n598088 , n70766 );
and ( n598091 , n595103 , n592486 );
and ( n70769 , n67636 , n592484 );
nor ( n598093 , n598091 , n70769 );
xnor ( n598094 , n598093 , n64990 );
and ( n70772 , n598090 , n598094 );
xor ( n70773 , n70231 , n70235 );
xor ( n598097 , n70773 , n597611 );
and ( n598098 , n598094 , n598097 );
and ( n70776 , n598090 , n598097 );
or ( n598100 , n70772 , n598098 , n70776 );
and ( n70778 , n67636 , n592486 );
and ( n598102 , n594952 , n592484 );
nor ( n70780 , n70778 , n598102 );
xnor ( n70781 , n70780 , n64990 );
and ( n70782 , n598100 , n70781 );
xor ( n70783 , n597614 , n70295 );
xor ( n70784 , n70783 , n70298 );
and ( n70785 , n70781 , n70784 );
and ( n70786 , n598100 , n70784 );
or ( n70787 , n70782 , n70785 , n70786 );
and ( n70788 , n594295 , n592683 );
and ( n598112 , n66967 , n592681 );
nor ( n598113 , n70788 , n598112 );
xnor ( n70791 , n598113 , n592475 );
and ( n598115 , n70787 , n70791 );
xor ( n70793 , n597624 , n70305 );
xor ( n70794 , n70793 , n597631 );
and ( n70795 , n70791 , n70794 );
and ( n598119 , n70787 , n70794 );
or ( n70797 , n598115 , n70795 , n598119 );
and ( n598121 , n66793 , n65592 );
and ( n598122 , n594124 , n592913 );
nor ( n598123 , n598121 , n598122 );
xnor ( n70801 , n598123 , n592638 );
and ( n598125 , n70797 , n70801 );
xor ( n70803 , n597732 , n597736 );
xor ( n70804 , n70803 , n70426 );
and ( n598128 , n70801 , n70804 );
and ( n70806 , n70797 , n70804 );
or ( n598130 , n598125 , n598128 , n70806 );
xor ( n70808 , n70551 , n70555 );
xor ( n598132 , n70808 , n70558 );
and ( n598133 , n598130 , n598132 );
xor ( n70811 , n70429 , n597756 );
xor ( n70812 , n70811 , n70446 );
and ( n598136 , n598132 , n70812 );
and ( n598137 , n598130 , n70812 );
or ( n70815 , n598133 , n598136 , n598137 );
and ( n598139 , n597950 , n70815 );
and ( n598140 , n65493 , n594441 );
and ( n70818 , n65384 , n67116 );
nor ( n598142 , n598140 , n70818 );
xnor ( n598143 , n598142 , n66190 );
and ( n598144 , n70815 , n598143 );
and ( n70822 , n597950 , n598143 );
or ( n598146 , n598139 , n598144 , n70822 );
and ( n598147 , n592645 , n594807 );
and ( n70825 , n592468 , n594804 );
nor ( n598149 , n598147 , n70825 );
xnor ( n598150 , n598149 , n66187 );
xor ( n70828 , n70561 , n70563 );
xor ( n70829 , n70828 , n70566 );
and ( n70830 , n598150 , n70829 );
xor ( n70831 , n70461 , n70465 );
xor ( n70832 , n70831 , n597801 );
and ( n70833 , n70829 , n70832 );
and ( n70834 , n598150 , n70832 );
or ( n70835 , n70830 , n70833 , n70834 );
and ( n70836 , n598146 , n70835 );
xor ( n70837 , n597816 , n597818 );
xor ( n598161 , n70837 , n597829 );
and ( n70839 , n70835 , n598161 );
and ( n70840 , n598146 , n598161 );
or ( n70841 , n70836 , n70839 , n70840 );
xor ( n598165 , n597812 , n597832 );
xor ( n598166 , n598165 , n70512 );
and ( n70844 , n70841 , n598166 );
xor ( n598168 , n70579 , n70583 );
xor ( n598169 , n598168 , n70586 );
and ( n70847 , n598166 , n598169 );
and ( n598171 , n70841 , n598169 );
or ( n598172 , n70844 , n70847 , n598171 );
and ( n598173 , n597924 , n598172 );
xor ( n70851 , n597924 , n598172 );
xor ( n598175 , n70841 , n598166 );
xor ( n70853 , n598175 , n598169 );
and ( n598177 , n596198 , n64744 );
and ( n70855 , n596193 , n64742 );
nor ( n70856 , n598177 , n70855 );
xnor ( n598180 , n70856 , n64623 );
and ( n598181 , n69283 , n64650 );
and ( n70859 , n596600 , n64648 );
nor ( n598183 , n598181 , n70859 );
xnor ( n598184 , n598183 , n591902 );
and ( n70862 , n598180 , n598184 );
xor ( n598186 , n70651 , n598072 );
xor ( n598187 , n598186 , n598075 );
and ( n70865 , n598184 , n598187 );
and ( n70866 , n598180 , n598187 );
or ( n598190 , n70862 , n70865 , n70866 );
and ( n598191 , n595521 , n592340 );
and ( n70869 , n68160 , n65015 );
nor ( n598193 , n598191 , n70869 );
xnor ( n598194 , n598193 , n64847 );
and ( n70872 , n598190 , n598194 );
xor ( n598196 , n597668 , n70349 );
xor ( n598197 , n598196 , n597675 );
and ( n70875 , n598194 , n598197 );
and ( n598199 , n598190 , n598197 );
or ( n70877 , n70872 , n70875 , n598199 );
and ( n598201 , n68160 , n592340 );
and ( n70879 , n67940 , n65015 );
nor ( n598203 , n598201 , n70879 );
xnor ( n70881 , n598203 , n64847 );
and ( n70882 , n70877 , n70881 );
xor ( n598206 , n597678 , n70359 );
xor ( n70884 , n598206 , n70364 );
and ( n598208 , n70881 , n70884 );
and ( n70886 , n70877 , n70884 );
or ( n598210 , n70882 , n598208 , n70886 );
and ( n598211 , n594710 , n592683 );
and ( n70889 , n594295 , n592681 );
nor ( n598213 , n598211 , n70889 );
xnor ( n598214 , n598213 , n592475 );
and ( n70892 , n598210 , n598214 );
xor ( n70893 , n597690 , n70371 );
xor ( n598217 , n70893 , n70386 );
and ( n598218 , n598214 , n598217 );
and ( n70896 , n598210 , n598217 );
or ( n598220 , n70892 , n598218 , n70896 );
and ( n598221 , n66951 , n65592 );
and ( n70899 , n66793 , n592913 );
nor ( n598223 , n598221 , n70899 );
xnor ( n598224 , n598223 , n592638 );
and ( n70902 , n598220 , n598224 );
xor ( n70903 , n70389 , n70393 );
xor ( n70904 , n70903 , n597729 );
and ( n70905 , n598224 , n70904 );
and ( n70906 , n598220 , n70904 );
or ( n70907 , n70902 , n70905 , n70906 );
and ( n70908 , n65844 , n594210 );
and ( n70909 , n65630 , n66885 );
nor ( n70910 , n70908 , n70909 );
xnor ( n70911 , n70910 , n593434 );
and ( n598235 , n70907 , n70911 );
and ( n598236 , n593437 , n66457 );
and ( n70914 , n593298 , n593778 );
nor ( n598238 , n598236 , n70914 );
xnor ( n70916 , n598238 , n593160 );
and ( n598240 , n70911 , n70916 );
and ( n70918 , n70907 , n70916 );
or ( n70919 , n598235 , n598240 , n70918 );
and ( n598243 , n65384 , n594807 );
and ( n598244 , n592645 , n594804 );
nor ( n70922 , n598243 , n598244 );
xnor ( n70923 , n70922 , n66187 );
and ( n70924 , n70919 , n70923 );
and ( n598248 , n592806 , n594441 );
and ( n70926 , n65493 , n67116 );
nor ( n598250 , n598248 , n70926 );
xnor ( n598251 , n598250 , n66190 );
and ( n70929 , n70923 , n598251 );
and ( n598253 , n70919 , n598251 );
or ( n598254 , n70924 , n70929 , n598253 );
and ( n70932 , n69581 , n64650 );
and ( n70933 , n69491 , n64648 );
nor ( n70934 , n70932 , n70933 );
xnor ( n598258 , n70934 , n591902 );
and ( n598259 , n597260 , n64559 );
and ( n70937 , n69739 , n591880 );
nor ( n70938 , n598259 , n70937 );
xnor ( n598262 , n70938 , n64521 );
and ( n598263 , n598258 , n598262 );
xor ( n70941 , n598042 , n70733 );
xor ( n70942 , n70941 , n70736 );
and ( n70943 , n598262 , n70942 );
and ( n598267 , n598258 , n70942 );
or ( n70945 , n598263 , n70943 , n598267 );
and ( n598269 , n596600 , n64744 );
and ( n598270 , n596198 , n64742 );
nor ( n70948 , n598269 , n598270 );
xnor ( n70949 , n70948 , n64623 );
and ( n70950 , n70945 , n70949 );
xor ( n598274 , n598062 , n70743 );
xor ( n598275 , n598274 , n70746 );
and ( n70953 , n70949 , n598275 );
and ( n598277 , n70945 , n598275 );
or ( n598278 , n70950 , n70953 , n598277 );
and ( n70956 , n595633 , n592340 );
and ( n70957 , n595521 , n65015 );
nor ( n70958 , n70956 , n70957 );
xnor ( n70959 , n70958 , n64847 );
and ( n598283 , n598278 , n70959 );
and ( n598284 , n596057 , n64862 );
and ( n70962 , n595827 , n64860 );
nor ( n598286 , n598284 , n70962 );
xnor ( n598287 , n598286 , n64764 );
and ( n598288 , n70959 , n598287 );
and ( n70966 , n598278 , n598287 );
or ( n70967 , n598283 , n598288 , n70966 );
and ( n598291 , n67940 , n592486 );
and ( n70969 , n595103 , n592484 );
nor ( n598293 , n598291 , n70969 );
xnor ( n598294 , n598293 , n64990 );
and ( n70972 , n70967 , n598294 );
xor ( n598296 , n70755 , n70759 );
xor ( n598297 , n598296 , n598087 );
and ( n70975 , n598294 , n598297 );
and ( n70976 , n70967 , n598297 );
or ( n70977 , n70972 , n70975 , n70976 );
and ( n598301 , n594952 , n592683 );
and ( n598302 , n594710 , n592681 );
nor ( n70980 , n598301 , n598302 );
xnor ( n70981 , n70980 , n592475 );
and ( n598305 , n70977 , n70981 );
xor ( n598306 , n598090 , n598094 );
xor ( n70984 , n598306 , n598097 );
and ( n70985 , n70981 , n70984 );
and ( n70986 , n70977 , n70984 );
or ( n598310 , n598305 , n70985 , n70986 );
and ( n70988 , n66967 , n65592 );
and ( n598312 , n66951 , n592913 );
nor ( n70990 , n70988 , n598312 );
xnor ( n598314 , n70990 , n592638 );
and ( n70992 , n598310 , n598314 );
xor ( n598316 , n598100 , n70781 );
xor ( n598317 , n598316 , n70784 );
and ( n70995 , n598314 , n598317 );
and ( n70996 , n598310 , n598317 );
or ( n598320 , n70992 , n70995 , n70996 );
and ( n70998 , n66104 , n66457 );
and ( n70999 , n593437 , n593778 );
nor ( n598323 , n70998 , n70999 );
xnor ( n71001 , n598323 , n593160 );
and ( n598325 , n598320 , n71001 );
and ( n598326 , n66507 , n66142 );
and ( n71004 , n593520 , n66140 );
nor ( n598328 , n598326 , n71004 );
xnor ( n71006 , n598328 , n592960 );
and ( n71007 , n71001 , n71006 );
and ( n598331 , n598320 , n71006 );
or ( n598332 , n598325 , n71007 , n598331 );
and ( n71010 , n65640 , n594441 );
and ( n598334 , n592806 , n67116 );
nor ( n71012 , n71010 , n598334 );
xnor ( n71013 , n71012 , n66190 );
and ( n598337 , n598332 , n71013 );
xor ( n71015 , n70605 , n597932 );
xor ( n598339 , n71015 , n597935 );
and ( n598340 , n71013 , n598339 );
and ( n71018 , n598332 , n598339 );
or ( n71019 , n598337 , n598340 , n71018 );
xor ( n71020 , n70615 , n70619 );
xor ( n598344 , n71020 , n70624 );
and ( n71022 , n71019 , n598344 );
xor ( n71023 , n598130 , n598132 );
xor ( n598347 , n71023 , n70812 );
and ( n598348 , n598344 , n598347 );
and ( n71026 , n71019 , n598347 );
or ( n71027 , n71022 , n598348 , n71026 );
and ( n598351 , n598254 , n71027 );
xor ( n598352 , n597950 , n70815 );
xor ( n71030 , n598352 , n598143 );
and ( n598354 , n71027 , n71030 );
and ( n598355 , n598254 , n71030 );
or ( n71033 , n598351 , n598354 , n598355 );
xor ( n598357 , n70569 , n597896 );
xor ( n71035 , n598357 , n597899 );
and ( n71036 , n71033 , n71035 );
xor ( n71037 , n598146 , n70835 );
xor ( n71038 , n71037 , n598161 );
and ( n598362 , n71035 , n71038 );
and ( n71040 , n71033 , n71038 );
or ( n598364 , n71036 , n598362 , n71040 );
and ( n71042 , n70853 , n598364 );
xor ( n71043 , n70853 , n598364 );
xor ( n598367 , n71033 , n71035 );
xor ( n598368 , n598367 , n71038 );
and ( n71046 , n593520 , n66457 );
and ( n598370 , n66104 , n593778 );
nor ( n598371 , n71046 , n598370 );
xnor ( n71049 , n598371 , n593160 );
and ( n598373 , n66606 , n66142 );
and ( n71051 , n66507 , n66140 );
nor ( n71052 , n598373 , n71051 );
xnor ( n71053 , n71052 , n592960 );
and ( n71054 , n71049 , n71053 );
xor ( n71055 , n598210 , n598214 );
xor ( n71056 , n71055 , n598217 );
and ( n598380 , n71053 , n71056 );
and ( n598381 , n71049 , n71056 );
or ( n71059 , n71054 , n598380 , n598381 );
and ( n598383 , n65630 , n594441 );
and ( n71061 , n65640 , n67116 );
nor ( n598385 , n598383 , n71061 );
xnor ( n71063 , n598385 , n66190 );
and ( n598387 , n71059 , n71063 );
and ( n598388 , n593298 , n594210 );
and ( n71066 , n65844 , n66885 );
nor ( n71067 , n598388 , n71066 );
xnor ( n71068 , n71067 , n593434 );
and ( n71069 , n71063 , n71068 );
and ( n71070 , n71059 , n71068 );
or ( n71071 , n598387 , n71069 , n71070 );
and ( n71072 , n594124 , n593256 );
and ( n71073 , n66606 , n593254 );
nor ( n71074 , n71072 , n71073 );
xnor ( n598398 , n71074 , n65490 );
xor ( n71076 , n70787 , n70791 );
xor ( n598400 , n71076 , n70794 );
and ( n71078 , n598398 , n598400 );
xor ( n71079 , n598220 , n598224 );
xor ( n71080 , n71079 , n70904 );
and ( n71081 , n598400 , n71080 );
and ( n598405 , n598398 , n71080 );
or ( n71083 , n71078 , n71081 , n598405 );
and ( n71084 , n71071 , n71083 );
xor ( n71085 , n70797 , n70801 );
xor ( n71086 , n71085 , n70804 );
and ( n71087 , n71083 , n71086 );
and ( n71088 , n71071 , n71086 );
or ( n598412 , n71084 , n71087 , n71088 );
and ( n598413 , n65493 , n594807 );
and ( n598414 , n65384 , n594804 );
nor ( n71092 , n598413 , n598414 );
xnor ( n598416 , n71092 , n66187 );
xor ( n71094 , n70907 , n70911 );
xor ( n71095 , n71094 , n70916 );
and ( n598419 , n598416 , n71095 );
xor ( n71097 , n598332 , n71013 );
xor ( n598421 , n71097 , n598339 );
and ( n71099 , n71095 , n598421 );
and ( n71100 , n598416 , n598421 );
or ( n71101 , n598419 , n71099 , n71100 );
and ( n598425 , n598412 , n71101 );
xor ( n598426 , n70919 , n70923 );
xor ( n71104 , n598426 , n598251 );
and ( n598428 , n71101 , n71104 );
and ( n598429 , n598412 , n71104 );
or ( n71107 , n598425 , n598428 , n598429 );
xor ( n598431 , n598254 , n71027 );
xor ( n598432 , n598431 , n71030 );
and ( n598433 , n71107 , n598432 );
xor ( n71111 , n598150 , n70829 );
xor ( n598435 , n71111 , n70832 );
and ( n598436 , n598432 , n598435 );
and ( n71114 , n71107 , n598435 );
or ( n598438 , n598433 , n598436 , n71114 );
and ( n598439 , n598368 , n598438 );
xor ( n71117 , n598368 , n598438 );
xor ( n598441 , n71107 , n598432 );
xor ( n71119 , n598441 , n598435 );
and ( n598443 , n596198 , n64862 );
and ( n71121 , n596193 , n64860 );
nor ( n71122 , n598443 , n71121 );
xnor ( n598446 , n71122 , n64764 );
and ( n71124 , n69283 , n64744 );
and ( n598448 , n596600 , n64742 );
nor ( n71126 , n71124 , n598448 );
xnor ( n71127 , n71126 , n64623 );
and ( n598451 , n598446 , n71127 );
xor ( n598452 , n597978 , n70660 );
and ( n71130 , n70652 , n64489 );
not ( n598454 , n71130 );
and ( n598455 , n598454 , n64448 );
and ( n71133 , n70652 , n64491 );
and ( n598457 , n597980 , n64489 );
nor ( n598458 , n71133 , n598457 );
xnor ( n598459 , n598458 , n64448 );
and ( n71137 , n598455 , n598459 );
and ( n598461 , n597980 , n64491 );
and ( n598462 , n70663 , n64489 );
nor ( n71140 , n598461 , n598462 );
xnor ( n598464 , n71140 , n64448 );
and ( n598465 , n71137 , n598464 );
and ( n71143 , n598464 , n70653 );
and ( n71144 , n71137 , n70653 );
or ( n71145 , n598465 , n71143 , n71144 );
and ( n598469 , n598452 , n71145 );
and ( n71147 , n70663 , n64491 );
and ( n598471 , n597996 , n64489 );
nor ( n71149 , n71147 , n598471 );
xnor ( n598473 , n71149 , n64448 );
and ( n71151 , n71145 , n598473 );
and ( n71152 , n598452 , n598473 );
or ( n71153 , n598469 , n71151 , n71152 );
and ( n71154 , n597996 , n64491 );
and ( n71155 , n70683 , n64489 );
nor ( n71156 , n71154 , n71155 );
xnor ( n598480 , n71156 , n64448 );
and ( n598481 , n71153 , n598480 );
xor ( n71159 , n597984 , n70666 );
xor ( n598483 , n71159 , n597991 );
and ( n598484 , n598480 , n598483 );
and ( n71162 , n71153 , n598483 );
or ( n598486 , n598481 , n598484 , n71162 );
and ( n71164 , n70683 , n64491 );
and ( n71165 , n70693 , n64489 );
nor ( n71166 , n71164 , n71165 );
xnor ( n598490 , n71166 , n64448 );
and ( n71168 , n598486 , n598490 );
xor ( n598492 , n70671 , n597999 );
xor ( n598493 , n598492 , n70678 );
and ( n71171 , n598490 , n598493 );
and ( n71172 , n598486 , n598493 );
or ( n598496 , n71168 , n71171 , n71172 );
and ( n71174 , n70693 , n64491 );
and ( n598498 , n70637 , n64489 );
nor ( n598499 , n71174 , n598498 );
xnor ( n71177 , n598499 , n64448 );
and ( n71178 , n598496 , n71177 );
xor ( n71179 , n598004 , n70686 );
xor ( n71180 , n71179 , n70688 );
and ( n71181 , n71177 , n71180 );
and ( n71182 , n598496 , n71180 );
or ( n71183 , n71178 , n71181 , n71182 );
and ( n71184 , n70637 , n64491 );
and ( n71185 , n70261 , n64489 );
nor ( n71186 , n71184 , n71185 );
xnor ( n71187 , n71186 , n64448 );
and ( n71188 , n71183 , n71187 );
xor ( n71189 , n598014 , n598019 );
xor ( n71190 , n71189 , n598021 );
and ( n71191 , n71187 , n71190 );
and ( n71192 , n71183 , n71190 );
or ( n71193 , n71188 , n71191 , n71192 );
and ( n71194 , n70261 , n64491 );
and ( n598518 , n70255 , n64489 );
nor ( n71196 , n71194 , n598518 );
xnor ( n71197 , n71196 , n64448 );
and ( n71198 , n71193 , n71197 );
xor ( n598522 , n70701 , n70705 );
xor ( n598523 , n598522 , n598030 );
and ( n71201 , n71197 , n598523 );
and ( n71202 , n71193 , n598523 );
or ( n71203 , n71198 , n71201 , n71202 );
and ( n598527 , n69739 , n64650 );
and ( n598528 , n69581 , n64648 );
nor ( n71206 , n598527 , n598528 );
xnor ( n71207 , n71206 , n591902 );
and ( n71208 , n71203 , n71207 );
xor ( n598532 , n70723 , n598050 );
xor ( n598533 , n598532 , n598053 );
and ( n71211 , n71207 , n598533 );
and ( n71212 , n71203 , n598533 );
or ( n71213 , n71208 , n71211 , n71212 );
and ( n598537 , n597402 , n64650 );
and ( n598538 , n597260 , n64648 );
nor ( n71216 , n598537 , n598538 );
xnor ( n598540 , n71216 , n591902 );
and ( n598541 , n70255 , n64559 );
and ( n71219 , n597569 , n591880 );
nor ( n598543 , n598541 , n71219 );
xnor ( n71221 , n598543 , n64521 );
and ( n71222 , n598540 , n71221 );
xor ( n598546 , n71183 , n71187 );
xor ( n598547 , n598546 , n71190 );
and ( n71225 , n71221 , n598547 );
and ( n598549 , n598540 , n598547 );
or ( n71227 , n71222 , n71225 , n598549 );
and ( n71228 , n597569 , n64559 );
and ( n71229 , n597402 , n591880 );
nor ( n598553 , n71228 , n71229 );
xnor ( n598554 , n598553 , n64521 );
and ( n71232 , n71227 , n598554 );
xor ( n598556 , n71193 , n71197 );
xor ( n71234 , n598556 , n598523 );
and ( n71235 , n598554 , n71234 );
and ( n71236 , n71227 , n71234 );
or ( n598560 , n71232 , n71235 , n71236 );
and ( n598561 , n69491 , n64744 );
and ( n71239 , n69283 , n64742 );
nor ( n598563 , n598561 , n71239 );
xnor ( n71241 , n598563 , n64623 );
and ( n71242 , n598560 , n71241 );
xor ( n71243 , n71203 , n71207 );
xor ( n598567 , n71243 , n598533 );
and ( n71245 , n71241 , n598567 );
and ( n598569 , n598560 , n598567 );
or ( n71247 , n71242 , n71245 , n598569 );
xor ( n71248 , n71213 , n71247 );
xor ( n598572 , n598258 , n598262 );
xor ( n598573 , n598572 , n70942 );
xor ( n71251 , n71248 , n598573 );
and ( n598575 , n71127 , n71251 );
and ( n71253 , n598446 , n71251 );
or ( n598577 , n598451 , n598575 , n71253 );
and ( n71255 , n595521 , n592486 );
and ( n71256 , n68160 , n592484 );
nor ( n598580 , n71255 , n71256 );
xnor ( n71258 , n598580 , n64990 );
and ( n598582 , n598577 , n71258 );
xor ( n71260 , n70945 , n70949 );
xor ( n71261 , n71260 , n598275 );
and ( n598585 , n71258 , n71261 );
and ( n598586 , n598577 , n71261 );
or ( n71264 , n598582 , n598585 , n598586 );
and ( n598588 , n595103 , n592683 );
and ( n598589 , n67636 , n592681 );
nor ( n71267 , n598588 , n598589 );
xnor ( n598591 , n71267 , n592475 );
and ( n598592 , n71264 , n598591 );
and ( n598593 , n68160 , n592486 );
and ( n71271 , n67940 , n592484 );
nor ( n598595 , n598593 , n71271 );
xnor ( n598596 , n598595 , n64990 );
and ( n71274 , n598591 , n598596 );
and ( n598598 , n71264 , n598596 );
or ( n598599 , n598592 , n71274 , n598598 );
and ( n598600 , n594710 , n65592 );
and ( n598601 , n594295 , n592913 );
nor ( n71279 , n598600 , n598601 );
xnor ( n598603 , n71279 , n592638 );
and ( n71281 , n598599 , n598603 );
xor ( n598605 , n70967 , n598294 );
xor ( n71283 , n598605 , n598297 );
and ( n71284 , n598603 , n71283 );
and ( n71285 , n598599 , n71283 );
or ( n71286 , n71281 , n71284 , n71285 );
and ( n71287 , n66951 , n593256 );
and ( n71288 , n66793 , n593254 );
nor ( n71289 , n71287 , n71288 );
xnor ( n71290 , n71289 , n65490 );
and ( n71291 , n71286 , n71290 );
xor ( n71292 , n70977 , n70981 );
xor ( n71293 , n71292 , n70984 );
and ( n71294 , n71290 , n71293 );
and ( n598618 , n71286 , n71293 );
or ( n71296 , n71291 , n71294 , n598618 );
and ( n598620 , n65844 , n594441 );
and ( n598621 , n65630 , n67116 );
nor ( n71299 , n598620 , n598621 );
xnor ( n598623 , n71299 , n66190 );
and ( n598624 , n71296 , n598623 );
and ( n71302 , n593437 , n594210 );
and ( n598626 , n593298 , n66885 );
nor ( n598627 , n71302 , n598626 );
xnor ( n598628 , n598627 , n593434 );
and ( n71306 , n598623 , n598628 );
and ( n598630 , n71296 , n598628 );
or ( n598631 , n598624 , n71306 , n598630 );
and ( n71309 , n66507 , n66457 );
and ( n598633 , n593520 , n593778 );
nor ( n71311 , n71309 , n598633 );
xnor ( n598635 , n71311 , n593160 );
and ( n71313 , n594124 , n66142 );
and ( n71314 , n66606 , n66140 );
nor ( n598638 , n71313 , n71314 );
xnor ( n71316 , n598638 , n592960 );
and ( n598640 , n598635 , n71316 );
and ( n598641 , n71213 , n71247 );
and ( n598642 , n71247 , n598573 );
and ( n598643 , n71213 , n598573 );
or ( n71321 , n598641 , n598642 , n598643 );
and ( n598645 , n595827 , n592340 );
and ( n598646 , n595633 , n65015 );
nor ( n71324 , n598645 , n598646 );
xnor ( n598648 , n71324 , n64847 );
and ( n598649 , n71321 , n598648 );
and ( n71327 , n596193 , n64862 );
and ( n71328 , n596057 , n64860 );
nor ( n598652 , n71327 , n71328 );
xnor ( n71330 , n598652 , n64764 );
and ( n71331 , n598648 , n71330 );
and ( n598655 , n71321 , n71330 );
or ( n598656 , n598649 , n71331 , n598655 );
xor ( n71334 , n598278 , n70959 );
xor ( n598658 , n71334 , n598287 );
and ( n598659 , n598656 , n598658 );
xor ( n71337 , n598180 , n598184 );
xor ( n598661 , n71337 , n598187 );
and ( n598662 , n598658 , n598661 );
and ( n71340 , n598656 , n598661 );
or ( n598664 , n598659 , n598662 , n71340 );
and ( n598665 , n67636 , n592683 );
and ( n598666 , n594952 , n592681 );
nor ( n71344 , n598665 , n598666 );
xnor ( n598668 , n71344 , n592475 );
and ( n598669 , n598664 , n598668 );
xor ( n71347 , n598190 , n598194 );
xor ( n71348 , n71347 , n598197 );
and ( n71349 , n598668 , n71348 );
and ( n71350 , n598664 , n71348 );
or ( n71351 , n598669 , n71349 , n71350 );
and ( n71352 , n594295 , n65592 );
and ( n71353 , n66967 , n592913 );
nor ( n71354 , n71352 , n71353 );
xnor ( n598678 , n71354 , n592638 );
xor ( n598679 , n71351 , n598678 );
xor ( n71357 , n70877 , n70881 );
xor ( n598681 , n71357 , n70884 );
xor ( n598682 , n598679 , n598681 );
and ( n71360 , n71316 , n598682 );
and ( n598684 , n598635 , n598682 );
or ( n598685 , n598640 , n71360 , n598684 );
and ( n71363 , n65640 , n594807 );
and ( n598687 , n592806 , n594804 );
nor ( n71365 , n71363 , n598687 );
xnor ( n598689 , n71365 , n66187 );
and ( n598690 , n598685 , n598689 );
and ( n71368 , n71351 , n598678 );
and ( n598692 , n598678 , n598681 );
and ( n598693 , n71351 , n598681 );
or ( n598694 , n71368 , n598692 , n598693 );
and ( n71372 , n66793 , n593256 );
and ( n598696 , n594124 , n593254 );
nor ( n71374 , n71372 , n598696 );
xnor ( n598698 , n71374 , n65490 );
xor ( n598699 , n598694 , n598698 );
xor ( n71377 , n598310 , n598314 );
xor ( n598701 , n71377 , n598317 );
xor ( n598702 , n598699 , n598701 );
and ( n71380 , n598689 , n598702 );
and ( n598704 , n598685 , n598702 );
or ( n598705 , n598690 , n71380 , n598704 );
and ( n71383 , n598631 , n598705 );
and ( n598707 , n592806 , n594807 );
and ( n71385 , n65493 , n594804 );
nor ( n598709 , n598707 , n71385 );
xnor ( n71387 , n598709 , n66187 );
and ( n71388 , n598705 , n71387 );
and ( n71389 , n598631 , n71387 );
or ( n598713 , n71383 , n71388 , n71389 );
and ( n598714 , n598694 , n598698 );
and ( n598715 , n598698 , n598701 );
and ( n71393 , n598694 , n598701 );
or ( n598717 , n598714 , n598715 , n71393 );
xor ( n598718 , n598320 , n71001 );
xor ( n71396 , n598718 , n71006 );
and ( n598720 , n598717 , n71396 );
xor ( n598721 , n598398 , n598400 );
xor ( n71399 , n598721 , n71080 );
and ( n71400 , n71396 , n71399 );
and ( n71401 , n598717 , n71399 );
or ( n598725 , n598720 , n71400 , n71401 );
and ( n71403 , n598713 , n598725 );
xor ( n71404 , n71071 , n71083 );
xor ( n71405 , n71404 , n71086 );
and ( n71406 , n598725 , n71405 );
and ( n71407 , n598713 , n71405 );
or ( n71408 , n71403 , n71406 , n71407 );
xor ( n71409 , n598412 , n71101 );
xor ( n71410 , n71409 , n71104 );
and ( n598734 , n71408 , n71410 );
xor ( n71412 , n71019 , n598344 );
xor ( n598736 , n71412 , n598347 );
and ( n71414 , n71410 , n598736 );
and ( n71415 , n71408 , n598736 );
or ( n71416 , n598734 , n71414 , n71415 );
and ( n71417 , n71119 , n71416 );
xor ( n71418 , n71119 , n71416 );
xor ( n71419 , n71408 , n71410 );
xor ( n71420 , n71419 , n598736 );
and ( n71421 , n69581 , n64744 );
and ( n71422 , n69491 , n64742 );
nor ( n71423 , n71421 , n71422 );
xnor ( n598747 , n71423 , n64623 );
and ( n71425 , n597260 , n64650 );
and ( n71426 , n69739 , n64648 );
nor ( n71427 , n71425 , n71426 );
xnor ( n71428 , n71427 , n591902 );
and ( n71429 , n598747 , n71428 );
xor ( n71430 , n71227 , n598554 );
xor ( n598754 , n71430 , n71234 );
and ( n71432 , n71428 , n598754 );
and ( n71433 , n598747 , n598754 );
or ( n71434 , n71429 , n71432 , n71433 );
and ( n71435 , n596600 , n64862 );
and ( n71436 , n596198 , n64860 );
nor ( n71437 , n71435 , n71436 );
xnor ( n598761 , n71437 , n64764 );
and ( n71439 , n71434 , n598761 );
xor ( n598763 , n598560 , n71241 );
xor ( n598764 , n598763 , n598567 );
and ( n71442 , n598761 , n598764 );
and ( n598766 , n71434 , n598764 );
or ( n598767 , n71439 , n71442 , n598766 );
and ( n71445 , n595633 , n592486 );
and ( n598769 , n595521 , n592484 );
nor ( n71447 , n71445 , n598769 );
xnor ( n71448 , n71447 , n64990 );
and ( n71449 , n598767 , n71448 );
and ( n71450 , n596057 , n592340 );
and ( n598774 , n595827 , n65015 );
nor ( n71452 , n71450 , n598774 );
xnor ( n598776 , n71452 , n64847 );
and ( n71454 , n71448 , n598776 );
and ( n71455 , n598767 , n598776 );
or ( n71456 , n71449 , n71454 , n71455 );
and ( n71457 , n67940 , n592683 );
and ( n71458 , n595103 , n592681 );
nor ( n71459 , n71457 , n71458 );
xnor ( n598783 , n71459 , n592475 );
and ( n598784 , n71456 , n598783 );
xor ( n71462 , n71321 , n598648 );
xor ( n598786 , n71462 , n71330 );
and ( n71464 , n598783 , n598786 );
and ( n71465 , n71456 , n598786 );
or ( n71466 , n598784 , n71464 , n71465 );
and ( n71467 , n594952 , n65592 );
and ( n71468 , n594710 , n592913 );
nor ( n71469 , n71467 , n71468 );
xnor ( n71470 , n71469 , n592638 );
and ( n71471 , n71466 , n71470 );
xor ( n71472 , n598656 , n598658 );
xor ( n71473 , n71472 , n598661 );
and ( n598797 , n71470 , n71473 );
and ( n598798 , n71466 , n71473 );
or ( n71476 , n71471 , n598797 , n598798 );
and ( n598800 , n66967 , n593256 );
and ( n71478 , n66951 , n593254 );
nor ( n71479 , n598800 , n71478 );
xnor ( n71480 , n71479 , n65490 );
and ( n71481 , n71476 , n71480 );
xor ( n71482 , n598664 , n598668 );
xor ( n71483 , n71482 , n71348 );
and ( n598807 , n71480 , n71483 );
and ( n71485 , n71476 , n71483 );
or ( n598809 , n71481 , n598807 , n71485 );
and ( n71487 , n66104 , n594210 );
and ( n598811 , n593437 , n66885 );
nor ( n71489 , n71487 , n598811 );
xnor ( n71490 , n71489 , n593434 );
and ( n71491 , n598809 , n71490 );
xor ( n71492 , n71286 , n71290 );
xor ( n71493 , n71492 , n71293 );
and ( n71494 , n71490 , n71493 );
and ( n598818 , n598809 , n71493 );
or ( n598819 , n71491 , n71494 , n598818 );
xor ( n71497 , n71296 , n598623 );
xor ( n598821 , n71497 , n598628 );
and ( n598822 , n598819 , n598821 );
xor ( n71500 , n71049 , n71053 );
xor ( n598824 , n71500 , n71056 );
and ( n598825 , n598821 , n598824 );
and ( n598826 , n598819 , n598824 );
or ( n71504 , n598822 , n598825 , n598826 );
xor ( n598828 , n71059 , n71063 );
xor ( n71506 , n598828 , n71068 );
and ( n71507 , n71504 , n71506 );
xor ( n598831 , n598717 , n71396 );
xor ( n71509 , n598831 , n71399 );
and ( n598833 , n71506 , n71509 );
and ( n71511 , n71504 , n71509 );
or ( n71512 , n71507 , n598833 , n71511 );
xor ( n71513 , n598416 , n71095 );
xor ( n71514 , n71513 , n598421 );
and ( n598838 , n71512 , n71514 );
xor ( n598839 , n598713 , n598725 );
xor ( n71517 , n598839 , n71405 );
and ( n598841 , n71514 , n71517 );
and ( n598842 , n71512 , n71517 );
or ( n71520 , n598838 , n598841 , n598842 );
and ( n598844 , n71420 , n71520 );
xor ( n598845 , n71420 , n71520 );
xor ( n71523 , n71512 , n71514 );
xor ( n598847 , n71523 , n71517 );
and ( n598848 , n66606 , n66457 );
and ( n598849 , n66507 , n593778 );
nor ( n598850 , n598848 , n598849 );
xnor ( n71528 , n598850 , n593160 );
and ( n71529 , n66793 , n66142 );
and ( n71530 , n594124 , n66140 );
nor ( n598854 , n71529 , n71530 );
xnor ( n598855 , n598854 , n592960 );
and ( n71533 , n71528 , n598855 );
xor ( n598857 , n598599 , n598603 );
xor ( n598858 , n598857 , n71283 );
and ( n71536 , n598855 , n598858 );
and ( n598860 , n71528 , n598858 );
or ( n598861 , n71533 , n71536 , n598860 );
and ( n71539 , n65630 , n594807 );
and ( n71540 , n65640 , n594804 );
nor ( n71541 , n71539 , n71540 );
xnor ( n598865 , n71541 , n66187 );
and ( n598866 , n598861 , n598865 );
and ( n71544 , n593298 , n594441 );
and ( n598868 , n65844 , n67116 );
nor ( n598869 , n71544 , n598868 );
xnor ( n71547 , n598869 , n66190 );
and ( n71548 , n598865 , n71547 );
and ( n71549 , n598861 , n71547 );
or ( n598873 , n598866 , n71548 , n71549 );
xor ( n598874 , n598455 , n598459 );
and ( n71552 , n70652 , n591880 );
not ( n598876 , n71552 );
and ( n598877 , n598876 , n64521 );
and ( n71555 , n70652 , n64559 );
and ( n71556 , n597980 , n591880 );
nor ( n598880 , n71555 , n71556 );
xnor ( n71558 , n598880 , n64521 );
and ( n598882 , n598877 , n71558 );
and ( n71560 , n597980 , n64559 );
and ( n71561 , n70663 , n591880 );
nor ( n598885 , n71560 , n71561 );
xnor ( n71563 , n598885 , n64521 );
and ( n71564 , n598882 , n71563 );
and ( n71565 , n71563 , n71130 );
and ( n598889 , n598882 , n71130 );
or ( n71567 , n71564 , n71565 , n598889 );
and ( n598891 , n598874 , n71567 );
and ( n598892 , n70663 , n64559 );
and ( n71570 , n597996 , n591880 );
nor ( n71571 , n598892 , n71570 );
xnor ( n598895 , n71571 , n64521 );
and ( n71573 , n71567 , n598895 );
and ( n598897 , n598874 , n598895 );
or ( n71575 , n598891 , n71573 , n598897 );
and ( n598899 , n597996 , n64559 );
and ( n598900 , n70683 , n591880 );
nor ( n71578 , n598899 , n598900 );
xnor ( n71579 , n71578 , n64521 );
and ( n598903 , n71575 , n71579 );
xor ( n71581 , n71137 , n598464 );
xor ( n598905 , n71581 , n70653 );
and ( n71583 , n71579 , n598905 );
and ( n598907 , n71575 , n598905 );
or ( n71585 , n598903 , n71583 , n598907 );
and ( n71586 , n70683 , n64559 );
and ( n598910 , n70693 , n591880 );
nor ( n598911 , n71586 , n598910 );
xnor ( n71589 , n598911 , n64521 );
and ( n598913 , n71585 , n71589 );
xor ( n598914 , n598452 , n71145 );
xor ( n71592 , n598914 , n598473 );
and ( n598916 , n71589 , n71592 );
and ( n598917 , n71585 , n71592 );
or ( n71595 , n598913 , n598916 , n598917 );
and ( n71596 , n70693 , n64559 );
and ( n598920 , n70637 , n591880 );
nor ( n598921 , n71596 , n598920 );
xnor ( n71599 , n598921 , n64521 );
and ( n598923 , n71595 , n71599 );
xor ( n598924 , n71153 , n598480 );
xor ( n71602 , n598924 , n598483 );
and ( n598926 , n71599 , n71602 );
and ( n598927 , n71595 , n71602 );
or ( n71605 , n598923 , n598926 , n598927 );
and ( n71606 , n70637 , n64559 );
and ( n598930 , n70261 , n591880 );
nor ( n598931 , n71606 , n598930 );
xnor ( n71609 , n598931 , n64521 );
and ( n598933 , n71605 , n71609 );
xor ( n71611 , n598486 , n598490 );
xor ( n598935 , n71611 , n598493 );
and ( n71613 , n71609 , n598935 );
and ( n598937 , n71605 , n598935 );
or ( n71615 , n598933 , n71613 , n598937 );
and ( n598939 , n70261 , n64559 );
and ( n598940 , n70255 , n591880 );
nor ( n71618 , n598939 , n598940 );
xnor ( n598942 , n71618 , n64521 );
and ( n598943 , n71615 , n598942 );
xor ( n71621 , n598496 , n71177 );
xor ( n71622 , n71621 , n71180 );
and ( n598946 , n598942 , n71622 );
and ( n71624 , n71615 , n71622 );
or ( n598948 , n598943 , n598946 , n71624 );
and ( n71626 , n69739 , n64744 );
and ( n598950 , n69581 , n64742 );
nor ( n598951 , n71626 , n598950 );
xnor ( n71629 , n598951 , n64623 );
and ( n598953 , n598948 , n71629 );
xor ( n598954 , n598540 , n71221 );
xor ( n71632 , n598954 , n598547 );
and ( n71633 , n71629 , n71632 );
and ( n598957 , n598948 , n71632 );
or ( n598958 , n598953 , n71633 , n598957 );
and ( n71636 , n597402 , n64744 );
and ( n598960 , n597260 , n64742 );
nor ( n598961 , n71636 , n598960 );
xnor ( n71639 , n598961 , n64623 );
and ( n598963 , n70255 , n64650 );
and ( n598964 , n597569 , n64648 );
nor ( n71642 , n598963 , n598964 );
xnor ( n71643 , n71642 , n591902 );
and ( n71644 , n71639 , n71643 );
xor ( n598968 , n71605 , n71609 );
xor ( n598969 , n598968 , n598935 );
and ( n71647 , n71643 , n598969 );
and ( n598971 , n71639 , n598969 );
or ( n598972 , n71644 , n71647 , n598971 );
and ( n71650 , n597569 , n64650 );
and ( n598974 , n597402 , n64648 );
nor ( n598975 , n71650 , n598974 );
xnor ( n71653 , n598975 , n591902 );
and ( n598977 , n598972 , n71653 );
xor ( n598978 , n71615 , n598942 );
xor ( n598979 , n598978 , n71622 );
and ( n71657 , n71653 , n598979 );
and ( n598981 , n598972 , n598979 );
or ( n71659 , n598977 , n71657 , n598981 );
and ( n598983 , n69491 , n64862 );
and ( n598984 , n69283 , n64860 );
nor ( n71662 , n598983 , n598984 );
xnor ( n598986 , n71662 , n64764 );
and ( n598987 , n71659 , n598986 );
xor ( n71665 , n598948 , n71629 );
xor ( n71666 , n71665 , n71632 );
and ( n598990 , n598986 , n71666 );
and ( n598991 , n71659 , n71666 );
or ( n71669 , n598987 , n598990 , n598991 );
and ( n71670 , n598958 , n71669 );
xor ( n598994 , n598747 , n71428 );
xor ( n71672 , n598994 , n598754 );
and ( n598996 , n71669 , n71672 );
and ( n71674 , n598958 , n71672 );
or ( n71675 , n71670 , n598996 , n71674 );
and ( n71676 , n595827 , n592486 );
and ( n599000 , n595633 , n592484 );
nor ( n599001 , n71676 , n599000 );
xnor ( n71679 , n599001 , n64990 );
and ( n599003 , n71675 , n71679 );
and ( n71681 , n596193 , n592340 );
and ( n71682 , n596057 , n65015 );
nor ( n599006 , n71681 , n71682 );
xnor ( n599007 , n599006 , n64847 );
and ( n599008 , n71679 , n599007 );
and ( n71686 , n71675 , n599007 );
or ( n599010 , n599003 , n599008 , n71686 );
and ( n71688 , n68160 , n592683 );
and ( n599012 , n67940 , n592681 );
nor ( n599013 , n71688 , n599012 );
xnor ( n71691 , n599013 , n592475 );
and ( n599015 , n599010 , n71691 );
xor ( n599016 , n598446 , n71127 );
xor ( n71694 , n599016 , n71251 );
and ( n599018 , n71691 , n71694 );
and ( n71696 , n599010 , n71694 );
or ( n599020 , n599015 , n599018 , n71696 );
and ( n71698 , n67636 , n65592 );
and ( n71699 , n594952 , n592913 );
nor ( n599023 , n71698 , n71699 );
xnor ( n71701 , n599023 , n592638 );
and ( n599025 , n599020 , n71701 );
xor ( n71703 , n598577 , n71258 );
xor ( n71704 , n71703 , n71261 );
and ( n599028 , n71701 , n71704 );
and ( n599029 , n599020 , n71704 );
or ( n71707 , n599025 , n599028 , n599029 );
and ( n599031 , n594295 , n593256 );
and ( n599032 , n66967 , n593254 );
nor ( n71710 , n599031 , n599032 );
xnor ( n599034 , n71710 , n65490 );
and ( n599035 , n71707 , n599034 );
xor ( n599036 , n71264 , n598591 );
xor ( n71714 , n599036 , n598596 );
and ( n599038 , n599034 , n71714 );
and ( n599039 , n71707 , n71714 );
or ( n71717 , n599035 , n599038 , n599039 );
and ( n599041 , n593437 , n594441 );
and ( n599042 , n593298 , n67116 );
nor ( n599043 , n599041 , n599042 );
xnor ( n71721 , n599043 , n66190 );
and ( n599045 , n71717 , n71721 );
and ( n71723 , n593520 , n594210 );
and ( n599047 , n66104 , n66885 );
nor ( n71725 , n71723 , n599047 );
xnor ( n71726 , n71725 , n593434 );
and ( n599050 , n71721 , n71726 );
and ( n71728 , n71717 , n71726 );
or ( n599052 , n599045 , n599050 , n71728 );
xor ( n71730 , n598635 , n71316 );
xor ( n599054 , n71730 , n598682 );
and ( n599055 , n599052 , n599054 );
xor ( n71733 , n598809 , n71490 );
xor ( n599057 , n71733 , n71493 );
and ( n599058 , n599054 , n599057 );
and ( n71736 , n599052 , n599057 );
or ( n71737 , n599055 , n599058 , n71736 );
and ( n599061 , n598873 , n71737 );
xor ( n599062 , n598685 , n598689 );
xor ( n71740 , n599062 , n598702 );
and ( n599064 , n71737 , n71740 );
and ( n599065 , n598873 , n71740 );
or ( n71743 , n599061 , n599064 , n599065 );
xor ( n599067 , n598631 , n598705 );
xor ( n599068 , n599067 , n71387 );
and ( n71746 , n71743 , n599068 );
xor ( n599070 , n71504 , n71506 );
xor ( n599071 , n599070 , n71509 );
and ( n71749 , n599068 , n599071 );
and ( n599073 , n71743 , n599071 );
or ( n71751 , n71746 , n71749 , n599073 );
and ( n599075 , n598847 , n71751 );
xor ( n71753 , n598847 , n71751 );
xor ( n71754 , n71743 , n599068 );
xor ( n599078 , n71754 , n599071 );
and ( n71756 , n65844 , n594807 );
and ( n599080 , n65630 , n594804 );
nor ( n71758 , n71756 , n599080 );
xnor ( n71759 , n71758 , n66187 );
xor ( n599083 , n71717 , n71721 );
xor ( n599084 , n599083 , n71726 );
and ( n71762 , n71759 , n599084 );
xor ( n599086 , n71528 , n598855 );
xor ( n599087 , n599086 , n598858 );
and ( n71765 , n599084 , n599087 );
and ( n599089 , n71759 , n599087 );
or ( n599090 , n71762 , n71765 , n599089 );
and ( n599091 , n69581 , n64862 );
and ( n71769 , n69491 , n64860 );
nor ( n599093 , n599091 , n71769 );
xnor ( n599094 , n599093 , n64764 );
and ( n71772 , n597260 , n64744 );
and ( n599096 , n69739 , n64742 );
nor ( n599097 , n71772 , n599096 );
xnor ( n71775 , n599097 , n64623 );
and ( n71776 , n599094 , n71775 );
xor ( n71777 , n598972 , n71653 );
xor ( n599101 , n71777 , n598979 );
and ( n71779 , n71775 , n599101 );
and ( n71780 , n599094 , n599101 );
or ( n71781 , n71776 , n71779 , n71780 );
and ( n71782 , n596193 , n592486 );
and ( n71783 , n596057 , n592484 );
nor ( n71784 , n71782 , n71783 );
xnor ( n599108 , n71784 , n64990 );
and ( n71786 , n71781 , n599108 );
xor ( n599110 , n71659 , n598986 );
xor ( n599111 , n599110 , n71666 );
and ( n71789 , n599108 , n599111 );
and ( n599113 , n71781 , n599111 );
or ( n71791 , n71786 , n71789 , n599113 );
and ( n71792 , n595633 , n592683 );
and ( n71793 , n595521 , n592681 );
nor ( n71794 , n71792 , n71793 );
xnor ( n599118 , n71794 , n592475 );
and ( n71796 , n71791 , n599118 );
and ( n599120 , n596057 , n592486 );
and ( n71798 , n595827 , n592484 );
nor ( n599122 , n599120 , n71798 );
xnor ( n71800 , n599122 , n64990 );
and ( n599124 , n599118 , n71800 );
and ( n599125 , n71791 , n71800 );
or ( n599126 , n71796 , n599124 , n599125 );
and ( n599127 , n67940 , n65592 );
and ( n71805 , n595103 , n592913 );
nor ( n599129 , n599127 , n71805 );
xnor ( n599130 , n599129 , n592638 );
and ( n71808 , n599126 , n599130 );
xor ( n599132 , n71675 , n71679 );
xor ( n599133 , n599132 , n599007 );
and ( n71811 , n599130 , n599133 );
and ( n71812 , n599126 , n599133 );
or ( n71813 , n71808 , n71811 , n71812 );
and ( n599137 , n594952 , n593256 );
and ( n599138 , n594710 , n593254 );
nor ( n71816 , n599137 , n599138 );
xnor ( n599140 , n71816 , n65490 );
and ( n71818 , n71813 , n599140 );
xor ( n71819 , n599010 , n71691 );
xor ( n71820 , n71819 , n71694 );
and ( n599144 , n599140 , n71820 );
and ( n71822 , n71813 , n71820 );
or ( n71823 , n71818 , n599144 , n71822 );
and ( n71824 , n66967 , n66142 );
and ( n71825 , n66951 , n66140 );
nor ( n71826 , n71824 , n71825 );
xnor ( n71827 , n71826 , n592960 );
and ( n71828 , n71823 , n71827 );
xor ( n599152 , n599020 , n71701 );
xor ( n599153 , n599152 , n71704 );
and ( n71831 , n71827 , n599153 );
and ( n71832 , n71823 , n599153 );
or ( n71833 , n71828 , n71831 , n71832 );
and ( n71834 , n66104 , n594441 );
and ( n599158 , n593437 , n67116 );
nor ( n599159 , n71834 , n599158 );
xnor ( n71837 , n599159 , n66190 );
and ( n71838 , n71833 , n71837 );
and ( n71839 , n66507 , n594210 );
and ( n71840 , n593520 , n66885 );
nor ( n71841 , n71839 , n71840 );
xnor ( n599165 , n71841 , n593434 );
and ( n599166 , n71837 , n599165 );
and ( n599167 , n71833 , n599165 );
or ( n71845 , n71838 , n599166 , n599167 );
and ( n599169 , n596198 , n592340 );
and ( n71847 , n596193 , n65015 );
nor ( n71848 , n599169 , n71847 );
xnor ( n599172 , n71848 , n64847 );
and ( n71850 , n69283 , n64862 );
and ( n599174 , n596600 , n64860 );
nor ( n71852 , n71850 , n599174 );
xnor ( n71853 , n71852 , n64764 );
and ( n599177 , n599172 , n71853 );
xor ( n71855 , n598958 , n71669 );
xor ( n599179 , n71855 , n71672 );
and ( n599180 , n71853 , n599179 );
and ( n599181 , n599172 , n599179 );
or ( n71859 , n599177 , n599180 , n599181 );
and ( n599183 , n595521 , n592683 );
and ( n599184 , n68160 , n592681 );
nor ( n71862 , n599183 , n599184 );
xnor ( n599186 , n71862 , n592475 );
and ( n599187 , n71859 , n599186 );
xor ( n599188 , n71434 , n598761 );
xor ( n71866 , n599188 , n598764 );
and ( n599190 , n599186 , n71866 );
and ( n599191 , n71859 , n71866 );
or ( n71869 , n599187 , n599190 , n599191 );
and ( n599193 , n595103 , n65592 );
and ( n599194 , n67636 , n592913 );
nor ( n71872 , n599193 , n599194 );
xnor ( n599196 , n71872 , n592638 );
and ( n71874 , n71869 , n599196 );
xor ( n599198 , n598767 , n71448 );
xor ( n71876 , n599198 , n598776 );
and ( n71877 , n599196 , n71876 );
and ( n599201 , n71869 , n71876 );
or ( n599202 , n71874 , n71877 , n599201 );
and ( n71880 , n594710 , n593256 );
and ( n599204 , n594295 , n593254 );
nor ( n599205 , n71880 , n599204 );
xnor ( n71883 , n599205 , n65490 );
and ( n599207 , n599202 , n71883 );
xor ( n599208 , n71456 , n598783 );
xor ( n71886 , n599208 , n598786 );
and ( n71887 , n71883 , n71886 );
and ( n599211 , n599202 , n71886 );
or ( n599212 , n599207 , n71887 , n599211 );
and ( n71890 , n66951 , n66142 );
and ( n599214 , n66793 , n66140 );
nor ( n599215 , n71890 , n599214 );
xnor ( n71893 , n599215 , n592960 );
and ( n599217 , n599212 , n71893 );
xor ( n71895 , n71466 , n71470 );
xor ( n599219 , n71895 , n71473 );
and ( n71897 , n71893 , n599219 );
and ( n599221 , n599212 , n599219 );
or ( n71899 , n599217 , n71897 , n599221 );
and ( n71900 , n71845 , n71899 );
xor ( n599224 , n71476 , n71480 );
xor ( n71902 , n599224 , n71483 );
and ( n599226 , n71899 , n71902 );
and ( n71904 , n71845 , n71902 );
or ( n599228 , n71900 , n599226 , n71904 );
and ( n599229 , n599090 , n599228 );
xor ( n71907 , n598861 , n598865 );
xor ( n71908 , n71907 , n71547 );
and ( n599232 , n599228 , n71908 );
and ( n599233 , n599090 , n71908 );
or ( n71911 , n599229 , n599232 , n599233 );
xor ( n599235 , n598819 , n598821 );
xor ( n599236 , n599235 , n598824 );
and ( n71914 , n71911 , n599236 );
xor ( n599238 , n598873 , n71737 );
xor ( n599239 , n599238 , n71740 );
and ( n599240 , n599236 , n599239 );
and ( n71918 , n71911 , n599239 );
or ( n599242 , n71914 , n599240 , n71918 );
and ( n599243 , n599078 , n599242 );
xor ( n71921 , n599078 , n599242 );
xor ( n599245 , n598877 , n71558 );
and ( n71923 , n70652 , n64648 );
not ( n599247 , n71923 );
and ( n71925 , n599247 , n591902 );
and ( n599249 , n70652 , n64650 );
and ( n599250 , n597980 , n64648 );
nor ( n71928 , n599249 , n599250 );
xnor ( n71929 , n71928 , n591902 );
and ( n71930 , n71925 , n71929 );
and ( n71931 , n597980 , n64650 );
and ( n599255 , n70663 , n64648 );
nor ( n599256 , n71931 , n599255 );
xnor ( n71934 , n599256 , n591902 );
and ( n599258 , n71930 , n71934 );
and ( n71936 , n71934 , n71552 );
and ( n71937 , n71930 , n71552 );
or ( n599261 , n599258 , n71936 , n71937 );
and ( n599262 , n599245 , n599261 );
and ( n71940 , n70663 , n64650 );
and ( n599264 , n597996 , n64648 );
nor ( n599265 , n71940 , n599264 );
xnor ( n71943 , n599265 , n591902 );
and ( n599267 , n599261 , n71943 );
and ( n599268 , n599245 , n71943 );
or ( n71946 , n599262 , n599267 , n599268 );
and ( n599270 , n597996 , n64650 );
and ( n71948 , n70683 , n64648 );
nor ( n599272 , n599270 , n71948 );
xnor ( n599273 , n599272 , n591902 );
and ( n599274 , n71946 , n599273 );
xor ( n71952 , n598882 , n71563 );
xor ( n599276 , n71952 , n71130 );
and ( n71954 , n599273 , n599276 );
and ( n599278 , n71946 , n599276 );
or ( n599279 , n599274 , n71954 , n599278 );
and ( n71957 , n70683 , n64650 );
and ( n599281 , n70693 , n64648 );
nor ( n599282 , n71957 , n599281 );
xnor ( n71960 , n599282 , n591902 );
and ( n599284 , n599279 , n71960 );
xor ( n71962 , n598874 , n71567 );
xor ( n599286 , n71962 , n598895 );
and ( n71964 , n71960 , n599286 );
and ( n599288 , n599279 , n599286 );
or ( n71966 , n599284 , n71964 , n599288 );
and ( n71967 , n70693 , n64650 );
and ( n599291 , n70637 , n64648 );
nor ( n599292 , n71967 , n599291 );
xnor ( n71970 , n599292 , n591902 );
and ( n599294 , n71966 , n71970 );
xor ( n599295 , n71575 , n71579 );
xor ( n71973 , n599295 , n598905 );
and ( n599297 , n71970 , n71973 );
and ( n599298 , n71966 , n71973 );
or ( n71976 , n599294 , n599297 , n599298 );
and ( n71977 , n70637 , n64650 );
and ( n599301 , n70261 , n64648 );
nor ( n599302 , n71977 , n599301 );
xnor ( n71980 , n599302 , n591902 );
and ( n599304 , n71976 , n71980 );
xor ( n599305 , n71585 , n71589 );
xor ( n71983 , n599305 , n71592 );
and ( n599307 , n71980 , n71983 );
and ( n599308 , n71976 , n71983 );
or ( n71986 , n599304 , n599307 , n599308 );
and ( n599310 , n70261 , n64650 );
and ( n599311 , n70255 , n64648 );
nor ( n71989 , n599310 , n599311 );
xnor ( n599313 , n71989 , n591902 );
and ( n71991 , n71986 , n599313 );
xor ( n599315 , n71595 , n71599 );
xor ( n71993 , n599315 , n71602 );
and ( n599317 , n599313 , n71993 );
and ( n71995 , n71986 , n71993 );
or ( n71996 , n71991 , n599317 , n71995 );
and ( n599320 , n69739 , n64862 );
and ( n599321 , n69581 , n64860 );
nor ( n71999 , n599320 , n599321 );
xnor ( n599323 , n71999 , n64764 );
and ( n599324 , n71996 , n599323 );
xor ( n72002 , n71639 , n71643 );
xor ( n599326 , n72002 , n598969 );
and ( n599327 , n599323 , n599326 );
and ( n72005 , n71996 , n599326 );
or ( n72006 , n599324 , n599327 , n72005 );
and ( n599330 , n69283 , n592340 );
and ( n599331 , n596600 , n65015 );
nor ( n72009 , n599330 , n599331 );
xnor ( n599333 , n72009 , n64847 );
and ( n599334 , n72006 , n599333 );
xor ( n72012 , n599094 , n71775 );
xor ( n599336 , n72012 , n599101 );
and ( n599337 , n599333 , n599336 );
and ( n72015 , n72006 , n599336 );
or ( n599339 , n599334 , n599337 , n72015 );
and ( n599340 , n595827 , n592683 );
and ( n72018 , n595633 , n592681 );
nor ( n72019 , n599340 , n72018 );
xnor ( n599343 , n72019 , n592475 );
and ( n72021 , n599339 , n599343 );
and ( n599345 , n596600 , n592340 );
and ( n599346 , n596198 , n65015 );
nor ( n599347 , n599345 , n599346 );
xnor ( n72025 , n599347 , n64847 );
and ( n599349 , n599343 , n72025 );
and ( n599350 , n599339 , n72025 );
or ( n72028 , n72021 , n599349 , n599350 );
and ( n599352 , n595103 , n593256 );
and ( n599353 , n67636 , n593254 );
nor ( n72031 , n599352 , n599353 );
xnor ( n72032 , n72031 , n65490 );
and ( n72033 , n72028 , n72032 );
xor ( n72034 , n599172 , n71853 );
xor ( n599358 , n72034 , n599179 );
and ( n599359 , n72032 , n599358 );
and ( n72037 , n72028 , n599358 );
or ( n599361 , n72033 , n599359 , n72037 );
and ( n599362 , n67636 , n593256 );
and ( n72040 , n594952 , n593254 );
nor ( n599364 , n599362 , n72040 );
xnor ( n72042 , n599364 , n65490 );
and ( n599366 , n599361 , n72042 );
xor ( n72044 , n71859 , n599186 );
xor ( n72045 , n72044 , n71866 );
and ( n599369 , n72042 , n72045 );
and ( n72047 , n599361 , n72045 );
or ( n599371 , n599366 , n599369 , n72047 );
and ( n72049 , n594295 , n66142 );
and ( n72050 , n66967 , n66140 );
nor ( n599374 , n72049 , n72050 );
xnor ( n599375 , n599374 , n592960 );
and ( n72053 , n599371 , n599375 );
xor ( n599377 , n71869 , n599196 );
xor ( n599378 , n599377 , n71876 );
and ( n72056 , n599375 , n599378 );
and ( n599380 , n599371 , n599378 );
or ( n599381 , n72053 , n72056 , n599380 );
and ( n599382 , n593437 , n594807 );
and ( n72060 , n593298 , n594804 );
nor ( n599384 , n599382 , n72060 );
xnor ( n599385 , n599384 , n66187 );
and ( n72063 , n599381 , n599385 );
and ( n599387 , n66793 , n66457 );
and ( n599388 , n594124 , n593778 );
nor ( n72066 , n599387 , n599388 );
xnor ( n72067 , n72066 , n593160 );
and ( n72068 , n599385 , n72067 );
and ( n72069 , n599381 , n72067 );
or ( n599393 , n72063 , n72068 , n72069 );
and ( n599394 , n593520 , n594441 );
and ( n72072 , n66104 , n67116 );
nor ( n599396 , n599394 , n72072 );
xnor ( n72074 , n599396 , n66190 );
and ( n599398 , n66606 , n594210 );
and ( n599399 , n66507 , n66885 );
nor ( n599400 , n599398 , n599399 );
xnor ( n72078 , n599400 , n593434 );
and ( n599402 , n72074 , n72078 );
xor ( n72080 , n599202 , n71883 );
xor ( n72081 , n72080 , n71886 );
and ( n599405 , n72078 , n72081 );
and ( n72083 , n72074 , n72081 );
or ( n599407 , n599402 , n599405 , n72083 );
and ( n72085 , n599393 , n599407 );
and ( n72086 , n593298 , n594807 );
and ( n599410 , n65844 , n594804 );
nor ( n72088 , n72086 , n599410 );
xnor ( n599412 , n72088 , n66187 );
and ( n599413 , n599407 , n599412 );
and ( n599414 , n599393 , n599412 );
or ( n72092 , n72085 , n599413 , n599414 );
and ( n599416 , n594124 , n66457 );
and ( n599417 , n66606 , n593778 );
nor ( n72095 , n599416 , n599417 );
xnor ( n599419 , n72095 , n593160 );
xor ( n599420 , n71707 , n599034 );
xor ( n599421 , n599420 , n71714 );
and ( n72099 , n599419 , n599421 );
xor ( n599423 , n599212 , n71893 );
xor ( n599424 , n599423 , n599219 );
and ( n72102 , n599421 , n599424 );
and ( n599426 , n599419 , n599424 );
or ( n599427 , n72099 , n72102 , n599426 );
and ( n72105 , n72092 , n599427 );
xor ( n599429 , n71845 , n71899 );
xor ( n72107 , n599429 , n71902 );
and ( n599431 , n599427 , n72107 );
and ( n72109 , n72092 , n72107 );
or ( n72110 , n72105 , n599431 , n72109 );
xor ( n599434 , n599090 , n599228 );
xor ( n72112 , n599434 , n71908 );
and ( n72113 , n72110 , n72112 );
xor ( n599437 , n599052 , n599054 );
xor ( n72115 , n599437 , n599057 );
and ( n72116 , n72112 , n72115 );
and ( n72117 , n72110 , n72115 );
or ( n599441 , n72113 , n72116 , n72117 );
xor ( n72119 , n71911 , n599236 );
xor ( n72120 , n72119 , n599239 );
and ( n599444 , n599441 , n72120 );
xor ( n599445 , n599441 , n72120 );
xor ( n599446 , n72110 , n72112 );
xor ( n72124 , n599446 , n72115 );
and ( n599448 , n66507 , n594441 );
and ( n599449 , n593520 , n67116 );
nor ( n72127 , n599448 , n599449 );
xnor ( n599451 , n72127 , n66190 );
and ( n599452 , n594124 , n594210 );
and ( n72130 , n66606 , n66885 );
nor ( n599454 , n599452 , n72130 );
xnor ( n599455 , n599454 , n593434 );
and ( n72133 , n599451 , n599455 );
xor ( n599457 , n599371 , n599375 );
xor ( n599458 , n599457 , n599378 );
and ( n599459 , n599455 , n599458 );
and ( n72137 , n599451 , n599458 );
or ( n599461 , n72133 , n599459 , n72137 );
and ( n72139 , n597402 , n64862 );
and ( n72140 , n597260 , n64860 );
nor ( n599464 , n72139 , n72140 );
xnor ( n599465 , n599464 , n64764 );
and ( n72143 , n70255 , n64744 );
and ( n599467 , n597569 , n64742 );
nor ( n72145 , n72143 , n599467 );
xnor ( n599469 , n72145 , n64623 );
and ( n599470 , n599465 , n599469 );
xor ( n72148 , n71976 , n71980 );
xor ( n599472 , n72148 , n71983 );
and ( n599473 , n599469 , n599472 );
and ( n72151 , n599465 , n599472 );
or ( n72152 , n599470 , n599473 , n72151 );
and ( n72153 , n597569 , n64744 );
and ( n72154 , n597402 , n64742 );
nor ( n599478 , n72153 , n72154 );
xnor ( n599479 , n599478 , n64623 );
and ( n72157 , n72152 , n599479 );
xor ( n599481 , n71986 , n599313 );
xor ( n72159 , n599481 , n71993 );
and ( n72160 , n599479 , n72159 );
and ( n599484 , n72152 , n72159 );
or ( n72162 , n72157 , n72160 , n599484 );
and ( n599486 , n69491 , n592340 );
and ( n599487 , n69283 , n65015 );
nor ( n72165 , n599486 , n599487 );
xnor ( n72166 , n72165 , n64847 );
and ( n72167 , n72162 , n72166 );
xor ( n72168 , n71996 , n599323 );
xor ( n72169 , n72168 , n599326 );
and ( n72170 , n72166 , n72169 );
and ( n72171 , n72162 , n72169 );
or ( n599495 , n72167 , n72170 , n72171 );
and ( n72173 , n596198 , n592486 );
and ( n72174 , n596193 , n592484 );
nor ( n72175 , n72173 , n72174 );
xnor ( n72176 , n72175 , n64990 );
and ( n599500 , n599495 , n72176 );
xor ( n599501 , n72006 , n599333 );
xor ( n72179 , n599501 , n599336 );
and ( n599503 , n72176 , n72179 );
and ( n72181 , n599495 , n72179 );
or ( n599505 , n599500 , n599503 , n72181 );
and ( n599506 , n595521 , n65592 );
and ( n72184 , n68160 , n592913 );
nor ( n599508 , n599506 , n72184 );
xnor ( n72186 , n599508 , n592638 );
and ( n599510 , n599505 , n72186 );
xor ( n72188 , n71781 , n599108 );
xor ( n599512 , n72188 , n599111 );
and ( n599513 , n72186 , n599512 );
and ( n72191 , n599505 , n599512 );
or ( n599515 , n599510 , n599513 , n72191 );
and ( n599516 , n68160 , n65592 );
and ( n72194 , n67940 , n592913 );
nor ( n599518 , n599516 , n72194 );
xnor ( n599519 , n599518 , n592638 );
and ( n72197 , n599515 , n599519 );
xor ( n599521 , n71791 , n599118 );
xor ( n599522 , n599521 , n71800 );
and ( n72200 , n599519 , n599522 );
and ( n599524 , n599515 , n599522 );
or ( n72202 , n72197 , n72200 , n599524 );
and ( n72203 , n594710 , n66142 );
and ( n72204 , n594295 , n66140 );
nor ( n72205 , n72203 , n72204 );
xnor ( n599529 , n72205 , n592960 );
and ( n72207 , n72202 , n599529 );
xor ( n72208 , n599126 , n599130 );
xor ( n72209 , n72208 , n599133 );
and ( n72210 , n599529 , n72209 );
and ( n72211 , n72202 , n72209 );
or ( n72212 , n72207 , n72210 , n72211 );
and ( n72213 , n66951 , n66457 );
and ( n72214 , n66793 , n593778 );
nor ( n72215 , n72213 , n72214 );
xnor ( n72216 , n72215 , n593160 );
and ( n599540 , n72212 , n72216 );
xor ( n599541 , n71813 , n599140 );
xor ( n72219 , n599541 , n71820 );
and ( n599543 , n72216 , n72219 );
and ( n599544 , n72212 , n72219 );
or ( n72222 , n599540 , n599543 , n599544 );
and ( n72223 , n599461 , n72222 );
xor ( n72224 , n71823 , n71827 );
xor ( n72225 , n72224 , n599153 );
and ( n72226 , n72222 , n72225 );
and ( n599550 , n599461 , n72225 );
or ( n599551 , n72223 , n72226 , n599550 );
xor ( n72229 , n71833 , n71837 );
xor ( n72230 , n72229 , n599165 );
and ( n72231 , n599551 , n72230 );
xor ( n72232 , n599419 , n599421 );
xor ( n72233 , n72232 , n599424 );
and ( n599557 , n72230 , n72233 );
and ( n72235 , n599551 , n72233 );
or ( n599559 , n72231 , n599557 , n72235 );
xor ( n599560 , n71759 , n599084 );
xor ( n599561 , n599560 , n599087 );
and ( n72239 , n599559 , n599561 );
xor ( n599563 , n72092 , n599427 );
xor ( n72241 , n599563 , n72107 );
and ( n72242 , n599561 , n72241 );
and ( n599566 , n599559 , n72241 );
or ( n72244 , n72239 , n72242 , n599566 );
and ( n599568 , n72124 , n72244 );
xor ( n599569 , n72124 , n72244 );
xor ( n72247 , n599559 , n599561 );
xor ( n599571 , n72247 , n72241 );
and ( n599572 , n69581 , n592340 );
and ( n72250 , n69491 , n65015 );
nor ( n72251 , n599572 , n72250 );
xnor ( n599575 , n72251 , n64847 );
and ( n599576 , n597260 , n64862 );
and ( n72254 , n69739 , n64860 );
nor ( n599578 , n599576 , n72254 );
xnor ( n599579 , n599578 , n64764 );
and ( n72257 , n599575 , n599579 );
xor ( n599581 , n72152 , n599479 );
xor ( n599582 , n599581 , n72159 );
and ( n599583 , n599579 , n599582 );
and ( n72261 , n599575 , n599582 );
or ( n599585 , n72257 , n599583 , n72261 );
and ( n72263 , n596600 , n592486 );
and ( n599587 , n596198 , n592484 );
nor ( n72265 , n72263 , n599587 );
xnor ( n599589 , n72265 , n64990 );
and ( n599590 , n599585 , n599589 );
xor ( n72268 , n72162 , n72166 );
xor ( n72269 , n72268 , n72169 );
and ( n599593 , n599589 , n72269 );
and ( n599594 , n599585 , n72269 );
or ( n72272 , n599590 , n599593 , n599594 );
and ( n599596 , n595633 , n65592 );
and ( n599597 , n595521 , n592913 );
nor ( n72275 , n599596 , n599597 );
xnor ( n599599 , n72275 , n592638 );
and ( n599600 , n72272 , n599599 );
and ( n72278 , n596057 , n592683 );
and ( n72279 , n595827 , n592681 );
nor ( n599603 , n72278 , n72279 );
xnor ( n599604 , n599603 , n592475 );
and ( n72282 , n599599 , n599604 );
and ( n599606 , n72272 , n599604 );
or ( n599607 , n599600 , n72282 , n599606 );
and ( n72285 , n67940 , n593256 );
and ( n599609 , n595103 , n593254 );
nor ( n599610 , n72285 , n599609 );
xnor ( n72288 , n599610 , n65490 );
and ( n599612 , n599607 , n72288 );
xor ( n599613 , n599339 , n599343 );
xor ( n72291 , n599613 , n72025 );
and ( n599615 , n72288 , n72291 );
and ( n72293 , n599607 , n72291 );
or ( n599617 , n599612 , n599615 , n72293 );
and ( n599618 , n594952 , n66142 );
and ( n599619 , n594710 , n66140 );
nor ( n72297 , n599618 , n599619 );
xnor ( n599621 , n72297 , n592960 );
and ( n599622 , n599617 , n599621 );
xor ( n72300 , n72028 , n72032 );
xor ( n599624 , n72300 , n599358 );
and ( n599625 , n599621 , n599624 );
and ( n72303 , n599617 , n599624 );
or ( n599627 , n599622 , n599625 , n72303 );
and ( n599628 , n66967 , n66457 );
and ( n72306 , n66951 , n593778 );
nor ( n599630 , n599628 , n72306 );
xnor ( n72308 , n599630 , n593160 );
and ( n599632 , n599627 , n72308 );
xor ( n599633 , n599361 , n72042 );
xor ( n72311 , n599633 , n72045 );
and ( n599635 , n72308 , n72311 );
and ( n599636 , n599627 , n72311 );
or ( n599637 , n599632 , n599635 , n599636 );
and ( n72315 , n66104 , n594807 );
and ( n599639 , n593437 , n594804 );
nor ( n72317 , n72315 , n599639 );
xnor ( n72318 , n72317 , n66187 );
and ( n599642 , n599637 , n72318 );
xor ( n72320 , n72212 , n72216 );
xor ( n599644 , n72320 , n72219 );
and ( n72322 , n72318 , n599644 );
and ( n72323 , n599637 , n599644 );
or ( n72324 , n599642 , n72322 , n72323 );
xor ( n72325 , n599381 , n599385 );
xor ( n599649 , n72325 , n72067 );
and ( n72327 , n72324 , n599649 );
xor ( n599651 , n72074 , n72078 );
xor ( n599652 , n599651 , n72081 );
and ( n599653 , n599649 , n599652 );
and ( n72331 , n72324 , n599652 );
or ( n599655 , n72327 , n599653 , n72331 );
xor ( n599656 , n599393 , n599407 );
xor ( n72334 , n599656 , n599412 );
and ( n599658 , n599655 , n72334 );
xor ( n599659 , n599551 , n72230 );
xor ( n72337 , n599659 , n72233 );
and ( n599661 , n72334 , n72337 );
and ( n72339 , n599655 , n72337 );
or ( n599663 , n599658 , n599661 , n72339 );
and ( n72341 , n599571 , n599663 );
xor ( n72342 , n599571 , n599663 );
xor ( n599666 , n599655 , n72334 );
xor ( n599667 , n599666 , n72337 );
xor ( n72345 , n71925 , n71929 );
and ( n72346 , n70652 , n64742 );
not ( n599670 , n72346 );
and ( n72348 , n599670 , n64623 );
and ( n72349 , n70652 , n64744 );
and ( n599673 , n597980 , n64742 );
nor ( n599674 , n72349 , n599673 );
xnor ( n599675 , n599674 , n64623 );
and ( n72353 , n72348 , n599675 );
and ( n599677 , n597980 , n64744 );
and ( n599678 , n70663 , n64742 );
nor ( n72356 , n599677 , n599678 );
xnor ( n599680 , n72356 , n64623 );
and ( n599681 , n72353 , n599680 );
and ( n72359 , n599680 , n71923 );
and ( n599683 , n72353 , n71923 );
or ( n599684 , n599681 , n72359 , n599683 );
and ( n72362 , n72345 , n599684 );
and ( n599686 , n70663 , n64744 );
and ( n72364 , n597996 , n64742 );
nor ( n599688 , n599686 , n72364 );
xnor ( n72366 , n599688 , n64623 );
and ( n599690 , n599684 , n72366 );
and ( n599691 , n72345 , n72366 );
or ( n72369 , n72362 , n599690 , n599691 );
and ( n599693 , n597996 , n64744 );
and ( n599694 , n70683 , n64742 );
nor ( n599695 , n599693 , n599694 );
xnor ( n72373 , n599695 , n64623 );
and ( n599697 , n72369 , n72373 );
xor ( n72375 , n71930 , n71934 );
xor ( n72376 , n72375 , n71552 );
and ( n72377 , n72373 , n72376 );
and ( n72378 , n72369 , n72376 );
or ( n72379 , n599697 , n72377 , n72378 );
and ( n72380 , n70683 , n64744 );
and ( n72381 , n70693 , n64742 );
nor ( n599705 , n72380 , n72381 );
xnor ( n599706 , n599705 , n64623 );
and ( n599707 , n72379 , n599706 );
xor ( n72385 , n599245 , n599261 );
xor ( n72386 , n72385 , n71943 );
and ( n72387 , n599706 , n72386 );
and ( n72388 , n72379 , n72386 );
or ( n72389 , n599707 , n72387 , n72388 );
and ( n599713 , n70693 , n64744 );
and ( n72391 , n70637 , n64742 );
nor ( n72392 , n599713 , n72391 );
xnor ( n599716 , n72392 , n64623 );
and ( n599717 , n72389 , n599716 );
xor ( n72395 , n71946 , n599273 );
xor ( n599719 , n72395 , n599276 );
and ( n599720 , n599716 , n599719 );
and ( n72398 , n72389 , n599719 );
or ( n599722 , n599717 , n599720 , n72398 );
and ( n599723 , n70637 , n64744 );
and ( n72401 , n70261 , n64742 );
nor ( n72402 , n599723 , n72401 );
xnor ( n72403 , n72402 , n64623 );
and ( n72404 , n599722 , n72403 );
xor ( n72405 , n599279 , n71960 );
xor ( n599729 , n72405 , n599286 );
and ( n599730 , n72403 , n599729 );
and ( n72408 , n599722 , n599729 );
or ( n72409 , n72404 , n599730 , n72408 );
and ( n72410 , n70261 , n64744 );
and ( n599734 , n70255 , n64742 );
nor ( n599735 , n72410 , n599734 );
xnor ( n599736 , n599735 , n64623 );
and ( n72414 , n72409 , n599736 );
xor ( n599738 , n71966 , n71970 );
xor ( n72416 , n599738 , n71973 );
and ( n72417 , n599736 , n72416 );
and ( n599741 , n72409 , n72416 );
or ( n72419 , n72414 , n72417 , n599741 );
and ( n599743 , n69739 , n592340 );
and ( n72421 , n69581 , n65015 );
nor ( n72422 , n599743 , n72421 );
xnor ( n599746 , n72422 , n64847 );
and ( n72424 , n72419 , n599746 );
xor ( n599748 , n599465 , n599469 );
xor ( n599749 , n599748 , n599472 );
and ( n72427 , n599746 , n599749 );
and ( n599751 , n72419 , n599749 );
or ( n599752 , n72424 , n72427 , n599751 );
and ( n72430 , n69283 , n592486 );
and ( n599754 , n596600 , n592484 );
nor ( n72432 , n72430 , n599754 );
xnor ( n599756 , n72432 , n64990 );
and ( n599757 , n599752 , n599756 );
xor ( n72435 , n599575 , n599579 );
xor ( n599759 , n72435 , n599582 );
and ( n72437 , n599756 , n599759 );
and ( n599761 , n599752 , n599759 );
or ( n599762 , n599757 , n72437 , n599761 );
and ( n72440 , n595827 , n65592 );
and ( n72441 , n595633 , n592913 );
nor ( n599765 , n72440 , n72441 );
xnor ( n72443 , n599765 , n592638 );
and ( n599767 , n599762 , n72443 );
and ( n599768 , n596193 , n592683 );
and ( n599769 , n596057 , n592681 );
nor ( n72447 , n599768 , n599769 );
xnor ( n599771 , n72447 , n592475 );
and ( n72449 , n72443 , n599771 );
and ( n599773 , n599762 , n599771 );
or ( n599774 , n599767 , n72449 , n599773 );
xor ( n72452 , n72272 , n599599 );
xor ( n599776 , n72452 , n599604 );
and ( n599777 , n599774 , n599776 );
xor ( n599778 , n599495 , n72176 );
xor ( n72456 , n599778 , n72179 );
and ( n599780 , n599776 , n72456 );
and ( n72458 , n599774 , n72456 );
or ( n599782 , n599777 , n599780 , n72458 );
and ( n599783 , n67636 , n66142 );
and ( n72461 , n594952 , n66140 );
nor ( n72462 , n599783 , n72461 );
xnor ( n599786 , n72462 , n592960 );
and ( n72464 , n599782 , n599786 );
xor ( n599788 , n599505 , n72186 );
xor ( n599789 , n599788 , n599512 );
and ( n599790 , n599786 , n599789 );
and ( n72468 , n599782 , n599789 );
or ( n599792 , n72464 , n599790 , n72468 );
and ( n72470 , n594295 , n66457 );
and ( n599794 , n66967 , n593778 );
nor ( n599795 , n72470 , n599794 );
xnor ( n72473 , n599795 , n593160 );
and ( n599797 , n599792 , n72473 );
xor ( n599798 , n599515 , n599519 );
xor ( n72476 , n599798 , n599522 );
and ( n599800 , n72473 , n72476 );
and ( n72478 , n599792 , n72476 );
or ( n599802 , n599797 , n599800 , n72478 );
and ( n72480 , n66793 , n594210 );
and ( n72481 , n594124 , n66885 );
nor ( n599805 , n72480 , n72481 );
xnor ( n72483 , n599805 , n593434 );
and ( n599807 , n599802 , n72483 );
xor ( n72485 , n72202 , n599529 );
xor ( n72486 , n72485 , n72209 );
and ( n599810 , n72483 , n72486 );
and ( n72488 , n599802 , n72486 );
or ( n599812 , n599807 , n599810 , n72488 );
and ( n72490 , n593520 , n594807 );
and ( n599814 , n66104 , n594804 );
nor ( n599815 , n72490 , n599814 );
xnor ( n72493 , n599815 , n66187 );
and ( n599817 , n66606 , n594441 );
and ( n599818 , n66507 , n67116 );
nor ( n599819 , n599817 , n599818 );
xnor ( n72497 , n599819 , n66190 );
and ( n599821 , n72493 , n72497 );
xor ( n599822 , n599627 , n72308 );
xor ( n72500 , n599822 , n72311 );
and ( n599824 , n72497 , n72500 );
and ( n72502 , n72493 , n72500 );
or ( n72503 , n599821 , n599824 , n72502 );
and ( n72504 , n599812 , n72503 );
xor ( n72505 , n599451 , n599455 );
xor ( n72506 , n72505 , n599458 );
and ( n599830 , n72503 , n72506 );
and ( n72508 , n599812 , n72506 );
or ( n599832 , n72504 , n599830 , n72508 );
xor ( n72510 , n72324 , n599649 );
xor ( n72511 , n72510 , n599652 );
and ( n599835 , n599832 , n72511 );
xor ( n599836 , n599461 , n72222 );
xor ( n72514 , n599836 , n72225 );
and ( n72515 , n72511 , n72514 );
and ( n599839 , n599832 , n72514 );
or ( n72517 , n599835 , n72515 , n599839 );
and ( n72518 , n599667 , n72517 );
xor ( n72519 , n599667 , n72517 );
and ( n599843 , n66507 , n594807 );
and ( n72521 , n593520 , n594804 );
nor ( n599845 , n599843 , n72521 );
xnor ( n599846 , n599845 , n66187 );
and ( n72524 , n594124 , n594441 );
and ( n599848 , n66606 , n67116 );
nor ( n72526 , n72524 , n599848 );
xnor ( n72527 , n72526 , n66190 );
and ( n599851 , n599846 , n72527 );
xor ( n72529 , n599792 , n72473 );
xor ( n599853 , n72529 , n72476 );
and ( n72531 , n72527 , n599853 );
and ( n72532 , n599846 , n599853 );
or ( n599856 , n599851 , n72531 , n72532 );
and ( n599857 , n597402 , n592340 );
and ( n72535 , n597260 , n65015 );
nor ( n599859 , n599857 , n72535 );
xnor ( n72537 , n599859 , n64847 );
and ( n599861 , n70255 , n64862 );
and ( n599862 , n597569 , n64860 );
nor ( n72540 , n599861 , n599862 );
xnor ( n599864 , n72540 , n64764 );
and ( n599865 , n72537 , n599864 );
xor ( n599866 , n599722 , n72403 );
xor ( n72544 , n599866 , n599729 );
and ( n599868 , n599864 , n72544 );
and ( n72546 , n72537 , n72544 );
or ( n72547 , n599865 , n599868 , n72546 );
and ( n599871 , n597569 , n64862 );
and ( n72549 , n597402 , n64860 );
nor ( n599873 , n599871 , n72549 );
xnor ( n72551 , n599873 , n64764 );
and ( n72552 , n72547 , n72551 );
xor ( n599876 , n72409 , n599736 );
xor ( n72554 , n599876 , n72416 );
and ( n599878 , n72551 , n72554 );
and ( n599879 , n72547 , n72554 );
or ( n599880 , n72552 , n599878 , n599879 );
and ( n72558 , n69491 , n592486 );
and ( n599882 , n69283 , n592484 );
nor ( n599883 , n72558 , n599882 );
xnor ( n72561 , n599883 , n64990 );
and ( n599885 , n599880 , n72561 );
xor ( n599886 , n72419 , n599746 );
xor ( n599887 , n599886 , n599749 );
and ( n72565 , n72561 , n599887 );
and ( n599889 , n599880 , n599887 );
or ( n599890 , n599885 , n72565 , n599889 );
and ( n72568 , n596198 , n592683 );
and ( n599892 , n596193 , n592681 );
nor ( n599893 , n72568 , n599892 );
xnor ( n599894 , n599893 , n592475 );
and ( n72572 , n599890 , n599894 );
xor ( n599896 , n599752 , n599756 );
xor ( n72574 , n599896 , n599759 );
and ( n599898 , n599894 , n72574 );
and ( n72576 , n599890 , n72574 );
or ( n72577 , n72572 , n599898 , n72576 );
and ( n599901 , n595521 , n593256 );
and ( n72579 , n68160 , n593254 );
nor ( n599903 , n599901 , n72579 );
xnor ( n599904 , n599903 , n65490 );
and ( n599905 , n72577 , n599904 );
xor ( n72583 , n599585 , n599589 );
xor ( n599907 , n72583 , n72269 );
and ( n599908 , n599904 , n599907 );
and ( n72586 , n72577 , n599907 );
or ( n599910 , n599905 , n599908 , n72586 );
and ( n599911 , n595103 , n66142 );
and ( n72589 , n67636 , n66140 );
nor ( n72590 , n599911 , n72589 );
xnor ( n599914 , n72590 , n592960 );
and ( n599915 , n599910 , n599914 );
and ( n72593 , n68160 , n593256 );
and ( n599917 , n67940 , n593254 );
nor ( n599918 , n72593 , n599917 );
xnor ( n72596 , n599918 , n65490 );
and ( n599920 , n599914 , n72596 );
and ( n599921 , n599910 , n72596 );
or ( n72599 , n599915 , n599920 , n599921 );
and ( n599923 , n594710 , n66457 );
and ( n72601 , n594295 , n593778 );
nor ( n599925 , n599923 , n72601 );
xnor ( n72603 , n599925 , n593160 );
and ( n72604 , n72599 , n72603 );
xor ( n599928 , n599607 , n72288 );
xor ( n72606 , n599928 , n72291 );
and ( n599930 , n72603 , n72606 );
and ( n72608 , n72599 , n72606 );
or ( n599932 , n72604 , n599930 , n72608 );
and ( n599933 , n66951 , n594210 );
and ( n72611 , n66793 , n66885 );
nor ( n72612 , n599933 , n72611 );
xnor ( n599936 , n72612 , n593434 );
and ( n599937 , n599932 , n599936 );
xor ( n72615 , n599617 , n599621 );
xor ( n599939 , n72615 , n599624 );
and ( n599940 , n599936 , n599939 );
and ( n72618 , n599932 , n599939 );
or ( n599942 , n599937 , n599940 , n72618 );
and ( n599943 , n599856 , n599942 );
xor ( n599944 , n599802 , n72483 );
xor ( n72622 , n599944 , n72486 );
and ( n599946 , n599942 , n72622 );
and ( n599947 , n599856 , n72622 );
or ( n72625 , n599943 , n599946 , n599947 );
xor ( n599949 , n599812 , n72503 );
xor ( n599950 , n599949 , n72506 );
and ( n72628 , n72625 , n599950 );
xor ( n599952 , n599637 , n72318 );
xor ( n599953 , n599952 , n599644 );
and ( n72631 , n599950 , n599953 );
and ( n72632 , n72625 , n599953 );
or ( n72633 , n72628 , n72631 , n72632 );
xor ( n599957 , n599832 , n72511 );
xor ( n599958 , n599957 , n72514 );
and ( n72636 , n72633 , n599958 );
xor ( n72637 , n72633 , n599958 );
xor ( n72638 , n72625 , n599950 );
xor ( n599962 , n72638 , n599953 );
and ( n599963 , n66606 , n594807 );
and ( n72641 , n66507 , n594804 );
nor ( n72642 , n599963 , n72641 );
xnor ( n72643 , n72642 , n66187 );
and ( n72644 , n66793 , n594441 );
and ( n599968 , n594124 , n67116 );
nor ( n599969 , n72644 , n599968 );
xnor ( n599970 , n599969 , n66190 );
and ( n72648 , n72643 , n599970 );
xor ( n599972 , n72599 , n72603 );
xor ( n72650 , n599972 , n72606 );
and ( n72651 , n599970 , n72650 );
and ( n599975 , n72643 , n72650 );
or ( n599976 , n72648 , n72651 , n599975 );
and ( n72654 , n69581 , n592486 );
and ( n72655 , n69491 , n592484 );
nor ( n599979 , n72654 , n72655 );
xnor ( n72657 , n599979 , n64990 );
and ( n72658 , n597260 , n592340 );
and ( n599982 , n69739 , n65015 );
nor ( n599983 , n72658 , n599982 );
xnor ( n599984 , n599983 , n64847 );
and ( n72662 , n72657 , n599984 );
xor ( n599986 , n72547 , n72551 );
xor ( n599987 , n599986 , n72554 );
and ( n72665 , n599984 , n599987 );
and ( n599989 , n72657 , n599987 );
or ( n599990 , n72662 , n72665 , n599989 );
and ( n599991 , n596193 , n65592 );
and ( n72669 , n596057 , n592913 );
nor ( n599993 , n599991 , n72669 );
xnor ( n72671 , n599993 , n592638 );
and ( n72672 , n599990 , n72671 );
xor ( n599996 , n599880 , n72561 );
xor ( n72674 , n599996 , n599887 );
and ( n599998 , n72671 , n72674 );
and ( n72676 , n599990 , n72674 );
or ( n72677 , n72672 , n599998 , n72676 );
and ( n600001 , n596057 , n65592 );
and ( n600002 , n595827 , n592913 );
nor ( n72680 , n600001 , n600002 );
xnor ( n600004 , n72680 , n592638 );
and ( n600005 , n72677 , n600004 );
xor ( n72683 , n599890 , n599894 );
xor ( n600007 , n72683 , n72574 );
and ( n600008 , n600004 , n600007 );
and ( n600009 , n72677 , n600007 );
or ( n72687 , n600005 , n600008 , n600009 );
and ( n600011 , n67940 , n66142 );
and ( n600012 , n595103 , n66140 );
nor ( n72690 , n600011 , n600012 );
xnor ( n600014 , n72690 , n592960 );
and ( n600015 , n72687 , n600014 );
xor ( n72693 , n599762 , n72443 );
xor ( n600017 , n72693 , n599771 );
and ( n72695 , n600014 , n600017 );
and ( n600019 , n72687 , n600017 );
or ( n72697 , n600015 , n72695 , n600019 );
and ( n600021 , n594952 , n66457 );
and ( n72699 , n594710 , n593778 );
nor ( n72700 , n600021 , n72699 );
xnor ( n600024 , n72700 , n593160 );
and ( n600025 , n72697 , n600024 );
xor ( n72703 , n599774 , n599776 );
xor ( n600027 , n72703 , n72456 );
and ( n600028 , n600024 , n600027 );
and ( n72706 , n72697 , n600027 );
or ( n600030 , n600025 , n600028 , n72706 );
and ( n600031 , n66967 , n594210 );
and ( n72709 , n66951 , n66885 );
nor ( n72710 , n600031 , n72709 );
xnor ( n600034 , n72710 , n593434 );
and ( n600035 , n600030 , n600034 );
xor ( n72713 , n599782 , n599786 );
xor ( n600037 , n72713 , n599789 );
and ( n600038 , n600034 , n600037 );
and ( n72716 , n600030 , n600037 );
or ( n600040 , n600035 , n600038 , n72716 );
and ( n600041 , n599976 , n600040 );
xor ( n72719 , n599932 , n599936 );
xor ( n600043 , n72719 , n599939 );
and ( n600044 , n600040 , n600043 );
and ( n72722 , n599976 , n600043 );
or ( n72723 , n600041 , n600044 , n72722 );
xor ( n72724 , n599856 , n599942 );
xor ( n72725 , n72724 , n72622 );
and ( n600049 , n72723 , n72725 );
xor ( n600050 , n72493 , n72497 );
xor ( n72728 , n600050 , n72500 );
and ( n600052 , n72725 , n72728 );
and ( n72730 , n72723 , n72728 );
or ( n72731 , n600049 , n600052 , n72730 );
and ( n600055 , n599962 , n72731 );
xor ( n600056 , n599962 , n72731 );
xor ( n72734 , n72723 , n72725 );
xor ( n600058 , n72734 , n72728 );
xor ( n72736 , n72348 , n599675 );
and ( n600060 , n70652 , n64860 );
not ( n600061 , n600060 );
and ( n72739 , n600061 , n64764 );
and ( n600063 , n70652 , n64862 );
and ( n600064 , n597980 , n64860 );
nor ( n72742 , n600063 , n600064 );
xnor ( n600066 , n72742 , n64764 );
and ( n72744 , n72739 , n600066 );
and ( n600068 , n597980 , n64862 );
and ( n600069 , n70663 , n64860 );
nor ( n72747 , n600068 , n600069 );
xnor ( n72748 , n72747 , n64764 );
and ( n600072 , n72744 , n72748 );
and ( n600073 , n72748 , n72346 );
and ( n72751 , n72744 , n72346 );
or ( n72752 , n600072 , n600073 , n72751 );
and ( n600076 , n72736 , n72752 );
and ( n600077 , n70663 , n64862 );
and ( n72755 , n597996 , n64860 );
nor ( n600079 , n600077 , n72755 );
xnor ( n600080 , n600079 , n64764 );
and ( n600081 , n72752 , n600080 );
and ( n72759 , n72736 , n600080 );
or ( n600083 , n600076 , n600081 , n72759 );
and ( n72761 , n597996 , n64862 );
and ( n72762 , n70683 , n64860 );
nor ( n600086 , n72761 , n72762 );
xnor ( n72764 , n600086 , n64764 );
and ( n600088 , n600083 , n72764 );
xor ( n72766 , n72353 , n599680 );
xor ( n72767 , n72766 , n71923 );
and ( n600091 , n72764 , n72767 );
and ( n600092 , n600083 , n72767 );
or ( n72770 , n600088 , n600091 , n600092 );
and ( n600094 , n70683 , n64862 );
and ( n600095 , n70693 , n64860 );
nor ( n72773 , n600094 , n600095 );
xnor ( n600097 , n72773 , n64764 );
and ( n600098 , n72770 , n600097 );
xor ( n600099 , n72345 , n599684 );
xor ( n72777 , n600099 , n72366 );
and ( n600101 , n600097 , n72777 );
and ( n600102 , n72770 , n72777 );
or ( n72780 , n600098 , n600101 , n600102 );
and ( n600104 , n70693 , n64862 );
and ( n600105 , n70637 , n64860 );
nor ( n72783 , n600104 , n600105 );
xnor ( n600107 , n72783 , n64764 );
and ( n72785 , n72780 , n600107 );
xor ( n600109 , n72369 , n72373 );
xor ( n72787 , n600109 , n72376 );
and ( n72788 , n600107 , n72787 );
and ( n600112 , n72780 , n72787 );
or ( n72790 , n72785 , n72788 , n600112 );
and ( n600114 , n70637 , n64862 );
and ( n72792 , n70261 , n64860 );
nor ( n72793 , n600114 , n72792 );
xnor ( n600117 , n72793 , n64764 );
and ( n72795 , n72790 , n600117 );
xor ( n600119 , n72379 , n599706 );
xor ( n600120 , n600119 , n72386 );
and ( n600121 , n600117 , n600120 );
and ( n72799 , n72790 , n600120 );
or ( n600123 , n72795 , n600121 , n72799 );
and ( n600124 , n70261 , n64862 );
and ( n72802 , n70255 , n64860 );
nor ( n600126 , n600124 , n72802 );
xnor ( n600127 , n600126 , n64764 );
and ( n600128 , n600123 , n600127 );
xor ( n72806 , n72389 , n599716 );
xor ( n600130 , n72806 , n599719 );
and ( n600131 , n600127 , n600130 );
and ( n72809 , n600123 , n600130 );
or ( n600133 , n600128 , n600131 , n72809 );
and ( n600134 , n69739 , n592486 );
and ( n72812 , n69581 , n592484 );
nor ( n600136 , n600134 , n72812 );
xnor ( n600137 , n600136 , n64990 );
and ( n72815 , n600133 , n600137 );
xor ( n600139 , n72537 , n599864 );
xor ( n600140 , n600139 , n72544 );
and ( n72818 , n600137 , n600140 );
and ( n600142 , n600133 , n600140 );
or ( n72820 , n72815 , n72818 , n600142 );
and ( n72821 , n597402 , n592486 );
and ( n72822 , n597260 , n592484 );
nor ( n600146 , n72821 , n72822 );
xnor ( n600147 , n600146 , n64990 );
and ( n72825 , n70255 , n592340 );
and ( n600149 , n597569 , n65015 );
nor ( n72827 , n72825 , n600149 );
xnor ( n72828 , n72827 , n64847 );
and ( n72829 , n600147 , n72828 );
xor ( n72830 , n72790 , n600117 );
xor ( n72831 , n72830 , n600120 );
and ( n72832 , n72828 , n72831 );
and ( n600156 , n600147 , n72831 );
or ( n72834 , n72829 , n72832 , n600156 );
and ( n72835 , n597569 , n592340 );
and ( n72836 , n597402 , n65015 );
nor ( n72837 , n72835 , n72836 );
xnor ( n600161 , n72837 , n64847 );
and ( n72839 , n72834 , n600161 );
xor ( n600163 , n600123 , n600127 );
xor ( n72841 , n600163 , n600130 );
and ( n72842 , n600161 , n72841 );
and ( n600166 , n72834 , n72841 );
or ( n72844 , n72839 , n72842 , n600166 );
and ( n600168 , n69491 , n592683 );
and ( n72846 , n69283 , n592681 );
nor ( n72847 , n600168 , n72846 );
xnor ( n72848 , n72847 , n592475 );
and ( n72849 , n72844 , n72848 );
xor ( n72850 , n600133 , n600137 );
xor ( n72851 , n72850 , n600140 );
and ( n72852 , n72848 , n72851 );
and ( n72853 , n72844 , n72851 );
or ( n72854 , n72849 , n72852 , n72853 );
and ( n600178 , n72820 , n72854 );
xor ( n600179 , n72657 , n599984 );
xor ( n72857 , n600179 , n599987 );
and ( n600181 , n72854 , n72857 );
and ( n72859 , n72820 , n72857 );
or ( n72860 , n600178 , n600181 , n72859 );
and ( n72861 , n596600 , n592683 );
and ( n72862 , n596198 , n592681 );
nor ( n72863 , n72861 , n72862 );
xnor ( n72864 , n72863 , n592475 );
and ( n72865 , n72860 , n72864 );
xor ( n72866 , n599990 , n72671 );
xor ( n72867 , n72866 , n72674 );
and ( n72868 , n72864 , n72867 );
and ( n72869 , n72860 , n72867 );
or ( n72870 , n72865 , n72868 , n72869 );
and ( n600194 , n68160 , n66142 );
and ( n600195 , n67940 , n66140 );
nor ( n72873 , n600194 , n600195 );
xnor ( n600197 , n72873 , n592960 );
and ( n72875 , n72870 , n600197 );
and ( n72876 , n595633 , n593256 );
and ( n72877 , n595521 , n593254 );
nor ( n72878 , n72876 , n72877 );
xnor ( n600202 , n72878 , n65490 );
and ( n72880 , n600197 , n600202 );
and ( n600204 , n72870 , n600202 );
or ( n600205 , n72875 , n72880 , n600204 );
and ( n72883 , n67636 , n66457 );
and ( n600207 , n594952 , n593778 );
nor ( n72885 , n72883 , n600207 );
xnor ( n600209 , n72885 , n593160 );
and ( n600210 , n600205 , n600209 );
xor ( n72888 , n72577 , n599904 );
xor ( n600212 , n72888 , n599907 );
and ( n72890 , n600209 , n600212 );
and ( n72891 , n600205 , n600212 );
or ( n600215 , n600210 , n72890 , n72891 );
and ( n72893 , n594295 , n594210 );
and ( n600217 , n66967 , n66885 );
nor ( n72895 , n72893 , n600217 );
xnor ( n600219 , n72895 , n593434 );
and ( n600220 , n600215 , n600219 );
xor ( n72898 , n599910 , n599914 );
xor ( n600222 , n72898 , n72596 );
and ( n72900 , n600219 , n600222 );
and ( n72901 , n600215 , n600222 );
or ( n72902 , n600220 , n72900 , n72901 );
and ( n72903 , n596198 , n65592 );
and ( n72904 , n596193 , n592913 );
nor ( n72905 , n72903 , n72904 );
xnor ( n72906 , n72905 , n592638 );
and ( n600230 , n69283 , n592683 );
and ( n72908 , n596600 , n592681 );
nor ( n600232 , n600230 , n72908 );
xnor ( n72910 , n600232 , n592475 );
and ( n72911 , n72906 , n72910 );
xor ( n600235 , n72820 , n72854 );
xor ( n600236 , n600235 , n72857 );
and ( n72914 , n72910 , n600236 );
and ( n600238 , n72906 , n600236 );
or ( n600239 , n72911 , n72914 , n600238 );
and ( n72917 , n595521 , n66142 );
and ( n600241 , n68160 , n66140 );
nor ( n600242 , n72917 , n600241 );
xnor ( n600243 , n600242 , n592960 );
and ( n72921 , n600239 , n600243 );
and ( n600245 , n595827 , n593256 );
and ( n72923 , n595633 , n593254 );
nor ( n600247 , n600245 , n72923 );
xnor ( n72925 , n600247 , n65490 );
and ( n72926 , n600243 , n72925 );
and ( n72927 , n600239 , n72925 );
or ( n600251 , n72921 , n72926 , n72927 );
and ( n72929 , n595103 , n66457 );
and ( n600253 , n67636 , n593778 );
nor ( n72931 , n72929 , n600253 );
xnor ( n72932 , n72931 , n593160 );
and ( n600256 , n600251 , n72932 );
xor ( n72934 , n72677 , n600004 );
xor ( n72935 , n72934 , n600007 );
and ( n600259 , n72932 , n72935 );
and ( n600260 , n600251 , n72935 );
or ( n72938 , n600256 , n600259 , n600260 );
and ( n600262 , n594710 , n594210 );
and ( n600263 , n594295 , n66885 );
nor ( n72941 , n600262 , n600263 );
xnor ( n600265 , n72941 , n593434 );
and ( n600266 , n72938 , n600265 );
xor ( n72944 , n72687 , n600014 );
xor ( n600268 , n72944 , n600017 );
and ( n72946 , n600265 , n600268 );
and ( n600270 , n72938 , n600268 );
or ( n72948 , n600266 , n72946 , n600270 );
and ( n72949 , n66951 , n594441 );
and ( n600273 , n66793 , n67116 );
nor ( n72951 , n72949 , n600273 );
xnor ( n600275 , n72951 , n66190 );
and ( n72953 , n72948 , n600275 );
xor ( n72954 , n72697 , n600024 );
xor ( n600278 , n72954 , n600027 );
and ( n600279 , n600275 , n600278 );
and ( n72957 , n72948 , n600278 );
or ( n600281 , n72953 , n600279 , n72957 );
and ( n600282 , n72902 , n600281 );
xor ( n72960 , n600030 , n600034 );
xor ( n600284 , n72960 , n600037 );
and ( n600285 , n600281 , n600284 );
and ( n600286 , n72902 , n600284 );
or ( n72964 , n600282 , n600285 , n600286 );
xor ( n600288 , n599846 , n72527 );
xor ( n600289 , n600288 , n599853 );
and ( n72967 , n72964 , n600289 );
xor ( n600291 , n599976 , n600040 );
xor ( n600292 , n600291 , n600043 );
and ( n72970 , n600289 , n600292 );
and ( n600294 , n72964 , n600292 );
or ( n72972 , n72967 , n72970 , n600294 );
and ( n600296 , n600058 , n72972 );
xor ( n72974 , n600058 , n72972 );
xor ( n600298 , n72964 , n600289 );
xor ( n600299 , n600298 , n600292 );
and ( n72977 , n69581 , n592683 );
and ( n72978 , n69491 , n592681 );
nor ( n600302 , n72977 , n72978 );
xnor ( n72980 , n600302 , n592475 );
and ( n72981 , n597260 , n592486 );
and ( n600305 , n69739 , n592484 );
nor ( n72983 , n72981 , n600305 );
xnor ( n72984 , n72983 , n64990 );
and ( n72985 , n72980 , n72984 );
xor ( n72986 , n72834 , n600161 );
xor ( n600310 , n72986 , n72841 );
and ( n600311 , n72984 , n600310 );
and ( n72989 , n72980 , n600310 );
or ( n72990 , n72985 , n600311 , n72989 );
and ( n600314 , n596193 , n593256 );
and ( n600315 , n596057 , n593254 );
nor ( n72993 , n600314 , n600315 );
xnor ( n600317 , n72993 , n65490 );
and ( n600318 , n72990 , n600317 );
xor ( n600319 , n72844 , n72848 );
xor ( n72997 , n600319 , n72851 );
and ( n600321 , n600317 , n72997 );
and ( n72999 , n72990 , n72997 );
or ( n600323 , n600318 , n600321 , n72999 );
and ( n73001 , n596057 , n593256 );
and ( n73002 , n595827 , n593254 );
nor ( n600326 , n73001 , n73002 );
xnor ( n600327 , n600326 , n65490 );
and ( n73005 , n600323 , n600327 );
xor ( n600329 , n72906 , n72910 );
xor ( n600330 , n600329 , n600236 );
and ( n73008 , n600327 , n600330 );
and ( n600332 , n600323 , n600330 );
or ( n600333 , n73005 , n73008 , n600332 );
and ( n73011 , n67940 , n66457 );
and ( n73012 , n595103 , n593778 );
nor ( n600336 , n73011 , n73012 );
xnor ( n600337 , n600336 , n593160 );
and ( n73015 , n600333 , n600337 );
xor ( n600339 , n72860 , n72864 );
xor ( n600340 , n600339 , n72867 );
and ( n73018 , n600337 , n600340 );
and ( n600342 , n600333 , n600340 );
or ( n600343 , n73015 , n73018 , n600342 );
and ( n73021 , n594952 , n594210 );
and ( n73022 , n594710 , n66885 );
nor ( n73023 , n73021 , n73022 );
xnor ( n73024 , n73023 , n593434 );
and ( n600348 , n600343 , n73024 );
xor ( n73026 , n72870 , n600197 );
xor ( n600350 , n73026 , n600202 );
and ( n73028 , n73024 , n600350 );
and ( n73029 , n600343 , n600350 );
or ( n600353 , n600348 , n73028 , n73029 );
and ( n600354 , n66967 , n594441 );
and ( n73032 , n66951 , n67116 );
nor ( n600356 , n600354 , n73032 );
xnor ( n600357 , n600356 , n66190 );
and ( n73035 , n600353 , n600357 );
xor ( n600359 , n600205 , n600209 );
xor ( n73037 , n600359 , n600212 );
and ( n73038 , n600357 , n73037 );
and ( n600362 , n600353 , n73037 );
or ( n73040 , n73035 , n73038 , n600362 );
and ( n600364 , n594124 , n594807 );
and ( n600365 , n66606 , n594804 );
nor ( n73043 , n600364 , n600365 );
xnor ( n73044 , n73043 , n66187 );
and ( n73045 , n73040 , n73044 );
xor ( n73046 , n600215 , n600219 );
xor ( n600370 , n73046 , n600222 );
and ( n600371 , n73044 , n600370 );
and ( n73049 , n73040 , n600370 );
or ( n600373 , n73045 , n600371 , n73049 );
xor ( n73051 , n72643 , n599970 );
xor ( n600375 , n73051 , n72650 );
and ( n73053 , n600373 , n600375 );
xor ( n73054 , n72902 , n600281 );
xor ( n600378 , n73054 , n600284 );
and ( n73056 , n600375 , n600378 );
and ( n600380 , n600373 , n600378 );
or ( n73058 , n73053 , n73056 , n600380 );
and ( n73059 , n600299 , n73058 );
xor ( n600383 , n600299 , n73058 );
xor ( n73061 , n600373 , n600375 );
xor ( n600385 , n73061 , n600378 );
xor ( n73063 , n72739 , n600066 );
and ( n600387 , n70652 , n65015 );
not ( n600388 , n600387 );
and ( n73066 , n600388 , n64847 );
and ( n600390 , n70652 , n592340 );
and ( n600391 , n597980 , n65015 );
nor ( n600392 , n600390 , n600391 );
xnor ( n73070 , n600392 , n64847 );
and ( n600394 , n73066 , n73070 );
and ( n600395 , n597980 , n592340 );
and ( n73073 , n70663 , n65015 );
nor ( n600397 , n600395 , n73073 );
xnor ( n600398 , n600397 , n64847 );
and ( n73076 , n600394 , n600398 );
and ( n600400 , n600398 , n600060 );
and ( n73078 , n600394 , n600060 );
or ( n600402 , n73076 , n600400 , n73078 );
and ( n73080 , n73063 , n600402 );
and ( n600404 , n70663 , n592340 );
and ( n73082 , n597996 , n65015 );
nor ( n73083 , n600404 , n73082 );
xnor ( n600407 , n73083 , n64847 );
and ( n73085 , n600402 , n600407 );
and ( n600409 , n73063 , n600407 );
or ( n73087 , n73080 , n73085 , n600409 );
and ( n73088 , n597996 , n592340 );
and ( n600412 , n70683 , n65015 );
nor ( n73090 , n73088 , n600412 );
xnor ( n600414 , n73090 , n64847 );
and ( n600415 , n73087 , n600414 );
xor ( n73093 , n72744 , n72748 );
xor ( n600417 , n73093 , n72346 );
and ( n600418 , n600414 , n600417 );
and ( n600419 , n73087 , n600417 );
or ( n73097 , n600415 , n600418 , n600419 );
and ( n600421 , n70683 , n592340 );
and ( n600422 , n70693 , n65015 );
nor ( n73100 , n600421 , n600422 );
xnor ( n600424 , n73100 , n64847 );
and ( n600425 , n73097 , n600424 );
xor ( n600426 , n72736 , n72752 );
xor ( n73104 , n600426 , n600080 );
and ( n600428 , n600424 , n73104 );
and ( n600429 , n73097 , n73104 );
or ( n73107 , n600425 , n600428 , n600429 );
and ( n600431 , n70693 , n592340 );
and ( n73109 , n70637 , n65015 );
nor ( n73110 , n600431 , n73109 );
xnor ( n600434 , n73110 , n64847 );
and ( n73112 , n73107 , n600434 );
xor ( n600436 , n600083 , n72764 );
xor ( n73114 , n600436 , n72767 );
and ( n73115 , n600434 , n73114 );
and ( n73116 , n73107 , n73114 );
or ( n600440 , n73112 , n73115 , n73116 );
and ( n73118 , n70637 , n592340 );
and ( n600442 , n70261 , n65015 );
nor ( n73120 , n73118 , n600442 );
xnor ( n73121 , n73120 , n64847 );
and ( n600445 , n600440 , n73121 );
xor ( n73123 , n72770 , n600097 );
xor ( n600447 , n73123 , n72777 );
and ( n73125 , n73121 , n600447 );
and ( n600449 , n600440 , n600447 );
or ( n600450 , n600445 , n73125 , n600449 );
and ( n73128 , n70261 , n592340 );
and ( n600452 , n70255 , n65015 );
nor ( n73130 , n73128 , n600452 );
xnor ( n73131 , n73130 , n64847 );
and ( n600455 , n600450 , n73131 );
xor ( n73133 , n72780 , n600107 );
xor ( n600457 , n73133 , n72787 );
and ( n73135 , n73131 , n600457 );
and ( n600459 , n600450 , n600457 );
or ( n73137 , n600455 , n73135 , n600459 );
and ( n73138 , n69739 , n592683 );
and ( n73139 , n69581 , n592681 );
nor ( n73140 , n73138 , n73139 );
xnor ( n73141 , n73140 , n592475 );
and ( n73142 , n73137 , n73141 );
xor ( n600466 , n600147 , n72828 );
xor ( n73144 , n600466 , n72831 );
and ( n600468 , n73141 , n73144 );
and ( n600469 , n73137 , n73144 );
or ( n73147 , n73142 , n600468 , n600469 );
and ( n600471 , n69283 , n65592 );
and ( n600472 , n596600 , n592913 );
nor ( n73150 , n600471 , n600472 );
xnor ( n73151 , n73150 , n592638 );
and ( n600475 , n73147 , n73151 );
xor ( n600476 , n72980 , n72984 );
xor ( n73154 , n600476 , n600310 );
and ( n600478 , n73151 , n73154 );
and ( n600479 , n73147 , n73154 );
or ( n73157 , n600475 , n600478 , n600479 );
and ( n600481 , n595827 , n66142 );
and ( n600482 , n595633 , n66140 );
nor ( n73160 , n600481 , n600482 );
xnor ( n600484 , n73160 , n592960 );
and ( n600485 , n73157 , n600484 );
and ( n600486 , n596600 , n65592 );
and ( n73164 , n596198 , n592913 );
nor ( n600488 , n600486 , n73164 );
xnor ( n73166 , n600488 , n592638 );
and ( n600490 , n600484 , n73166 );
and ( n600491 , n73157 , n73166 );
or ( n73169 , n600485 , n600490 , n600491 );
and ( n73170 , n595103 , n594210 );
and ( n600494 , n67636 , n66885 );
nor ( n600495 , n73170 , n600494 );
xnor ( n73173 , n600495 , n593434 );
and ( n600497 , n73169 , n73173 );
and ( n73175 , n595633 , n66142 );
and ( n600499 , n595521 , n66140 );
nor ( n600500 , n73175 , n600499 );
xnor ( n73178 , n600500 , n592960 );
and ( n600502 , n73173 , n73178 );
and ( n600503 , n73169 , n73178 );
or ( n73181 , n600497 , n600502 , n600503 );
and ( n600505 , n67636 , n594210 );
and ( n73183 , n594952 , n66885 );
nor ( n600507 , n600505 , n73183 );
xnor ( n600508 , n600507 , n593434 );
and ( n600509 , n73181 , n600508 );
xor ( n73187 , n600239 , n600243 );
xor ( n600511 , n73187 , n72925 );
and ( n600512 , n600508 , n600511 );
and ( n73190 , n73181 , n600511 );
or ( n73191 , n600509 , n600512 , n73190 );
and ( n600515 , n594295 , n594441 );
and ( n600516 , n66967 , n67116 );
nor ( n73194 , n600515 , n600516 );
xnor ( n600518 , n73194 , n66190 );
and ( n73196 , n73191 , n600518 );
xor ( n73197 , n600251 , n72932 );
xor ( n600521 , n73197 , n72935 );
and ( n73199 , n600518 , n600521 );
and ( n600523 , n73191 , n600521 );
or ( n73201 , n73196 , n73199 , n600523 );
and ( n73202 , n66793 , n594807 );
and ( n600526 , n594124 , n594804 );
nor ( n600527 , n73202 , n600526 );
xnor ( n73205 , n600527 , n66187 );
and ( n600529 , n73201 , n73205 );
xor ( n73207 , n72938 , n600265 );
xor ( n600531 , n73207 , n600268 );
and ( n600532 , n73205 , n600531 );
and ( n73210 , n73201 , n600531 );
or ( n600534 , n600529 , n600532 , n73210 );
xor ( n600535 , n73040 , n73044 );
xor ( n600536 , n600535 , n600370 );
and ( n73214 , n600534 , n600536 );
xor ( n600538 , n72948 , n600275 );
xor ( n73216 , n600538 , n600278 );
and ( n73217 , n600536 , n73216 );
and ( n600541 , n600534 , n73216 );
or ( n73219 , n73214 , n73217 , n600541 );
and ( n600543 , n600385 , n73219 );
xor ( n73221 , n600385 , n73219 );
and ( n73222 , n597402 , n592683 );
and ( n600546 , n597260 , n592681 );
nor ( n600547 , n73222 , n600546 );
xnor ( n73225 , n600547 , n592475 );
and ( n600549 , n70255 , n592486 );
and ( n600550 , n597569 , n592484 );
nor ( n73228 , n600549 , n600550 );
xnor ( n600552 , n73228 , n64990 );
and ( n600553 , n73225 , n600552 );
xor ( n600554 , n600440 , n73121 );
xor ( n73232 , n600554 , n600447 );
and ( n600556 , n600552 , n73232 );
and ( n600557 , n73225 , n73232 );
or ( n73235 , n600553 , n600556 , n600557 );
and ( n600559 , n597569 , n592486 );
and ( n600560 , n597402 , n592484 );
nor ( n73238 , n600559 , n600560 );
xnor ( n600562 , n73238 , n64990 );
and ( n73240 , n73235 , n600562 );
xor ( n600564 , n600450 , n73131 );
xor ( n73242 , n600564 , n600457 );
and ( n73243 , n600562 , n73242 );
and ( n600567 , n73235 , n73242 );
or ( n73245 , n73240 , n73243 , n600567 );
and ( n600569 , n69491 , n65592 );
and ( n73247 , n69283 , n592913 );
nor ( n73248 , n600569 , n73247 );
xnor ( n600572 , n73248 , n592638 );
and ( n600573 , n73245 , n600572 );
xor ( n73251 , n73137 , n73141 );
xor ( n600575 , n73251 , n73144 );
and ( n600576 , n600572 , n600575 );
and ( n73254 , n73245 , n600575 );
or ( n600578 , n600573 , n600576 , n73254 );
and ( n600579 , n596198 , n593256 );
and ( n600580 , n596193 , n593254 );
nor ( n73258 , n600579 , n600580 );
xnor ( n600582 , n73258 , n65490 );
and ( n600583 , n600578 , n600582 );
xor ( n73261 , n73147 , n73151 );
xor ( n600585 , n73261 , n73154 );
and ( n600586 , n600582 , n600585 );
and ( n73264 , n600578 , n600585 );
or ( n600588 , n600583 , n600586 , n73264 );
and ( n73266 , n595521 , n66457 );
and ( n600590 , n68160 , n593778 );
nor ( n73268 , n73266 , n600590 );
xnor ( n600592 , n73268 , n593160 );
and ( n73270 , n600588 , n600592 );
xor ( n73271 , n72990 , n600317 );
xor ( n600595 , n73271 , n72997 );
and ( n73273 , n600592 , n600595 );
and ( n600597 , n600588 , n600595 );
or ( n73275 , n73270 , n73273 , n600597 );
and ( n73276 , n68160 , n66457 );
and ( n600600 , n67940 , n593778 );
nor ( n600601 , n73276 , n600600 );
xnor ( n73279 , n600601 , n593160 );
and ( n600603 , n73275 , n73279 );
xor ( n600604 , n600323 , n600327 );
xor ( n73282 , n600604 , n600330 );
and ( n600606 , n73279 , n73282 );
and ( n600607 , n73275 , n73282 );
or ( n600608 , n600603 , n600606 , n600607 );
and ( n73286 , n594710 , n594441 );
and ( n600610 , n594295 , n67116 );
nor ( n600611 , n73286 , n600610 );
xnor ( n73289 , n600611 , n66190 );
and ( n600613 , n600608 , n73289 );
xor ( n73291 , n600333 , n600337 );
xor ( n73292 , n73291 , n600340 );
and ( n73293 , n73289 , n73292 );
and ( n73294 , n600608 , n73292 );
or ( n600618 , n600613 , n73293 , n73294 );
and ( n73296 , n66951 , n594807 );
and ( n600620 , n66793 , n594804 );
nor ( n600621 , n73296 , n600620 );
xnor ( n73299 , n600621 , n66187 );
and ( n600623 , n600618 , n73299 );
xor ( n73301 , n600343 , n73024 );
xor ( n600625 , n73301 , n600350 );
and ( n600626 , n73299 , n600625 );
and ( n73304 , n600618 , n600625 );
or ( n600628 , n600623 , n600626 , n73304 );
xor ( n600629 , n73201 , n73205 );
xor ( n73307 , n600629 , n600531 );
and ( n600631 , n600628 , n73307 );
xor ( n73309 , n600353 , n600357 );
xor ( n600633 , n73309 , n73037 );
and ( n600634 , n73307 , n600633 );
and ( n73312 , n600628 , n600633 );
or ( n600636 , n600631 , n600634 , n73312 );
xor ( n600637 , n600534 , n600536 );
xor ( n73315 , n600637 , n73216 );
and ( n73316 , n600636 , n73315 );
xor ( n600640 , n600636 , n73315 );
xor ( n600641 , n600628 , n73307 );
xor ( n73319 , n600641 , n600633 );
and ( n600643 , n69581 , n65592 );
and ( n600644 , n69491 , n592913 );
nor ( n73322 , n600643 , n600644 );
xnor ( n600646 , n73322 , n592638 );
and ( n600647 , n597260 , n592683 );
and ( n73325 , n69739 , n592681 );
nor ( n600649 , n600647 , n73325 );
xnor ( n73327 , n600649 , n592475 );
and ( n73328 , n600646 , n73327 );
xor ( n73329 , n73235 , n600562 );
xor ( n73330 , n73329 , n73242 );
and ( n73331 , n73327 , n73330 );
and ( n73332 , n600646 , n73330 );
or ( n600656 , n73328 , n73331 , n73332 );
and ( n600657 , n596600 , n593256 );
and ( n600658 , n596198 , n593254 );
nor ( n600659 , n600657 , n600658 );
xnor ( n73337 , n600659 , n65490 );
and ( n600661 , n600656 , n73337 );
xor ( n73339 , n73245 , n600572 );
xor ( n73340 , n73339 , n600575 );
and ( n73341 , n73337 , n73340 );
and ( n73342 , n600656 , n73340 );
or ( n73343 , n600661 , n73341 , n73342 );
and ( n73344 , n595633 , n66457 );
and ( n73345 , n595521 , n593778 );
nor ( n600669 , n73344 , n73345 );
xnor ( n73347 , n600669 , n593160 );
and ( n73348 , n73343 , n73347 );
and ( n600672 , n596057 , n66142 );
and ( n73350 , n595827 , n66140 );
nor ( n600674 , n600672 , n73350 );
xnor ( n73352 , n600674 , n592960 );
and ( n73353 , n73347 , n73352 );
and ( n600677 , n73343 , n73352 );
or ( n600678 , n73348 , n73353 , n600677 );
and ( n73356 , n67940 , n594210 );
and ( n600680 , n595103 , n66885 );
nor ( n73358 , n73356 , n600680 );
xnor ( n600682 , n73358 , n593434 );
and ( n73360 , n600678 , n600682 );
xor ( n73361 , n73157 , n600484 );
xor ( n600685 , n73361 , n73166 );
and ( n600686 , n600682 , n600685 );
and ( n73364 , n600678 , n600685 );
or ( n600688 , n73360 , n600686 , n73364 );
and ( n600689 , n594952 , n594441 );
and ( n73367 , n594710 , n67116 );
nor ( n600691 , n600689 , n73367 );
xnor ( n600692 , n600691 , n66190 );
and ( n73370 , n600688 , n600692 );
xor ( n73371 , n73169 , n73173 );
xor ( n600695 , n73371 , n73178 );
and ( n600696 , n600692 , n600695 );
and ( n73374 , n600688 , n600695 );
or ( n600698 , n73370 , n600696 , n73374 );
and ( n600699 , n66967 , n594807 );
and ( n73377 , n66951 , n594804 );
nor ( n600701 , n600699 , n73377 );
xnor ( n600702 , n600701 , n66187 );
and ( n73380 , n600698 , n600702 );
xor ( n73381 , n73181 , n600508 );
xor ( n73382 , n73381 , n600511 );
and ( n73383 , n600702 , n73382 );
and ( n73384 , n600698 , n73382 );
or ( n600708 , n73380 , n73383 , n73384 );
xor ( n73386 , n600618 , n73299 );
xor ( n73387 , n73386 , n600625 );
and ( n600711 , n600708 , n73387 );
xor ( n600712 , n73191 , n600518 );
xor ( n73390 , n600712 , n600521 );
and ( n600714 , n73387 , n73390 );
and ( n600715 , n600708 , n73390 );
or ( n73393 , n600711 , n600714 , n600715 );
and ( n600717 , n73319 , n73393 );
xor ( n73395 , n73319 , n73393 );
xor ( n600719 , n73066 , n73070 );
and ( n73397 , n70652 , n592484 );
not ( n600721 , n73397 );
and ( n73399 , n600721 , n64990 );
and ( n73400 , n70652 , n592486 );
and ( n73401 , n597980 , n592484 );
nor ( n73402 , n73400 , n73401 );
xnor ( n73403 , n73402 , n64990 );
and ( n600727 , n73399 , n73403 );
and ( n600728 , n597980 , n592486 );
and ( n73406 , n70663 , n592484 );
nor ( n600730 , n600728 , n73406 );
xnor ( n73408 , n600730 , n64990 );
and ( n600732 , n600727 , n73408 );
and ( n600733 , n73408 , n600387 );
and ( n73411 , n600727 , n600387 );
or ( n600735 , n600732 , n600733 , n73411 );
and ( n600736 , n600719 , n600735 );
and ( n73414 , n70663 , n592486 );
and ( n600738 , n597996 , n592484 );
nor ( n600739 , n73414 , n600738 );
xnor ( n73417 , n600739 , n64990 );
and ( n600741 , n600735 , n73417 );
and ( n73419 , n600719 , n73417 );
or ( n600743 , n600736 , n600741 , n73419 );
and ( n73421 , n597996 , n592486 );
and ( n600745 , n70683 , n592484 );
nor ( n600746 , n73421 , n600745 );
xnor ( n73424 , n600746 , n64990 );
and ( n73425 , n600743 , n73424 );
xor ( n600749 , n600394 , n600398 );
xor ( n73427 , n600749 , n600060 );
and ( n73428 , n73424 , n73427 );
and ( n600752 , n600743 , n73427 );
or ( n600753 , n73425 , n73428 , n600752 );
and ( n73431 , n70683 , n592486 );
and ( n73432 , n70693 , n592484 );
nor ( n73433 , n73431 , n73432 );
xnor ( n73434 , n73433 , n64990 );
and ( n73435 , n600753 , n73434 );
xor ( n73436 , n73063 , n600402 );
xor ( n73437 , n73436 , n600407 );
and ( n73438 , n73434 , n73437 );
and ( n73439 , n600753 , n73437 );
or ( n600763 , n73435 , n73438 , n73439 );
and ( n73441 , n70693 , n592486 );
and ( n600765 , n70637 , n592484 );
nor ( n73443 , n73441 , n600765 );
xnor ( n73444 , n73443 , n64990 );
and ( n600768 , n600763 , n73444 );
xor ( n600769 , n73087 , n600414 );
xor ( n73447 , n600769 , n600417 );
and ( n600771 , n73444 , n73447 );
and ( n73449 , n600763 , n73447 );
or ( n73450 , n600768 , n600771 , n73449 );
and ( n600774 , n70637 , n592486 );
and ( n600775 , n70261 , n592484 );
nor ( n73453 , n600774 , n600775 );
xnor ( n600777 , n73453 , n64990 );
and ( n73455 , n73450 , n600777 );
xor ( n73456 , n73097 , n600424 );
xor ( n73457 , n73456 , n73104 );
and ( n73458 , n600777 , n73457 );
and ( n73459 , n73450 , n73457 );
or ( n73460 , n73455 , n73458 , n73459 );
and ( n73461 , n70261 , n592486 );
and ( n600785 , n70255 , n592484 );
nor ( n600786 , n73461 , n600785 );
xnor ( n73464 , n600786 , n64990 );
and ( n600788 , n73460 , n73464 );
xor ( n73466 , n73107 , n600434 );
xor ( n73467 , n73466 , n73114 );
and ( n600791 , n73464 , n73467 );
and ( n73469 , n73460 , n73467 );
or ( n600793 , n600788 , n600791 , n73469 );
and ( n600794 , n69739 , n65592 );
and ( n73472 , n69581 , n592913 );
nor ( n600796 , n600794 , n73472 );
xnor ( n73474 , n600796 , n592638 );
and ( n600798 , n600793 , n73474 );
xor ( n73476 , n73225 , n600552 );
xor ( n600800 , n73476 , n73232 );
and ( n600801 , n73474 , n600800 );
and ( n73479 , n600793 , n600800 );
or ( n600803 , n600798 , n600801 , n73479 );
and ( n73481 , n597402 , n65592 );
and ( n600805 , n597260 , n592913 );
nor ( n73483 , n73481 , n600805 );
xnor ( n73484 , n73483 , n592638 );
and ( n73485 , n70255 , n592683 );
and ( n73486 , n597569 , n592681 );
nor ( n73487 , n73485 , n73486 );
xnor ( n73488 , n73487 , n592475 );
and ( n73489 , n73484 , n73488 );
xor ( n73490 , n73450 , n600777 );
xor ( n73491 , n73490 , n73457 );
and ( n73492 , n73488 , n73491 );
and ( n73493 , n73484 , n73491 );
or ( n73494 , n73489 , n73492 , n73493 );
and ( n73495 , n597569 , n592683 );
and ( n73496 , n597402 , n592681 );
nor ( n73497 , n73495 , n73496 );
xnor ( n73498 , n73497 , n592475 );
and ( n73499 , n73494 , n73498 );
xor ( n73500 , n73460 , n73464 );
xor ( n73501 , n73500 , n73467 );
and ( n73502 , n73498 , n73501 );
and ( n73503 , n73494 , n73501 );
or ( n73504 , n73499 , n73502 , n73503 );
and ( n73505 , n69491 , n593256 );
and ( n600829 , n69283 , n593254 );
nor ( n73507 , n73505 , n600829 );
xnor ( n73508 , n73507 , n65490 );
and ( n73509 , n73504 , n73508 );
xor ( n73510 , n600793 , n73474 );
xor ( n73511 , n73510 , n600800 );
and ( n73512 , n73508 , n73511 );
and ( n73513 , n73504 , n73511 );
or ( n73514 , n73509 , n73512 , n73513 );
and ( n73515 , n600803 , n73514 );
xor ( n73516 , n600646 , n73327 );
xor ( n73517 , n73516 , n73330 );
and ( n73518 , n73514 , n73517 );
and ( n73519 , n600803 , n73517 );
or ( n73520 , n73515 , n73518 , n73519 );
and ( n73521 , n595827 , n66457 );
and ( n73522 , n595633 , n593778 );
nor ( n73523 , n73521 , n73522 );
xnor ( n73524 , n73523 , n593160 );
and ( n73525 , n73520 , n73524 );
and ( n600849 , n596193 , n66142 );
and ( n73527 , n596057 , n66140 );
nor ( n600851 , n600849 , n73527 );
xnor ( n600852 , n600851 , n592960 );
and ( n600853 , n73524 , n600852 );
and ( n73531 , n73520 , n600852 );
or ( n600855 , n73525 , n600853 , n73531 );
and ( n600856 , n595103 , n594441 );
and ( n73534 , n67636 , n67116 );
nor ( n600858 , n600856 , n73534 );
xnor ( n600859 , n600858 , n66190 );
and ( n600860 , n600855 , n600859 );
xor ( n73538 , n600578 , n600582 );
xor ( n600862 , n73538 , n600585 );
and ( n600863 , n600859 , n600862 );
and ( n73541 , n600855 , n600862 );
or ( n600865 , n600860 , n600863 , n73541 );
and ( n600866 , n67636 , n594441 );
and ( n73544 , n594952 , n67116 );
nor ( n600868 , n600866 , n73544 );
xnor ( n73546 , n600868 , n66190 );
and ( n73547 , n600865 , n73546 );
xor ( n73548 , n600588 , n600592 );
xor ( n73549 , n73548 , n600595 );
and ( n73550 , n73546 , n73549 );
and ( n73551 , n600865 , n73549 );
or ( n600875 , n73547 , n73550 , n73551 );
and ( n73553 , n594295 , n594807 );
and ( n600877 , n66967 , n594804 );
nor ( n73555 , n73553 , n600877 );
xnor ( n600879 , n73555 , n66187 );
and ( n600880 , n600875 , n600879 );
xor ( n73558 , n73275 , n73279 );
xor ( n600882 , n73558 , n73282 );
and ( n600883 , n600879 , n600882 );
and ( n73561 , n600875 , n600882 );
or ( n600885 , n600880 , n600883 , n73561 );
xor ( n600886 , n600698 , n600702 );
xor ( n73564 , n600886 , n73382 );
and ( n600888 , n600885 , n73564 );
xor ( n600889 , n600608 , n73289 );
xor ( n73567 , n600889 , n73292 );
and ( n600891 , n73564 , n73567 );
and ( n73569 , n600885 , n73567 );
or ( n73570 , n600888 , n600891 , n73569 );
xor ( n73571 , n600708 , n73387 );
xor ( n73572 , n73571 , n73390 );
and ( n73573 , n73570 , n73572 );
xor ( n73574 , n73570 , n73572 );
xor ( n73575 , n600885 , n73564 );
xor ( n73576 , n73575 , n73567 );
and ( n73577 , n596198 , n66142 );
and ( n73578 , n596193 , n66140 );
nor ( n73579 , n73577 , n73578 );
xnor ( n73580 , n73579 , n592960 );
and ( n73581 , n69283 , n593256 );
and ( n600905 , n596600 , n593254 );
nor ( n73583 , n73581 , n600905 );
xnor ( n600907 , n73583 , n65490 );
and ( n600908 , n73580 , n600907 );
xor ( n73586 , n600803 , n73514 );
xor ( n73587 , n73586 , n73517 );
and ( n73588 , n600907 , n73587 );
and ( n73589 , n73580 , n73587 );
or ( n600913 , n600908 , n73588 , n73589 );
and ( n73591 , n595521 , n594210 );
and ( n600915 , n68160 , n66885 );
nor ( n73593 , n73591 , n600915 );
xnor ( n600917 , n73593 , n593434 );
and ( n600918 , n600913 , n600917 );
xor ( n73596 , n600656 , n73337 );
xor ( n73597 , n73596 , n73340 );
and ( n600921 , n600917 , n73597 );
and ( n73599 , n600913 , n73597 );
or ( n73600 , n600918 , n600921 , n73599 );
and ( n600924 , n68160 , n594210 );
and ( n73602 , n67940 , n66885 );
nor ( n600926 , n600924 , n73602 );
xnor ( n600927 , n600926 , n593434 );
and ( n73605 , n73600 , n600927 );
xor ( n600929 , n73343 , n73347 );
xor ( n600930 , n600929 , n73352 );
and ( n73608 , n600927 , n600930 );
and ( n73609 , n73600 , n600930 );
or ( n600933 , n73605 , n73608 , n73609 );
and ( n600934 , n594710 , n594807 );
and ( n73612 , n594295 , n594804 );
nor ( n600936 , n600934 , n73612 );
xnor ( n600937 , n600936 , n66187 );
and ( n73615 , n600933 , n600937 );
xor ( n600939 , n600678 , n600682 );
xor ( n73617 , n600939 , n600685 );
and ( n73618 , n600937 , n73617 );
and ( n73619 , n600933 , n73617 );
or ( n73620 , n73615 , n73618 , n73619 );
xor ( n73621 , n600688 , n600692 );
xor ( n73622 , n73621 , n600695 );
and ( n73623 , n73620 , n73622 );
xor ( n73624 , n600875 , n600879 );
xor ( n73625 , n73624 , n600882 );
and ( n73626 , n73622 , n73625 );
and ( n600950 , n73620 , n73625 );
or ( n73628 , n73623 , n73626 , n600950 );
and ( n600952 , n73576 , n73628 );
xor ( n73630 , n73576 , n73628 );
xor ( n600954 , n73620 , n73622 );
xor ( n600955 , n600954 , n73625 );
and ( n73633 , n69581 , n593256 );
and ( n600957 , n69491 , n593254 );
nor ( n600958 , n73633 , n600957 );
xnor ( n73636 , n600958 , n65490 );
and ( n73637 , n597260 , n65592 );
and ( n600961 , n69739 , n592913 );
nor ( n73639 , n73637 , n600961 );
xnor ( n600963 , n73639 , n592638 );
and ( n73641 , n73636 , n600963 );
xor ( n600965 , n73494 , n73498 );
xor ( n600966 , n600965 , n73501 );
and ( n73644 , n600963 , n600966 );
and ( n600968 , n73636 , n600966 );
or ( n73646 , n73641 , n73644 , n600968 );
and ( n73647 , n596600 , n66142 );
and ( n73648 , n596198 , n66140 );
nor ( n600972 , n73647 , n73648 );
xnor ( n73650 , n600972 , n592960 );
and ( n600974 , n73646 , n73650 );
xor ( n73652 , n73504 , n73508 );
xor ( n600976 , n73652 , n73511 );
and ( n73654 , n73650 , n600976 );
and ( n73655 , n73646 , n600976 );
or ( n600979 , n600974 , n73654 , n73655 );
and ( n600980 , n595633 , n594210 );
and ( n73658 , n595521 , n66885 );
nor ( n600982 , n600980 , n73658 );
xnor ( n600983 , n600982 , n593434 );
and ( n73661 , n600979 , n600983 );
and ( n600985 , n596057 , n66457 );
and ( n600986 , n595827 , n593778 );
nor ( n600987 , n600985 , n600986 );
xnor ( n73665 , n600987 , n593160 );
and ( n73666 , n600983 , n73665 );
and ( n600990 , n600979 , n73665 );
or ( n73668 , n73661 , n73666 , n600990 );
and ( n600992 , n67940 , n594441 );
and ( n73670 , n595103 , n67116 );
nor ( n73671 , n600992 , n73670 );
xnor ( n600995 , n73671 , n66190 );
and ( n600996 , n73668 , n600995 );
xor ( n73674 , n73520 , n73524 );
xor ( n600998 , n73674 , n600852 );
and ( n600999 , n600995 , n600998 );
and ( n73677 , n73668 , n600998 );
or ( n601001 , n600996 , n600999 , n73677 );
and ( n73679 , n594952 , n594807 );
and ( n601003 , n594710 , n594804 );
nor ( n73681 , n73679 , n601003 );
xnor ( n601005 , n73681 , n66187 );
and ( n601006 , n601001 , n601005 );
xor ( n73684 , n600855 , n600859 );
xor ( n601008 , n73684 , n600862 );
and ( n601009 , n601005 , n601008 );
and ( n73687 , n601001 , n601008 );
or ( n73688 , n601006 , n601009 , n73687 );
xor ( n601012 , n600933 , n600937 );
xor ( n73690 , n601012 , n73617 );
and ( n601014 , n73688 , n73690 );
xor ( n73692 , n600865 , n73546 );
xor ( n73693 , n73692 , n73549 );
and ( n601017 , n73690 , n73693 );
and ( n73695 , n73688 , n73693 );
or ( n601019 , n601014 , n601017 , n73695 );
and ( n73697 , n600955 , n601019 );
xor ( n601021 , n600955 , n601019 );
xor ( n73699 , n73399 , n73403 );
and ( n73700 , n70652 , n592681 );
not ( n601024 , n73700 );
and ( n73702 , n601024 , n592475 );
and ( n601026 , n70652 , n592683 );
and ( n73704 , n597980 , n592681 );
nor ( n601028 , n601026 , n73704 );
xnor ( n601029 , n601028 , n592475 );
and ( n73707 , n73702 , n601029 );
and ( n601031 , n597980 , n592683 );
and ( n601032 , n70663 , n592681 );
nor ( n73710 , n601031 , n601032 );
xnor ( n73711 , n73710 , n592475 );
and ( n73712 , n73707 , n73711 );
and ( n73713 , n73711 , n73397 );
and ( n73714 , n73707 , n73397 );
or ( n73715 , n73712 , n73713 , n73714 );
and ( n73716 , n73699 , n73715 );
and ( n601040 , n70663 , n592683 );
and ( n601041 , n597996 , n592681 );
nor ( n73719 , n601040 , n601041 );
xnor ( n601043 , n73719 , n592475 );
and ( n601044 , n73715 , n601043 );
and ( n73722 , n73699 , n601043 );
or ( n601046 , n73716 , n601044 , n73722 );
and ( n601047 , n597996 , n592683 );
and ( n73725 , n70683 , n592681 );
nor ( n601049 , n601047 , n73725 );
xnor ( n601050 , n601049 , n592475 );
and ( n73728 , n601046 , n601050 );
xor ( n601052 , n600727 , n73408 );
xor ( n73730 , n601052 , n600387 );
and ( n601054 , n601050 , n73730 );
and ( n73732 , n601046 , n73730 );
or ( n601056 , n73728 , n601054 , n73732 );
and ( n73734 , n70683 , n592683 );
and ( n601058 , n70693 , n592681 );
nor ( n73736 , n73734 , n601058 );
xnor ( n73737 , n73736 , n592475 );
and ( n601061 , n601056 , n73737 );
xor ( n601062 , n600719 , n600735 );
xor ( n73740 , n601062 , n73417 );
and ( n601064 , n73737 , n73740 );
and ( n601065 , n601056 , n73740 );
or ( n73743 , n601061 , n601064 , n601065 );
and ( n601067 , n70693 , n592683 );
and ( n73745 , n70637 , n592681 );
nor ( n73746 , n601067 , n73745 );
xnor ( n601070 , n73746 , n592475 );
and ( n73748 , n73743 , n601070 );
xor ( n601072 , n600743 , n73424 );
xor ( n73750 , n601072 , n73427 );
and ( n73751 , n601070 , n73750 );
and ( n601075 , n73743 , n73750 );
or ( n601076 , n73748 , n73751 , n601075 );
and ( n73754 , n70637 , n592683 );
and ( n601078 , n70261 , n592681 );
nor ( n601079 , n73754 , n601078 );
xnor ( n73757 , n601079 , n592475 );
and ( n601081 , n601076 , n73757 );
xor ( n73759 , n600753 , n73434 );
xor ( n73760 , n73759 , n73437 );
and ( n601084 , n73757 , n73760 );
and ( n73762 , n601076 , n73760 );
or ( n73763 , n601081 , n601084 , n73762 );
and ( n73764 , n70261 , n592683 );
and ( n601088 , n70255 , n592681 );
nor ( n73766 , n73764 , n601088 );
xnor ( n73767 , n73766 , n592475 );
and ( n601091 , n73763 , n73767 );
xor ( n601092 , n600763 , n73444 );
xor ( n601093 , n601092 , n73447 );
and ( n73771 , n73767 , n601093 );
and ( n601095 , n73763 , n601093 );
or ( n601096 , n601091 , n73771 , n601095 );
and ( n73774 , n69739 , n593256 );
and ( n73775 , n69581 , n593254 );
nor ( n73776 , n73774 , n73775 );
xnor ( n73777 , n73776 , n65490 );
and ( n601101 , n601096 , n73777 );
xor ( n73779 , n73484 , n73488 );
xor ( n601103 , n73779 , n73491 );
and ( n73781 , n73777 , n601103 );
and ( n601105 , n601096 , n601103 );
or ( n601106 , n601101 , n73781 , n601105 );
and ( n73784 , n597402 , n593256 );
and ( n73785 , n597260 , n593254 );
nor ( n601109 , n73784 , n73785 );
xnor ( n601110 , n601109 , n65490 );
and ( n73788 , n70255 , n65592 );
and ( n601112 , n597569 , n592913 );
nor ( n601113 , n73788 , n601112 );
xnor ( n73791 , n601113 , n592638 );
and ( n601115 , n601110 , n73791 );
xor ( n601116 , n601076 , n73757 );
xor ( n73794 , n601116 , n73760 );
and ( n73795 , n73791 , n73794 );
and ( n601119 , n601110 , n73794 );
or ( n73797 , n601115 , n73795 , n601119 );
and ( n601121 , n597569 , n65592 );
and ( n73799 , n597402 , n592913 );
nor ( n73800 , n601121 , n73799 );
xnor ( n601124 , n73800 , n592638 );
and ( n73802 , n73797 , n601124 );
xor ( n601126 , n73763 , n73767 );
xor ( n73804 , n601126 , n601093 );
and ( n601128 , n601124 , n73804 );
and ( n601129 , n73797 , n73804 );
or ( n73807 , n73802 , n601128 , n601129 );
and ( n601131 , n69491 , n66142 );
and ( n601132 , n69283 , n66140 );
nor ( n601133 , n601131 , n601132 );
xnor ( n73811 , n601133 , n592960 );
and ( n601135 , n73807 , n73811 );
xor ( n601136 , n601096 , n73777 );
xor ( n73814 , n601136 , n601103 );
and ( n601138 , n73811 , n73814 );
and ( n601139 , n73807 , n73814 );
or ( n73817 , n601135 , n601138 , n601139 );
and ( n601141 , n601106 , n73817 );
xor ( n601142 , n73636 , n600963 );
xor ( n73820 , n601142 , n600966 );
and ( n601144 , n73817 , n73820 );
and ( n73822 , n601106 , n73820 );
or ( n601146 , n601141 , n601144 , n73822 );
and ( n601147 , n596193 , n66457 );
and ( n73825 , n596057 , n593778 );
nor ( n601149 , n601147 , n73825 );
xnor ( n73827 , n601149 , n593160 );
and ( n601151 , n601146 , n73827 );
xor ( n73829 , n73646 , n73650 );
xor ( n73830 , n73829 , n600976 );
and ( n601154 , n73827 , n73830 );
and ( n73832 , n601146 , n73830 );
or ( n601156 , n601151 , n601154 , n73832 );
and ( n73834 , n68160 , n594441 );
and ( n601158 , n67940 , n67116 );
nor ( n601159 , n73834 , n601158 );
xnor ( n73837 , n601159 , n66190 );
and ( n601161 , n601156 , n73837 );
xor ( n601162 , n73580 , n600907 );
xor ( n73840 , n601162 , n73587 );
and ( n73841 , n73837 , n73840 );
and ( n73842 , n601156 , n73840 );
or ( n73843 , n601161 , n73841 , n73842 );
and ( n73844 , n67636 , n594807 );
and ( n601168 , n594952 , n594804 );
nor ( n73846 , n73844 , n601168 );
xnor ( n601170 , n73846 , n66187 );
and ( n73848 , n73843 , n601170 );
xor ( n601172 , n600913 , n600917 );
xor ( n73850 , n601172 , n73597 );
and ( n601174 , n601170 , n73850 );
and ( n601175 , n73843 , n73850 );
or ( n73853 , n73848 , n601174 , n601175 );
xor ( n601177 , n73600 , n600927 );
xor ( n601178 , n601177 , n600930 );
and ( n73856 , n73853 , n601178 );
xor ( n601180 , n601001 , n601005 );
xor ( n601181 , n601180 , n601008 );
and ( n73859 , n601178 , n601181 );
and ( n601183 , n73853 , n601181 );
or ( n601184 , n73856 , n73859 , n601183 );
xor ( n73862 , n73688 , n73690 );
xor ( n73863 , n73862 , n73693 );
and ( n601187 , n601184 , n73863 );
xor ( n601188 , n601184 , n73863 );
xor ( n73866 , n73853 , n601178 );
xor ( n601190 , n73866 , n601181 );
and ( n73868 , n596198 , n66457 );
and ( n601192 , n596193 , n593778 );
nor ( n73870 , n73868 , n601192 );
xnor ( n601194 , n73870 , n593160 );
and ( n73872 , n69283 , n66142 );
and ( n73873 , n596600 , n66140 );
nor ( n601197 , n73872 , n73873 );
xnor ( n601198 , n601197 , n592960 );
and ( n73876 , n601194 , n601198 );
xor ( n601200 , n601106 , n73817 );
xor ( n601201 , n601200 , n73820 );
and ( n73879 , n601198 , n601201 );
and ( n601203 , n601194 , n601201 );
or ( n601204 , n73876 , n73879 , n601203 );
and ( n73882 , n595521 , n594441 );
and ( n73883 , n68160 , n67116 );
nor ( n601207 , n73882 , n73883 );
xnor ( n73885 , n601207 , n66190 );
and ( n601209 , n601204 , n73885 );
and ( n73887 , n595827 , n594210 );
and ( n73888 , n595633 , n66885 );
nor ( n601212 , n73887 , n73888 );
xnor ( n601213 , n601212 , n593434 );
and ( n73891 , n73885 , n601213 );
and ( n601215 , n601204 , n601213 );
or ( n601216 , n601209 , n73891 , n601215 );
and ( n73894 , n595103 , n594807 );
and ( n601218 , n67636 , n594804 );
nor ( n601219 , n73894 , n601218 );
xnor ( n601220 , n601219 , n66187 );
and ( n73898 , n601216 , n601220 );
xor ( n601222 , n600979 , n600983 );
xor ( n601223 , n601222 , n73665 );
and ( n73901 , n601220 , n601223 );
and ( n601225 , n601216 , n601223 );
or ( n601226 , n73898 , n73901 , n601225 );
xor ( n73904 , n73668 , n600995 );
xor ( n601228 , n73904 , n600998 );
and ( n601229 , n601226 , n601228 );
xor ( n73907 , n73843 , n601170 );
xor ( n601231 , n73907 , n73850 );
and ( n601232 , n601228 , n601231 );
and ( n73910 , n601226 , n601231 );
or ( n601234 , n601229 , n601232 , n73910 );
and ( n73912 , n601190 , n601234 );
xor ( n601236 , n601190 , n601234 );
xor ( n73914 , n601226 , n601228 );
xor ( n601238 , n73914 , n601231 );
and ( n73916 , n69581 , n66142 );
and ( n73917 , n69491 , n66140 );
nor ( n601241 , n73916 , n73917 );
xnor ( n601242 , n601241 , n592960 );
and ( n73920 , n597260 , n593256 );
and ( n601244 , n69739 , n593254 );
nor ( n601245 , n73920 , n601244 );
xnor ( n73923 , n601245 , n65490 );
and ( n601247 , n601242 , n73923 );
xor ( n601248 , n73797 , n601124 );
xor ( n73926 , n601248 , n73804 );
and ( n73927 , n73923 , n73926 );
and ( n601251 , n601242 , n73926 );
or ( n73929 , n601247 , n73927 , n601251 );
and ( n601253 , n596600 , n66457 );
and ( n73931 , n596198 , n593778 );
nor ( n73932 , n601253 , n73931 );
xnor ( n601256 , n73932 , n593160 );
and ( n601257 , n73929 , n601256 );
xor ( n73935 , n73807 , n73811 );
xor ( n601259 , n73935 , n73814 );
and ( n601260 , n601256 , n601259 );
and ( n73938 , n73929 , n601259 );
or ( n601262 , n601257 , n601260 , n73938 );
and ( n601263 , n595633 , n594441 );
and ( n601264 , n595521 , n67116 );
nor ( n73942 , n601263 , n601264 );
xnor ( n601266 , n73942 , n66190 );
and ( n601267 , n601262 , n601266 );
and ( n73945 , n596057 , n594210 );
and ( n601269 , n595827 , n66885 );
nor ( n601270 , n73945 , n601269 );
xnor ( n73948 , n601270 , n593434 );
and ( n601272 , n601266 , n73948 );
and ( n73950 , n601262 , n73948 );
or ( n73951 , n601267 , n601272 , n73950 );
and ( n601275 , n67940 , n594807 );
and ( n601276 , n595103 , n594804 );
nor ( n73954 , n601275 , n601276 );
xnor ( n601278 , n73954 , n66187 );
and ( n601279 , n73951 , n601278 );
xor ( n73957 , n601146 , n73827 );
xor ( n601281 , n73957 , n73830 );
and ( n601282 , n601278 , n601281 );
and ( n73960 , n73951 , n601281 );
or ( n601284 , n601279 , n601282 , n73960 );
xor ( n601285 , n601216 , n601220 );
xor ( n73963 , n601285 , n601223 );
and ( n601287 , n601284 , n73963 );
xor ( n73965 , n601156 , n73837 );
xor ( n73966 , n73965 , n73840 );
and ( n601290 , n73963 , n73966 );
and ( n73968 , n601284 , n73966 );
or ( n601292 , n601287 , n601290 , n73968 );
and ( n73970 , n601238 , n601292 );
xor ( n73971 , n601238 , n601292 );
xor ( n73972 , n73702 , n601029 );
and ( n601296 , n70652 , n592913 );
not ( n601297 , n601296 );
and ( n73975 , n601297 , n592638 );
and ( n601299 , n70652 , n65592 );
and ( n601300 , n597980 , n592913 );
nor ( n73978 , n601299 , n601300 );
xnor ( n601302 , n73978 , n592638 );
and ( n601303 , n73975 , n601302 );
and ( n601304 , n597980 , n65592 );
and ( n73982 , n70663 , n592913 );
nor ( n73983 , n601304 , n73982 );
xnor ( n601307 , n73983 , n592638 );
and ( n73985 , n601303 , n601307 );
and ( n601309 , n601307 , n73700 );
and ( n73987 , n601303 , n73700 );
or ( n601311 , n73985 , n601309 , n73987 );
and ( n73989 , n73972 , n601311 );
and ( n73990 , n70663 , n65592 );
and ( n601314 , n597996 , n592913 );
nor ( n73992 , n73990 , n601314 );
xnor ( n601316 , n73992 , n592638 );
and ( n601317 , n601311 , n601316 );
and ( n601318 , n73972 , n601316 );
or ( n73996 , n73989 , n601317 , n601318 );
and ( n601320 , n597996 , n65592 );
and ( n73998 , n70683 , n592913 );
nor ( n601322 , n601320 , n73998 );
xnor ( n601323 , n601322 , n592638 );
and ( n74001 , n73996 , n601323 );
xor ( n601325 , n73707 , n73711 );
xor ( n601326 , n601325 , n73397 );
and ( n74004 , n601323 , n601326 );
and ( n74005 , n73996 , n601326 );
or ( n601329 , n74001 , n74004 , n74005 );
and ( n74007 , n70683 , n65592 );
and ( n74008 , n70693 , n592913 );
nor ( n601332 , n74007 , n74008 );
xnor ( n601333 , n601332 , n592638 );
and ( n74011 , n601329 , n601333 );
xor ( n601335 , n73699 , n73715 );
xor ( n601336 , n601335 , n601043 );
and ( n601337 , n601333 , n601336 );
and ( n74015 , n601329 , n601336 );
or ( n601339 , n74011 , n601337 , n74015 );
and ( n601340 , n70693 , n65592 );
and ( n74018 , n70637 , n592913 );
nor ( n74019 , n601340 , n74018 );
xnor ( n74020 , n74019 , n592638 );
and ( n74021 , n601339 , n74020 );
xor ( n74022 , n601046 , n601050 );
xor ( n74023 , n74022 , n73730 );
and ( n74024 , n74020 , n74023 );
and ( n74025 , n601339 , n74023 );
or ( n74026 , n74021 , n74024 , n74025 );
and ( n74027 , n70637 , n65592 );
and ( n74028 , n70261 , n592913 );
nor ( n74029 , n74027 , n74028 );
xnor ( n74030 , n74029 , n592638 );
and ( n74031 , n74026 , n74030 );
xor ( n74032 , n601056 , n73737 );
xor ( n74033 , n74032 , n73740 );
and ( n74034 , n74030 , n74033 );
and ( n74035 , n74026 , n74033 );
or ( n74036 , n74031 , n74034 , n74035 );
and ( n74037 , n70261 , n65592 );
and ( n74038 , n70255 , n592913 );
nor ( n74039 , n74037 , n74038 );
xnor ( n74040 , n74039 , n592638 );
and ( n74041 , n74036 , n74040 );
xor ( n74042 , n73743 , n601070 );
xor ( n74043 , n74042 , n73750 );
and ( n74044 , n74040 , n74043 );
and ( n74045 , n74036 , n74043 );
or ( n74046 , n74041 , n74044 , n74045 );
and ( n74047 , n69739 , n66142 );
and ( n74048 , n69581 , n66140 );
nor ( n74049 , n74047 , n74048 );
xnor ( n74050 , n74049 , n592960 );
and ( n74051 , n74046 , n74050 );
xor ( n74052 , n601110 , n73791 );
xor ( n74053 , n74052 , n73794 );
and ( n74054 , n74050 , n74053 );
and ( n74055 , n74046 , n74053 );
or ( n74056 , n74051 , n74054 , n74055 );
and ( n601380 , n69283 , n66457 );
and ( n74058 , n596600 , n593778 );
nor ( n601382 , n601380 , n74058 );
xnor ( n74060 , n601382 , n593160 );
and ( n74061 , n74056 , n74060 );
xor ( n74062 , n601242 , n73923 );
xor ( n74063 , n74062 , n73926 );
and ( n74064 , n74060 , n74063 );
and ( n74065 , n74056 , n74063 );
or ( n74066 , n74061 , n74064 , n74065 );
and ( n74067 , n596193 , n594210 );
and ( n74068 , n596057 , n66885 );
nor ( n74069 , n74067 , n74068 );
xnor ( n74070 , n74069 , n593434 );
and ( n74071 , n74066 , n74070 );
xor ( n74072 , n73929 , n601256 );
xor ( n74073 , n74072 , n601259 );
and ( n74074 , n74070 , n74073 );
and ( n74075 , n74066 , n74073 );
or ( n74076 , n74071 , n74074 , n74075 );
and ( n74077 , n68160 , n594807 );
and ( n74078 , n67940 , n594804 );
nor ( n74079 , n74077 , n74078 );
xnor ( n601403 , n74079 , n66187 );
and ( n74081 , n74076 , n601403 );
xor ( n601405 , n601194 , n601198 );
xor ( n601406 , n601405 , n601201 );
and ( n74084 , n601403 , n601406 );
and ( n601408 , n74076 , n601406 );
or ( n601409 , n74081 , n74084 , n601408 );
xor ( n601410 , n601204 , n73885 );
xor ( n74088 , n601410 , n601213 );
and ( n601412 , n601409 , n74088 );
xor ( n74090 , n73951 , n601278 );
xor ( n74091 , n74090 , n601281 );
and ( n74092 , n74088 , n74091 );
and ( n601416 , n601409 , n74091 );
or ( n74094 , n601412 , n74092 , n601416 );
xor ( n601418 , n601284 , n73963 );
xor ( n74096 , n601418 , n73966 );
and ( n601420 , n74094 , n74096 );
xor ( n74098 , n74094 , n74096 );
xor ( n601422 , n601409 , n74088 );
xor ( n74100 , n601422 , n74091 );
and ( n601424 , n597402 , n66142 );
and ( n601425 , n597260 , n66140 );
nor ( n74103 , n601424 , n601425 );
xnor ( n74104 , n74103 , n592960 );
and ( n74105 , n70255 , n593256 );
and ( n601429 , n597569 , n593254 );
nor ( n74107 , n74105 , n601429 );
xnor ( n601431 , n74107 , n65490 );
and ( n601432 , n74104 , n601431 );
xor ( n74110 , n74026 , n74030 );
xor ( n74111 , n74110 , n74033 );
and ( n601435 , n601431 , n74111 );
and ( n74113 , n74104 , n74111 );
or ( n601437 , n601432 , n601435 , n74113 );
and ( n601438 , n597569 , n593256 );
and ( n74116 , n597402 , n593254 );
nor ( n74117 , n601438 , n74116 );
xnor ( n601441 , n74117 , n65490 );
and ( n74119 , n601437 , n601441 );
xor ( n74120 , n74036 , n74040 );
xor ( n601444 , n74120 , n74043 );
and ( n601445 , n601441 , n601444 );
and ( n74123 , n601437 , n601444 );
or ( n601447 , n74119 , n601445 , n74123 );
and ( n601448 , n69491 , n66457 );
and ( n74126 , n69283 , n593778 );
nor ( n601450 , n601448 , n74126 );
xnor ( n601451 , n601450 , n593160 );
and ( n74129 , n601447 , n601451 );
xor ( n74130 , n74046 , n74050 );
xor ( n601454 , n74130 , n74053 );
and ( n74132 , n601451 , n601454 );
and ( n601456 , n601447 , n601454 );
or ( n601457 , n74129 , n74132 , n601456 );
and ( n74135 , n596198 , n594210 );
and ( n601459 , n596193 , n66885 );
nor ( n601460 , n74135 , n601459 );
xnor ( n601461 , n601460 , n593434 );
and ( n74139 , n601457 , n601461 );
xor ( n601463 , n74056 , n74060 );
xor ( n601464 , n601463 , n74063 );
and ( n74142 , n601461 , n601464 );
and ( n601466 , n601457 , n601464 );
or ( n601467 , n74139 , n74142 , n601466 );
and ( n601468 , n595521 , n594807 );
and ( n74146 , n68160 , n594804 );
nor ( n601470 , n601468 , n74146 );
xnor ( n601471 , n601470 , n66187 );
and ( n74149 , n601467 , n601471 );
and ( n601473 , n595827 , n594441 );
and ( n601474 , n595633 , n67116 );
nor ( n74152 , n601473 , n601474 );
xnor ( n601476 , n74152 , n66190 );
and ( n601477 , n601471 , n601476 );
and ( n601478 , n601467 , n601476 );
or ( n74156 , n74149 , n601477 , n601478 );
xor ( n601480 , n601262 , n601266 );
xor ( n74158 , n601480 , n73948 );
and ( n601482 , n74156 , n74158 );
xor ( n74160 , n74076 , n601403 );
xor ( n74161 , n74160 , n601406 );
and ( n601485 , n74158 , n74161 );
and ( n601486 , n74156 , n74161 );
or ( n74164 , n601482 , n601485 , n601486 );
and ( n601488 , n74100 , n74164 );
xor ( n601489 , n74100 , n74164 );
xor ( n74167 , n74156 , n74158 );
xor ( n601491 , n74167 , n74161 );
and ( n601492 , n69581 , n66457 );
and ( n74170 , n69491 , n593778 );
nor ( n74171 , n601492 , n74170 );
xnor ( n601495 , n74171 , n593160 );
and ( n74173 , n597260 , n66142 );
and ( n601497 , n69739 , n66140 );
nor ( n74175 , n74173 , n601497 );
xnor ( n74176 , n74175 , n592960 );
and ( n601500 , n601495 , n74176 );
xor ( n601501 , n601437 , n601441 );
xor ( n74179 , n601501 , n601444 );
and ( n601503 , n74176 , n74179 );
and ( n601504 , n601495 , n74179 );
or ( n74182 , n601500 , n601503 , n601504 );
and ( n601506 , n596193 , n594441 );
and ( n601507 , n596057 , n67116 );
nor ( n601508 , n601506 , n601507 );
xnor ( n74186 , n601508 , n66190 );
and ( n601510 , n74182 , n74186 );
xor ( n601511 , n601447 , n601451 );
xor ( n74189 , n601511 , n601454 );
and ( n601513 , n74186 , n74189 );
and ( n601514 , n74182 , n74189 );
or ( n74192 , n601510 , n601513 , n601514 );
and ( n601516 , n595633 , n594807 );
and ( n74194 , n595521 , n594804 );
nor ( n74195 , n601516 , n74194 );
xnor ( n74196 , n74195 , n66187 );
and ( n74197 , n74192 , n74196 );
and ( n74198 , n596057 , n594441 );
and ( n601522 , n595827 , n67116 );
nor ( n74200 , n74198 , n601522 );
xnor ( n74201 , n74200 , n66190 );
and ( n601525 , n74196 , n74201 );
and ( n601526 , n74192 , n74201 );
or ( n74204 , n74197 , n601525 , n601526 );
xor ( n601528 , n601467 , n601471 );
xor ( n601529 , n601528 , n601476 );
and ( n74207 , n74204 , n601529 );
xor ( n601531 , n74066 , n74070 );
xor ( n601532 , n601531 , n74073 );
and ( n74210 , n601529 , n601532 );
and ( n601534 , n74204 , n601532 );
or ( n74212 , n74207 , n74210 , n601534 );
and ( n601536 , n601491 , n74212 );
xor ( n74214 , n601491 , n74212 );
xor ( n601538 , n73975 , n601302 );
and ( n601539 , n70652 , n593254 );
not ( n601540 , n601539 );
and ( n74218 , n601540 , n65490 );
and ( n601542 , n70652 , n593256 );
and ( n74220 , n597980 , n593254 );
nor ( n601544 , n601542 , n74220 );
xnor ( n74222 , n601544 , n65490 );
and ( n74223 , n74218 , n74222 );
and ( n601547 , n597980 , n593256 );
and ( n74225 , n70663 , n593254 );
nor ( n601549 , n601547 , n74225 );
xnor ( n74227 , n601549 , n65490 );
and ( n601551 , n74223 , n74227 );
and ( n601552 , n74227 , n601296 );
and ( n74230 , n74223 , n601296 );
or ( n601554 , n601551 , n601552 , n74230 );
and ( n601555 , n601538 , n601554 );
and ( n74233 , n70663 , n593256 );
and ( n74234 , n597996 , n593254 );
nor ( n601558 , n74233 , n74234 );
xnor ( n601559 , n601558 , n65490 );
and ( n74237 , n601554 , n601559 );
and ( n601561 , n601538 , n601559 );
or ( n601562 , n601555 , n74237 , n601561 );
and ( n74240 , n597996 , n593256 );
and ( n601564 , n70683 , n593254 );
nor ( n601565 , n74240 , n601564 );
xnor ( n74243 , n601565 , n65490 );
and ( n601567 , n601562 , n74243 );
xor ( n74245 , n601303 , n601307 );
xor ( n601569 , n74245 , n73700 );
and ( n74247 , n74243 , n601569 );
and ( n601571 , n601562 , n601569 );
or ( n601572 , n601567 , n74247 , n601571 );
and ( n74250 , n70683 , n593256 );
and ( n74251 , n70693 , n593254 );
nor ( n601575 , n74250 , n74251 );
xnor ( n74253 , n601575 , n65490 );
and ( n74254 , n601572 , n74253 );
xor ( n601578 , n73972 , n601311 );
xor ( n601579 , n601578 , n601316 );
and ( n74257 , n74253 , n601579 );
and ( n74258 , n601572 , n601579 );
or ( n601582 , n74254 , n74257 , n74258 );
and ( n74260 , n70693 , n593256 );
and ( n601584 , n70637 , n593254 );
nor ( n74262 , n74260 , n601584 );
xnor ( n601586 , n74262 , n65490 );
and ( n74264 , n601582 , n601586 );
xor ( n601588 , n73996 , n601323 );
xor ( n74266 , n601588 , n601326 );
and ( n601590 , n601586 , n74266 );
and ( n74268 , n601582 , n74266 );
or ( n601592 , n74264 , n601590 , n74268 );
and ( n601593 , n70637 , n593256 );
and ( n601594 , n70261 , n593254 );
nor ( n74272 , n601593 , n601594 );
xnor ( n601596 , n74272 , n65490 );
and ( n74274 , n601592 , n601596 );
xor ( n601598 , n601329 , n601333 );
xor ( n74276 , n601598 , n601336 );
and ( n74277 , n601596 , n74276 );
and ( n601601 , n601592 , n74276 );
or ( n74279 , n74274 , n74277 , n601601 );
and ( n601603 , n70261 , n593256 );
and ( n74281 , n70255 , n593254 );
nor ( n601605 , n601603 , n74281 );
xnor ( n601606 , n601605 , n65490 );
and ( n74284 , n74279 , n601606 );
xor ( n74285 , n601339 , n74020 );
xor ( n601609 , n74285 , n74023 );
and ( n601610 , n601606 , n601609 );
and ( n74288 , n74279 , n601609 );
or ( n601612 , n74284 , n601610 , n74288 );
and ( n601613 , n69739 , n66457 );
and ( n74291 , n69581 , n593778 );
nor ( n601615 , n601613 , n74291 );
xnor ( n601616 , n601615 , n593160 );
and ( n601617 , n601612 , n601616 );
xor ( n74295 , n74104 , n601431 );
xor ( n601619 , n74295 , n74111 );
and ( n601620 , n601616 , n601619 );
and ( n74298 , n601612 , n601619 );
or ( n601622 , n601617 , n601620 , n74298 );
and ( n601623 , n69283 , n594210 );
and ( n74301 , n596600 , n66885 );
nor ( n601625 , n601623 , n74301 );
xnor ( n74303 , n601625 , n593434 );
and ( n601627 , n601622 , n74303 );
xor ( n74305 , n601495 , n74176 );
xor ( n601629 , n74305 , n74179 );
and ( n74307 , n74303 , n601629 );
and ( n601631 , n601622 , n601629 );
or ( n74309 , n601627 , n74307 , n601631 );
and ( n74310 , n595827 , n594807 );
and ( n601634 , n595633 , n594804 );
nor ( n74312 , n74310 , n601634 );
xnor ( n601636 , n74312 , n66187 );
and ( n601637 , n74309 , n601636 );
and ( n601638 , n596600 , n594210 );
and ( n74316 , n596198 , n66885 );
nor ( n601640 , n601638 , n74316 );
xnor ( n74318 , n601640 , n593434 );
and ( n601642 , n601636 , n74318 );
and ( n74320 , n74309 , n74318 );
or ( n601644 , n601637 , n601642 , n74320 );
xor ( n74322 , n74192 , n74196 );
xor ( n74323 , n74322 , n74201 );
and ( n601647 , n601644 , n74323 );
xor ( n74325 , n601457 , n601461 );
xor ( n601649 , n74325 , n601464 );
and ( n601650 , n74323 , n601649 );
and ( n74328 , n601644 , n601649 );
or ( n601652 , n601647 , n601650 , n74328 );
xor ( n74330 , n74204 , n601529 );
xor ( n74331 , n74330 , n601532 );
and ( n601655 , n601652 , n74331 );
xor ( n74333 , n601652 , n74331 );
xor ( n601657 , n601644 , n74323 );
xor ( n74335 , n601657 , n601649 );
and ( n74336 , n597402 , n66457 );
and ( n601660 , n597260 , n593778 );
nor ( n601661 , n74336 , n601660 );
xnor ( n74339 , n601661 , n593160 );
and ( n601663 , n70255 , n66142 );
and ( n74341 , n597569 , n66140 );
nor ( n74342 , n601663 , n74341 );
xnor ( n601666 , n74342 , n592960 );
and ( n601667 , n74339 , n601666 );
xor ( n74345 , n601592 , n601596 );
xor ( n601669 , n74345 , n74276 );
and ( n601670 , n601666 , n601669 );
and ( n74348 , n74339 , n601669 );
or ( n601672 , n601667 , n601670 , n74348 );
and ( n601673 , n597569 , n66142 );
and ( n74351 , n597402 , n66140 );
nor ( n601675 , n601673 , n74351 );
xnor ( n601676 , n601675 , n592960 );
and ( n74354 , n601672 , n601676 );
xor ( n601678 , n74279 , n601606 );
xor ( n601679 , n601678 , n601609 );
and ( n74357 , n601676 , n601679 );
and ( n601681 , n601672 , n601679 );
or ( n74359 , n74354 , n74357 , n601681 );
and ( n601683 , n69491 , n594210 );
and ( n601684 , n69283 , n66885 );
nor ( n74362 , n601683 , n601684 );
xnor ( n601686 , n74362 , n593434 );
and ( n601687 , n74359 , n601686 );
xor ( n74365 , n601612 , n601616 );
xor ( n74366 , n74365 , n601619 );
and ( n601690 , n601686 , n74366 );
and ( n601691 , n74359 , n74366 );
or ( n74369 , n601687 , n601690 , n601691 );
and ( n74370 , n596198 , n594441 );
and ( n601694 , n596193 , n67116 );
nor ( n74372 , n74370 , n601694 );
xnor ( n74373 , n74372 , n66190 );
and ( n74374 , n74369 , n74373 );
xor ( n74375 , n601622 , n74303 );
xor ( n74376 , n74375 , n601629 );
and ( n74377 , n74373 , n74376 );
and ( n74378 , n74369 , n74376 );
or ( n74379 , n74374 , n74377 , n74378 );
xor ( n601703 , n74309 , n601636 );
xor ( n74381 , n601703 , n74318 );
and ( n601705 , n74379 , n74381 );
xor ( n601706 , n74182 , n74186 );
xor ( n601707 , n601706 , n74189 );
and ( n74385 , n74381 , n601707 );
and ( n601709 , n74379 , n601707 );
or ( n74387 , n601705 , n74385 , n601709 );
and ( n74388 , n74335 , n74387 );
xor ( n74389 , n74335 , n74387 );
xor ( n74390 , n74379 , n74381 );
xor ( n601714 , n74390 , n601707 );
and ( n74392 , n69581 , n594210 );
and ( n601716 , n69491 , n66885 );
nor ( n601717 , n74392 , n601716 );
xnor ( n74395 , n601717 , n593434 );
and ( n601719 , n597260 , n66457 );
and ( n74397 , n69739 , n593778 );
nor ( n601721 , n601719 , n74397 );
xnor ( n601722 , n601721 , n593160 );
and ( n74400 , n74395 , n601722 );
xor ( n74401 , n601672 , n601676 );
xor ( n601725 , n74401 , n601679 );
and ( n601726 , n601722 , n601725 );
and ( n74404 , n74395 , n601725 );
or ( n74405 , n74400 , n601726 , n74404 );
and ( n601729 , n596193 , n594807 );
and ( n74407 , n596057 , n594804 );
nor ( n601731 , n601729 , n74407 );
xnor ( n601732 , n601731 , n66187 );
and ( n74410 , n74405 , n601732 );
xor ( n74411 , n74359 , n601686 );
xor ( n601735 , n74411 , n74366 );
and ( n601736 , n601732 , n601735 );
and ( n601737 , n74405 , n601735 );
or ( n74415 , n74410 , n601736 , n601737 );
and ( n74416 , n596057 , n594807 );
and ( n601740 , n595827 , n594804 );
nor ( n601741 , n74416 , n601740 );
xnor ( n74419 , n601741 , n66187 );
and ( n601743 , n74415 , n74419 );
xor ( n601744 , n74369 , n74373 );
xor ( n74422 , n601744 , n74376 );
and ( n74423 , n74419 , n74422 );
and ( n601747 , n74415 , n74422 );
or ( n74425 , n601743 , n74423 , n601747 );
and ( n601749 , n601714 , n74425 );
xor ( n74427 , n601714 , n74425 );
and ( n74428 , n597569 , n66457 );
and ( n601752 , n597402 , n593778 );
nor ( n601753 , n74428 , n601752 );
xnor ( n74431 , n601753 , n593160 );
and ( n74432 , n70261 , n66142 );
and ( n601756 , n70255 , n66140 );
nor ( n601757 , n74432 , n601756 );
xnor ( n74435 , n601757 , n592960 );
and ( n74436 , n74431 , n74435 );
xor ( n601760 , n601582 , n601586 );
xor ( n601761 , n601760 , n74266 );
and ( n601762 , n74435 , n601761 );
and ( n601763 , n74431 , n601761 );
or ( n74441 , n74436 , n601762 , n601763 );
and ( n601765 , n69739 , n594210 );
and ( n74443 , n69581 , n66885 );
nor ( n74444 , n601765 , n74443 );
xnor ( n601768 , n74444 , n593434 );
and ( n74446 , n74441 , n601768 );
xor ( n74447 , n74339 , n601666 );
xor ( n601771 , n74447 , n601669 );
and ( n601772 , n601768 , n601771 );
and ( n74450 , n74441 , n601771 );
or ( n601774 , n74446 , n601772 , n74450 );
and ( n601775 , n69283 , n594441 );
and ( n74453 , n596600 , n67116 );
nor ( n601777 , n601775 , n74453 );
xnor ( n601778 , n601777 , n66190 );
and ( n74456 , n601774 , n601778 );
xor ( n601780 , n74395 , n601722 );
xor ( n74458 , n601780 , n601725 );
and ( n601782 , n601778 , n74458 );
and ( n601783 , n601774 , n74458 );
or ( n74461 , n74456 , n601782 , n601783 );
and ( n601785 , n596600 , n594441 );
and ( n74463 , n596198 , n67116 );
nor ( n74464 , n601785 , n74463 );
xnor ( n74465 , n74464 , n66190 );
and ( n74466 , n74461 , n74465 );
xor ( n74467 , n74405 , n601732 );
xor ( n74468 , n74467 , n601735 );
and ( n74469 , n74465 , n74468 );
and ( n74470 , n74461 , n74468 );
or ( n74471 , n74466 , n74469 , n74470 );
xor ( n74472 , n74415 , n74419 );
xor ( n74473 , n74472 , n74422 );
and ( n74474 , n74471 , n74473 );
xor ( n74475 , n74471 , n74473 );
xor ( n74476 , n74461 , n74465 );
xor ( n74477 , n74476 , n74468 );
xor ( n74478 , n74218 , n74222 );
and ( n74479 , n70652 , n66140 );
not ( n74480 , n74479 );
and ( n74481 , n74480 , n592960 );
and ( n74482 , n70652 , n66142 );
and ( n601806 , n597980 , n66140 );
nor ( n601807 , n74482 , n601806 );
xnor ( n74485 , n601807 , n592960 );
and ( n601809 , n74481 , n74485 );
and ( n74487 , n597980 , n66142 );
and ( n74488 , n70663 , n66140 );
nor ( n74489 , n74487 , n74488 );
xnor ( n74490 , n74489 , n592960 );
and ( n74491 , n601809 , n74490 );
and ( n74492 , n74490 , n601539 );
and ( n74493 , n601809 , n601539 );
or ( n74494 , n74491 , n74492 , n74493 );
and ( n74495 , n74478 , n74494 );
and ( n74496 , n70663 , n66142 );
and ( n74497 , n597996 , n66140 );
nor ( n74498 , n74496 , n74497 );
xnor ( n74499 , n74498 , n592960 );
and ( n74500 , n74494 , n74499 );
and ( n74501 , n74478 , n74499 );
or ( n74502 , n74495 , n74500 , n74501 );
and ( n74503 , n597996 , n66142 );
and ( n74504 , n70683 , n66140 );
nor ( n74505 , n74503 , n74504 );
xnor ( n74506 , n74505 , n592960 );
and ( n74507 , n74502 , n74506 );
xor ( n74508 , n74223 , n74227 );
xor ( n74509 , n74508 , n601296 );
and ( n74510 , n74506 , n74509 );
and ( n74511 , n74502 , n74509 );
or ( n74512 , n74507 , n74510 , n74511 );
and ( n74513 , n70683 , n66142 );
and ( n74514 , n70693 , n66140 );
nor ( n74515 , n74513 , n74514 );
xnor ( n74516 , n74515 , n592960 );
and ( n74517 , n74512 , n74516 );
xor ( n74518 , n601538 , n601554 );
xor ( n74519 , n74518 , n601559 );
and ( n74520 , n74516 , n74519 );
and ( n74521 , n74512 , n74519 );
or ( n74522 , n74517 , n74520 , n74521 );
and ( n74523 , n70693 , n66142 );
and ( n74524 , n70637 , n66140 );
nor ( n74525 , n74523 , n74524 );
xnor ( n601849 , n74525 , n592960 );
and ( n74527 , n74522 , n601849 );
xor ( n601851 , n601562 , n74243 );
xor ( n74529 , n601851 , n601569 );
and ( n74530 , n601849 , n74529 );
and ( n601854 , n74522 , n74529 );
or ( n74532 , n74527 , n74530 , n601854 );
and ( n74533 , n70637 , n66142 );
and ( n601857 , n70261 , n66140 );
nor ( n74535 , n74533 , n601857 );
xnor ( n74536 , n74535 , n592960 );
and ( n601860 , n74532 , n74536 );
xor ( n601861 , n601572 , n74253 );
xor ( n74539 , n601861 , n601579 );
and ( n601863 , n74536 , n74539 );
and ( n601864 , n74532 , n74539 );
or ( n74542 , n601860 , n601863 , n601864 );
and ( n601866 , n597402 , n594210 );
and ( n601867 , n597260 , n66885 );
nor ( n601868 , n601866 , n601867 );
xnor ( n74546 , n601868 , n593434 );
and ( n601870 , n70255 , n66457 );
and ( n601871 , n597569 , n593778 );
nor ( n74549 , n601870 , n601871 );
xnor ( n601873 , n74549 , n593160 );
and ( n74551 , n74546 , n601873 );
xor ( n74552 , n74532 , n74536 );
xor ( n74553 , n74552 , n74539 );
and ( n601877 , n601873 , n74553 );
and ( n74555 , n74546 , n74553 );
or ( n601879 , n74551 , n601877 , n74555 );
and ( n74557 , n74542 , n601879 );
xor ( n601881 , n74431 , n74435 );
xor ( n74559 , n601881 , n601761 );
and ( n74560 , n601879 , n74559 );
and ( n601884 , n74542 , n74559 );
or ( n601885 , n74557 , n74560 , n601884 );
and ( n74563 , n69491 , n594441 );
and ( n601887 , n69283 , n67116 );
nor ( n601888 , n74563 , n601887 );
xnor ( n74566 , n601888 , n66190 );
and ( n601890 , n601885 , n74566 );
xor ( n74568 , n74441 , n601768 );
xor ( n601892 , n74568 , n601771 );
and ( n74570 , n74566 , n601892 );
and ( n601894 , n601885 , n601892 );
or ( n601895 , n601890 , n74570 , n601894 );
and ( n74573 , n596198 , n594807 );
and ( n74574 , n596193 , n594804 );
nor ( n601898 , n74573 , n74574 );
xnor ( n74576 , n601898 , n66187 );
and ( n601900 , n601895 , n74576 );
xor ( n601901 , n601774 , n601778 );
xor ( n74579 , n601901 , n74458 );
and ( n74580 , n74576 , n74579 );
and ( n601904 , n601895 , n74579 );
or ( n601905 , n601900 , n74580 , n601904 );
and ( n601906 , n74477 , n601905 );
xor ( n74584 , n74477 , n601905 );
and ( n74585 , n69581 , n594441 );
and ( n74586 , n69491 , n67116 );
nor ( n74587 , n74585 , n74586 );
xnor ( n74588 , n74587 , n66190 );
and ( n74589 , n597260 , n594210 );
and ( n601913 , n69739 , n66885 );
nor ( n74591 , n74589 , n601913 );
xnor ( n74592 , n74591 , n593434 );
and ( n601916 , n74588 , n74592 );
xor ( n74594 , n74542 , n601879 );
xor ( n601918 , n74594 , n74559 );
and ( n74596 , n74592 , n601918 );
and ( n74597 , n74588 , n601918 );
or ( n601921 , n601916 , n74596 , n74597 );
and ( n601922 , n596600 , n594807 );
and ( n74600 , n596198 , n594804 );
nor ( n601924 , n601922 , n74600 );
xnor ( n601925 , n601924 , n66187 );
and ( n74603 , n601921 , n601925 );
xor ( n601927 , n601885 , n74566 );
xor ( n601928 , n601927 , n601892 );
and ( n601929 , n601925 , n601928 );
and ( n74607 , n601921 , n601928 );
or ( n601931 , n74603 , n601929 , n74607 );
xor ( n601932 , n601895 , n74576 );
xor ( n74610 , n601932 , n74579 );
and ( n601934 , n601931 , n74610 );
xor ( n601935 , n601931 , n74610 );
xor ( n74613 , n601921 , n601925 );
xor ( n74614 , n74613 , n601928 );
and ( n74615 , n597569 , n594210 );
and ( n74616 , n597402 , n66885 );
nor ( n74617 , n74615 , n74616 );
xnor ( n74618 , n74617 , n593434 );
and ( n74619 , n70261 , n66457 );
and ( n74620 , n70255 , n593778 );
nor ( n601944 , n74619 , n74620 );
xnor ( n74622 , n601944 , n593160 );
and ( n601946 , n74618 , n74622 );
xor ( n74624 , n74522 , n601849 );
xor ( n74625 , n74624 , n74529 );
and ( n601949 , n74622 , n74625 );
and ( n601950 , n74618 , n74625 );
or ( n74628 , n601946 , n601949 , n601950 );
and ( n601952 , n69739 , n594441 );
and ( n601953 , n69581 , n67116 );
nor ( n74631 , n601952 , n601953 );
xnor ( n601955 , n74631 , n66190 );
and ( n601956 , n74628 , n601955 );
xor ( n601957 , n74546 , n601873 );
xor ( n74635 , n601957 , n74553 );
and ( n601959 , n601955 , n74635 );
and ( n74637 , n74628 , n74635 );
or ( n74638 , n601956 , n601959 , n74637 );
xor ( n74639 , n74481 , n74485 );
and ( n74640 , n70652 , n593778 );
not ( n74641 , n74640 );
and ( n74642 , n74641 , n593160 );
and ( n74643 , n70652 , n66457 );
and ( n74644 , n597980 , n593778 );
nor ( n74645 , n74643 , n74644 );
xnor ( n74646 , n74645 , n593160 );
and ( n74647 , n74642 , n74646 );
and ( n601971 , n597980 , n66457 );
and ( n601972 , n70663 , n593778 );
nor ( n601973 , n601971 , n601972 );
xnor ( n74651 , n601973 , n593160 );
and ( n74652 , n74647 , n74651 );
and ( n601976 , n74651 , n74479 );
and ( n74654 , n74647 , n74479 );
or ( n74655 , n74652 , n601976 , n74654 );
and ( n601979 , n74639 , n74655 );
and ( n601980 , n70663 , n66457 );
and ( n74658 , n597996 , n593778 );
nor ( n601982 , n601980 , n74658 );
xnor ( n601983 , n601982 , n593160 );
and ( n74661 , n74655 , n601983 );
and ( n601985 , n74639 , n601983 );
or ( n74663 , n601979 , n74661 , n601985 );
and ( n74664 , n597996 , n66457 );
and ( n601988 , n70683 , n593778 );
nor ( n74666 , n74664 , n601988 );
xnor ( n601990 , n74666 , n593160 );
and ( n74668 , n74663 , n601990 );
xor ( n74669 , n601809 , n74490 );
xor ( n74670 , n74669 , n601539 );
and ( n74671 , n601990 , n74670 );
and ( n601995 , n74663 , n74670 );
or ( n601996 , n74668 , n74671 , n601995 );
and ( n74674 , n70683 , n66457 );
and ( n74675 , n70693 , n593778 );
nor ( n601999 , n74674 , n74675 );
xnor ( n602000 , n601999 , n593160 );
and ( n74678 , n601996 , n602000 );
xor ( n74679 , n74478 , n74494 );
xor ( n74680 , n74679 , n74499 );
and ( n74681 , n602000 , n74680 );
and ( n74682 , n601996 , n74680 );
or ( n74683 , n74678 , n74681 , n74682 );
and ( n74684 , n70693 , n66457 );
and ( n74685 , n70637 , n593778 );
nor ( n74686 , n74684 , n74685 );
xnor ( n602010 , n74686 , n593160 );
and ( n74688 , n74683 , n602010 );
xor ( n602012 , n74502 , n74506 );
xor ( n74690 , n602012 , n74509 );
and ( n602014 , n602010 , n74690 );
and ( n74692 , n74683 , n74690 );
or ( n602016 , n74688 , n602014 , n74692 );
and ( n602017 , n70637 , n66457 );
and ( n74695 , n70261 , n593778 );
nor ( n74696 , n602017 , n74695 );
xnor ( n602020 , n74696 , n593160 );
and ( n602021 , n602016 , n602020 );
xor ( n74699 , n74512 , n74516 );
xor ( n602023 , n74699 , n74519 );
and ( n602024 , n602020 , n602023 );
and ( n74702 , n602016 , n602023 );
or ( n602026 , n602021 , n602024 , n74702 );
and ( n602027 , n597402 , n594441 );
and ( n74705 , n597260 , n67116 );
nor ( n74706 , n602027 , n74705 );
xnor ( n602030 , n74706 , n66190 );
and ( n74708 , n70255 , n594210 );
and ( n602032 , n597569 , n66885 );
nor ( n74710 , n74708 , n602032 );
xnor ( n74711 , n74710 , n593434 );
and ( n602035 , n602030 , n74711 );
xor ( n74713 , n602016 , n602020 );
xor ( n74714 , n74713 , n602023 );
and ( n74715 , n74711 , n74714 );
and ( n74716 , n602030 , n74714 );
or ( n74717 , n602035 , n74715 , n74716 );
and ( n74718 , n602026 , n74717 );
xor ( n74719 , n74618 , n74622 );
xor ( n74720 , n74719 , n74625 );
and ( n74721 , n74717 , n74720 );
and ( n74722 , n602026 , n74720 );
or ( n74723 , n74718 , n74721 , n74722 );
and ( n74724 , n69491 , n594807 );
and ( n74725 , n69283 , n594804 );
nor ( n74726 , n74724 , n74725 );
xnor ( n74727 , n74726 , n66187 );
and ( n74728 , n74723 , n74727 );
xor ( n74729 , n74628 , n601955 );
xor ( n602053 , n74729 , n74635 );
and ( n74731 , n74727 , n602053 );
and ( n74732 , n74723 , n602053 );
or ( n602056 , n74728 , n74731 , n74732 );
and ( n602057 , n74638 , n602056 );
xor ( n74735 , n74588 , n74592 );
xor ( n602059 , n74735 , n601918 );
and ( n602060 , n602056 , n602059 );
and ( n74738 , n74638 , n602059 );
or ( n602062 , n602057 , n602060 , n74738 );
and ( n602063 , n74614 , n602062 );
xor ( n602064 , n74614 , n602062 );
and ( n74742 , n69283 , n594807 );
and ( n602066 , n596600 , n594804 );
nor ( n602067 , n74742 , n602066 );
xnor ( n74745 , n602067 , n66187 );
xor ( n602069 , n74638 , n602056 );
xor ( n602070 , n602069 , n602059 );
and ( n74748 , n74745 , n602070 );
xor ( n74749 , n74745 , n602070 );
xor ( n74750 , n74723 , n74727 );
xor ( n74751 , n74750 , n602053 );
and ( n74752 , n69581 , n594807 );
and ( n74753 , n69491 , n594804 );
nor ( n74754 , n74752 , n74753 );
xnor ( n74755 , n74754 , n66187 );
and ( n74756 , n597260 , n594441 );
and ( n74757 , n69739 , n67116 );
nor ( n74758 , n74756 , n74757 );
xnor ( n74759 , n74758 , n66190 );
and ( n74760 , n74755 , n74759 );
xor ( n74761 , n602026 , n74717 );
xor ( n74762 , n74761 , n74720 );
and ( n74763 , n74759 , n74762 );
and ( n74764 , n74755 , n74762 );
or ( n74765 , n74760 , n74763 , n74764 );
and ( n74766 , n74751 , n74765 );
xor ( n74767 , n74751 , n74765 );
xor ( n74768 , n74642 , n74646 );
and ( n74769 , n70652 , n66885 );
not ( n74770 , n74769 );
and ( n74771 , n74770 , n593434 );
and ( n74772 , n70652 , n594210 );
and ( n74773 , n597980 , n66885 );
nor ( n74774 , n74772 , n74773 );
xnor ( n74775 , n74774 , n593434 );
and ( n602099 , n74771 , n74775 );
and ( n74777 , n597980 , n594210 );
and ( n602101 , n70663 , n66885 );
nor ( n74779 , n74777 , n602101 );
xnor ( n74780 , n74779 , n593434 );
and ( n602104 , n602099 , n74780 );
and ( n74782 , n74780 , n74640 );
and ( n602106 , n602099 , n74640 );
or ( n74784 , n602104 , n74782 , n602106 );
and ( n74785 , n74768 , n74784 );
and ( n74786 , n70663 , n594210 );
and ( n74787 , n597996 , n66885 );
nor ( n74788 , n74786 , n74787 );
xnor ( n74789 , n74788 , n593434 );
and ( n74790 , n74784 , n74789 );
and ( n74791 , n74768 , n74789 );
or ( n74792 , n74785 , n74790 , n74791 );
and ( n74793 , n597996 , n594210 );
and ( n74794 , n70683 , n66885 );
nor ( n74795 , n74793 , n74794 );
xnor ( n74796 , n74795 , n593434 );
and ( n602120 , n74792 , n74796 );
xor ( n74798 , n74647 , n74651 );
xor ( n74799 , n74798 , n74479 );
and ( n74800 , n74796 , n74799 );
and ( n74801 , n74792 , n74799 );
or ( n74802 , n602120 , n74800 , n74801 );
and ( n74803 , n70683 , n594210 );
and ( n74804 , n70693 , n66885 );
nor ( n74805 , n74803 , n74804 );
xnor ( n74806 , n74805 , n593434 );
and ( n74807 , n74802 , n74806 );
xor ( n74808 , n74639 , n74655 );
xor ( n74809 , n74808 , n601983 );
and ( n602133 , n74806 , n74809 );
and ( n74811 , n74802 , n74809 );
or ( n602135 , n74807 , n602133 , n74811 );
and ( n74813 , n70693 , n594210 );
and ( n74814 , n70637 , n66885 );
nor ( n74815 , n74813 , n74814 );
xnor ( n602139 , n74815 , n593434 );
and ( n74817 , n602135 , n602139 );
xor ( n74818 , n74663 , n601990 );
xor ( n74819 , n74818 , n74670 );
and ( n602143 , n602139 , n74819 );
and ( n602144 , n602135 , n74819 );
or ( n74822 , n74817 , n602143 , n602144 );
and ( n602146 , n70637 , n594210 );
and ( n602147 , n70261 , n66885 );
nor ( n74825 , n602146 , n602147 );
xnor ( n602149 , n74825 , n593434 );
and ( n602150 , n74822 , n602149 );
xor ( n602151 , n601996 , n602000 );
xor ( n74829 , n602151 , n74680 );
and ( n602153 , n602149 , n74829 );
and ( n602154 , n74822 , n74829 );
or ( n74832 , n602150 , n602153 , n602154 );
and ( n602156 , n70261 , n594210 );
and ( n74834 , n70255 , n66885 );
nor ( n74835 , n602156 , n74834 );
xnor ( n74836 , n74835 , n593434 );
and ( n74837 , n74832 , n74836 );
xor ( n602161 , n74683 , n602010 );
xor ( n74839 , n602161 , n74690 );
and ( n74840 , n74836 , n74839 );
and ( n74841 , n74832 , n74839 );
or ( n602165 , n74837 , n74840 , n74841 );
and ( n74843 , n69739 , n594807 );
and ( n602167 , n69581 , n594804 );
nor ( n74845 , n74843 , n602167 );
xnor ( n74846 , n74845 , n66187 );
and ( n74847 , n602165 , n74846 );
xor ( n74848 , n602030 , n74711 );
xor ( n74849 , n74848 , n74714 );
and ( n74850 , n74846 , n74849 );
and ( n602174 , n602165 , n74849 );
or ( n74852 , n74847 , n74850 , n602174 );
xor ( n74853 , n74755 , n74759 );
xor ( n602177 , n74853 , n74762 );
and ( n602178 , n74852 , n602177 );
xor ( n74856 , n74852 , n602177 );
xor ( n602180 , n602165 , n74846 );
xor ( n602181 , n602180 , n74849 );
and ( n74859 , n597402 , n594807 );
and ( n602183 , n597260 , n594804 );
nor ( n74861 , n74859 , n602183 );
xnor ( n602185 , n74861 , n66187 );
and ( n74863 , n70255 , n594441 );
and ( n602187 , n597569 , n67116 );
nor ( n602188 , n74863 , n602187 );
xnor ( n74866 , n602188 , n66190 );
and ( n602190 , n602185 , n74866 );
xor ( n602191 , n74822 , n602149 );
xor ( n74869 , n602191 , n74829 );
and ( n602193 , n74866 , n74869 );
and ( n602194 , n602185 , n74869 );
or ( n74872 , n602190 , n602193 , n602194 );
and ( n74873 , n597569 , n594441 );
and ( n74874 , n597402 , n67116 );
nor ( n74875 , n74873 , n74874 );
xnor ( n602199 , n74875 , n66190 );
and ( n602200 , n74872 , n602199 );
xor ( n74878 , n74832 , n74836 );
xor ( n602202 , n74878 , n74839 );
and ( n74880 , n602199 , n602202 );
and ( n602204 , n74872 , n602202 );
or ( n74882 , n602200 , n74880 , n602204 );
and ( n74883 , n602181 , n74882 );
xor ( n602207 , n602181 , n74882 );
and ( n602208 , n597260 , n594807 );
and ( n74886 , n69739 , n594804 );
nor ( n602210 , n602208 , n74886 );
xnor ( n602211 , n602210 , n66187 );
xor ( n74889 , n74872 , n602199 );
xor ( n602213 , n74889 , n602202 );
and ( n602214 , n602211 , n602213 );
xor ( n74892 , n602211 , n602213 );
xor ( n74893 , n602185 , n74866 );
xor ( n602217 , n74893 , n74869 );
xor ( n602218 , n74771 , n74775 );
and ( n74896 , n70652 , n67116 );
not ( n602220 , n74896 );
and ( n602221 , n602220 , n66190 );
and ( n74899 , n70652 , n594441 );
and ( n602223 , n597980 , n67116 );
nor ( n602224 , n74899 , n602223 );
xnor ( n602225 , n602224 , n66190 );
and ( n74903 , n602221 , n602225 );
and ( n74904 , n597980 , n594441 );
and ( n74905 , n70663 , n67116 );
nor ( n74906 , n74904 , n74905 );
xnor ( n74907 , n74906 , n66190 );
and ( n602231 , n74903 , n74907 );
and ( n74909 , n74907 , n74769 );
and ( n74910 , n74903 , n74769 );
or ( n602234 , n602231 , n74909 , n74910 );
and ( n74912 , n602218 , n602234 );
and ( n602236 , n70663 , n594441 );
and ( n74914 , n597996 , n67116 );
nor ( n74915 , n602236 , n74914 );
xnor ( n602239 , n74915 , n66190 );
and ( n74917 , n602234 , n602239 );
and ( n602241 , n602218 , n602239 );
or ( n74919 , n74912 , n74917 , n602241 );
and ( n602243 , n597996 , n594441 );
and ( n602244 , n70683 , n67116 );
nor ( n74922 , n602243 , n602244 );
xnor ( n602246 , n74922 , n66190 );
and ( n602247 , n74919 , n602246 );
xor ( n602248 , n602099 , n74780 );
xor ( n74926 , n602248 , n74640 );
and ( n602250 , n602246 , n74926 );
and ( n602251 , n74919 , n74926 );
or ( n74929 , n602247 , n602250 , n602251 );
and ( n602253 , n70683 , n594441 );
and ( n602254 , n70693 , n67116 );
nor ( n74932 , n602253 , n602254 );
xnor ( n602256 , n74932 , n66190 );
and ( n74934 , n74929 , n602256 );
xor ( n602258 , n74768 , n74784 );
xor ( n74936 , n602258 , n74789 );
and ( n602260 , n602256 , n74936 );
and ( n74938 , n74929 , n74936 );
or ( n74939 , n74934 , n602260 , n74938 );
and ( n602263 , n70693 , n594441 );
and ( n602264 , n70637 , n67116 );
nor ( n74942 , n602263 , n602264 );
xnor ( n602266 , n74942 , n66190 );
and ( n602267 , n74939 , n602266 );
xor ( n74945 , n74792 , n74796 );
xor ( n602269 , n74945 , n74799 );
and ( n602270 , n602266 , n602269 );
and ( n74948 , n74939 , n602269 );
or ( n74949 , n602267 , n602270 , n74948 );
and ( n602273 , n70637 , n594441 );
and ( n602274 , n70261 , n67116 );
nor ( n74952 , n602273 , n602274 );
xnor ( n602276 , n74952 , n66190 );
and ( n602277 , n74949 , n602276 );
xor ( n74955 , n74802 , n74806 );
xor ( n602279 , n74955 , n74809 );
and ( n602280 , n602276 , n602279 );
and ( n74958 , n74949 , n602279 );
or ( n602282 , n602277 , n602280 , n74958 );
and ( n602283 , n70261 , n594441 );
and ( n74961 , n70255 , n67116 );
nor ( n602285 , n602283 , n74961 );
xnor ( n74963 , n602285 , n66190 );
and ( n602287 , n602282 , n74963 );
xor ( n74965 , n602135 , n602139 );
xor ( n74966 , n74965 , n74819 );
and ( n602290 , n74963 , n74966 );
and ( n74968 , n602282 , n74966 );
or ( n602292 , n602287 , n602290 , n74968 );
and ( n74970 , n602217 , n602292 );
xor ( n602294 , n602217 , n602292 );
and ( n602295 , n597569 , n594807 );
and ( n74973 , n597402 , n594804 );
nor ( n602297 , n602295 , n74973 );
xnor ( n602298 , n602297 , n66187 );
xor ( n74976 , n602282 , n74963 );
xor ( n74977 , n74976 , n74966 );
and ( n74978 , n602298 , n74977 );
xor ( n602302 , n602298 , n74977 );
and ( n74980 , n70255 , n594807 );
and ( n602304 , n597569 , n594804 );
nor ( n602305 , n74980 , n602304 );
xnor ( n602306 , n602305 , n66187 );
xor ( n74984 , n74949 , n602276 );
xor ( n602308 , n74984 , n602279 );
and ( n602309 , n602306 , n602308 );
xor ( n74987 , n602306 , n602308 );
and ( n602311 , n70261 , n594807 );
and ( n602312 , n70255 , n594804 );
nor ( n602313 , n602311 , n602312 );
xnor ( n74991 , n602313 , n66187 );
xor ( n602315 , n74939 , n602266 );
xor ( n74993 , n602315 , n602269 );
and ( n602317 , n74991 , n74993 );
xor ( n74995 , n74991 , n74993 );
and ( n602319 , n70637 , n594807 );
and ( n602320 , n70261 , n594804 );
nor ( n74998 , n602319 , n602320 );
xnor ( n74999 , n74998 , n66187 );
xor ( n602323 , n74929 , n602256 );
xor ( n602324 , n602323 , n74936 );
and ( n75002 , n74999 , n602324 );
xor ( n602326 , n74999 , n602324 );
and ( n602327 , n70693 , n594807 );
and ( n75005 , n70637 , n594804 );
nor ( n602329 , n602327 , n75005 );
xnor ( n602330 , n602329 , n66187 );
xor ( n75008 , n74919 , n602246 );
xor ( n75009 , n75008 , n74926 );
and ( n602333 , n602330 , n75009 );
xor ( n602334 , n602330 , n75009 );
and ( n75012 , n70683 , n594807 );
and ( n602336 , n70693 , n594804 );
nor ( n602337 , n75012 , n602336 );
xnor ( n75015 , n602337 , n66187 );
xor ( n602339 , n602218 , n602234 );
xor ( n602340 , n602339 , n602239 );
and ( n75018 , n75015 , n602340 );
xor ( n75019 , n75015 , n602340 );
and ( n75020 , n597996 , n594807 );
and ( n75021 , n70683 , n594804 );
nor ( n75022 , n75020 , n75021 );
xnor ( n75023 , n75022 , n66187 );
xor ( n75024 , n74903 , n74907 );
xor ( n75025 , n75024 , n74769 );
and ( n75026 , n75023 , n75025 );
xor ( n75027 , n75023 , n75025 );
and ( n75028 , n70663 , n594807 );
and ( n75029 , n597996 , n594804 );
nor ( n75030 , n75028 , n75029 );
xnor ( n75031 , n75030 , n66187 );
xor ( n75032 , n602221 , n602225 );
and ( n75033 , n75031 , n75032 );
xor ( n75034 , n75031 , n75032 );
and ( n75035 , n597980 , n594807 );
and ( n602359 , n70663 , n594804 );
nor ( n75037 , n75035 , n602359 );
xnor ( n602361 , n75037 , n66187 );
and ( n75039 , n602361 , n74896 );
xor ( n602363 , n602361 , n74896 );
and ( n75041 , n70652 , n594807 );
and ( n602365 , n597980 , n594804 );
nor ( n75043 , n75041 , n602365 );
xnor ( n602367 , n75043 , n66187 );
and ( n602368 , n70652 , n594804 );
not ( n75046 , n602368 );
and ( n75047 , n75046 , n66187 );
and ( n602371 , n602367 , n75047 );
and ( n75049 , n602363 , n602371 );
or ( n602373 , n75039 , n75049 );
and ( n602374 , n75034 , n602373 );
or ( n602375 , n75033 , n602374 );
and ( n75053 , n75027 , n602375 );
or ( n602377 , n75026 , n75053 );
and ( n602378 , n75019 , n602377 );
or ( n75056 , n75018 , n602378 );
and ( n602380 , n602334 , n75056 );
or ( n602381 , n602333 , n602380 );
and ( n75059 , n602326 , n602381 );
or ( n75060 , n75002 , n75059 );
and ( n602384 , n74995 , n75060 );
or ( n602385 , n602317 , n602384 );
and ( n75063 , n74987 , n602385 );
or ( n602387 , n602309 , n75063 );
and ( n602388 , n602302 , n602387 );
or ( n75066 , n74978 , n602388 );
and ( n602390 , n602294 , n75066 );
or ( n602391 , n74970 , n602390 );
and ( n75069 , n74892 , n602391 );
or ( n75070 , n602214 , n75069 );
and ( n75071 , n602207 , n75070 );
or ( n75072 , n74883 , n75071 );
and ( n75073 , n74856 , n75072 );
or ( n75074 , n602178 , n75073 );
and ( n75075 , n74767 , n75074 );
or ( n75076 , n74766 , n75075 );
and ( n602400 , n74749 , n75076 );
or ( n75078 , n74748 , n602400 );
and ( n602402 , n602064 , n75078 );
or ( n602403 , n602063 , n602402 );
and ( n75081 , n601935 , n602403 );
or ( n75082 , n601934 , n75081 );
and ( n75083 , n74584 , n75082 );
or ( n602407 , n601906 , n75083 );
and ( n602408 , n74475 , n602407 );
or ( n602409 , n74474 , n602408 );
and ( n75087 , n74427 , n602409 );
or ( n602411 , n601749 , n75087 );
and ( n75089 , n74389 , n602411 );
or ( n602413 , n74388 , n75089 );
and ( n75091 , n74333 , n602413 );
or ( n75092 , n601655 , n75091 );
and ( n602416 , n74214 , n75092 );
or ( n602417 , n601536 , n602416 );
and ( n75095 , n601489 , n602417 );
or ( n602419 , n601488 , n75095 );
and ( n602420 , n74098 , n602419 );
or ( n75098 , n601420 , n602420 );
and ( n602422 , n73971 , n75098 );
or ( n602423 , n73970 , n602422 );
and ( n75101 , n601236 , n602423 );
or ( n75102 , n73912 , n75101 );
and ( n602426 , n601188 , n75102 );
or ( n602427 , n601187 , n602426 );
and ( n75105 , n601021 , n602427 );
or ( n602429 , n73697 , n75105 );
and ( n602430 , n73630 , n602429 );
or ( n75108 , n600952 , n602430 );
and ( n602432 , n73574 , n75108 );
or ( n602433 , n73573 , n602432 );
and ( n75111 , n73395 , n602433 );
or ( n602435 , n600717 , n75111 );
and ( n75113 , n600640 , n602435 );
or ( n602437 , n73316 , n75113 );
and ( n75115 , n73221 , n602437 );
or ( n602439 , n600543 , n75115 );
and ( n75117 , n600383 , n602439 );
or ( n75118 , n73059 , n75117 );
and ( n602442 , n72974 , n75118 );
or ( n602443 , n600296 , n602442 );
and ( n75121 , n600056 , n602443 );
or ( n602445 , n600055 , n75121 );
and ( n602446 , n72637 , n602445 );
or ( n75124 , n72636 , n602446 );
and ( n602448 , n72519 , n75124 );
or ( n602449 , n72518 , n602448 );
and ( n75127 , n72342 , n602449 );
or ( n75128 , n72341 , n75127 );
and ( n602452 , n599569 , n75128 );
or ( n602453 , n599568 , n602452 );
and ( n75131 , n599445 , n602453 );
or ( n602455 , n599444 , n75131 );
and ( n602456 , n71921 , n602455 );
or ( n75134 , n599243 , n602456 );
and ( n602458 , n71753 , n75134 );
or ( n602459 , n599075 , n602458 );
and ( n75137 , n598845 , n602459 );
or ( n602461 , n598844 , n75137 );
and ( n602462 , n71418 , n602461 );
or ( n602463 , n71417 , n602462 );
and ( n75141 , n71117 , n602463 );
or ( n602465 , n598439 , n75141 );
and ( n75143 , n71043 , n602465 );
or ( n602467 , n71042 , n75143 );
and ( n75145 , n70851 , n602467 );
or ( n75146 , n598173 , n75145 );
and ( n602470 , n70599 , n75146 );
or ( n602471 , n70598 , n602470 );
and ( n75149 , n597868 , n602471 );
or ( n602473 , n70544 , n75149 );
and ( n602474 , n70225 , n602473 );
or ( n75152 , n597547 , n602474 );
and ( n602476 , n70069 , n75152 );
or ( n602477 , n70068 , n602476 );
and ( n75155 , n597232 , n602477 );
or ( n75156 , n597231 , n75155 );
and ( n602480 , n69859 , n75156 );
or ( n602481 , n597181 , n602480 );
and ( n75159 , n597010 , n602481 );
or ( n602483 , n69686 , n75159 );
and ( n602484 , n69435 , n602483 );
or ( n75162 , n69434 , n602484 );
and ( n602486 , n69240 , n75162 );
or ( n602487 , n69239 , n602486 );
and ( n75165 , n69038 , n602487 );
or ( n75166 , n69037 , n75165 );
and ( n75167 , n68866 , n75166 );
or ( n602491 , n596188 , n75167 );
and ( n75169 , n68704 , n602491 );
or ( n602493 , n596026 , n75169 );
and ( n75171 , n595985 , n602493 );
or ( n602495 , n68661 , n75171 );
and ( n75173 , n595787 , n602495 );
or ( n602497 , n68463 , n75173 );
and ( n75175 , n595625 , n602497 );
or ( n75176 , n595624 , n75175 );
and ( n602500 , n68100 , n75176 );
or ( n75178 , n68099 , n602500 );
and ( n602502 , n67918 , n75178 );
or ( n602503 , n67917 , n602502 );
and ( n602504 , n67878 , n602503 );
or ( n75182 , n67877 , n602504 );
and ( n602506 , n67558 , n75182 );
or ( n602507 , n67557 , n602506 );
and ( n75185 , n67379 , n602507 );
or ( n602509 , n67378 , n75185 );
and ( n602510 , n67291 , n602509 );
or ( n75188 , n594613 , n602510 );
and ( n75189 , n594409 , n75188 );
or ( n602513 , n594408 , n75189 );
and ( n602514 , n594267 , n602513 );
or ( n75192 , n66943 , n602514 );
and ( n602516 , n66747 , n75192 );
or ( n602517 , n66746 , n602516 );
and ( n75195 , n593922 , n602517 );
or ( n602519 , n66598 , n75195 );
and ( n75197 , n593750 , n602519 );
or ( n75198 , n593749 , n75197 );
and ( n75199 , n66286 , n75198 );
or ( n75200 , n593608 , n75199 );
and ( n75201 , n593424 , n75200 );
or ( n75202 , n66100 , n75201 );
and ( n75203 , n593286 , n75202 );
or ( n75204 , n65962 , n75203 );
and ( n75205 , n65821 , n75204 );
or ( n602529 , n593143 , n75205 );
and ( n75207 , n592950 , n602529 );
or ( n75208 , n592949 , n75207 );
and ( n75209 , n65572 , n75208 );
or ( n75210 , n65571 , n75209 );
and ( n75211 , n65452 , n75210 );
or ( n602535 , n592774 , n75211 );
and ( n602536 , n592631 , n602535 );
or ( n75214 , n592630 , n602536 );
and ( n602538 , n65243 , n75214 );
or ( n602539 , n65242 , n602538 );
and ( n75217 , n592465 , n602539 );
or ( n602541 , n592464 , n75217 );
and ( n602542 , n65053 , n602541 );
or ( n75220 , n65052 , n602542 );
and ( n602544 , n64963 , n75220 );
or ( n602545 , n592285 , n602544 );
and ( n75223 , n64892 , n602545 );
or ( n75224 , n592214 , n75223 );
and ( n602548 , n592135 , n75224 );
or ( n75226 , n592134 , n602548 );
and ( n602550 , n592038 , n75226 );
or ( n75228 , n592037 , n602550 );
and ( n602552 , n592003 , n75228 );
or ( n602553 , n64679 , n602552 );
and ( n75231 , n64618 , n602553 );
or ( n75232 , n64617 , n75231 );
and ( n602556 , n64553 , n75232 );
or ( n602557 , n64552 , n602556 );
and ( n75235 , n64514 , n602557 );
or ( n602559 , n64513 , n75235 );
xor ( n602560 , n64485 , n602559 );
buf ( n602561 , n602560 );
xor ( n602562 , n64514 , n602557 );
buf ( n602563 , n602562 );
xor ( n602564 , n64553 , n75232 );
buf ( n602565 , n602564 );
xor ( n75243 , n64618 , n602553 );
buf ( n602567 , n75243 );
xor ( n602568 , n592003 , n75228 );
buf ( n602569 , n602568 );
xor ( n602570 , n592038 , n75226 );
buf ( n602571 , n602570 );
xor ( n602572 , n592135 , n75224 );
buf ( n602573 , n602572 );
xor ( n75251 , n64892 , n602545 );
buf ( n602575 , n75251 );
xor ( n75253 , n64963 , n75220 );
buf ( n602577 , n75253 );
xor ( n75255 , n65053 , n602541 );
buf ( n602579 , n75255 );
xor ( n75257 , n592465 , n602539 );
buf ( n602581 , n75257 );
xor ( n75259 , n65243 , n75214 );
buf ( n602583 , n75259 );
xor ( n75261 , n592631 , n602535 );
buf ( n602585 , n75261 );
xor ( n75263 , n65452 , n75210 );
buf ( n602587 , n75263 );
xor ( n602588 , n65572 , n75208 );
buf ( n602589 , n602588 );
xor ( n75267 , n592950 , n602529 );
buf ( n602591 , n75267 );
xor ( n75269 , n65821 , n75204 );
buf ( n602593 , n75269 );
xor ( n75271 , n593286 , n75202 );
buf ( n602595 , n75271 );
xor ( n75273 , n593424 , n75200 );
buf ( n602597 , n75273 );
xor ( n75275 , n66286 , n75198 );
buf ( n602599 , n75275 );
xor ( n602600 , n593750 , n602519 );
buf ( n602601 , n602600 );
xor ( n75279 , n593922 , n602517 );
buf ( n602603 , n75279 );
xor ( n602604 , n66747 , n75192 );
buf ( n602605 , n602604 );
xor ( n602606 , n594267 , n602513 );
buf ( n602607 , n602606 );
xor ( n75285 , n594409 , n75188 );
buf ( n602609 , n75285 );
xor ( n75287 , n67291 , n602509 );
buf ( n602611 , n75287 );
xor ( n602612 , n67379 , n602507 );
buf ( n602613 , n602612 );
xor ( n602614 , n67558 , n75182 );
buf ( n602615 , n602614 );
xor ( n75293 , n67878 , n602503 );
buf ( n602617 , n75293 );
xor ( n75295 , n67918 , n75178 );
buf ( n602619 , n75295 );
xor ( n75297 , n68100 , n75176 );
buf ( n602621 , n75297 );
xor ( n75299 , n595625 , n602497 );
buf ( n602623 , n75299 );
xor ( n75301 , n595787 , n602495 );
buf ( n602625 , n75301 );
xor ( n75303 , n595985 , n602493 );
buf ( n602627 , n75303 );
xor ( n602628 , n68704 , n602491 );
buf ( n602629 , n602628 );
xor ( n602630 , n68866 , n75166 );
buf ( n602631 , n602630 );
xor ( n75309 , n69038 , n602487 );
buf ( n602633 , n75309 );
xor ( n602634 , n69240 , n75162 );
buf ( n602635 , n602634 );
xor ( n602636 , n69435 , n602483 );
buf ( n602637 , n602636 );
xor ( n75315 , n597010 , n602481 );
buf ( n602639 , n75315 );
xor ( n602640 , n69859 , n75156 );
buf ( n602641 , n602640 );
xor ( n75319 , n597232 , n602477 );
buf ( n602643 , n75319 );
xor ( n75321 , n70069 , n75152 );
buf ( n602645 , n75321 );
xor ( n75323 , n70225 , n602473 );
buf ( n602647 , n75323 );
xor ( n75325 , n597868 , n602471 );
buf ( n602649 , n75325 );
xor ( n75327 , n70599 , n75146 );
buf ( n602651 , n75327 );
xor ( n75329 , n70851 , n602467 );
buf ( n602653 , n75329 );
xor ( n602654 , n71043 , n602465 );
buf ( n602655 , n602654 );
xor ( n602656 , n71117 , n602463 );
buf ( n602657 , n602656 );
xor ( n75335 , n71418 , n602461 );
buf ( n602659 , n75335 );
xor ( n602660 , n598845 , n602459 );
buf ( n602661 , n602660 );
xor ( n75339 , n71753 , n75134 );
buf ( n602663 , n75339 );
xor ( n602664 , n71921 , n602455 );
buf ( n602665 , n602664 );
xor ( n75343 , n599445 , n602453 );
buf ( n602667 , n75343 );
xor ( n602668 , n599569 , n75128 );
buf ( n602669 , n602668 );
xor ( n75347 , n72342 , n602449 );
buf ( n602671 , n75347 );
xor ( n75349 , n72519 , n75124 );
buf ( n602673 , n75349 );
xor ( n602674 , n72637 , n602445 );
buf ( n602675 , n602674 );
xor ( n75353 , n600056 , n602443 );
buf ( n602677 , n75353 );
xor ( n75355 , n72974 , n75118 );
buf ( n602679 , n75355 );
xor ( n75357 , n600383 , n602439 );
buf ( n602681 , n75357 );
xor ( n602682 , n73221 , n602437 );
buf ( n602683 , n602682 );
xor ( n75361 , n600640 , n602435 );
buf ( n602685 , n75361 );
xor ( n602686 , n73395 , n602433 );
buf ( n602687 , n602686 );
xor ( n602688 , n73574 , n75108 );
buf ( n602689 , n602688 );
xor ( n602690 , n73630 , n602429 );
buf ( n602691 , n602690 );
xor ( n602692 , n601021 , n602427 );
buf ( n602693 , n602692 );
xor ( n75371 , n601188 , n75102 );
buf ( n602695 , n75371 );
xor ( n75373 , n601236 , n602423 );
buf ( n602697 , n75373 );
xor ( n75375 , n73971 , n75098 );
buf ( n602699 , n75375 );
xor ( n75377 , n74098 , n602419 );
buf ( n602701 , n75377 );
xor ( n75379 , n601489 , n602417 );
buf ( n602703 , n75379 );
xor ( n75381 , n74214 , n75092 );
buf ( n602705 , n75381 );
xor ( n602706 , n74333 , n602413 );
buf ( n602707 , n602706 );
xor ( n602708 , n74389 , n602411 );
buf ( n602709 , n602708 );
xor ( n75387 , n74427 , n602409 );
buf ( n602711 , n75387 );
xor ( n602712 , n74475 , n602407 );
buf ( n602713 , n602712 );
xor ( n602714 , n74584 , n75082 );
buf ( n602715 , n602714 );
xor ( n75393 , n601935 , n602403 );
buf ( n602717 , n75393 );
xor ( n602718 , n602064 , n75078 );
buf ( n602719 , n602718 );
xor ( n75397 , n74749 , n75076 );
buf ( n602721 , n75397 );
xor ( n602722 , n74767 , n75074 );
buf ( n602723 , n602722 );
xor ( n602724 , n74856 , n75072 );
buf ( n602725 , n602724 );
xor ( n75403 , n602207 , n75070 );
buf ( n602727 , n75403 );
xor ( n602728 , n74892 , n602391 );
buf ( n602729 , n602728 );
xor ( n602730 , n602294 , n75066 );
buf ( n602731 , n602730 );
xor ( n602732 , n602302 , n602387 );
buf ( n602733 , n602732 );
xor ( n602734 , n74987 , n602385 );
buf ( n602735 , n602734 );
xor ( n75413 , n74995 , n75060 );
buf ( n602737 , n75413 );
xor ( n602738 , n602326 , n602381 );
buf ( n602739 , n602738 );
xor ( n602740 , n602334 , n75056 );
buf ( n602741 , n602740 );
xor ( n75419 , n75019 , n602377 );
buf ( n602743 , n75419 );
xor ( n602744 , n75027 , n602375 );
buf ( n602745 , n602744 );
xor ( n75423 , n75034 , n602373 );
buf ( n602747 , n75423 );
xor ( n602748 , n602363 , n602371 );
buf ( n602749 , n602748 );
xor ( n75427 , n602367 , n75047 );
buf ( n602751 , n75427 );
buf ( n602752 , n602368 );
buf ( n602753 , n602752 );
buf ( n602754 , 1'b0 );
buf ( n602755 , 1'b0 );
buf ( n602756 , 1'b0 );
buf ( n602757 , 1'b0 );
buf ( n75435 , 1'b0 );
buf ( n75436 , 1'b0 );
buf ( n602760 , 1'b0 );
buf ( n75438 , 1'b0 );
buf ( n602762 , 1'b0 );
buf ( n602763 , 1'b0 );
buf ( n75441 , 1'b0 );
buf ( n75442 , 1'b0 );
buf ( n602766 , 1'b0 );
buf ( n75444 , 1'b0 );
buf ( n75445 , 1'b0 );
buf ( n75446 , 1'b0 );
buf ( n602770 , 1'b0 );
buf ( n75448 , 1'b0 );
buf ( n602772 , 1'b0 );
buf ( n75450 , 1'b0 );
buf ( n75451 , 1'b0 );
buf ( n75452 , 1'b0 );
buf ( n602776 , 1'b0 );
buf ( n75454 , 1'b0 );
buf ( n602778 , 1'b0 );
buf ( n75456 , 1'b0 );
buf ( n75457 , 1'b0 );
buf ( n602781 , 1'b0 );
buf ( n75459 , 1'b0 );
buf ( n602783 , 1'b0 );
buf ( n602784 , 1'b0 );
buf ( n75462 , 1'b0 );
buf ( n75463 , 1'b0 );
buf ( n75464 , 1'b0 );
buf ( n75465 , 1'b0 );
buf ( n75466 , 1'b0 );
buf ( n75467 , 1'b0 );
buf ( n75468 , 1'b0 );
buf ( n75469 , 1'b0 );
buf ( n75470 , 1'b0 );
buf ( n75471 , 1'b0 );
buf ( n75472 , 1'b0 );
buf ( n602796 , 1'b0 );
buf ( n75474 , 1'b0 );
buf ( n602798 , 1'b0 );
buf ( n75476 , 1'b0 );
buf ( n75477 , 1'b0 );
buf ( n75478 , 1'b0 );
buf ( n602802 , 1'b0 );
buf ( n602803 , 1'b0 );
buf ( n75481 , 1'b0 );
buf ( n602805 , 1'b0 );
buf ( n75483 , 1'b0 );
buf ( n602807 , 1'b0 );
buf ( n75485 , 1'b0 );
buf ( n602809 , 1'b0 );
buf ( n602810 , 1'b0 );
buf ( n602811 , 1'b0 );
buf ( n602812 , 1'b0 );
buf ( n75490 , 1'b0 );
buf ( n602814 , 1'b0 );
buf ( n602815 , 1'b0 );
buf ( n75493 , 1'b0 );
buf ( n602817 , 1'b0 );
buf ( n602818 , 1'b0 );
buf ( n602819 , 1'b1 );
buf ( n75497 , 1'b1 );
buf ( n602821 , 1'b1 );
buf ( n75499 , 1'b1 );
buf ( n75500 , 1'b1 );
buf ( n75501 , 1'b1 );
buf ( n75502 , 1'b1 );
buf ( n75503 , 1'b1 );
endmodule

