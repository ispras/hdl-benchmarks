module lt_10_4(a, b, c);
  input [9:0] a;
  input [3:0] b;
  output c;

  assign c = (a < b);

endmodule
