// IWLS benchmark module "dalu" printed on Wed May 29 16:31:30 2002
module dalu(inA15, inA14, inA13, inA12, inA11, inA10, inA9, inA8, inA7, inA6, inA5, inA4, inA3, inA2, inA1, inA0, inB15, inB14, inB13, inB12, inB11, inB10, inB9, inB8, inB7, inB6, inB5, inB4, inB3, inB2, inB1, inB0, inC15, inC14, inC13, inC12, inC11, inC10, inC9, inC8, inC7, inC6, inC5, inC4, inC3, inC2, inC1, inC0, inD15, inD14, inD13, inD12, inD11, inD10, inD9, inD8, inD7, inD6, inD5, inD4, inD3, inD2, inD1, inD0, opsel3, opsel2, opsel1, opsel0, musel4, musel3, musel2, musel1, sh2, sh1, sh0, O15, O14, O13, O12, O11, O10, O9, O8, O7, O6, O5, O4, O3, O2, O1, O0);
input
  inA10,
  inA11,
  inA12,
  inA13,
  inA14,
  inA15,
  inB10,
  inB11,
  inB12,
  inB13,
  inB14,
  inB15,
  inC10,
  inC11,
  inC12,
  inC13,
  inC14,
  inC15,
  inD10,
  inD11,
  inD12,
  inD13,
  inD14,
  inD15,
  inA0,
  inA1,
  inA2,
  inA3,
  inA4,
  inA5,
  inA6,
  inA7,
  inA8,
  inA9,
  inB0,
  inB1,
  inB2,
  inB3,
  inB4,
  inB5,
  inB6,
  inB7,
  inB8,
  inB9,
  inC0,
  inC1,
  inC2,
  inC3,
  inC4,
  inC5,
  inC6,
  inC7,
  inC8,
  inC9,
  inD0,
  inD1,
  inD2,
  inD3,
  inD4,
  inD5,
  inD6,
  inD7,
  inD8,
  inD9,
  sh0,
  sh1,
  sh2,
  musel1,
  musel2,
  musel3,
  musel4,
  opsel0,
  opsel1,
  opsel2,
  opsel3;
output
  O0,
  O1,
  O2,
  O3,
  O4,
  O5,
  O6,
  O7,
  O8,
  O9,
  O10,
  O11,
  O12,
  O13,
  O14,
  O15;
wire
  \[5893] ,
  \[378] ,
  \[189] ,
  \[5894] ,
  \[569] ,
  \[8520] ,
  \[6055] ,
  \[9880] ,
  \[6056] ,
  \[4349] ,
  \[5897] ,
  \[5898] ,
  \[10744] ,
  \[8335] ,
  \[9883] ,
  \[8905] ,
  \[10556] ,
  \[190] ,
  \[570] ,
  \[950] ,
  \[381] ,
  \[8908] ,
  \[382] ,
  \[11100] ,
  \[2642] ,
  \[10372] ,
  \[193] ,
  \[383] ,
  \[4540] ,
  \[194] ,
  \[384] ,
  \[4352] ,
  \[2645] ,
  \[575] ,
  \[576] ,
  \[6061] ,
  \[197] ,
  \[6062] ,
  \[198] ,
  \[6063] ,
  \[199] ,
  \[8911] ,
  \[6065] ,
  \[6066] ,
  \[10944] ,
  \[8914] ,
  \[0] ,
  \[10946] ,
  \[1] ,
  \[2] ,
  \[8917] ,
  \[10570] ,
  \[391] ,
  \[581] ,
  \[3] ,
  \[582] ,
  \[4] ,
  \[1105] ,
  \[5] ,
  \[11302] ,
  \[6] ,
  \[1107] ,
  \[7] ,
  \[8] ,
  \[6071] ,
  \[587] ,
  \[9] ,
  \[6072] ,
  \[588] ,
  \[6073] ,
  \[399] ,
  \[8540] ,
  \[969] ,
  \[8920] ,
  \[6074] ,
  \[11308] ,
  \[6075] ,
  \[8923] ,
  \[10764] ,
  \[8926] ,
  \[10960] ,
  \[11310] ,
  \[782] ,
  \[8929] ,
  \[1115] ,
  \[593] ,
  \[594] ,
  \[6080] ,
  \[6081] ,
  \[6082] ,
  \[10588] ,
  \[8360] ,
  \[599] ,
  \[11318] ,
  \[8932] ,
  \[6086] ,
  \[6087] ,
  \[8935] ,
  \[10396] ,
  \[1501] ,
  \[1312] ,
  \[11316] ,
  \[1502] ,
  \[11506] ,
  \[8938] ,
  \[3404] ,
  \[4954] ,
  \[6092] ,
  \[5304] ,
  \[6093] ,
  \[10978] ,
  \[799] ,
  \[6094] ,
  \[8181] ,
  \[8941] ,
  \[8562] ,
  \[6097] ,
  \[8944] ,
  \[6098] ,
  \[1130] ,
  \[11324] ,
  \[10786] ,
  \[1511] ,
  \[2490] ,
  \[11326] ,
  \[1512] ,
  \[8947] ,
  \[3600] ,
  G3,
  \[2493] ,
  \[1136] ,
  \[11332] ,
  \[4392] ,
  \[1517] ,
  \[1329] ,
  \[1519] ,
  \[4965] ,
  \[3228] ,
  \[8950] ,
  \[11908] ,
  \[4968] ,
  \[9301] ,
  \[8953] ,
  \[11334] ,
  \[1520] ,
  \[1331] ,
  \[8956] ,
  \[11146] ,
  \[1332] ,
  \[8388] ,
  \[9117] ,
  \[3231] ,
  \[11340] ,
  \[8959] ,
  \[11910] ,
  \[4780] ,
  \[1525] ,
  \[9119] ,
  \[11342] ,
  \[1526] ,
  \[1337] ,
  \[5701] ,
  \[1338] ,
  \[5514] ,
  \[5704] ,
  \[10998] ,
  \[11348] ,
  \[11728] ,
  \[5517] ,
  \[8962] ,
  b0,
  b1,
  b2,
  b3,
  b4,
  b5,
  b6,
  b7,
  b8,
  b9,
  \[9314] ,
  \[8965] ,
  \[1910] ,
  \[8586] ,
  e0,
  e1,
  e2,
  e3,
  e5,
  e6,
  e7,
  \[8777] ,
  e9,
  \[11726] ,
  \[8968] ,
  \[1913] ,
  \[9507] ,
  \[11350] ,
  \[11920] ,
  \[1535] ,
  \[11922] ,
  \[5900] ,
  \[1347] ,
  \[1537] ,
  \[1538] ,
  \[5712] ,
  \[1349] ,
  \[3626] ,
  \[5713] ,
  \[5903] ,
  \[5904] ,
  \[5905] ,
  \[11358] ,
  \[3629] ,
  \[8971] ,
  \[9511] ,
  \[9132] ,
  \[5908] ,
  \[8974] ,
  \[5719] ,
  \[9513] ,
  \[5909] ,
  \[1350] ,
  \[11544] ,
  \[11166] ,
  \[11356] ,
  \[11546] ,
  \[8977] ,
  \[1353] ,
  \[1543] ,
  \[202] ,
  \[9707] ,
  \[1354] ,
  \[1544] ,
  \[203] ,
  \[204] ,
  \[1356] ,
  \[1167] ,
  \[5911] ,
  \[5722] ,
  \[207] ,
  \[5533] ,
  \[208] ,
  \[5913] ,
  \[209] ,
  \[8980] ,
  \[5156] ,
  \[5536] ,
  \[5916] ,
  \[9331] ,
  \[5917] ,
  \[9711] ,
  \[9901] ,
  b10,
  b11,
  b12,
  \[8983] ,
  b13,
  b14,
  b15,
  \[5918] ,
  \[9523] ,
  \[9713] ,
  \[11364] ,
  \[1361] ,
  \[9145] ,
  \[9335] ,
  \[8986] ,
  \[210] ,
  \[9905] ,
  \[11366] ,
  \[1363] ,
  \[1553] ,
  \[9337] ,
  \[9527] ,
  \[11180] ,
  \[1364] ,
  \[8989] ,
  \[213] ,
  \[1555] ,
  \[9529] ,
  \[214] ,
  \[9719] ,
  \[11372] ,
  \[1556] ,
  \[5730] ,
  \[5731] ,
  \[5921] ,
  \[5542] ,
  \[217] ,
  \[5922] ,
  \[3076] ,
  \[1369] ,
  \[5543] ,
  \[218] ,
  \[219] ,
  \[5924] ,
  \[3079] ,
  \[8992] ,
  \[5737] ,
  \[5927] ,
  \[9721] ,
  \[9911] ,
  \[10204] ,
  \[5928] ,
  \[10013] ,
  \[5929] ,
  \[9913] ,
  \[1370] ,
  \[11374] ,
  \[10015] ,
  \[1561] ,
  \[600] ,
  \[1562] ,
  \[10400] ,
  \[411] ,
  \[3270] ,
  \[9347] ,
  \[222] ,
  \[11380] ,
  \[11760] ,
  \[223] ,
  \[9728] ,
  \[9539] ,
  \[224] ,
  \[11382] ,
  \[11762] ,
  \[5740] ,
  \[605] ,
  \[1567] ,
  \[5551] ,
  \[606] ,
  \[1568] ,
  \[227] ,
  \[5932] ,
  \[1379] ,
  \[228] ,
  \[5933] ,
  \[5554] ,
  \[229] ,
  \[5555] ,
  \[5935] ,
  \[11388] ,
  \[11578] ,
  \[9920] ,
  \[10029] ,
  \[9351] ,
  \[9731] ,
  \[5748] ,
  \[9353] ,
  \[5749] ,
  \[9543] ,
  \[5939] ,
  \[1190] ,
  \[9923] ,
  \[1381] ,
  \[9165] ,
  \[9545] ,
  \[230] ,
  \[11196] ,
  \[1382] ,
  \[611] ,
  \[612] ,
  \[11390] ,
  \[11580] ,
  \[233] ,
  \[423] ,
  \[10031] ,
  \[234] ,
  \[424] ,
  \[11772] ,
  \[425] ,
  \[1387] ,
  \[1577] ,
  \[426] ,
  \[1388] ,
  \[237] ,
  \[617] ,
  \[1579] ,
  \[5563] ,
  \[238] ,
  \[618] ,
  \[5564] ,
  \[6103] ,
  \[239] ,
  \[10608] ,
  \[6104] ,
  \[5755] ,
  \[5945] ,
  \[11398] ,
  \[6105] ,
  \[9740] ,
  \[9171] ,
  \[5378] ,
  e10,
  \[10224] ,
  e11,
  e13,
  \[6107] ,
  \[10414] ,
  e14,
  \[5758] ,
  e15,
  \[9932] ,
  \[9363] ,
  \[6108] ,
  \[9743] ,
  \[1580] ,
  \[11774] ,
  \[9555] ,
  \[9935] ,
  \[11396] ,
  \[1772] ,
  \[9367] ,
  \[242] ,
  \[432] ,
  \[243] ,
  \[623] ,
  \[1775] ,
  \[9369] ,
  \[9559] ,
  \[244] ,
  \[9749] ,
  \[624] ,
  \[5570] ,
  \[5760] ,
  \[5950] ,
  \[1397] ,
  \[5951] ,
  \[247] ,
  \[5952] ,
  \[1399] ,
  \[1589] ,
  \[5573] ,
  \[5763] ,
  \[248] ,
  \[438] ,
  \[10048] ,
  \[6113] ,
  \[249] ,
  \[6114] ,
  \[5955] ,
  \[6115] ,
  \[11978] ,
  \[5956] ,
  \[9561] ,
  \[5957] ,
  \[9941] ,
  \[10044] ,
  \[6117] ,
  \[9753] ,
  \[10046] ,
  \[9184] ,
  pgx3,
  \[1591] ,
  \[9755] ,
  \[9945] ,
  \[10050] ,
  \[1592] ,
  \[11976] ,
  \[441] ,
  \[631] ,
  \[252] ,
  \[9757] ,
  \[9947] ,
  \[10432] ,
  \[9379] ,
  \[9949] ,
  \[4222] ,
  \[255] ,
  \[1597] ,
  \[5581] ,
  \[5771] ,
  \[256] ,
  \[1598] ,
  \[5582] ,
  \[5772] ,
  \[5962] ,
  \[258] ,
  \[5963] ,
  \[10058] ,
  \[11988] ,
  \[5966] ,
  \[9760] ,
  \[9571] ,
  \[5967] ,
  \[10244] ,
  \[5588] ,
  \[5778] ,
  \[9952] ,
  \[9383] ,
  \[5969] ,
  \[9763] ,
  \[10056] ,
  \[9385] ,
  \[9575] ,
  \[9955] ,
  \[10060] ,
  \[10630] ,
  \[9766] ,
  \[9197] ,
  \[9577] ,
  \[10062] ,
  \[11990] ,
  \[263] ,
  \[10632] ,
  \[9958] ,
  \[264] ,
  \[5970] ,
  \[835] ,
  \[5591] ,
  \[5781] ,
  \[266] ,
  \[10068] ,
  \[10258] ,
  \[5975] ,
  \[5976] ,
  \[5977] ,
  \[5978] ,
  \[9772] ,
  \[5599] ,
  \[5789] ,
  \[5979] ,
  \[9964] ,
  \[9395] ,
  \[10070] ,
  \[271] ,
  \[9776] ,
  \[8418] ,
  \[10830] ,
  \[272] ,
  \[10072] ,
  \[10452] ,
  \[9968] ,
  \[9399] ,
  \[274] ,
  \[9779] ,
  \[464] ,
  \[5790] ,
  \[5980] ,
  \[465] ,
  \[5981] ,
  \[466] ,
  \[5982] ,
  \[467] ,
  \[468] ,
  \[279] ,
  \[8611] ,
  \[5796] ,
  \[5987] ,
  \[9971] ,
  \[10074] ,
  \[5988] ,
  \[5799] ,
  \[10646] ,
  \[280] ,
  \[10080] ,
  \[661] ,
  \[2352] ,
  \[282] ,
  \[10082] ,
  \[2355] ,
  \[5990] ,
  \[287] ,
  \[5992] ,
  \[667] ,
  \[288] ,
  \[5993] ,
  \[10468] ,
  \[5994] ,
  \[10084] ,
  \[5998] ,
  \[10086] ,
  \[10276] ,
  \[290] ,
  \[480] ,
  \[10850] ,
  \[10092] ,
  \[1005] ,
  \[483] ,
  \[4640] ,
  \[484] ,
  \[295] ,
  \[865] ,
  \[296] ,
  \[298] ,
  \[2938] ,
  \[10098] ,
  \[489] ,
  \[8440] ,
  \[11018] ,
  \[10094] ,
  \[10474] ,
  \[10664] ,
  \[11014] ,
  \[1200] ,
  \[11204] ,
  \[10096] ,
  \[10476] ,
  \[2941] ,
  \[11022] ,
  \[875] ,
  \[496] ,
  \[4466] ,
  \[10868] ,
  \[8263] ,
  \[5008] ,
  \[11024] ,
  \[1400] ,
  \[11404] ,
  \[10296] ,
  \[11026] ,
  \[11406] ,
  \[10870] ,
  \[1405] ,
  \[1406] ,
  \[11412] ,
  \[4663] ,
  \[697] ,
  \[4854] ,
  \[4666] ,
  \[11228] ,
  \[10684] ,
  \[8464] ,
  \[1221] ,
  \[1411] ,
  \[11226] ,
  \[1412] ,
  \[1603] ,
  \[11040] ,
  \[11420] ,
  \[1604] ,
  \[8849] ,
  \[1035] ,
  \[11612] ,
  \[10884] ,
  \[11424] ,
  \[11614] ,
  \[8286] ,
  \[1421] ,
  \[11806] ,
  \[1423] ,
  \[1613] ,
  \[1424] ,
  \[1045] ,
  \[1235] ,
  \[1615] ,
  \[3512] ,
  \[11242] ,
  \[12790] ,
  \[1616] ,
  \[5600] ,
  \[3515] ,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[5606] ,
  \[14] ,
  \[9401] ,
  \[15] ,
  \[5609] ,
  \[11434] ,
  \[11624] ,
  \[12799] ,
  \[1431] ,
  \[1432] ,
  \[11626] ,
  \[12793] ,
  \[9217] ,
  \[12796] ,
  \[1434] ,
  \[1627] ,
  \[1439] ,
  \[1629] ,
  \[11068] ,
  \[8491] ,
  \[5617] ,
  \[9411] ,
  \[5807] ,
  \[5618] ,
  \[5808] ,
  \[9223] ,
  \[11254] ,
  \[1630] ,
  \[1441] ,
  \[9415] ,
  \[9605] ,
  \[1442] ,
  \[9417] ,
  \[1635] ,
  \[9609] ,
  \[11262] ,
  \[1636] ,
  \[1447] ,
  \[1448] ,
  \[5624] ,
  \[5814] ,
  \[3348] ,
  \[5627] ,
  \[5817] ,
  \[9611] ,
  \[9615] ,
  \[11456] ,
  \[9236] ,
  \[9427] ,
  \[9617] ,
  \[9807] ,
  \[11840] ,
  \[303] ,
  \[1075] ,
  \[304] ,
  \[11842] ,
  \[1457] ,
  \[306] ,
  \[1459] ,
  \[3736] ,
  \[10108] ,
  \[5635] ,
  \[5825] ,
  \[5256] ,
  \[5636] ,
  \[5826] ,
  \[9431] ,
  \[9621] ,
  \[10104] ,
  \[9433] ,
  \[9623] ,
  \[1460] ,
  \[10106] ,
  \[11654] ,
  \[9815] ,
  \[10110] ,
  \[311] ,
  \[312] ,
  \[11090] ,
  \[9817] ,
  \[8899] ,
  \[503] ,
  \[1465] ,
  \[9249] ,
  \[9629] ,
  \[314] ,
  \[11282] ,
  \[1466] ,
  \[506] ,
  \[5642] ,
  \[5832] ,
  \[1089] ,
  \[507] ,
  \[508] ,
  \[10118] ,
  \[319] ,
  \[509] ,
  \[5645] ,
  \[5835] ,
  \[11288] ,
  \[5456] ,
  \[5837] ,
  \[9443] ,
  \[9823] ,
  \[10116] ,
  \[9635] ,
  \[320] ,
  \[9825] ,
  \[11286] ,
  \[10120] ,
  \[511] ,
  \[9447] ,
  \[322] ,
  \[11290] ,
  \[10122] ,
  \[9638] ,
  \[1475] ,
  \[12020] ,
  \[9449] ,
  \[514] ,
  \[5840] ,
  \[1477] ,
  \[6000] ,
  \[5082] ,
  \[1478] ,
  \[6001] ,
  \[327] ,
  \[517] ,
  \[707] ,
  \[5653] ,
  \[5843] ,
  \[328] ,
  \[10128] ,
  \[10318] ,
  \[5654] ,
  \[5844] ,
  \[11298] ,
  \[11488] ,
  \[5846] ,
  \[6006] ,
  \[9641] ,
  \[6007] ,
  \[9832] ,
  \[6008] ,
  \[5849] ,
  \[10316] ,
  \[330] ,
  \[9835] ,
  \[10130] ,
  \[10320] ,
  \[1483] ,
  \[9647] ,
  \[1484] ,
  \[11490] ,
  \[10132] ,
  \[9269] ,
  \[3762] ,
  \[9459] ,
  \[5660] ,
  \[5850] ,
  \[335] ,
  \[905] ,
  \[336] ,
  \[6011] ,
  \[3765] ,
  \[1489] ,
  \[6012] ,
  \[5663] ,
  \[5853] ,
  \[338] ,
  \[5854] ,
  \[10708] ,
  \[3388] ,
  \[5855] ,
  \[4308] ,
  \[10134] ,
  \[6017] ,
  \[5858] ,
  \[10704] ,
  \[6018] ,
  \[9463] ,
  \[5859] ,
  \[9653] ,
  \[1490] ,
  \[6019] ,
  \[11874] ,
  \[10516] ,
  \[9844] ,
  \[9275] ,
  \[9465] ,
  \[9655] ,
  \[11496] ,
  \[10140] ,
  \[11876] ,
  \[10710] ,
  \[9847] ,
  \[3391] ,
  \[10142] ,
  \[343] ,
  \[10712] ,
  \[10902] ,
  \[344] ,
  \[11692] ,
  \[5671] ,
  \[5861] ,
  \[346] ,
  \[12802] ,
  \[6021] ,
  \[5672] ,
  \[1499] ,
  \[2228] ,
  \[6022] ,
  \[5864] ,
  \[919] ,
  \[5865] ,
  \[5866] ,
  \[12048] ,
  \[9661] ,
  \[12808] ,
  \[10144] ,
  \[6027] ,
  \[10334] ,
  \[5678] ,
  \[6028] ,
  \[5869] ,
  \[9853] ,
  \[10146] ,
  \[11694] ,
  \[6029] ,
  \[9664] ,
  \[9475] ,
  \[2231] ,
  \[351] ,
  \[352] ,
  \[9857] ,
  \[10152] ,
  \[9288] ,
  \[12805] ,
  \[12050] ,
  \[3592] ,
  \[9479] ,
  \[354] ,
  \[9859] ,
  \[5870] ,
  \[6030] ,
  \[5681] ,
  \[5871] ,
  \[6031] ,
  \[5682] ,
  \[12811] ,
  \[737] ,
  \[10158] ,
  \[5874] ,
  \[359] ,
  \[4706] ,
  \[5875] ,
  \[9670] ,
  \[6036] ,
  \[9481] ,
  \[5877] ,
  \[8313] ,
  \[9861] ,
  \[10154] ,
  \[6037] ,
  \[6038] ,
  \[10156] ,
  \[6039] ,
  \[10536] ,
  \[9674] ,
  \[10726] ,
  \[9864] ,
  \[360] ,
  \[9677] ,
  \[362] ,
  \[9867] ,
  \[10352] ,
  \[173] ,
  \[10922] ,
  \[2814] ,
  \[5880] ,
  \[555] ,
  \[5881] ,
  \[556] ,
  \[177] ,
  \[5882] ,
  \[367] ,
  \[2817] ,
  \[178] ,
  \[368] ,
  \[10168] ,
  \[5694] ,
  \[179] ,
  \[6044] ,
  \[5695] ,
  \[5885] ,
  \[6045] ,
  \[4338] ,
  \[5886] ,
  \[9870] ,
  \[9491] ,
  \[10164] ,
  \[5888] ,
  \[5889] ,
  \[10166] ,
  \[9495] ,
  \[370] ,
  \[10170] ,
  \[9876] ,
  \[561] ,
  \[751] ,
  \[2062] ,
  \[9497] ,
  \[182] ,
  \[562] ,
  \[10172] ,
  \[183] ,
  \[563] ,
  \[184] ,
  \[564] ,
  \[2065] ,
  \[375] ,
  \[6050] ,
  \[376] ,
  \[6051] ,
  \[187] ,
  \[5892] ,
  \[6052] ,
  \[188] ;
assign
  \[5893]  = (~\[5892]  & \[5849] ) | ~\[11358] ,
  \[378]  = (~inB0 & ~\[1772] ) | ((~inB0 & ~musel1) | ((~\[9575]  & ~\[1772] ) | (~\[9575]  & ~musel1))),
  \[189]  = (~\[8911]  & ~\[8956] ) | ((~\[8911]  & ~opsel2) | (~\[8956]  & opsel2)),
  \[5894]  = ~inC10 | ~musel2,
  \[569]  = (~\[10060]  & ~\[10056] ) | ((~\[10060]  & ~sh1) | (~\[10056]  & sh1)),
  \[8520]  = (~\[6071]  & ~\[346] ) | ~\[10536] ,
  \[6055]  = ~\[5886]  | (~\[5881]  | ~\[12790] ),
  \[9880]  = ~\[5681]  | \[5671] ,
  \[6056]  = ~opsel2 | ~\[8929] ,
  \[4349]  = (\[5835]  & \[5817] ) | ((\[5835]  & ~\[5807] ) | ((~\[5825]  & \[5817] ) | (~\[5825]  & ~\[5807] ))),
  \[5897]  = ~\[9417]  | (musel3 | ~musel4),
  \[5898]  = (~\[5897]  & \[5849] ) | ~\[11350] ,
  \[10744]  = ~sh2 | ~\[8440] ,
  \[8335]  = (~\[5987]  & ~\[290] ) | ~\[11068] ,
  \[9883]  = \[5681]  | ~\[5671] ,
  \[8905]  = (~\[5955]  & ~\[5854] ) | ~\[11242] ,
  \[10556]  = ~\[9249]  | (opsel2 | ~opsel3),
  \[190]  = (~\[9165]  & \[5979] ) | ((~\[9165]  & ~\[8956] ) | ((~\[8899]  & \[5979] ) | (~\[8899]  & ~\[8956] ))),
  \[570]  = (~\[10062]  & ~\[10058] ) | ((~\[10062]  & ~sh1) | (~\[10058]  & sh1)),
  \[950]  = (~\[6038]  & ~\[10786] ) | (~\[6038]  & ~\[9740] ),
  \[381]  = ~\[1421]  & (~opsel0 & ~\[5778] ),
  \[8908]  = (~\[5969]  & ~\[5859] ) | ~\[11180] ,
  \[382]  = ~\[1397]  & (~opsel0 & ~\[5796] ),
  \[11100]  = \[5627]  | \[5617] ,
  \[2642]  = musel2 & inD6,
  \[10372]  = ~\[2065]  | (musel3 | (~musel4 | ~inD2)),
  \[193]  = (~\[1089]  & \[194] ) | (~\[1089]  & ~\[5992] ),
  \[383]  = ~\[1379]  & (~opsel0 & ~\[5814] ),
  \[4540]  = musel2 & inC2,
  \[194]  = (~\[8914]  & ~\[8959] ) | ((~\[8914]  & ~opsel2) | (~\[8959]  & opsel2)),
  \[384]  = ~\[1361]  & (~opsel0 & ~\[5832] ),
  \[4352]  = (\[5799]  & \[5781] ) | ((\[5799]  & ~\[5771] ) | ((~\[5789]  & \[5781] ) | (~\[5789]  & ~\[5771] ))),
  \[2645]  = ~musel1 & ~musel2,
  \[575]  = (~\[10072]  & ~\[10068] ) | ((~\[10072]  & ~sh1) | (~\[10068]  & sh1)),
  \[576]  = (~\[10074]  & ~\[10070] ) | ((~\[10074]  & ~sh1) | (~\[10070]  & sh1)),
  \[6061]  = ~musel3 | musel4,
  \[197]  = (~opsel0 & ~opsel1) | (opsel0 & opsel1),
  \[6062]  = opsel0 | opsel1,
  \[198]  = (~\[1045]  & \[199] ) | (~\[1045]  & ~\[6007] ),
  \[6063]  = (~\[5740]  & ~\[5730] ) | (\[5740]  & \[5730] ),
  \[199]  = (~\[8917]  & ~\[8962] ) | ((~\[8917]  & ~opsel2) | (~\[8962]  & opsel2)),
  \[8911]  = (~pgx3 & \[5865] ) | (pgx3 & ~\[5865] ),
  \[6065]  = ~\[12790]  | ~\[5886] ,
  \[6066]  = ~opsel2 | ~\[8932] ,
  \[10944]  = ~\[9883]  | ~\[5994] ,
  \[8914]  = (~\[6000]  & ~\[5893] ) | ~\[11040] ,
  \[0]  = (~\[173]  & ~opsel3) | ~\[11290] ,
  \[10946]  = ~\[9184]  | (opsel2 | ~opsel3),
  \[1]  = (~\[178]  & ~opsel3) | ~\[11228] ,
  \[2]  = (~\[183]  & ~opsel3) | ~\[11166] ,
  \[8917]  = (~\[6011]  & ~\[5898] ) | ~\[10960] ,
  \[10570]  = ~\[6065]  | ~\[5881] ,
  \[391]  = (~\[1356]  & ~\[4338] ) | (~\[1356]  & ~\[9605] ),
  \[581]  = (~\[10084]  & ~\[10080] ) | ((~\[10084]  & ~sh1) | (~\[10080]  & sh1)),
  \[3]  = (~\[188]  & ~opsel3) | (~\[5981]  & ~\[190] ),
  \[582]  = (~\[10086]  & ~\[10082] ) | ((~\[10086]  & ~sh1) | (~\[10082]  & sh1)),
  \[4]  = (~\[193]  & ~opsel3) | ~\[11026] ,
  \[1105]  = \[8286]  & sh1,
  \[5]  = (~\[198]  & ~opsel3) | ~\[10946] ,
  \[11302]  = ~\[5932]  | \[5849] ,
  \[6]  = (~\[203]  & ~opsel3) | ~\[10870] ,
  \[1107]  = \[8263]  & ~sh2,
  \[7]  = (~\[208]  & ~opsel3) | (~\[6030]  & ~\[210] ),
  \[8]  = (~\[213]  & ~opsel3) | ~\[10712] ,
  \[6071]  = ~musel3 | musel4,
  \[587]  = (~\[10096]  & ~\[10092] ) | ((~\[10096]  & ~sh1) | (~\[10092]  & sh1)),
  \[9]  = (~\[218]  & ~opsel3) | ~\[10632] ,
  \[6072]  = opsel0 | opsel1,
  \[588]  = (~\[10098]  & ~\[10094] ) | ((~\[10098]  & ~sh1) | (~\[10094]  & sh1)),
  \[6073]  = (~\[5758]  & ~\[5748] ) | (\[5758]  & \[5748] ),
  \[399]  = (~\[12799]  & ~\[9623] ) | (~\[12799]  & ~\[5840] ),
  \[8540]  = (~\[6080]  & ~\[354] ) | ~\[10452] ,
  \[969]  = ~\[6031]  & ~\[6028] ,
  \[8920]  = (~\[6021]  & ~\[5904] ) | ~\[10884] ,
  \[6074]  = opsel2 | ~opsel3,
  \[11308]  = ~musel1 | (musel2 | ~inA0),
  \[6075]  = ~opsel2 | ~\[8935] ,
  \[8923]  = (~\[5998]  & ~\[5909] ) | (\[5998]  & \[5909] ),
  \[10764]  = ~\[2817]  | (musel3 | (~musel4 | ~inD7)),
  \[8926]  = (~\[6044]  & ~\[5870] ) | ~\[10726] ,
  \[10960]  = ~\[6011]  | ~\[5898] ,
  \[11310]  = ~\[5927]  | \[5849] ,
  \[782]  = (~\[6082]  & ~\[10474] ) | (~\[6082]  & ~\[9638] ),
  \[8929]  = (~\[6055]  & ~\[5875] ) | ~\[10646] ,
  \[1115]  = (~\[5993]  & ~\[11090] ) | (~\[5993]  & ~\[9844] ),
  \[593]  = (~\[10108]  & ~\[10104] ) | ((~\[10108]  & ~sh1) | (~\[10104]  & sh1)),
  \[594]  = (~\[10110]  & ~\[10106] ) | ((~\[10110]  & ~sh1) | (~\[10106]  & sh1)),
  \[6080]  = ~musel3 | musel4,
  \[6081]  = opsel0 | opsel1,
  \[6082]  = (~\[5781]  & ~\[5771] ) | (\[5781]  & \[5771] ),
  \[10588]  = ~sh2 | ~\[8491] ,
  \[8360]  = (~\[6006]  & ~\[298] ) | ~\[10998] ,
  \[599]  = (~\[10120]  & ~\[10116] ) | ((~\[10120]  & ~sh1) | (~\[10116]  & sh1)),
  \[11318]  = ~\[5921]  | \[5849] ,
  \[8932]  = (~\[6065]  & ~\[5881] ) | ~\[10570] ,
  \[6086]  = ~\[5933]  | (~\[5928]  | (~\[5922]  | \[5849] )),
  \[6087]  = ~opsel2 | ~\[8938] ,
  \[8935]  = (~\[12790]  & \[5886] ) | (\[12790]  & ~\[5886] ),
  \[10396]  = ~\[9653]  | ~\[9664] ,
  \[1501]  = ~musel1 & (~musel2 & (~\[5695]  & ~musel3)),
  \[1312]  = (~\[5555]  & ~\[11456] ) | (~\[5555]  & ~\[9932] ),
  \[11316]  = ~musel1 | (musel2 | ~inA1),
  \[1502]  = ~\[320]  & (musel3 & ~musel4),
  \[11506]  = (~\[1354]  & ~\[1353] ) | ~\[9609] ,
  \[8938]  = (~\[6086]  & ~\[5917] ) | ~\[10414] ,
  \[3404]  = \[8181]  & sh2,
  \[4954]  = musel2 & inC7,
  \[6092]  = ~musel3 | musel4,
  \[5304]  = musel2 & inC13,
  \[6093]  = opsel0 | opsel1,
  \[10978]  = ~sh2 | ~\[8360] ,
  \[799]  = ~\[6075]  & ~\[6072] ,
  \[6094]  = (~\[5799]  & ~\[5789] ) | (\[5799]  & \[5789] ),
  \[8181]  = (~\[5533]  & ~\[258] ) | ~\[11434] ,
  \[8941]  = (~\[6097]  & ~\[5922] ) | ~\[10334] ,
  \[8562]  = (~\[6092]  & ~\[362] ) | ~\[10372] ,
  \[6097]  = ~\[5933]  | (~\[5928]  | \[5849] ),
  \[8944]  = (~\[6107]  & ~\[5928] ) | ~\[10258] ,
  \[6098]  = ~opsel2 | ~\[8941] ,
  \[1130]  = ~\[5843]  & ~\[5840] ,
  \[11324]  = ~musel1 | (musel2 | ~inA2),
  \[10786]  = ~\[9719]  | ~\[9743] ,
  \[1511]  = (~\[5682]  & \[5663] ) | (~\[5682]  & ~\[5653] ),
  \[2490]  = musel2 & inD5,
  \[11326]  = ~\[5916]  | \[5849] ,
  \[1512]  = \[5663]  & ~\[5653] ,
  \[8947]  = (~\[5933]  & ~\[5849] ) | (\[5933]  & \[5849] ),
  \[3600]  = ~sh1 & ~sh2,
  G3 = (~\[9807]  & ~\[5627] ) | ((~\[9807]  & \[5617] ) | ((~\[9815]  & ~\[5627] ) | (~\[9815]  & \[5617] ))),
  \[2493]  = ~musel1 & ~musel2,
  \[1136]  = ~\[5982]  & ~\[5979] ,
  \[11332]  = ~musel1 | (musel2 | ~inA3),
  \[4392]  = musel2 & inC0,
  \[1517]  = opsel2 & opsel3,
  \[1329]  = opsel2 & opsel3,
  \[1519]  = ~musel1 & (~musel2 & (~\[5672]  & ~musel3)),
  \[4965]  = (\[5681]  & \[5663] ) | ((\[5681]  & ~\[5653] ) | ((~\[5671]  & \[5663] ) | (~\[5671]  & ~\[5653] ))),
  \[3228]  = musel2 & inD10,
  \[8950]  = (~\[5950]  & \[8263] ) | ~\[11254] ,
  O0 = \[15] ,
  O1 = \[14] ,
  O2 = \[13] ,
  O3 = \[12] ,
  O4 = \[11] ,
  O5 = \[10] ,
  O6 = \[9] ,
  O7 = \[8] ,
  O8 = \[7] ,
  O9 = \[6] ,
  \[11908]  = musel2 | (~musel3 | ~inD10),
  \[4968]  = (\[5645]  & \[5627] ) | ((\[5645]  & ~\[5617] ) | ((~\[5635]  & \[5627] ) | (~\[5635]  & ~\[5617] ))),
  \[9301]  = (~\[247]  & ~e1) | (\[8989]  & ~\[6104] ),
  \[8953]  = (~\[5963]  & ~\[5957] ) | ~\[3592] ,
  \[11334]  = ~\[5908]  | \[5849] ,
  \[1520]  = ~\[312]  & (musel3 & ~musel4),
  \[1331]  = ~musel1 & (~musel2 & (~\[5600]  & ~musel3)),
  \[8956]  = (~\[556]  & ~sh2) | (~\[555]  & sh2),
  \[11146]  = ~\[3515]  | (musel3 | (~musel4 | ~inD12)),
  \[1332]  = ~\[280]  & (musel3 & ~musel4),
  \[8388]  = (~\[6017]  & ~\[306] ) | ~\[10922] ,
  \[9117]  = (~\[5939]  & ~opsel2) | ~\[11298] ,
  \[3231]  = ~musel1 & ~musel2,
  \[11340]  = ~musel1 | (musel2 | ~inA8),
  \[8959]  = (~\[5988]  & ~\[561] ) | ~\[3348] ,
  \[11910]  = ~musel2 | (musel3 | ~inB10),
  \[4780]  = musel2 & inC5,
  \[1525]  = ~\[311]  & (musel1 & ~musel3),
  \[9119]  = (~\[177]  & ~e15) | (\[8181]  & ~\[5536] ),
  \[11342]  = ~\[5903]  | \[5849] ,
  \[1526]  = (~musel1 & ~\[11842] ) | (~musel1 & ~\[11840] ),
  \[1337]  = ~\[279]  & (musel1 & ~musel3),
  \[5701]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[1338]  = (~musel1 & ~\[11490] ) | (~musel1 & ~\[11488] ),
  \[5514]  = musel2 & inD15,
  \[5704]  = (~\[423]  & ~b7) | (\[423]  & b7),
  \[10998]  = ~\[3231]  | (musel3 | (~musel4 | ~inD10)),
  \[11348]  = ~musel1 | (musel2 | ~inA9),
  \[11728]  = ~musel2 | (musel3 | ~inB5),
  \[5517]  = ~musel1 & ~musel2,
  \[8962]  = (~\[564]  & ~sh0) | (~\[563]  & sh0),
  b0 = ~\[1364]  & ~\[1363] ,
  b1 = ~\[1382]  & ~\[1381] ,
  b2 = ~\[1400]  & ~\[1399] ,
  b3 = ~\[1424]  & ~\[1423] ,
  b4 = ~\[1442]  & ~\[1441] ,
  b5 = ~\[1460]  & ~\[1459] ,
  b6 = ~\[1478]  & ~\[1477] ,
  b7 = ~\[1502]  & ~\[1501] ,
  b8 = ~\[1520]  & ~\[1519] ,
  b9 = ~\[1538]  & ~\[1537] ,
  \[9314]  = (~\[252]  & ~e0) | (\[8992]  & ~\[6114] ),
  \[8965]  = (~\[570]  & ~sh0) | (~\[569]  & sh0),
  \[1910]  = musel2 & inD1,
  \[8586]  = (~\[6103]  & ~\[370] ) | ~\[10296] ,
  e0 = (~\[661]  & ~\[6115] ) | (~\[661]  & ~\[5840] ),
  e1 = (~\[697]  & ~\[6105] ) | (~\[697]  & ~\[9670] ),
  e2 = (~\[737]  & ~\[6094] ) | (~\[737]  & ~\[9647] ),
  e3 = (~\[782]  & ~\[9611] ) | (~\[782]  & ~\[6082] ),
  e5 = (~\[865]  & ~\[6063] ) | (~\[865]  & ~\[9772] ),
  e6 = (~\[905]  & ~\[6052] ) | (~\[905]  & ~\[9749] ),
  e7 = (~\[950]  & ~\[9713] ) | (~\[950]  & ~\[6038] ),
  \[8777]  = (~\[6073]  & \[6039] ) | (\[6073]  & ~\[6039] ),
  e9 = (~\[1035]  & ~\[6019] ) | (~\[1035]  & ~\[9876] ),
  \[11726]  = musel2 | (~musel3 | ~inD5),
  \[8968]  = (~\[576]  & ~sh0) | (~\[575]  & sh0),
  \[1913]  = ~musel1 & ~musel2,
  \[9507]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[11350]  = ~\[5897]  | \[5849] ,
  \[11920]  = musel2 | (~musel3 | ~inD11),
  \[1535]  = opsel2 & opsel3,
  \[11922]  = ~musel2 | (musel3 | ~inB11),
  \[5900]  = ~inC9 | ~musel2,
  \[1347]  = ~\[5843]  & ~\[5840] ,
  \[1537]  = ~musel1 & (~musel2 & (~\[5654]  & ~musel3)),
  \[1538]  = ~\[304]  & (musel3 & ~musel4),
  \[5712]  = (~\[1484]  & ~\[1483] ) | musel4,
  \[1349]  = ~opsel1 & (~opsel2 & opsel3),
  \[3626]  = musel2 & inD13,
  \[5713]  = ~inC6 | ~musel4,
  \[5903]  = ~\[9433]  | (musel3 | ~musel4),
  \[5904]  = (~\[5903]  & \[5849] ) | ~\[11342] ,
  \[5905]  = ~inC8 | ~musel2,
  \[11358]  = ~\[5892]  | \[5849] ,
  \[3629]  = ~musel1 & ~musel2,
  \[8971]  = (~\[582]  & ~sh0) | (~\[581]  & sh0),
  \[9511]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[9132]  = (~\[182]  & ~e14) | (\[8950]  & ~\[5951] ),
  \[5908]  = ~\[9449]  | (musel3 | ~musel4),
  \[8974]  = (~\[588]  & ~sh0) | (~\[587]  & sh0),
  \[5719]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[9513]  = (~\[5882]  & ~musel1) | ~\[11372] ,
  \[5909]  = (~\[5908]  & \[5849] ) | ~\[11334] ,
  \[1350]  = opsel1 & (opsel2 & ~opsel3),
  \[11544]  = musel2 | (~musel3 | ~inD0),
  \[11166]  = ~\[9145]  | (opsel2 | ~opsel3),
  \[11356]  = ~musel1 | (musel2 | ~inA10),
  \[11546]  = ~musel2 | (musel3 | ~inB0),
  \[8977]  = (~\[594]  & ~sh0) | (~\[593]  & sh0),
  \[1353]  = (~\[391]  & \[5799] ) | (~\[391]  & ~\[5789] ),
  \[1543]  = ~\[303]  & (musel1 & ~musel3),
  \[202]  = (~opsel0 & ~opsel1) | (opsel0 & opsel1),
  \[9707]  = \[5740]  | ~\[5730] ,
  \[1354]  = \[5799]  & ~\[5789] ,
  \[1544]  = (~musel1 & ~\[11876] ) | (~musel1 & ~\[11874] ),
  \[203]  = (~\[1005]  & \[204] ) | (~\[1005]  & ~\[6018] ),
  \[204]  = (~\[8920]  & ~\[8965] ) | ((~\[8920]  & ~opsel2) | (~\[8965]  & opsel2)),
  \[1356]  = \[5817]  & ~\[5807] ,
  \[1167]  = ~\[5970]  & ~\[5966] ,
  \[5911]  = ~\[5909]  | (~\[5904]  | (~\[5898]  | ~\[5893] )),
  \[5722]  = (~\[424]  & ~b6) | (\[424]  & b6),
  \[207]  = (~opsel0 & ~opsel1) | (opsel0 & opsel1),
  \[5533]  = ~musel3 | musel4,
  \[208]  = (~\[969]  & \[209] ) | (~\[969]  & ~\[6028] ),
  \[5913]  = ~inC3 | ~musel2,
  \[209]  = (~\[8923]  & ~\[8968] ) | ((~\[8923]  & ~opsel2) | (~\[8968]  & opsel2)),
  \[8980]  = (~\[600]  & ~sh0) | (~\[599]  & sh0),
  \[5156]  = musel2 & inC10,
  \[5536]  = opsel0 | opsel1,
  \[5916]  = ~\[9529]  | (musel3 | ~musel4),
  \[9331]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[5917]  = (~\[5916]  & \[5849] ) | ~\[11326] ,
  \[9711]  = \[5704]  | ~\[5694] ,
  \[9901]  = (~\[5763]  & ~\[511] ) | \[5760] ,
  b10 = ~\[1556]  & ~\[1555] ,
  b11 = ~\[1580]  & ~\[1579] ,
  b12 = ~\[1332]  & ~\[1331] ,
  \[8983]  = (~\[606]  & ~sh0) | (~\[605]  & sh0),
  b13 = ~\[1592]  & ~\[1591] ,
  b14 = ~\[1616]  & ~\[1615] ,
  b15 = ~\[1630]  & ~\[1629] ,
  \[5918]  = ~inC2 | ~musel2,
  \[9523]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[9713]  = (~\[438]  & \[9740] ) | ~\[9743] ,
  \[11364]  = ~musel1 | (musel2 | ~inA11),
  \[1361]  = opsel2 & opsel3,
  \[9145]  = (~\[187]  & ~e13) | (\[8953]  & ~\[5966] ),
  \[9335]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[8986]  = (~\[612]  & ~sh0) | (~\[611]  & sh0),
  \[210]  = (~\[9217]  & \[6028] ) | ((~\[9217]  & ~\[8968] ) | ((~\[8849]  & \[6028] ) | (~\[8849]  & ~\[8968] ))),
  \[9905]  = (~\[514]  & \[9932] ) | ~\[9935] ,
  \[11366]  = ~\[5885]  | \[5849] ,
  \[1363]  = ~musel1 & (~musel2 & (~\[5826]  & ~musel3)),
  \[1553]  = opsel2 & opsel3,
  \[9337]  = (~\[5846]  & ~musel1) | ~\[11424] ,
  \[9527]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[11180]  = ~\[5969]  | ~\[5859] ,
  \[1364]  = ~\[376]  & (musel3 & ~musel4),
  \[8989]  = (~\[618]  & ~sh0) | (~\[617]  & sh0),
  \[213]  = (~\[919]  & \[214] ) | (~\[919]  & ~\[6037] ),
  \[1555]  = ~musel1 & (~musel2 & (~\[5636]  & ~musel3)),
  \[9529]  = (~\[5913]  & ~musel1) | ~\[11332] ,
  \[214]  = (~\[8926]  & ~\[8971] ) | ((~\[8926]  & ~opsel2) | (~\[8971]  & opsel2)),
  \[9719]  = (~\[441]  & ~\[12805] ) | ~\[9731] ,
  \[11372]  = ~musel1 | (musel2 | ~inA4),
  \[1556]  = ~\[296]  & (musel3 & ~musel4),
  \[5730]  = (~\[1466]  & ~\[1465] ) | musel4,
  \[5731]  = ~inC5 | ~musel4,
  \[5921]  = ~\[9545]  | (musel3 | ~musel4),
  \[5542]  = (~\[1636]  & ~\[1635] ) | musel4,
  \[217]  = (~opsel0 & ~opsel1) | (opsel0 & opsel1),
  \[5922]  = (~\[5921]  & \[5849] ) | ~\[11318] ,
  \[3076]  = musel2 & inD9,
  \[1369]  = ~\[375]  & (musel1 & ~musel3),
  \[5543]  = ~inC15 | ~musel4,
  \[218]  = (~\[875]  & \[219] ) | (~\[875]  & ~\[6051] ),
  \[219]  = (~\[8929]  & ~\[8974] ) | ((~\[8929]  & ~opsel2) | (~\[8974]  & opsel2)),
  \[5924]  = ~inC1 | ~musel2,
  \[3079]  = ~musel1 & ~musel2,
  \[8992]  = (~\[624]  & ~sh0) | (~\[623]  & sh0),
  \[5737]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[5927]  = ~\[9561]  | (musel3 | ~musel4),
  \[9721]  = (~\[6039]  & ~\[12808] ) | ~\[9728] ,
  \[9911]  = (~\[517]  & ~\[12793] ) | ~\[9923] ,
  \[10204]  = ~sh2 | ~\[8611] ,
  \[5928]  = (~\[5927]  & \[5849] ) | ~\[11310] ,
  \[10013]  = (~sh1 & sh2) | ~\[11196] ,
  \[5929]  = ~inC0 | ~musel2,
  \[9913]  = (~\[5844]  & ~\[12796] ) | ~\[9920] ,
  \[1370]  = (~musel1 & ~\[11546] ) | (~musel1 & ~\[11544] ),
  \[11374]  = ~\[5880]  | \[5849] ,
  \[10015]  = (\[8286]  & ~sh0) | (\[8263]  & sh0),
  \[1561]  = ~\[295]  & (musel1 & ~musel3),
  \[600]  = (~\[10122]  & ~\[10118] ) | ((~\[10122]  & ~sh1) | (~\[10118]  & sh1)),
  \[1562]  = (~musel1 & ~\[11910] ) | (~musel1 & ~\[11908] ),
  \[10400]  = ~\[9275]  | (opsel2 | ~opsel3),
  \[411]  = (~\[12802]  & ~\[9655] ) | (~\[12802]  & ~\[5840] ),
  \[3270]  = ~\[5935]  & ~\[5911] ,
  \[9347]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[222]  = (~opsel0 & ~opsel1) | (opsel0 & opsel1),
  \[11380]  = ~musel1 | (musel2 | ~inA5),
  \[11760]  = musel2 | (~musel3 | ~inD6),
  \[223]  = (~\[835]  & \[224] ) | (~\[835]  & ~\[6062] ),
  \[9728]  = \[5758]  | ~\[5748] ,
  \[9539]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[224]  = (~\[8932]  & ~\[8977] ) | ((~\[8932]  & ~opsel2) | (~\[8977]  & opsel2)),
  \[11382]  = ~\[5874]  | \[5849] ,
  \[11762]  = ~musel2 | (musel3 | ~inB6),
  \[5740]  = (~\[425]  & ~b5) | (\[425]  & b5),
  \[605]  = (~\[10132]  & ~\[10128] ) | ((~\[10132]  & ~sh1) | (~\[10128]  & sh1)),
  \[1567]  = ~\[287]  & (musel1 & ~musel3),
  \[5551]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[606]  = (~\[10134]  & ~\[10130] ) | ((~\[10134]  & ~sh1) | (~\[10130]  & sh1)),
  \[1568]  = (~musel1 & ~\[11922] ) | (~musel1 & ~\[11920] ),
  \[227]  = (~opsel0 & ~opsel1) | (opsel0 & opsel1),
  \[5932]  = ~\[9577]  | (musel3 | ~musel4),
  \[1379]  = opsel2 & opsel3,
  \[228]  = (~\[799]  & \[229] ) | (~\[799]  & ~\[6072] ),
  \[5933]  = (~\[5932]  & \[5849] ) | ~\[11302] ,
  \[5554]  = (~\[506]  & ~b15) | (\[506]  & b15),
  \[229]  = (~\[8935]  & ~\[8980] ) | ((~\[8935]  & ~opsel2) | (~\[8980]  & opsel2)),
  \[5555]  = (~\[5554]  & ~\[5542] ) | ~\[12020] ,
  \[5935]  = ~\[5933]  | (~\[5928]  | (~\[5922]  | ~\[5917] )),
  \[11388]  = ~musel1 | (musel2 | ~inA6),
  \[11578]  = musel2 | (~musel3 | ~inD1),
  \[9920]  = ~\[5599]  | \[5609] ,
  \[10029]  = (\[8313]  & ~sh1) | (\[8263]  & sh1),
  \[9351]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[9731]  = ~\[5740]  | \[5730] ,
  \[5748]  = (~\[1448]  & ~\[1447] ) | musel4,
  \[9353]  = (~\[5850]  & ~musel1) | ~\[11420] ,
  \[5749]  = ~inC4 | ~musel4,
  \[9543]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[5939]  = ~pgx3 | (~\[5865]  | (~\[5859]  | ~\[5854] )),
  \[1190]  = (~\[5967]  & ~\[11226] ) | (~\[5967]  & ~\[9968] ),
  \[9923]  = \[5581]  | ~\[5591] ,
  \[1381]  = ~musel1 & (~musel2 & (~\[5808]  & ~musel3)),
  \[9165]  = (~opsel0 & opsel1) | (opsel0 & ~opsel1),
  \[9545]  = (~\[5918]  & ~musel1) | ~\[11324] ,
  \[230]  = (~\[9269]  & \[6072] ) | ((~\[9269]  & ~\[8980] ) | ((~\[8777]  & \[6072] ) | (~\[8777]  & ~\[8980] ))),
  \[11196]  = ~sh1 | ~\[5957] ,
  \[1382]  = ~\[368]  & (musel3 & ~musel4),
  \[611]  = (~\[10144]  & ~\[10140] ) | ((~\[10144]  & ~sh1) | (~\[10140]  & sh1)),
  \[612]  = (~\[10146]  & ~\[10142] ) | ((~\[10146]  & ~sh1) | (~\[10142]  & sh1)),
  \[11390]  = ~\[5869]  | \[5849] ,
  \[11580]  = ~musel2 | (musel3 | ~inB1),
  \[233]  = (~\[751]  & \[234] ) | (~\[751]  & ~\[6081] ),
  \[423]  = ~\[1499]  & (~opsel0 & ~\[5701] ),
  \[10031]  = (~\[562]  & ~sh0) | (~\[5990]  & \[8313] ),
  \[234]  = (~\[8938]  & ~\[8983] ) | ((~\[8938]  & ~opsel2) | (~\[8983]  & opsel2)),
  \[424]  = ~\[1475]  & (~opsel0 & ~\[5719] ),
  \[11772]  = musel2 | (~musel3 | ~inD7),
  \[425]  = ~\[1457]  & (~opsel0 & ~\[5737] ),
  \[1387]  = ~\[367]  & (musel1 & ~musel3),
  \[1577]  = opsel2 & opsel3,
  \[426]  = ~\[1439]  & (~opsel0 & ~\[5755] ),
  \[1388]  = (~musel1 & ~\[11580] ) | (~musel1 & ~\[11578] ),
  \[237]  = (~opsel0 & ~opsel1) | (opsel0 & opsel1),
  \[617]  = (~\[10156]  & ~\[10152] ) | ((~\[10156]  & ~sh1) | (~\[10152]  & sh1)),
  \[1579]  = ~musel1 & (~musel2 & (~\[5618]  & ~musel3)),
  \[5563]  = (~\[1604]  & ~\[1603] ) | musel4,
  \[238]  = (~\[707]  & \[239] ) | (~\[707]  & ~\[6093] ),
  \[618]  = (~\[10158]  & ~\[10154] ) | ((~\[10158]  & ~sh1) | (~\[10154]  & sh1)),
  \[5564]  = ~inC14 | ~musel4,
  \[6103]  = ~musel3 | musel4,
  \[239]  = (~\[8941]  & ~\[8986] ) | ((~\[8941]  & ~opsel2) | (~\[8986]  & opsel2)),
  \[10608]  = ~\[2493]  | (musel3 | (~musel4 | ~inD5)),
  \[6104]  = opsel0 | opsel1,
  \[5755]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[5945]  = ~musel3 | musel4,
  \[11398]  = ~\[5864]  | \[5849] ,
  \[6105]  = (~\[5817]  & ~\[5807] ) | (\[5817]  & \[5807] ),
  \[9740]  = ~\[5722]  | \[5712] ,
  \[9171]  = (~\[197]  & ~e11) | (\[8959]  & ~\[5992] ),
  \[5378]  = musel2 & inC14,
  e10 = (~\[1075]  & ~\[6008] ) | (~\[1075]  & ~\[9853] ),
  \[10224]  = ~\[1775]  | (musel3 | (~musel4 | ~inD0)),
  e11 = (~\[1115]  & ~\[9817] ) | (~\[1115]  & ~\[5993] ),
  e13 = (~\[1190]  & ~\[5967] ) | (~\[1190]  & ~\[9964] ),
  \[6107]  = ~\[5933]  | \[5849] ,
  \[10414]  = ~\[6086]  | ~\[5917] ,
  e14 = (~\[1221]  & ~\[5952] ) | (~\[1221]  & ~\[9941] ),
  \[5758]  = (~\[426]  & ~b4) | (\[426]  & b4),
  e15 = (~\[1312]  & ~\[9905] ) | (~\[1312]  & ~\[5555] ),
  \[9932]  = \[5563]  | ~\[5573] ,
  \[9363]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[6108]  = ~opsel2 | ~\[8944] ,
  \[9743]  = \[5722]  | ~\[5712] ,
  \[1580]  = ~\[288]  & (musel3 & ~musel4),
  \[11774]  = ~musel2 | (musel3 | ~inB7),
  \[9555]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[9935]  = ~\[5563]  | \[5573] ,
  \[11396]  = ~musel1 | (musel2 | ~inA7),
  \[1772]  = musel2 & inD0,
  \[9367]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[242]  = (~opsel0 & ~opsel1) | (opsel0 & opsel1),
  \[432]  = (~\[1434]  & ~\[4308] ) | (~\[1434]  & ~\[9707] ),
  \[243]  = (~\[667]  & \[244] ) | (~\[667]  & ~\[6104] ),
  \[623]  = (~\[10168]  & ~\[10164] ) | ((~\[10168]  & ~sh1) | (~\[10164]  & sh1)),
  \[1775]  = ~musel1 & ~musel2,
  \[9369]  = (~\[5855]  & ~musel1) | ~\[11412] ,
  \[9559]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[244]  = (~\[8944]  & ~\[8989] ) | ((~\[8944]  & ~opsel2) | (~\[8989]  & opsel2)),
  \[9749]  = ~\[10704]  | ~\[9766] ,
  \[624]  = (~\[10170]  & ~\[10166] ) | ((~\[10170]  & ~sh1) | (~\[10166]  & sh1)),
  \[5570]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[5760]  = (\[5704]  & ~\[5694] ) | ~\[11654] ,
  \[5950]  = (sh1 & ~sh2) | ~\[3736] ,
  \[1397]  = opsel2 & opsel3,
  \[5951]  = opsel0 | opsel1,
  \[247]  = (~opsel0 & ~opsel1) | (opsel0 & opsel1),
  \[5952]  = (~\[5563]  & ~\[5573] ) | (\[5563]  & \[5573] ),
  \[1399]  = ~musel1 & (~musel2 & (~\[5790]  & ~musel3)),
  \[1589]  = opsel2 & opsel3,
  \[5573]  = (~\[507]  & ~b14) | (\[507]  & b14),
  \[5763]  = ~\[4663]  | ~\[4666] ,
  \[248]  = (~\[631]  & \[249] ) | (~\[631]  & ~\[6114] ),
  \[438]  = (~\[12805]  & ~\[9721] ) | (~\[12805]  & ~\[9731] ),
  \[10048]  = (\[8335]  & ~sh2) | (\[8181]  & sh2),
  \[6113]  = ~musel3 | musel4,
  \[249]  = (~\[8947]  & ~\[8992] ) | ((~\[8947]  & ~opsel2) | (~\[8992]  & opsel2)),
  \[6114]  = opsel0 | opsel1,
  \[5955]  = ~\[5865]  | (~\[5859]  | ~pgx3),
  \[6115]  = (~\[5835]  & ~\[5825] ) | (\[5835]  & \[5825] ),
  \[11978]  = ~musel2 | (musel3 | ~inB13),
  \[5956]  = ~opsel2 | ~\[8905] ,
  \[9561]  = (~\[5924]  & ~musel1) | ~\[11316] ,
  \[5957]  = ~sh0 | ~sh2,
  \[9941]  = ~\[11282]  | ~\[9958] ,
  \[10044]  = (\[8286]  & ~sh2) | ~\[10978] ,
  \[6117]  = ~opsel2 | ~\[8947] ,
  \[9753]  = (\[9757]  & ~\[6039] ) | ~\[9760] ,
  \[10046]  = (\[8313]  & ~sh2) | (\[8181]  & sh2),
  \[9184]  = (~\[202]  & ~e10) | (\[8962]  & ~\[6007] ),
  pgx3 = ~\[5935]  & (~\[5849]  & (~\[5911]  & ~\[5888] )),
  \[1591]  = ~musel1 & (~musel2 & (~\[5582]  & ~musel3)),
  \[9755]  = ~\[10710]  | ~\[9757] ,
  \[9945]  = (\[9949]  & ~\[5844] ) | ~\[9952] ,
  \[10050]  = (\[8360]  & ~sh2) | (\[8263]  & sh2),
  \[1592]  = ~\[272]  & (musel3 & ~musel4),
  \[11976]  = musel2 | (~musel3 | ~inD13),
  \[441]  = (~\[12808]  & ~\[9728] ) | (~\[12808]  & ~\[6039] ),
  \[631]  = ~\[6117]  & ~\[6114] ,
  \[252]  = (~opsel0 & ~opsel1) | (opsel0 & opsel1),
  \[9757]  = ~\[5758]  | \[5748] ,
  \[9947]  = ~\[11288]  | ~\[9949] ,
  \[10432]  = ~sh2 | ~\[8540] ,
  \[9379]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[9949]  = \[5599]  | ~\[5609] ,
  \[4222]  = musel2 & inC12,
  \[255]  = (~musel2 & ~inA15) | ((musel2 & ~inC15) | (~inC15 & ~inA15)),
  \[1597]  = ~\[271]  & (musel1 & ~musel3),
  \[5581]  = (~\[1598]  & ~\[1597] ) | musel4,
  \[5771]  = (~\[1412]  & ~\[1411] ) | musel4,
  \[256]  = (~inA15 & ~\[5456] ) | ((~inA15 & ~musel1) | ((~\[9331]  & ~\[5456] ) | (~\[9331]  & ~musel1))),
  \[1598]  = (~musel1 & ~\[11978] ) | (~musel1 & ~\[11976] ),
  \[5582]  = ~inC13 | ~musel4,
  \[5772]  = ~inC3 | ~musel4,
  \[5962]  = ~musel3 | musel4,
  \[258]  = (~inB15 & ~\[5514] ) | ((~inB15 & ~musel1) | ((~\[9335]  & ~\[5514] ) | (~\[9335]  & ~musel1))),
  \[5963]  = ~sh1 | ~\[8286] ,
  \[10058]  = (\[8335]  & ~sh2) | (\[8181]  & sh2),
  \[11988]  = musel2 | (~musel3 | ~inD14),
  \[5966]  = opsel0 | opsel1,
  \[9760]  = \[5758]  | ~\[5748] ,
  \[9571]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[5967]  = (~\[5581]  & ~\[5591] ) | (\[5581]  & \[5591] ),
  \[10244]  = ~\[9301]  | (opsel2 | ~opsel3),
  \[5588]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[5778]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[9952]  = ~\[5599]  | \[5609] ,
  \[9383]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[5969]  = ~pgx3 | ~\[5865] ,
  \[9763]  = ~\[5740]  | \[5730] ,
  \[10056]  = (\[8313]  & ~sh2) | ~\[10902] ,
  \[9385]  = (~\[5861]  & ~musel1) | ~\[11404] ,
  \[9575]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[9955]  = \[5581]  | ~\[5591] ,
  \[10060]  = (\[8360]  & ~sh2) | (\[8263]  & sh2),
  \[10630]  = ~\[9779]  | ~\[6039] ,
  \[9766]  = \[5740]  | ~\[5730] ,
  \[9197]  = (~\[207]  & ~e9) | (\[8965]  & ~\[6018] ),
  \[9577]  = (~\[5929]  & ~musel1) | ~\[11308] ,
  \[10062]  = (\[8388]  & ~sh2) | (\[8286]  & sh2),
  \[11990]  = ~musel2 | (musel3 | ~inB14),
  \[263]  = (~musel2 & ~inA14) | ((musel2 & ~inC14) | (~inC14 & ~inA14)),
  \[10632]  = ~\[9236]  | (opsel2 | ~opsel3),
  \[9958]  = ~\[5581]  | \[5591] ,
  \[264]  = (~inA14 & ~\[5378] ) | ((~inA14 & ~musel1) | ((~\[9347]  & ~\[5378] ) | (~\[9347]  & ~musel1))),
  \[5970]  = ~opsel2 | ~\[8908] ,
  \[835]  = ~\[6066]  & ~\[6062] ,
  \[5591]  = (~\[508]  & ~b13) | (\[508]  & b13),
  \[5781]  = (~\[381]  & ~b3) | (\[381]  & b3),
  \[266]  = (~inB14 & ~\[3762] ) | ((~inB14 & ~musel1) | ((~\[9351]  & ~\[3762] ) | (~\[9351]  & ~musel1))),
  \[10068]  = (\[8335]  & ~sh2) | ~\[10830] ,
  \[10258]  = ~\[6107]  | ~\[5928] ,
  \[5975]  = ~musel3 | musel4,
  \[5976]  = ~sh0 | ~sh1,
  \[5977]  = ~sh0 | sh1,
  \[5978]  = (~\[5977]  & \[8286] ) | (~\[5976]  & \[8181] ),
  \[9772]  = (\[9776]  & ~\[6039] ) | ~\[9779] ,
  \[5599]  = (~\[1338]  & ~\[1337] ) | musel4,
  \[5789]  = (~\[1406]  & ~\[1405] ) | musel4,
  \[5979]  = opsel0 | opsel1,
  \[9964]  = (\[9968]  & ~\[5844] ) | ~\[9971] ,
  \[9395]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[10070]  = (\[8360]  & ~sh2) | (\[8181]  & sh2),
  \[271]  = (~musel2 & ~inA13) | ((musel2 & ~inC13) | (~inC13 & ~inA13)),
  \[9776]  = ~\[5758]  | \[5748] ,
  \[8418]  = (~\[6027]  & ~\[314] ) | ~\[10850] ,
  \[10830]  = ~sh2 | ~\[8418] ,
  \[272]  = (~inA13 & ~\[5304] ) | ((~inA13 & ~musel1) | ((~\[9363]  & ~\[5304] ) | (~\[9363]  & ~musel1))),
  \[10072]  = (\[8388]  & ~sh2) | (\[8286]  & sh2),
  \[10452]  = ~\[2231]  | (musel3 | (~musel4 | ~inD3)),
  \[9968]  = \[5599]  | ~\[5609] ,
  \[9399]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[274]  = (~inB13 & ~\[3626] ) | ((~inB13 & ~musel1) | ((~\[9367]  & ~\[3626] ) | (~\[9367]  & ~musel1))),
  \[9779]  = \[5758]  | ~\[5748] ,
  \[464]  = ~\[1577]  & (~opsel0 & ~\[5624] ),
  \[5790]  = ~inC2 | ~musel4,
  \[5980]  = (~\[5599]  & ~\[5609] ) | (\[5599]  & \[5609] ),
  \[465]  = ~\[1553]  & (~opsel0 & ~\[5642] ),
  \[5981]  = opsel2 | ~opsel3,
  \[466]  = ~\[1535]  & (~opsel0 & ~\[5660] ),
  \[5982]  = ~opsel2 | ~\[8911] ,
  \[467]  = ~\[1517]  & (~opsel0 & ~\[5678] ),
  \[468]  = ~\[5837]  & ~\[1130] ,
  \[279]  = (~musel2 & ~inA12) | ((musel2 & ~inC12) | (~inC12 & ~inA12)),
  \[8611]  = (~\[6113]  & ~\[378] ) | ~\[10224] ,
  \[5796]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[5987]  = ~musel3 | musel4,
  \[9971]  = ~\[5599]  | \[5609] ,
  \[10074]  = (\[8418]  & ~sh2) | (\[8313]  & sh2),
  \[5988]  = ~sh0 | ~sh1,
  \[5799]  = (~\[382]  & ~b2) | (\[382]  & b2),
  \[10646]  = ~\[6055]  | ~\[5875] ,
  \[280]  = (~inA12 & ~\[4222] ) | ((~inA12 & ~musel1) | ((~\[9379]  & ~\[4222] ) | (~\[9379]  & ~musel1))),
  \[10080]  = (\[8360]  & ~sh2) | ~\[10744] ,
  \[661]  = ~\[6115]  & ~\[5840] ,
  \[2352]  = musel2 & inD4,
  \[282]  = (~inB12 & ~\[3512] ) | ((~inB12 & ~musel1) | ((~\[9383]  & ~\[3512] ) | (~\[9383]  & ~musel1))),
  \[10082]  = (\[8388]  & ~sh2) | (\[8181]  & sh2),
  \[2355]  = ~musel1 & ~musel2,
  \[5990]  = ~sh0 | sh1,
  \[287]  = (~musel2 & ~inA11) | ((musel2 & ~inC11) | (~inC11 & ~inA11)),
  \[5992]  = opsel0 | opsel1,
  \[667]  = ~\[6108]  & ~\[6104] ,
  \[288]  = (~inA11 & ~\[5256] ) | ((~inA11 & ~musel1) | ((~\[9395]  & ~\[5256] ) | (~\[9395]  & ~musel1))),
  \[5993]  = (\[5627]  & \[5617] ) | ~\[11100] ,
  \[10468]  = ~\[9615]  | ~\[9638] ,
  \[5994]  = (~\[468]  & ~\[5763] ) | \[5760] ,
  \[10084]  = (\[8418]  & ~sh2) | (\[8313]  & sh2),
  \[5998]  = ~\[3270]  | \[5849] ,
  \[10086]  = (\[8440]  & ~sh2) | (\[8335]  & sh2),
  \[10276]  = ~sh2 | ~\[8586] ,
  \[290]  = (~inB11 & ~\[3388] ) | ((~inB11 & ~musel1) | ((~\[9399]  & ~\[3388] ) | (~\[9399]  & ~musel1))),
  \[480]  = (~\[12811]  & ~\[9825] ) | (~\[12811]  & ~\[9835] ),
  \[10850]  = ~\[2941]  | (musel3 | (~musel4 | ~inD8)),
  \[10092]  = (\[8388]  & ~sh2) | ~\[10664] ,
  \[1005]  = ~\[6022]  & ~\[6018] ,
  \[483]  = (~\[484]  & ~\[9832] ) | (~\[484]  & ~\[5994] ),
  \[4640]  = musel2 & inC3,
  \[484]  = \[5681]  & ~\[5671] ,
  \[295]  = (~musel2 & ~inA10) | ((musel2 & ~inC10) | (~inC10 & ~inA10)),
  \[865]  = (~\[6063]  & ~\[10630] ) | (~\[6063]  & ~\[9776] ),
  \[296]  = (~inA10 & ~\[5156] ) | ((~inA10 & ~musel1) | ((~\[9411]  & ~\[5156] ) | (~\[9411]  & ~musel1))),
  \[298]  = (~inB10 & ~\[3228] ) | ((~inB10 & ~musel1) | ((~\[9415]  & ~\[3228] ) | (~\[9415]  & ~musel1))),
  \[2938]  = musel2 & inD8,
  \[10098]  = (\[8464]  & ~sh2) | (\[8360]  & sh2),
  \[489]  = \[5645]  & ~\[5635] ,
  \[8440]  = (~\[6036]  & ~\[322] ) | ~\[10764] ,
  \[11018]  = ~\[9857]  | ~\[9867] ,
  \[10094]  = (\[8418]  & ~sh2) | (\[8263]  & sh2),
  \[10474]  = ~\[9617]  | ~\[9641] ,
  \[10664]  = ~sh2 | ~\[8464] ,
  \[11014]  = \[5645]  | \[5635] ,
  \[1200]  = ~\[5956]  & ~\[5951] ,
  \[11204]  = ~\[3629]  | (musel3 | (~musel4 | ~inD13)),
  \[10096]  = (\[8440]  & ~sh2) | (\[8335]  & sh2),
  \[10476]  = ~\[9621]  | ~\[9635] ,
  \[2941]  = ~musel1 & ~musel2,
  \[11022]  = ~\[9859]  | ~\[9870] ,
  \[875]  = ~\[6056]  & ~\[6051] ,
  \[496]  = \[5681]  & ~\[5671] ,
  \[4466]  = musel2 & inC1,
  \[10868]  = \[5681]  | \[5671] ,
  \[8263]  = (~\[5945]  & ~\[266] ) | ~\[11262] ,
  \[5008]  = musel2 & inC8,
  \[11024]  = ~\[9864]  | ~\[5994] ,
  \[1400]  = ~\[360]  & (musel3 & ~musel4),
  \[11404]  = ~musel1 | (musel2 | ~inA12),
  \[10296]  = ~\[1913]  | (musel3 | (~musel4 | ~inD1)),
  \[11026]  = ~\[9171]  | (opsel2 | ~opsel3),
  \[11406]  = ~\[5858]  | \[5849] ,
  \[10870]  = ~\[9197]  | (opsel2 | ~opsel3),
  \[1405]  = ~\[359]  & (musel1 & ~musel3),
  \[1406]  = (~musel1 & ~\[11614] ) | (~musel1 & ~\[11612] ),
  \[11412]  = ~musel1 | (musel2 | ~inA13),
  \[4663]  = (\[5758]  & \[5740] ) | ((\[5758]  & ~\[5730] ) | ((~\[5748]  & \[5740] ) | (~\[5748]  & ~\[5730] ))),
  \[697]  = (~\[6105]  & ~\[10318] ) | (~\[6105]  & ~\[9674] ),
  \[4854]  = musel2 & inC6,
  \[4666]  = (\[5722]  & \[5704] ) | ((\[5722]  & ~\[5694] ) | ((~\[5712]  & \[5704] ) | (~\[5712]  & ~\[5694] ))),
  \[11228]  = ~\[9132]  | (opsel2 | ~opsel3),
  \[10684]  = ~\[2645]  | (musel3 | (~musel4 | ~inD6)),
  \[8464]  = (~\[6050]  & ~\[330] ) | ~\[10684] ,
  \[1221]  = (~\[5952]  & ~\[11286] ) | (~\[5952]  & ~\[9955] ),
  \[1411]  = ~\[351]  & (musel1 & ~musel3),
  \[11226]  = ~\[9971]  | ~\[5844] ,
  \[1412]  = (~musel1 & ~\[11626] ) | (~musel1 & ~\[11624] ),
  \[1603]  = ~\[263]  & (musel1 & ~musel3),
  \[11040]  = ~\[6000]  | ~\[5893] ,
  \[11420]  = ~musel1 | (musel2 | ~inA14),
  \[1604]  = (~musel1 & ~\[11990] ) | (~musel1 & ~\[11988] ),
  \[8849]  = (~\[6029]  & \[5994] ) | (\[6029]  & ~\[5994] ),
  \[1035]  = (~\[6019]  & ~\[10944] ) | (~\[6019]  & ~\[9880] ),
  \[11612]  = musel2 | (~musel3 | ~inD2),
  O10 = \[5] ,
  O11 = \[4] ,
  O12 = \[3] ,
  O13 = \[2] ,
  O14 = \[1] ,
  O15 = \[0] ,
  \[10884]  = ~\[6021]  | ~\[5904] ,
  \[11424]  = ~musel1 | (musel2 | ~inA15),
  \[11614]  = ~musel2 | (musel3 | ~inB2),
  \[8286]  = (~\[5962]  & ~\[274] ) | ~\[11204] ,
  \[1421]  = opsel2 & opsel3,
  \[11806]  = (~\[1512]  & ~\[1511] ) | (~\[5645]  & \[5635] ),
  \[1423]  = ~musel1 & (~musel2 & (~\[5772]  & ~musel3)),
  \[1613]  = opsel2 & opsel3,
  \[1424]  = ~\[352]  & (musel3 & ~musel4),
  \[1045]  = ~\[6012]  & ~\[6007] ,
  \[1235]  = ~\[5939]  & (~\[5536]  & opsel2),
  \[1615]  = ~musel1 & (~musel2 & (~\[5564]  & ~musel3)),
  \[3512]  = musel2 & inD12,
  \[11242]  = ~\[5955]  | ~\[5854] ,
  \[12790]  = ~\[5935]  & ~\[5849] ,
  \[1616]  = ~\[264]  & (musel3 & ~musel4),
  \[5600]  = ~inC12 | ~musel4,
  \[3515]  = ~musel1 & ~musel2,
  \[10]  = (~\[223]  & ~opsel3) | ~\[10556] ,
  \[11]  = (~\[228]  & ~opsel3) | (~\[6074]  & ~\[230] ),
  \[12]  = (~\[233]  & ~opsel3) | ~\[10400] ,
  \[13]  = (~\[238]  & ~opsel3) | ~\[10320] ,
  \[5606]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[14]  = (~\[243]  & ~opsel3) | ~\[10244] ,
  \[9401]  = (~\[5889]  & ~musel1) | ~\[11364] ,
  \[15]  = (~\[248]  & ~opsel3) | ~\[10172] ,
  \[5609]  = (~\[509]  & ~b12) | (\[509]  & b12),
  \[11434]  = ~\[5517]  | (musel3 | (~musel4 | ~inD15)),
  \[11624]  = musel2 | (~musel3 | ~inD3),
  \[12799]  = ~\[5835]  & \[5825] ,
  \[1431]  = (~\[432]  & \[5722] ) | (~\[432]  & ~\[5712] ),
  \[1432]  = \[5722]  & ~\[5712] ,
  \[11626]  = ~musel2 | (musel3 | ~inB3),
  \[12793]  = \[5581]  & ~\[5591] ,
  \[9217]  = (~opsel0 & opsel1) | (opsel0 & ~opsel1),
  \[12796]  = ~\[5599]  & \[5609] ,
  \[1434]  = \[5740]  & ~\[5730] ,
  \[1627]  = opsel2 & opsel3,
  \[1439]  = opsel2 & opsel3,
  \[1629]  = ~musel1 & (~musel2 & (~\[5543]  & ~musel3)),
  \[11068]  = ~\[3391]  | (musel3 | (~musel4 | ~inD11)),
  \[8491]  = (~\[6061]  & ~\[338] ) | ~\[10608] ,
  \[5617]  = (~\[1568]  & ~\[1567] ) | musel4,
  \[9411]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[5807]  = (~\[1388]  & ~\[1387] ) | musel4,
  \[5618]  = ~inC11 | ~musel4,
  \[5808]  = ~inC1 | ~musel4,
  \[9223]  = (~\[217]  & ~e7) | (\[8971]  & ~\[6037] ),
  \[11254]  = ~\[5950]  | ~\[8181] ,
  \[1630]  = ~\[256]  & (musel3 & ~musel4),
  \[1441]  = ~musel1 & (~musel2 & (~\[5749]  & ~musel3)),
  \[9415]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[9605]  = \[5817]  | ~\[5807] ,
  \[1442]  = ~\[344]  & (musel3 & ~musel4),
  \[9417]  = (~\[5894]  & ~musel1) | ~\[11356] ,
  \[1635]  = ~\[255]  & (musel1 & ~musel3),
  \[9609]  = \[5781]  | ~\[5771] ,
  \[11262]  = ~\[3765]  | (musel3 | (~musel4 | ~inD14)),
  \[1636]  = (~musel1 & ~\[12050] ) | (~musel1 & ~\[12048] ),
  \[1447]  = ~\[343]  & (musel1 & ~musel3),
  \[1448]  = (~musel1 & ~\[11694] ) | (~musel1 & ~\[11692] ),
  \[5624]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[5814]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[3348]  = (~\[10031]  & ~\[3404] ) | ((~\[10031]  & ~\[5988] ) | ((~\[3404]  & sh2) | (~\[5988]  & sh2))),
  \[5627]  = (~\[464]  & ~b11) | (\[464]  & b11),
  \[5817]  = (~\[383]  & ~b1) | (\[383]  & b1),
  \[9611]  = ~\[10468]  | ~\[9641] ,
  \[9615]  = (~\[399]  & \[9629] ) | ~\[9635] ,
  \[11456]  = ~\[9911]  | ~\[9935] ,
  \[9236]  = (~\[222]  & ~e6) | (\[8974]  & ~\[6051] ),
  \[9427]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[9617]  = ~\[10476]  | ~\[9629] ,
  \[9807]  = (\[5645]  & ~\[5635] ) | ~\[11806] ,
  \[11840]  = musel2 | (~musel3 | ~inD8),
  \[303]  = (~musel2 & ~inA9) | ((musel2 & ~inC9) | (~inC9 & ~inA9)),
  \[1075]  = (~\[6008]  & ~\[11022] ) | (~\[6008]  & ~\[9867] ),
  \[304]  = (~inA9 & ~\[5082] ) | ((~inA9 & ~musel1) | ((~\[9427]  & ~\[5082] ) | (~\[9427]  & ~musel1))),
  \[11842]  = ~musel2 | (musel3 | ~inB8),
  \[1457]  = opsel2 & opsel3,
  \[306]  = (~inB9 & ~\[3076] ) | ((~inB9 & ~musel1) | ((~\[9431]  & ~\[3076] ) | (~\[9431]  & ~musel1))),
  \[1459]  = ~musel1 & (~musel2 & (~\[5731]  & ~musel3)),
  \[3736]  = (~sh0 & ~sh2) | ((sh0 & sh1) | (sh1 & ~sh2)),
  \[10108]  = (\[8464]  & ~sh2) | (\[8360]  & sh2),
  \[5635]  = (~\[1562]  & ~\[1561] ) | musel4,
  \[5825]  = (~\[1370]  & ~\[1369] ) | musel4,
  \[5256]  = musel2 & inC11,
  \[5636]  = ~inC10 | ~musel4,
  \[5826]  = ~inC0 | ~musel4,
  \[9431]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[9621]  = (~\[5840]  & ~\[12799] ) | ~\[9623] ,
  \[10104]  = (\[8418]  & ~sh2) | ~\[10588] ,
  \[9433]  = (~\[5900]  & ~musel1) | ~\[11348] ,
  \[9623]  = ~\[5835]  | \[5825] ,
  \[1460]  = ~\[336]  & (musel3 & ~musel4),
  \[10106]  = (\[8440]  & ~sh2) | (\[8286]  & sh2),
  \[11654]  = (~\[1432]  & ~\[1431] ) | ~\[9711] ,
  \[9815]  = \[5627]  | ~\[5617] ,
  \[10110]  = (\[8491]  & ~sh2) | (\[8388]  & sh2),
  \[311]  = (~musel2 & ~inA8) | ((musel2 & ~inC8) | (~inC8 & ~inA8)),
  \[312]  = (~inA8 & ~\[5008] ) | ((~inA8 & ~musel1) | ((~\[9443]  & ~\[5008] ) | (~\[9443]  & ~musel1))),
  \[11090]  = ~\[9823]  | ~\[9847] ,
  \[9817]  = (~\[480]  & ~\[489] ) | ~\[9847] ,
  \[8899]  = (~\[5980]  & \[5844] ) | (\[5980]  & ~\[5844] ),
  \[503]  = \[5681]  & ~\[5671] ,
  \[1465]  = ~\[335]  & (musel1 & ~musel3),
  \[9249]  = (~\[227]  & ~e5) | (\[8977]  & ~\[6062] ),
  \[9629]  = ~\[5817]  | \[5807] ,
  \[314]  = (~inB8 & ~\[2938] ) | ((~inB8 & ~musel1) | ((~\[9447]  & ~\[2938] ) | (~\[9447]  & ~musel1))),
  \[11282]  = ~\[9945]  | ~\[9955] ,
  \[1466]  = (~musel1 & ~\[11728] ) | (~musel1 & ~\[11726] ),
  \[506]  = ~\[1627]  & (~opsel0 & ~\[5551] ),
  \[5642]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[5832]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[1089]  = ~\[6001]  & ~\[5992] ,
  \[507]  = ~\[1613]  & (~opsel0 & ~\[5570] ),
  \[508]  = ~\[1589]  & (~opsel0 & ~\[5588] ),
  \[10118]  = (\[8464]  & ~sh2) | (\[8313]  & sh2),
  \[319]  = (~musel2 & ~inA7) | ((musel2 & ~inC7) | (~inC7 & ~inA7)),
  \[509]  = ~\[1329]  & (~opsel0 & ~\[5606] ),
  \[5645]  = (~\[465]  & ~b10) | (\[465]  & b10),
  \[5835]  = (~\[384]  & ~b0) | (\[384]  & b0),
  \[11288]  = ~\[9952]  | ~\[5844] ,
  \[5456]  = musel2 & inC15,
  \[5837]  = (\[5781]  & ~\[5771] ) | ~\[11506] ,
  \[9443]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[9823]  = (~\[483]  & ~\[12811] ) | ~\[9835] ,
  \[10116]  = (\[8440]  & ~sh2) | ~\[10516] ,
  \[9635]  = \[5817]  | ~\[5807] ,
  \[320]  = (~inA7 & ~\[4954] ) | ((~inA7 & ~musel1) | ((~\[9459]  & ~\[4954] ) | (~\[9459]  & ~musel1))),
  \[9825]  = (~\[5994]  & ~\[484] ) | ~\[9832] ,
  \[11286]  = ~\[9947]  | ~\[9958] ,
  \[10120]  = (\[8491]  & ~sh2) | (\[8388]  & sh2),
  \[511]  = ~\[5837]  & ~\[1347] ,
  \[9447]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[322]  = (~inB7 & ~\[2814] ) | ((~inB7 & ~musel1) | ((~\[9463]  & ~\[2814] ) | (~\[9463]  & ~musel1))),
  \[11290]  = ~\[9119]  | (opsel2 | ~opsel3),
  \[10122]  = (\[8520]  & ~sh2) | (\[8418]  & sh2),
  \[9638]  = ~\[5799]  | \[5789] ,
  \[1475]  = opsel2 & opsel3,
  \[12020]  = ~\[5554]  | ~\[5542] ,
  \[9449]  = (~\[5905]  & ~musel1) | ~\[11340] ,
  \[514]  = (~\[12793]  & ~\[9913] ) | (~\[12793]  & ~\[9923] ),
  \[5840]  = (~\[1350]  & ~\[1349] ) | opsel0,
  \[1477]  = ~musel1 & (~musel2 & (~\[5713]  & ~musel3)),
  \[6000]  = \[5998]  | (~\[5909]  | (~\[5904]  | ~\[5898] )),
  \[5082]  = musel2 & inC9,
  \[1478]  = ~\[328]  & (musel3 & ~musel4),
  \[6001]  = ~opsel2 | ~\[8914] ,
  \[327]  = (~musel2 & ~inA6) | ((musel2 & ~inC6) | (~inC6 & ~inA6)),
  \[517]  = (~\[12796]  & ~\[9920] ) | (~\[12796]  & ~\[5844] ),
  \[707]  = ~\[6098]  & ~\[6093] ,
  \[5653]  = (~\[1544]  & ~\[1543] ) | musel4,
  \[5843]  = ~\[4349]  | ~\[4352] ,
  \[328]  = (~inA6 & ~\[4854] ) | ((~inA6 & ~musel1) | ((~\[9475]  & ~\[4854] ) | (~\[9475]  & ~musel1))),
  \[10128]  = (\[8464]  & ~sh2) | ~\[10432] ,
  \[10318]  = ~\[9677]  | \[5840] ,
  \[5654]  = ~inC9 | ~musel4,
  \[5844]  = ~G3 | ~\[11496] ,
  \[11298]  = ~opsel2 | ~\[8181] ,
  \[11488]  = musel2 | (~musel3 | ~inD12),
  \[5846]  = ~inC15 | ~musel2,
  \[6006]  = ~musel3 | musel4,
  \[9641]  = \[5799]  | ~\[5789] ,
  \[6007]  = opsel0 | opsel1,
  \[9832]  = \[5681]  | ~\[5671] ,
  \[6008]  = (\[5645]  & \[5635] ) | ~\[11014] ,
  \[5849]  = ~\[9337]  | (musel3 | ~musel4),
  \[10316]  = ~\[9674]  | ~\[5840] ,
  \[330]  = (~inB6 & ~\[2642] ) | ((~inB6 & ~musel1) | ((~\[9479]  & ~\[2642] ) | (~\[9479]  & ~musel1))),
  \[9835]  = ~\[5663]  | \[5653] ,
  \[10130]  = (\[8491]  & ~sh2) | (\[8335]  & sh2),
  \[10320]  = ~\[9288]  | (opsel2 | ~opsel3),
  \[1483]  = ~\[327]  & (musel1 & ~musel3),
  \[9647]  = (~\[411]  & \[9661] ) | ~\[9664] ,
  \[1484]  = (~musel1 & ~\[11762] ) | (~musel1 & ~\[11760] ),
  \[11490]  = ~musel2 | (musel3 | ~inB12),
  \[10132]  = (\[8520]  & ~sh2) | (\[8418]  & sh2),
  \[9269]  = (~opsel0 & opsel1) | (opsel0 & ~opsel1),
  \[3762]  = musel2 & inD14,
  \[9459]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[5660]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[5850]  = ~inC14 | ~musel2,
  \[335]  = (~musel2 & ~inA5) | ((musel2 & ~inC5) | (~inC5 & ~inA5)),
  \[905]  = (~\[6052]  & ~\[10708] ) | (~\[6052]  & ~\[9763] ),
  \[336]  = (~inA5 & ~\[4780] ) | ((~inA5 & ~musel1) | ((~\[9491]  & ~\[4780] ) | (~\[9491]  & ~musel1))),
  \[6011]  = \[5998]  | (~\[5909]  | ~\[5904] ),
  \[3765]  = ~musel1 & ~musel2,
  \[1489]  = ~\[319]  & (musel1 & ~musel3),
  \[6012]  = ~opsel2 | ~\[8917] ,
  \[5663]  = (~\[466]  & ~b9) | (\[466]  & b9),
  \[5853]  = ~\[9353]  | (musel3 | ~musel4),
  \[338]  = (~inB5 & ~\[2490] ) | ((~inB5 & ~musel1) | ((~\[9495]  & ~\[2490] ) | (~\[9495]  & ~musel1))),
  \[5854]  = (~\[5849]  & \[5853] ) | (\[5849]  & ~\[5853] ),
  \[10708]  = ~\[9755]  | ~\[9766] ,
  \[3388]  = musel2 & inD11,
  \[5855]  = ~inC13 | ~musel2,
  \[4308]  = \[5758]  & ~\[5748] ,
  \[10134]  = (\[8540]  & ~sh2) | (\[8440]  & sh2),
  \[6017]  = ~musel3 | musel4,
  \[5858]  = ~\[9369]  | (musel3 | ~musel4),
  \[10704]  = ~\[9753]  | ~\[9763] ,
  \[6018]  = opsel0 | opsel1,
  \[9463]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[5859]  = (~\[5858]  & \[5849] ) | ~\[11406] ,
  \[9653]  = (~\[5840]  & ~\[12802] ) | ~\[9655] ,
  \[1490]  = (~musel1 & ~\[11774] ) | (~musel1 & ~\[11772] ),
  \[6019]  = (~\[5663]  & ~\[5653] ) | (\[5663]  & \[5653] ),
  \[11874]  = musel2 | (~musel3 | ~inD9),
  \[10516]  = ~sh2 | ~\[8520] ,
  \[9844]  = ~\[5645]  | \[5635] ,
  \[9275]  = (~\[237]  & ~e3) | (\[8983]  & ~\[6081] ),
  \[9465]  = (~\[5866]  & ~musel1) | ~\[11396] ,
  \[9655]  = ~\[5835]  | \[5825] ,
  \[11496]  = ~\[4965]  | (~\[4968]  | ~\[9901] ),
  \[10140]  = (\[8491]  & ~sh2) | ~\[10352] ,
  \[11876]  = ~musel2 | (musel3 | ~inB9),
  \[10710]  = ~\[9760]  | ~\[6039] ,
  \[9847]  = \[5645]  | ~\[5635] ,
  \[3391]  = ~musel1 & ~musel2,
  \[10142]  = (\[8520]  & ~sh2) | (\[8360]  & sh2),
  \[343]  = (~musel2 & ~inA4) | ((musel2 & ~inC4) | (~inC4 & ~inA4)),
  \[10712]  = ~\[9223]  | (opsel2 | ~opsel3),
  \[10902]  = ~sh2 | ~\[8388] ,
  \[344]  = (~inA4 & ~\[4706] ) | ((~inA4 & ~musel1) | ((~\[9507]  & ~\[4706] ) | (~\[9507]  & ~musel1))),
  \[11692]  = musel2 | (~musel3 | ~inD4),
  \[5671]  = (~\[1526]  & ~\[1525] ) | musel4,
  \[5861]  = ~inC12 | ~musel2,
  \[346]  = (~inB4 & ~\[2352] ) | ((~inB4 & ~musel1) | ((~\[9511]  & ~\[2352] ) | (~\[9511]  & ~musel1))),
  \[12802]  = ~\[5835]  & \[5825] ,
  \[6021]  = \[5998]  | ~\[5909] ,
  \[5672]  = ~inC8 | ~musel4,
  \[1499]  = opsel2 & opsel3,
  \[2228]  = musel2 & inD3,
  \[6022]  = ~opsel2 | ~\[8920] ,
  \[5864]  = ~\[9385]  | (musel3 | ~musel4),
  \[919]  = ~\[6045]  & ~\[6037] ,
  \[5865]  = (~\[5864]  & \[5849] ) | ~\[11398] ,
  \[5866]  = ~inC7 | ~musel2,
  \[12048]  = musel2 | (~musel3 | ~inD15),
  \[9661]  = ~\[5817]  | \[5807] ,
  \[12808]  = \[5758]  & ~\[5748] ,
  \[10144]  = (\[8540]  & ~sh2) | (\[8440]  & sh2),
  \[6027]  = ~musel3 | musel4,
  \[10334]  = ~\[6097]  | ~\[5922] ,
  \[5678]  = (~opsel1 & ~opsel3) | (opsel1 & ~opsel2),
  \[6028]  = opsel0 | opsel1,
  \[5869]  = ~\[9465]  | (musel3 | ~musel4),
  \[9853]  = ~\[11018]  | ~\[9870] ,
  \[10146]  = (\[8562]  & ~sh2) | (\[8464]  & sh2),
  \[11694]  = ~musel2 | (musel3 | ~inB4),
  \[6029]  = (\[5681]  & \[5671] ) | ~\[10868] ,
  \[9664]  = \[5817]  | ~\[5807] ,
  \[9475]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[2231]  = ~musel1 & ~musel2,
  \[351]  = (~musel2 & ~inA3) | ((musel2 & ~inC3) | (~inC3 & ~inA3)),
  \[352]  = (~inA3 & ~\[4640] ) | ((~inA3 & ~musel1) | ((~\[9523]  & ~\[4640] ) | (~\[9523]  & ~musel1))),
  \[9857]  = (~\[5994]  & ~\[496] ) | ~\[9864] ,
  \[10152]  = (\[8520]  & ~sh2) | ~\[10276] ,
  \[9288]  = (~\[242]  & ~e2) | (\[8986]  & ~\[6093] ),
  \[12805]  = ~\[5740]  & \[5730] ,
  \[12050]  = ~musel2 | (musel3 | ~inB15),
  \[3592]  = (~\[3600]  & ~\[10013] ) | ((~\[3600]  & ~\[8181] ) | ((~\[10015]  & ~\[10013] ) | (~\[10015]  & ~\[8181] ))),
  \[9479]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[354]  = (~inB3 & ~\[2228] ) | ((~inB3 & ~musel1) | ((~\[9527]  & ~\[2228] ) | (~\[9527]  & ~musel1))),
  \[9859]  = ~\[11024]  | ~\[9861] ,
  \[5870]  = (~\[5869]  & \[5849] ) | ~\[11390] ,
  \[6030]  = opsel2 | ~opsel3,
  \[5681]  = (~\[467]  & ~b8) | (\[467]  & b8),
  \[5871]  = ~inC6 | ~musel2,
  \[6031]  = ~opsel2 | ~\[8923] ,
  \[5682]  = ~\[5681]  | \[5671] ,
  \[12811]  = ~\[5663]  & \[5653] ,
  \[737]  = (~\[6094]  & ~\[10396] ) | (~\[6094]  & ~\[9661] ),
  \[10158]  = (\[8586]  & ~sh2) | (\[8491]  & sh2),
  \[5874]  = ~\[9481]  | (musel3 | ~musel4),
  \[359]  = (~musel2 & ~inA2) | ((musel2 & ~inC2) | (~inC2 & ~inA2)),
  \[4706]  = musel2 & inC4,
  \[5875]  = (~\[5874]  & \[5849] ) | ~\[11382] ,
  \[9670]  = ~\[10316]  | ~\[9677] ,
  \[6036]  = ~musel3 | musel4,
  \[9481]  = (~\[5871]  & ~musel1) | ~\[11388] ,
  \[5877]  = ~inC5 | ~musel2,
  \[8313]  = (~\[5975]  & ~\[282] ) | ~\[11146] ,
  \[9861]  = ~\[5681]  | \[5671] ,
  \[10154]  = (\[8540]  & ~sh2) | (\[8388]  & sh2),
  \[6037]  = opsel0 | opsel1,
  \[6038]  = (~\[5704]  & ~\[5694] ) | (\[5704]  & \[5694] ),
  \[10156]  = (\[8562]  & ~sh2) | (\[8464]  & sh2),
  \[6039]  = (~\[5843]  & ~\[5840] ) | \[5837] ,
  \[10536]  = ~\[2355]  | (musel3 | (~musel4 | ~inD4)),
  \[9674]  = ~\[5835]  | \[5825] ,
  \[10726]  = ~\[6044]  | ~\[5870] ,
  \[9864]  = \[5681]  | ~\[5671] ,
  \[360]  = (~inA2 & ~\[4540] ) | ((~inA2 & ~musel1) | ((~\[9539]  & ~\[4540] ) | (~\[9539]  & ~musel1))),
  \[9677]  = \[5835]  | ~\[5825] ,
  \[362]  = (~inB2 & ~\[2062] ) | ((~inB2 & ~musel1) | ((~\[9543]  & ~\[2062] ) | (~\[9543]  & ~musel1))),
  \[9867]  = ~\[5663]  | \[5653] ,
  \[10352]  = ~sh2 | ~\[8562] ,
  \[173]  = (~\[1235]  & ~\[9117] ) | (~\[1235]  & ~\[5536] ),
  \[10922]  = ~\[3079]  | (musel3 | (~musel4 | ~inD9)),
  \[2814]  = musel2 & inD7,
  \[5880]  = ~\[9497]  | (musel3 | ~musel4),
  \[555]  = (~\[5976]  & ~\[8313] ) | ((\[5976]  & ~\[8181] ) | (~\[8313]  & ~\[8181] )),
  \[5881]  = (~\[5880]  & \[5849] ) | ~\[11374] ,
  \[556]  = (~\[5978]  & ~\[10029] ) | (~\[5978]  & sh0),
  \[177]  = (~opsel0 & ~opsel1) | (opsel0 & opsel1),
  \[5882]  = ~inC4 | ~musel2,
  \[367]  = (~musel2 & ~inA1) | ((musel2 & ~inC1) | (~inC1 & ~inA1)),
  \[2817]  = ~musel1 & ~musel2,
  \[178]  = (~\[1200]  & \[179] ) | (~\[1200]  & ~\[5951] ),
  \[368]  = (~inA1 & ~\[4466] ) | ((~inA1 & ~musel1) | ((~\[9555]  & ~\[4466] ) | (~\[9555]  & ~musel1))),
  \[10168]  = (\[8586]  & ~sh2) | (\[8491]  & sh2),
  \[5694]  = (~\[1490]  & ~\[1489] ) | musel4,
  \[179]  = (~\[8905]  & ~\[8950] ) | ((~\[8905]  & ~opsel2) | (~\[8950]  & opsel2)),
  \[6044]  = ~\[12790]  | (~\[5886]  | (~\[5881]  | ~\[5875] )),
  \[5695]  = ~inC7 | ~musel4,
  \[5885]  = ~\[9513]  | (musel3 | ~musel4),
  \[6045]  = ~opsel2 | ~\[8926] ,
  \[4338]  = \[5835]  & ~\[5825] ,
  \[5886]  = (~\[5885]  & \[5849] ) | ~\[11366] ,
  \[9870]  = \[5663]  | ~\[5653] ,
  \[9491]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[10164]  = (\[8540]  & ~sh2) | ~\[10204] ,
  \[5888]  = ~\[5886]  | (~\[5881]  | (~\[5875]  | ~\[5870] )),
  \[5889]  = ~inC11 | ~musel2,
  \[10166]  = (\[8562]  & ~sh2) | (\[8418]  & sh2),
  \[9495]  = (~musel1 & musel2) | (musel1 & ~musel2),
  \[370]  = (~inB1 & ~\[1910] ) | ((~inB1 & ~musel1) | ((~\[9559]  & ~\[1910] ) | (~\[9559]  & ~musel1))),
  \[10170]  = (\[8611]  & ~sh2) | (\[8520]  & sh2),
  \[9876]  = (~\[5994]  & ~\[503] ) | ~\[9883] ,
  \[561]  = (~\[1107]  & ~sh2) | (~\[1107]  & ~\[8335] ),
  \[751]  = ~\[6087]  & ~\[6081] ,
  \[2062]  = musel2 & inD2,
  \[9497]  = (~\[5877]  & ~musel1) | ~\[11380] ,
  \[182]  = (~opsel0 & ~opsel1) | (opsel0 & opsel1),
  \[562]  = (~\[1105]  & ~\[8335] ) | (~\[1105]  & sh1),
  \[10172]  = ~\[9314]  | (opsel2 | ~opsel3),
  \[183]  = (~\[1167]  & \[184] ) | (~\[1167]  & ~\[5966] ),
  \[563]  = (~\[10048]  & ~\[10044] ) | ((~\[10048]  & ~sh1) | (~\[10044]  & sh1)),
  \[184]  = (~\[8908]  & ~\[8953] ) | ((~\[8908]  & ~opsel2) | (~\[8953]  & opsel2)),
  \[564]  = (~\[10050]  & ~\[10046] ) | ((~\[10050]  & ~sh1) | (~\[10046]  & sh1)),
  \[2065]  = ~musel1 & ~musel2,
  \[375]  = (~musel2 & ~inA0) | ((musel2 & ~inC0) | (~inC0 & ~inA0)),
  \[6050]  = ~musel3 | musel4,
  \[376]  = (~inA0 & ~\[4392] ) | ((~inA0 & ~musel1) | ((~\[9571]  & ~\[4392] ) | (~\[9571]  & ~musel1))),
  \[6051]  = opsel0 | opsel1,
  \[187]  = (~opsel0 & ~opsel1) | (opsel0 & opsel1),
  \[5892]  = ~\[9401]  | (musel3 | ~musel4),
  \[6052]  = (~\[5722]  & ~\[5712] ) | (\[5722]  & \[5712] ),
  \[188]  = (~\[1136]  & \[189] ) | (~\[1136]  & ~\[5979] );
endmodule

