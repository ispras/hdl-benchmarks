//NOTE: no-implementation module stub

module EU (
    input DSPCLK,
    input T_RST,
    input GO_Ex,
    input GO_Cx,
    input EX_en,
    input EX_enc,
    input cdAM_E,
    input DIVQ_E,
    input DIVS_E,
    input Double_E,
    input MTAR_E,
    input MTAX0_E,
    input MTAX1_E,
    input MTAY0_E,
    input MTAY1_E,
    input Rbyp_Rg,
    input MFAR_E,
    input MFAX0_E,
    input MFAX1_E,
    input MFAY0_E,
    input MFAY1_E,
    input MFASTAT_E,
    input MTMX0_Eg,
    input MTMX1_Eg,
    input MTMY0_Eg,
    input MTMY1_Eg,
    input MTMR0_Eg,
    input MTMR1_Eg,
    input MTMR2_Eg,
    input MFMX0_E,
    input MFMX1_E,
    input MFMY0_E,
    input MFMY1_E,
    input MFMR0_E,
    input MFMR1_E,
    input MFMR2_E,
    input Ybyp_Rg,
    input MTASTAT_E,
    input MTSI_E,
    input MTSB_E,
    input MTSE_E,
    input MTSR0_E,
    input MTSR1_E,
    input MFSI_E,
    input MFSB_E,
    input MFSE_E,
    input MFSR1_E,
    input MFSR0_E,
    input imSHT_E,
    input Xbyp_Rg,
    input MFALU_E,
    input MFMAC_E,
    input MFSHT_E,
    input pMFALU_E,
    input pMFMAC_E,
    input pMFSHT_E,
    input accPM_E,
    input Squ_Rx,
    input GO_MAC,
    input updSR0_Eg,
    input updSR1_Eg,
    input SHTop_E,
    input satMR_Eg,
    input MACop_E,
    input updMF_E,
    input updMR_E,
    input ALUop_E,
    input updAR_E,
    input updAF_E,
    input ALUop_R,
    input type9,
    input updSR_E,
    input MACop_R,
    input DIVQ_R,
    input DIVS_R,
    input [17:0] IR,
    input [14:0] IRE,
    input [3:0] Term,
    input MSTAT,
    input CE,
    input VpopST_Eg,
    input [7:0] popASTATo,
    input RSTtext_h,
    input BIASRND,
    `ifdef FD_DFT
    input SCAN_TEST,
    `endif
    input [7:0] ASTAT,
    input Ctrue,
    input Ttrue,
    input [15:0] DMDid,
    output [15:0] euDMD_do,
    input [15:0] PMDin,
    output [15:0] euPMD_do
);

endmodule
