//NOTE: no-implementation module stub

module MREG16MC (
    input wire DSPCLK,
    input wire MMR_web,
    input wire SYSR_we,
    input wire [15:0] DMD,
    output reg [15:0] SYSR,
    input wire RST
);

endmodule
