//NOTE: no-implementation module stub

module REG12L (
    input wire DSPCLK,
    input wire CLKEMCOREenb,
    input wire GO_E,
    input wire [11:0] EMCOREdi,
    output reg [11:0] EMCOREdo
);

endmodule
