module logical_and_2_1(a, b, c);
  input [1:0] a;
  input b;
  output c;
  assign c = a && b;
endmodule
