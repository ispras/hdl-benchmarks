// IWLS benchmark module "MultiplierB_32" printed on Wed May 29 22:12:35 2002
module MultiplierB_32(\1 , \3 , \4 , \5 , \6 , \7 , \8 , \9 , \10 , \11 , \12 , \13 , \14 , \15 , \16 , \17 , \18 , \19 , \20 , \21 , \22 , \23 , \24 , \25 , \26 , \27 , \28 , \29 , \30 , \31 , \32 , \33 , \98 );
input
  \1 ,
  \3 ,
  \4 ,
  \5 ,
  \6 ,
  \7 ,
  \8 ,
  \9 ,
  \10 ,
  \11 ,
  \12 ,
  \13 ,
  \14 ,
  \15 ,
  \16 ,
  \17 ,
  \18 ,
  \19 ,
  \20 ,
  \21 ,
  \22 ,
  \23 ,
  \24 ,
  \25 ,
  \26 ,
  \27 ,
  \28 ,
  \29 ,
  \30 ,
  \31 ,
  \32 ,
  \33 ;
output
  \98 ;
reg
  \2 ,
  \34 ,
  \36 ,
  \37 ,
  \38 ,
  \39 ,
  \40 ,
  \41 ,
  \42 ,
  \43 ,
  \44 ,
  \45 ,
  \46 ,
  \47 ,
  \48 ,
  \49 ,
  \50 ,
  \51 ,
  \52 ,
  \53 ,
  \54 ,
  \55 ,
  \56 ,
  \57 ,
  \58 ,
  \59 ,
  \60 ,
  \61 ,
  \62 ,
  \63 ,
  \64 ,
  \65 ,
  \66 ,
  \67 ,
  \68 ,
  \69 ,
  \70 ,
  \71 ,
  \72 ,
  \73 ,
  \74 ,
  \75 ,
  \76 ,
  \77 ,
  \78 ,
  \79 ,
  \80 ,
  \81 ,
  \82 ,
  \83 ,
  \84 ,
  \85 ,
  \86 ,
  \87 ,
  \88 ,
  \89 ,
  \90 ,
  \91 ,
  \92 ,
  \93 ,
  \94 ,
  \95 ;
wire
  \[77] ,
  \[78] ,
  \[79] ,
  \[80] ,
  \[81] ,
  \[82] ,
  \[83] ,
  \[84] ,
  \[85] ,
  \[86] ,
  \[87] ,
  \[88] ,
  \[89] ,
  \[90] ,
  \[91] ,
  \[92] ,
  \[93] ,
  \[94] ,
  \[95] ,
  \[96] ,
  \[97] ,
  \[100] ,
  \[98] ,
  \[101] ,
  \[99] ,
  \[102] ,
  \[103] ,
  \[104] ,
  \[105] ,
  \[106] ,
  \[107] ,
  \[108] ,
  \[109] ,
  \[110] ,
  \[111] ,
  \[112] ,
  \[113] ,
  \[114] ,
  \[115] ,
  \[116] ,
  \[117] ,
  \[118] ,
  \[119] ,
  \96 ,
  \97 ,
  \[120] ,
  \[121] ,
  \[122] ,
  \[123] ,
  \[124] ,
  \160 ,
  \161 ,
  \162 ,
  \163 ,
  \164 ,
  \165 ,
  \166 ,
  \167 ,
  \168 ,
  \169 ,
  \170 ,
  \171 ,
  \172 ,
  \173 ,
  \174 ,
  \175 ,
  \176 ,
  \177 ,
  \178 ,
  \179 ,
  \180 ,
  \181 ,
  \182 ,
  \183 ,
  \184 ,
  \185 ,
  \186 ,
  \187 ,
  \188 ,
  \189 ,
  \190 ,
  \191 ,
  \192 ,
  \193 ,
  \194 ,
  \195 ,
  \196 ,
  \197 ,
  \198 ,
  \199 ,
  \200 ,
  \201 ,
  \202 ,
  \203 ,
  \204 ,
  \205 ,
  \206 ,
  \207 ,
  \208 ,
  \209 ,
  \210 ,
  \211 ,
  \212 ,
  \213 ,
  \214 ,
  \215 ,
  \216 ,
  \217 ,
  \218 ,
  \219 ,
  \220 ,
  \221 ,
  \222 ,
  \223 ,
  \224 ,
  \225 ,
  \226 ,
  \227 ,
  \228 ,
  \229 ,
  \230 ,
  \231 ,
  \232 ,
  \233 ,
  \234 ,
  \235 ,
  \236 ,
  \237 ,
  \238 ,
  \239 ,
  \240 ,
  \241 ,
  \242 ,
  \243 ,
  \244 ,
  \245 ,
  \246 ,
  \247 ,
  \248 ,
  \249 ,
  \250 ,
  \251 ,
  \252 ,
  \253 ,
  \254 ,
  \255 ,
  \256 ,
  \257 ,
  \258 ,
  \259 ,
  \260 ,
  \261 ,
  \262 ,
  \263 ,
  \264 ,
  \265 ,
  \266 ,
  \267 ,
  \268 ,
  \269 ,
  \270 ,
  \271 ,
  \272 ,
  \273 ,
  \274 ,
  \275 ,
  \276 ,
  \277 ,
  \278 ,
  \279 ,
  \280 ,
  \281 ,
  \282 ,
  \283 ,
  \284 ,
  \285 ,
  \286 ,
  \287 ,
  \288 ,
  \289 ,
  \290 ,
  \291 ,
  \292 ,
  \293 ,
  \294 ,
  \295 ,
  \296 ,
  \297 ,
  \298 ,
  \299 ,
  \300 ,
  \301 ,
  \302 ,
  \303 ,
  \304 ,
  \305 ,
  \306 ,
  \307 ,
  \308 ,
  \309 ,
  \310 ,
  \311 ,
  \312 ,
  \313 ,
  \314 ,
  \315 ,
  \316 ,
  \317 ,
  \318 ,
  \319 ,
  \320 ,
  \321 ,
  \322 ,
  \323 ,
  \324 ,
  \325 ,
  \326 ,
  \327 ,
  \328 ,
  \329 ,
  \330 ,
  \331 ,
  \332 ,
  \333 ,
  \334 ,
  \335 ,
  \336 ,
  \337 ,
  \338 ,
  \339 ,
  \340 ,
  \341 ,
  \342 ,
  \343 ,
  \344 ,
  \345 ,
  \346 ,
  \347 ,
  \348 ,
  \349 ,
  \350 ,
  \351 ,
  \352 ,
  \353 ,
  \354 ,
  \355 ,
  \356 ,
  \357 ,
  \358 ,
  \359 ,
  \360 ,
  \361 ,
  \362 ,
  \363 ,
  \364 ,
  \365 ,
  \366 ,
  \367 ,
  \368 ,
  \369 ,
  \370 ,
  \371 ,
  \372 ,
  \373 ,
  \374 ,
  \375 ,
  \376 ,
  \377 ,
  \378 ,
  \379 ,
  \380 ,
  \381 ,
  \382 ,
  \383 ,
  \384 ,
  \385 ,
  \386 ,
  \387 ,
  \388 ,
  \389 ,
  \390 ,
  \391 ,
  \392 ,
  \393 ,
  \394 ,
  \395 ,
  \396 ,
  \397 ,
  \398 ,
  \399 ,
  \400 ,
  \401 ,
  \402 ,
  \403 ,
  \404 ,
  \405 ,
  \406 ,
  \407 ,
  \408 ,
  \409 ,
  \410 ,
  \411 ,
  \412 ,
  \413 ,
  \414 ,
  \415 ,
  \416 ,
  \417 ,
  \418 ,
  \419 ,
  \420 ,
  \421 ,
  \422 ,
  \423 ,
  \424 ,
  \425 ,
  \426 ,
  \427 ,
  \428 ,
  \429 ,
  \430 ,
  \431 ,
  \432 ,
  \433 ,
  \434 ,
  \435 ,
  \436 ,
  \437 ,
  \438 ,
  \439 ,
  \440 ,
  \441 ,
  \442 ,
  \443 ,
  \444 ,
  \445 ,
  \446 ,
  \447 ,
  \448 ,
  \449 ,
  \450 ,
  \451 ,
  \452 ,
  \453 ,
  \454 ,
  \455 ,
  \456 ,
  \457 ,
  \458 ,
  \459 ,
  \460 ,
  \461 ,
  \462 ,
  \463 ,
  \464 ,
  \465 ,
  \466 ,
  \467 ,
  \468 ,
  \469 ,
  \470 ,
  \471 ,
  \472 ,
  \473 ,
  \474 ,
  \475 ,
  \476 ,
  \477 ,
  \478 ,
  \479 ,
  \480 ,
  \481 ,
  \482 ,
  \483 ,
  \484 ,
  \485 ,
  \486 ,
  \487 ,
  \488 ,
  \489 ,
  \490 ,
  \491 ,
  \492 ,
  \493 ,
  \494 ,
  \495 ,
  \496 ,
  \497 ,
  \498 ,
  \499 ,
  \500 ,
  \501 ,
  \502 ,
  \503 ,
  \504 ,
  \505 ,
  \506 ,
  \507 ,
  \508 ,
  \509 ,
  \510 ,
  \511 ,
  \512 ,
  \513 ,
  \514 ,
  \515 ,
  \516 ,
  \517 ,
  \518 ,
  \519 ,
  \520 ,
  \521 ,
  \522 ,
  \523 ,
  \524 ,
  \525 ,
  \526 ,
  \527 ,
  \528 ,
  \529 ,
  \530 ,
  \531 ,
  \532 ,
  \533 ,
  \534 ,
  \535 ,
  \536 ,
  \537 ,
  \538 ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[66] ,
  \[67] ,
  \[68] ,
  \[69] ,
  \[70] ,
  \[71] ,
  \[72] ,
  \[73] ,
  \[74] ,
  \[75] ,
  \[76] ;
assign
  \[77]  = \296 ,
  \[78]  = \301 ,
  \[79]  = \306 ,
  \[80]  = \311 ,
  \[81]  = \316 ,
  \[82]  = \321 ,
  \[83]  = \326 ,
  \[84]  = \331 ,
  \[85]  = \336 ,
  \[86]  = \341 ,
  \[87]  = \346 ,
  \[88]  = \351 ,
  \[89]  = \356 ,
  \[90]  = \361 ,
  \[91]  = \366 ,
  \[92]  = \371 ,
  \[93]  = \376 ,
  \[94]  = \230 ,
  \[95]  = \235 ,
  \[96]  = \240 ,
  \[97]  = \245 ,
  \[100]  = \260 ,
  \[98]  = \250 ,
  \[101]  = \265 ,
  \[99]  = \255 ,
  \[102]  = \270 ,
  \[103]  = \275 ,
  \[104]  = \280 ,
  \[105]  = \285 ,
  \[106]  = \290 ,
  \[107]  = \295 ,
  \[108]  = \300 ,
  \[109]  = \305 ,
  \[110]  = \310 ,
  \[111]  = \315 ,
  \[112]  = \320 ,
  \[113]  = \325 ,
  \[114]  = \330 ,
  \[115]  = \335 ,
  \[116]  = \340 ,
  \[117]  = \345 ,
  \[118]  = \350 ,
  \[119]  = \355 ,
  \96  = 0,
  \97  = \476  | \475 ,
  \98  = \226 ,
  \[120]  = \360 ,
  \[121]  = \365 ,
  \[122]  = \370 ,
  \[123]  = \375 ,
  \[124]  = \380 ,
  \160  = ~\161 ,
  \161  = (~\381  & ~\1 ) | (\381  & \1 ),
  \162  = \3 ,
  \163  = \4 ,
  \164  = \5 ,
  \165  = \6 ,
  \166  = \7 ,
  \167  = \8 ,
  \168  = \9 ,
  \169  = \10 ,
  \170  = \11 ,
  \171  = \12 ,
  \172  = \13 ,
  \173  = \14 ,
  \174  = \15 ,
  \175  = \16 ,
  \176  = \17 ,
  \177  = \18 ,
  \178  = \19 ,
  \179  = \20 ,
  \180  = \21 ,
  \181  = \22 ,
  \182  = \23 ,
  \183  = \24 ,
  \184  = \25 ,
  \185  = \26 ,
  \186  = \27 ,
  \187  = \28 ,
  \188  = \29 ,
  \189  = \30 ,
  \190  = \31 ,
  \191  = \32 ,
  \192  = \33 ,
  \193  = 0,
  \194  = 0,
  \195  = 0,
  \196  = 0,
  \197  = 0,
  \198  = 0,
  \199  = 0,
  \200  = 0,
  \201  = 0,
  \202  = 0,
  \203  = 0,
  \204  = 0,
  \205  = 0,
  \206  = 0,
  \207  = 0,
  \208  = 0,
  \209  = 0,
  \210  = 0,
  \211  = 0,
  \212  = 0,
  \213  = 0,
  \214  = 0,
  \215  = 0,
  \216  = 0,
  \217  = 0,
  \218  = 0,
  \219  = 0,
  \220  = 0,
  \221  = 0,
  \222  = 0,
  \223  = 0,
  \224  = \34 ,
  \225  = 0,
  \226  = (~\383  & \382 ) | (\383  & ~\382 ),
  \227  = \382  & \36 ,
  \228  = \382  & \66 ,
  \229  = \36  & \66 ,
  \230  = \384  | \229 ,
  \231  = (~\386  & \385 ) | (\386  & ~\385 ),
  \232  = \385  & \37 ,
  \233  = \385  & \67 ,
  \234  = \37  & \67 ,
  \235  = \387  | \234 ,
  \236  = (~\389  & \388 ) | (\389  & ~\388 ),
  \237  = \388  & \38 ,
  \238  = \388  & \68 ,
  \239  = \38  & \68 ,
  \240  = \390  | \239 ,
  \241  = (~\392  & \391 ) | (\392  & ~\391 ),
  \242  = \391  & \39 ,
  \243  = \391  & \69 ,
  \244  = \39  & \69 ,
  \245  = \393  | \244 ,
  \246  = (~\395  & \394 ) | (\395  & ~\394 ),
  \247  = \394  & \40 ,
  \248  = \394  & \70 ,
  \249  = \40  & \70 ,
  \250  = \396  | \249 ,
  \251  = (~\398  & \397 ) | (\398  & ~\397 ),
  \252  = \397  & \41 ,
  \253  = \397  & \71 ,
  \254  = \41  & \71 ,
  \255  = \399  | \254 ,
  \256  = (~\401  & \400 ) | (\401  & ~\400 ),
  \257  = \400  & \42 ,
  \258  = \400  & \72 ,
  \259  = \42  & \72 ,
  \260  = \402  | \259 ,
  \261  = (~\404  & \403 ) | (\404  & ~\403 ),
  \262  = \403  & \43 ,
  \263  = \403  & \73 ,
  \264  = \43  & \73 ,
  \265  = \405  | \264 ,
  \266  = (~\407  & \406 ) | (\407  & ~\406 ),
  \267  = \406  & \44 ,
  \268  = \406  & \74 ,
  \269  = \44  & \74 ,
  \270  = \408  | \269 ,
  \271  = (~\410  & \409 ) | (\410  & ~\409 ),
  \272  = \409  & \45 ,
  \273  = \409  & \75 ,
  \274  = \45  & \75 ,
  \275  = \411  | \274 ,
  \276  = (~\413  & \412 ) | (\413  & ~\412 ),
  \277  = \412  & \46 ,
  \278  = \412  & \76 ,
  \279  = \46  & \76 ,
  \280  = \414  | \279 ,
  \281  = (~\416  & \415 ) | (\416  & ~\415 ),
  \282  = \415  & \47 ,
  \283  = \415  & \77 ,
  \284  = \47  & \77 ,
  \285  = \417  | \284 ,
  \286  = (~\419  & \418 ) | (\419  & ~\418 ),
  \287  = \418  & \48 ,
  \288  = \418  & \78 ,
  \289  = \48  & \78 ,
  \290  = \420  | \289 ,
  \291  = (~\422  & \421 ) | (\422  & ~\421 ),
  \292  = \421  & \49 ,
  \293  = \421  & \79 ,
  \294  = \49  & \79 ,
  \295  = \423  | \294 ,
  \296  = (~\425  & \424 ) | (\425  & ~\424 ),
  \297  = \424  & \50 ,
  \298  = \424  & \80 ,
  \299  = \50  & \80 ,
  \300  = \426  | \299 ,
  \301  = (~\428  & \427 ) | (\428  & ~\427 ),
  \302  = \427  & \51 ,
  \303  = \427  & \81 ,
  \304  = \51  & \81 ,
  \305  = \429  | \304 ,
  \306  = (~\431  & \430 ) | (\431  & ~\430 ),
  \307  = \430  & \52 ,
  \308  = \430  & \82 ,
  \309  = \52  & \82 ,
  \310  = \432  | \309 ,
  \311  = (~\434  & \433 ) | (\434  & ~\433 ),
  \312  = \433  & \53 ,
  \313  = \433  & \83 ,
  \314  = \53  & \83 ,
  \315  = \435  | \314 ,
  \316  = (~\437  & \436 ) | (\437  & ~\436 ),
  \317  = \436  & \54 ,
  \318  = \436  & \84 ,
  \319  = \54  & \84 ,
  \320  = \438  | \319 ,
  \321  = (~\440  & \439 ) | (\440  & ~\439 ),
  \322  = \439  & \55 ,
  \323  = \439  & \85 ,
  \324  = \55  & \85 ,
  \325  = \441  | \324 ,
  \326  = (~\443  & \442 ) | (\443  & ~\442 ),
  \327  = \442  & \56 ,
  \328  = \442  & \86 ,
  \329  = \56  & \86 ,
  \330  = \444  | \329 ,
  \331  = (~\446  & \445 ) | (\446  & ~\445 ),
  \332  = \445  & \57 ,
  \333  = \445  & \87 ,
  \334  = \57  & \87 ,
  \335  = \447  | \334 ,
  \336  = (~\449  & \448 ) | (\449  & ~\448 ),
  \337  = \448  & \58 ,
  \338  = \448  & \88 ,
  \339  = \58  & \88 ,
  \340  = \450  | \339 ,
  \341  = (~\452  & \451 ) | (\452  & ~\451 ),
  \342  = \451  & \59 ,
  \343  = \451  & \89 ,
  \344  = \59  & \89 ,
  \345  = \453  | \344 ,
  \346  = (~\455  & \454 ) | (\455  & ~\454 ),
  \347  = \454  & \60 ,
  \348  = \454  & \90 ,
  \349  = \60  & \90 ,
  \350  = \456  | \349 ,
  \351  = (~\458  & \457 ) | (\458  & ~\457 ),
  \352  = \457  & \61 ,
  \353  = \457  & \91 ,
  \354  = \61  & \91 ,
  \355  = \459  | \354 ,
  \356  = (~\461  & \460 ) | (\461  & ~\460 ),
  \357  = \460  & \62 ,
  \358  = \460  & \92 ,
  \359  = \62  & \92 ,
  \360  = \462  | \359 ,
  \361  = (~\464  & \463 ) | (\464  & ~\463 ),
  \362  = \463  & \63 ,
  \363  = \463  & \93 ,
  \364  = \63  & \93 ,
  \365  = \465  | \364 ,
  \366  = (~\467  & \466 ) | (\467  & ~\466 ),
  \367  = \466  & \64 ,
  \368  = \466  & \94 ,
  \369  = \64  & \94 ,
  \370  = \468  | \369 ,
  \371  = (~\470  & \469 ) | (\470  & ~\469 ),
  \372  = \469  & \65 ,
  \373  = \469  & \95 ,
  \374  = \65  & \95 ,
  \375  = \471  | \374 ,
  \376  = (~\473  & \472 ) | (\473  & ~\472 ),
  \377  = \472  & \2 ,
  \378  = \472  & \96 ,
  \379  = \2  & \96 ,
  \380  = \474  | \379 ,
  \381  = 0,
  \382  = \538  | \537 ,
  \383  = (~\36  & \66 ) | (\36  & ~\66 ),
  \384  = \228  | \227 ,
  \385  = \536  | \535 ,
  \386  = (~\37  & \67 ) | (\37  & ~\67 ),
  \387  = \233  | \232 ,
  \388  = \534  | \533 ,
  \389  = (~\38  & \68 ) | (\38  & ~\68 ),
  \390  = \238  | \237 ,
  \391  = \532  | \531 ,
  \392  = (~\39  & \69 ) | (\39  & ~\69 ),
  \393  = \243  | \242 ,
  \394  = \530  | \529 ,
  \395  = (~\40  & \70 ) | (\40  & ~\70 ),
  \396  = \248  | \247 ,
  \397  = \528  | \527 ,
  \398  = (~\41  & \71 ) | (\41  & ~\71 ),
  \399  = \253  | \252 ,
  \400  = \526  | \525 ,
  \401  = (~\42  & \72 ) | (\42  & ~\72 ),
  \402  = \258  | \257 ,
  \403  = \524  | \523 ,
  \404  = (~\43  & \73 ) | (\43  & ~\73 ),
  \405  = \263  | \262 ,
  \406  = \522  | \521 ,
  \407  = (~\44  & \74 ) | (\44  & ~\74 ),
  \408  = \268  | \267 ,
  \409  = \520  | \519 ,
  \410  = (~\45  & \75 ) | (\45  & ~\75 ),
  \411  = \273  | \272 ,
  \412  = \518  | \517 ,
  \413  = (~\46  & \76 ) | (\46  & ~\76 ),
  \414  = \278  | \277 ,
  \415  = \516  | \515 ,
  \416  = (~\47  & \77 ) | (\47  & ~\77 ),
  \417  = \283  | \282 ,
  \418  = \514  | \513 ,
  \419  = (~\48  & \78 ) | (\48  & ~\78 ),
  \420  = \288  | \287 ,
  \421  = \512  | \511 ,
  \422  = (~\49  & \79 ) | (\49  & ~\79 ),
  \423  = \293  | \292 ,
  \424  = \510  | \509 ,
  \425  = (~\50  & \80 ) | (\50  & ~\80 ),
  \426  = \298  | \297 ,
  \427  = \508  | \507 ,
  \428  = (~\51  & \81 ) | (\51  & ~\81 ),
  \429  = \303  | \302 ,
  \430  = \506  | \505 ,
  \431  = (~\52  & \82 ) | (\52  & ~\82 ),
  \432  = \308  | \307 ,
  \433  = \504  | \503 ,
  \434  = (~\53  & \83 ) | (\53  & ~\83 ),
  \435  = \313  | \312 ,
  \436  = \502  | \501 ,
  \437  = (~\54  & \84 ) | (\54  & ~\84 ),
  \438  = \318  | \317 ,
  \439  = \500  | \499 ,
  \440  = (~\55  & \85 ) | (\55  & ~\85 ),
  \441  = \323  | \322 ,
  \442  = \498  | \497 ,
  \443  = (~\56  & \86 ) | (\56  & ~\86 ),
  \444  = \328  | \327 ,
  \445  = \496  | \495 ,
  \446  = (~\57  & \87 ) | (\57  & ~\87 ),
  \447  = \333  | \332 ,
  \448  = \494  | \493 ,
  \449  = (~\58  & \88 ) | (\58  & ~\88 ),
  \450  = \338  | \337 ,
  \451  = \492  | \491 ,
  \452  = (~\59  & \89 ) | (\59  & ~\89 ),
  \453  = \343  | \342 ,
  \454  = \490  | \489 ,
  \455  = (~\60  & \90 ) | (\60  & ~\90 ),
  \456  = \348  | \347 ,
  \457  = \488  | \487 ,
  \458  = (~\61  & \91 ) | (\61  & ~\91 ),
  \459  = \353  | \352 ,
  \460  = \486  | \485 ,
  \461  = (~\62  & \92 ) | (\62  & ~\92 ),
  \462  = \358  | \357 ,
  \463  = \484  | \483 ,
  \464  = (~\63  & \93 ) | (\63  & ~\93 ),
  \465  = \363  | \362 ,
  \466  = \482  | \481 ,
  \467  = (~\64  & \94 ) | (\64  & ~\94 ),
  \468  = \368  | \367 ,
  \469  = \480  | \479 ,
  \470  = (~\65  & \95 ) | (\65  & ~\95 ),
  \471  = \373  | \372 ,
  \472  = \478  | \477 ,
  \473  = (~\2  & \96 ) | (\2  & ~\96 ),
  \474  = \378  | \377 ,
  \475  = \224  & \160 ,
  \476  = \225  & \161 ,
  \477  = \192  & \160 ,
  \478  = \223  & \161 ,
  \479  = \191  & \160 ,
  \480  = \222  & \161 ,
  \481  = \190  & \160 ,
  \482  = \221  & \161 ,
  \483  = \189  & \160 ,
  \484  = \220  & \161 ,
  \485  = \188  & \160 ,
  \486  = \219  & \161 ,
  \487  = \187  & \160 ,
  \488  = \218  & \161 ,
  \489  = \186  & \160 ,
  \490  = \217  & \161 ,
  \491  = \185  & \160 ,
  \492  = \216  & \161 ,
  \493  = \184  & \160 ,
  \494  = \215  & \161 ,
  \495  = \183  & \160 ,
  \496  = \214  & \161 ,
  \497  = \182  & \160 ,
  \498  = \213  & \161 ,
  \499  = \181  & \160 ,
  \500  = \212  & \161 ,
  \501  = \180  & \160 ,
  \502  = \211  & \161 ,
  \503  = \179  & \160 ,
  \504  = \210  & \161 ,
  \505  = \178  & \160 ,
  \506  = \209  & \161 ,
  \507  = \177  & \160 ,
  \508  = \208  & \161 ,
  \509  = \176  & \160 ,
  \510  = \207  & \161 ,
  \511  = \175  & \160 ,
  \512  = \206  & \161 ,
  \513  = \174  & \160 ,
  \514  = \205  & \161 ,
  \515  = \173  & \160 ,
  \516  = \204  & \161 ,
  \517  = \172  & \160 ,
  \518  = \203  & \161 ,
  \519  = \171  & \160 ,
  \520  = \202  & \161 ,
  \521  = \170  & \160 ,
  \522  = \201  & \161 ,
  \523  = \169  & \160 ,
  \524  = \200  & \161 ,
  \525  = \168  & \160 ,
  \526  = \199  & \161 ,
  \527  = \167  & \160 ,
  \528  = \198  & \161 ,
  \529  = \166  & \160 ,
  \530  = \197  & \161 ,
  \531  = \165  & \160 ,
  \532  = \196  & \161 ,
  \533  = \164  & \160 ,
  \534  = \195  & \161 ,
  \535  = \163  & \160 ,
  \536  = \194  & \161 ,
  \537  = \162  & \160 ,
  \538  = \193  & \161 ,
  \[63]  = \97 ,
  \[64]  = \231 ,
  \[65]  = \236 ,
  \[66]  = \241 ,
  \[67]  = \246 ,
  \[68]  = \251 ,
  \[69]  = \256 ,
  \[70]  = \261 ,
  \[71]  = \266 ,
  \[72]  = \271 ,
  \[73]  = \276 ,
  \[74]  = \281 ,
  \[75]  = \286 ,
  \[76]  = \291 ;
always begin
  \2  = \[64] ;
  \34  = \[63] ;
  \36  = \[65] ;
  \37  = \[66] ;
  \38  = \[67] ;
  \39  = \[68] ;
  \40  = \[69] ;
  \41  = \[70] ;
  \42  = \[71] ;
  \43  = \[72] ;
  \44  = \[73] ;
  \45  = \[74] ;
  \46  = \[75] ;
  \47  = \[76] ;
  \48  = \[77] ;
  \49  = \[78] ;
  \50  = \[79] ;
  \51  = \[80] ;
  \52  = \[81] ;
  \53  = \[82] ;
  \54  = \[83] ;
  \55  = \[84] ;
  \56  = \[85] ;
  \57  = \[86] ;
  \58  = \[87] ;
  \59  = \[88] ;
  \60  = \[89] ;
  \61  = \[90] ;
  \62  = \[91] ;
  \63  = \[92] ;
  \64  = \[93] ;
  \65  = \[94] ;
  \66  = \[95] ;
  \67  = \[96] ;
  \68  = \[97] ;
  \69  = \[98] ;
  \70  = \[99] ;
  \71  = \[100] ;
  \72  = \[101] ;
  \73  = \[102] ;
  \74  = \[103] ;
  \75  = \[104] ;
  \76  = \[105] ;
  \77  = \[106] ;
  \78  = \[107] ;
  \79  = \[108] ;
  \80  = \[109] ;
  \81  = \[110] ;
  \82  = \[111] ;
  \83  = \[112] ;
  \84  = \[113] ;
  \85  = \[114] ;
  \86  = \[115] ;
  \87  = \[116] ;
  \88  = \[117] ;
  \89  = \[118] ;
  \90  = \[119] ;
  \91  = \[120] ;
  \92  = \[121] ;
  \93  = \[122] ;
  \94  = \[123] ;
  \95  = \[124] ;
end
initial begin
  \2  = 0;
  \34  = 0;
  \36  = 0;
  \37  = 0;
  \38  = 0;
  \39  = 0;
  \40  = 0;
  \41  = 0;
  \42  = 0;
  \43  = 0;
  \44  = 0;
  \45  = 0;
  \46  = 0;
  \47  = 0;
  \48  = 0;
  \49  = 0;
  \50  = 0;
  \51  = 0;
  \52  = 0;
  \53  = 0;
  \54  = 0;
  \55  = 0;
  \56  = 0;
  \57  = 0;
  \58  = 0;
  \59  = 0;
  \60  = 0;
  \61  = 0;
  \62  = 0;
  \63  = 0;
  \64  = 0;
  \65  = 0;
  \66  = 0;
  \67  = 0;
  \68  = 0;
  \69  = 0;
  \70  = 0;
  \71  = 0;
  \72  = 0;
  \73  = 0;
  \74  = 0;
  \75  = 0;
  \76  = 0;
  \77  = 0;
  \78  = 0;
  \79  = 0;
  \80  = 0;
  \81  = 0;
  \82  = 0;
  \83  = 0;
  \84  = 0;
  \85  = 0;
  \86  = 0;
  \87  = 0;
  \88  = 0;
  \89  = 0;
  \90  = 0;
  \91  = 0;
  \92  = 0;
  \93  = 0;
  \94  = 0;
  \95  = 0;
end
endmodule

