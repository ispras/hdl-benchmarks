module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 , g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 , g539 , g540 , g541 , g542 , g543 , g544 , g545 , g546 , g547 , g548 , g549 , g550 , g551 , g552 , g553 , g554 , g555 , g556 , g557 , g558 , g559 , g560 , g561 , g562 , g563 , g564 , g565 , g566 , g567 , g568 , g569 , g570 , g571 , g572 , g573 , g574 , g575 , g576 , g577 , g578 , g579 , g580 , g581 , g582 , g583 , g584 , g585 , g586 , g587 , g588 , g589 , g590 , g591 , g592 , g593 , g594 , g595 , g596 , g597 , g598 , g599 , g600 , g601 , g602 , g603 , g604 , g605 , g606 , g607 , g608 , g609 , g610 , g611 , g612 , g613 , g614 , g615 , g616 , g617 , g618 , g619 , g620 , g621 , g622 , g623 , g624 , g625 , g626 , g627 , g628 , g629 , g630 , g631 , g632 , g633 , g634 , g635 , g636 , g637 , g638 , g639 , g640 , g641 , g642 , g643 , g644 , g645 , g646 , g647 , g648 , g649 , g650 , g651 , g652 , g653 , g654 , g655 , g656 , g657 , g658 , g659 , g660 , g661 , g662 , g663 , g664 , g665 , g666 , g667 , g668 , g669 , g670 , g671 , g672 , g673 , g674 , g675 , g676 , g677 , g678 , g679 , g680 , g681 , g682 , g683 , g684 , g685 , g686 , g687 , g688 , g689 , g690 , g691 , g692 , g693 , g694 , g695 , g696 , g697 , g698 , g699 , g700 , g701 , g702 , g703 , g704 , g705 , g706 , g707 , g708 , g709 , g710 , g711 , g712 , g713 , g714 , g715 , g716 , g717 , g718 , g719 , g720 , g721 , g722 , g723 , g724 , g725 , g726 , g727 , g728 , g729 , g730 , g731 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 , g231 , g232 , g233 , g234 , g235 , g236 , g237 , g238 , g239 , g240 , g241 , g242 , g243 , g244 , g245 , g246 , g247 , g248 , g249 , g250 , g251 , g252 , g253 , g254 , g255 , g256 , g257 , g258 , g259 , g260 , g261 , g262 , g263 , g264 , g265 , g266 , g267 , g268 , g269 , g270 , g271 , g272 , g273 , g274 , g275 , g276 , g277 , g278 , g279 , g280 , g281 , g282 , g283 , g284 , g285 , g286 , g287 , g288 , g289 , g290 , g291 , g292 , g293 , g294 , g295 , g296 , g297 , g298 , g299 , g300 , g301 , g302 , g303 , g304 , g305 , g306 , g307 , g308 , g309 , g310 , g311 , g312 , g313 , g314 , g315 , g316 , g317 , g318 , g319 , g320 , g321 , g322 , g323 , g324 , g325 , g326 , g327 , g328 , g329 , g330 , g331 , g332 , g333 , g334 , g335 , g336 , g337 , g338 , g339 , g340 , g341 , g342 , g343 , g344 , g345 , g346 , g347 , g348 , g349 , g350 , g351 , g352 , g353 , g354 , g355 , g356 , g357 , g358 , g359 , g360 , g361 , g362 , g363 , g364 , g365 , g366 , g367 , g368 , g369 , g370 , g371 , g372 , g373 , g374 , g375 , g376 , g377 , g378 , g379 , g380 , g381 , g382 , g383 , g384 , g385 , g386 , g387 , g388 , g389 , g390 , g391 , g392 , g393 , g394 , g395 , g396 , g397 , g398 , g399 , g400 , g401 , g402 , g403 , g404 , g405 , g406 , g407 , g408 , g409 , g410 , g411 , g412 , g413 , g414 , g415 , g416 , g417 , g418 , g419 , g420 , g421 , g422 , g423 , g424 , g425 , g426 , g427 , g428 , g429 , g430 , g431 , g432 , g433 , g434 , g435 , g436 , g437 , g438 , g439 , g440 , g441 , g442 , g443 , g444 , g445 , g446 , g447 , g448 , g449 ;
output g450 , g451 , g452 , g453 , g454 , g455 , g456 , g457 , g458 , g459 , g460 , g461 , g462 , g463 , g464 , g465 , g466 , g467 , g468 , g469 , g470 , g471 , g472 , g473 , g474 , g475 , g476 , g477 , g478 , g479 , g480 , g481 , g482 , g483 , g484 , g485 , g486 , g487 , g488 , g489 , g490 , g491 , g492 , g493 , g494 , g495 , g496 , g497 , g498 , g499 , g500 , g501 , g502 , g503 , g504 , g505 , g506 , g507 , g508 , g509 , g510 , g511 , g512 , g513 , g514 , g515 , g516 , g517 , g518 , g519 , g520 , g521 , g522 , g523 , g524 , g525 , g526 , g527 , g528 , g529 , g530 , g531 , g532 , g533 , g534 , g535 , g536 , g537 , g538 , g539 , g540 , g541 , g542 , g543 , g544 , g545 , g546 , g547 , g548 , g549 , g550 , g551 , g552 , g553 , g554 , g555 , g556 , g557 , g558 , g559 , g560 , g561 , g562 , g563 , g564 , g565 , g566 , g567 , g568 , g569 , g570 , g571 , g572 , g573 , g574 , g575 , g576 , g577 , g578 , g579 , g580 , g581 , g582 , g583 , g584 , g585 , g586 , g587 , g588 , g589 , g590 , g591 , g592 , g593 , g594 , g595 , g596 , g597 , g598 , g599 , g600 , g601 , g602 , g603 , g604 , g605 , g606 , g607 , g608 , g609 , g610 , g611 , g612 , g613 , g614 , g615 , g616 , g617 , g618 , g619 , g620 , g621 , g622 , g623 , g624 , g625 , g626 , g627 , g628 , g629 , g630 , g631 , g632 , g633 , g634 , g635 , g636 , g637 , g638 , g639 , g640 , g641 , g642 , g643 , g644 , g645 , g646 , g647 , g648 , g649 , g650 , g651 , g652 , g653 , g654 , g655 , g656 , g657 , g658 , g659 , g660 , g661 , g662 , g663 , g664 , g665 , g666 , g667 , g668 , g669 , g670 , g671 , g672 , g673 , g674 , g675 , g676 , g677 , g678 , g679 , g680 , g681 , g682 , g683 , g684 , g685 , g686 , g687 , g688 , g689 , g690 , g691 , g692 , g693 , g694 , g695 , g696 , g697 , g698 , g699 , g700 , g701 , g702 , g703 , g704 , g705 , g706 , g707 , g708 , g709 , g710 , g711 , g712 , g713 , g714 , g715 , g716 , g717 , g718 , g719 , g720 , g721 , g722 , g723 , g724 , g725 , g726 , g727 , g728 , g729 , g730 , g731 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , 
     n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , 
     n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , 
     n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , 
     n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , 
     n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , 
     n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , 
     n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , 
     n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , 
     n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , 
     n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , 
     n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , 
     n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , 
     n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , 
     n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , 
     n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , 
     n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , 
     n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , 
     n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , 
     n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , 
     n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , 
     n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , 
     n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , 
     n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , 
     n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , 
     n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , 
     n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , 
     n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , 
     n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , 
     n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , 
     n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , 
     n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , 
     n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , 
     n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , 
     n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , 
     n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , 
     n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , 
     n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , 
     n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , 
     n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , 
     n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , 
     n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , 
     n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , 
     n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , 
     n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , 
     n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , 
     n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , 
     n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , 
     n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , 
     n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , 
     n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , 
     n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , 
     n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , 
     n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , 
     n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , 
     n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , 
     n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , 
     n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , 
     n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , 
     n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , 
     n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , 
     n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , 
     n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , 
     n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , 
     n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , 
     n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , 
     n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , 
     n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , 
     n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , 
     n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , 
     n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , 
     n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , 
     n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , 
     n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , 
     n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , 
     n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , 
     n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , 
     n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , 
     n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , 
     n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , 
     n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , 
     n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , 
     n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , 
     n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , 
     n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , 
     n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , 
     n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , 
     n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , 
     n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , 
     n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , 
     n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , 
     n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , 
     n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , 
     n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , 
     n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , 
     n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , 
     n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , 
     n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , 
     n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , 
     n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , 
     n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , 
     n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , 
     n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , 
     n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , 
     n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , 
     n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , 
     n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , 
     n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , 
     n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , 
     n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , 
     n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , 
     n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , 
     n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , 
     n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , 
     n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , 
     n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , 
     n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , 
     n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , 
     n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , 
     n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , 
     n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , 
     n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , 
     n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , 
     n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , 
     n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , 
     n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , 
     n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , 
     n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , 
     n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , 
     n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , 
     n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , 
     n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , 
     n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , 
     n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , 
     n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , 
     n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , 
     n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , 
     n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , 
     n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , 
     n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , 
     n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , 
     n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , 
     n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , 
     n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , 
     n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , 
     n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , 
     n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , 
     n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , 
     n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , 
     n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , 
     n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , 
     n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , 
     n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , 
     n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , 
     n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , 
     n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , 
     n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , 
     n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , 
     n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , 
     n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , 
     n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , 
     n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , 
     n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , 
     n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , 
     n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , 
     n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , 
     n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , 
     n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , 
     n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , 
     n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , 
     n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , 
     n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , 
     n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , 
     n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , 
     n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , 
     n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , 
     n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , 
     n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , 
     n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , 
     n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , 
     n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , 
     n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , 
     n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , 
     n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , 
     n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , 
     n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , 
     n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , 
     n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , 
     n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , 
     n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , 
     n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , 
     n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , 
     n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , 
     n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , 
     n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , 
     n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , 
     n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , 
     n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , 
     n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , 
     n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , 
     n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , 
     n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , 
     n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , 
     n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , 
     n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , 
     n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , 
     n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , 
     n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , 
     n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , 
     n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , 
     n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , 
     n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , 
     n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , 
     n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , 
     n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , 
     n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , 
     n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , 
     n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , 
     n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , 
     n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , 
     n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , 
     n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , 
     n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , 
     n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , 
     n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , 
     n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , 
     n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , 
     n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , 
     n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , 
     n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , 
     n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , 
     n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , 
     n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , 
     n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , 
     n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , 
     n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , 
     n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , 
     n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , 
     n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , 
     n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , 
     n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , 
     n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , 
     n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , 
     n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , 
     n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , 
     n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , 
     n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , 
     n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , 
     n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , 
     n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , 
     n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , 
     n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , 
     n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , 
     n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , 
     n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , 
     n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , 
     n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , 
     n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , 
     n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , 
     n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , 
     n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , 
     n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , 
     n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , 
     n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , 
     n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , 
     n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , 
     n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , 
     n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , 
     n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , 
     n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , 
     n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , 
     n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , 
     n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , 
     n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , 
     n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , 
     n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , 
     n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , 
     n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , 
     n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , 
     n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , 
     n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , 
     n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , 
     n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , 
     n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , 
     n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , 
     n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , 
     n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , 
     n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , 
     n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , 
     n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , 
     n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , 
     n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , 
     n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , 
     n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , 
     n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , 
     n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , 
     n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , 
     n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , 
     n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , 
     n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , 
     n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , 
     n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , 
     n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , 
     n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , 
     n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , 
     n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , 
     n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , 
     n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , 
     n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , 
     n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , 
     n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , 
     n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , 
     n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , 
     n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , 
     n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , 
     n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , 
     n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , 
     n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , 
     n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , 
     n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , 
     n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , 
     n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , 
     n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , 
     n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , 
     n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , 
     n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , 
     n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , 
     n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , 
     n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , 
     n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , 
     n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , 
     n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , 
     n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , 
     n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , 
     n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , 
     n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , 
     n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , 
     n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , 
     n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , 
     n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , 
     n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , 
     n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , 
     n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , 
     n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , 
     n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , 
     n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , 
     n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , 
     n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , 
     n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , 
     n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , 
     n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , 
     n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , 
     n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , 
     n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , 
     n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , 
     n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , 
     n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , 
     n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , 
     n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , 
     n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , 
     n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , 
     n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , 
     n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , 
     n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , 
     n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , 
     n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , 
     n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , 
     n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , 
     n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , 
     n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , 
     n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , 
     n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , 
     n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , 
     n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , 
     n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , 
     n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , 
     n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , 
     n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , 
     n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , 
     n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , 
     n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , 
     n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , 
     n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , 
     n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , 
     n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , 
     n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , 
     n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , 
     n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , 
     n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , 
     n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , 
     n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , 
     n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , 
     n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , 
     n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , 
     n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , 
     n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , 
     n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , 
     n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , 
     n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , 
     n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , 
     n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , 
     n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , 
     n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , 
     n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , 
     n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , 
     n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , 
     n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , 
     n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , 
     n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , 
     n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , 
     n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , 
     n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , 
     n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , 
     n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , 
     n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , 
     n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , 
     n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , 
     n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , 
     n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , 
     n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , 
     n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , 
     n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , 
     n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , 
     n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , 
     n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , 
     n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , 
     n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , 
     n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , 
     n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , 
     n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , 
     n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , 
     n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , 
     n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , 
     n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , 
     n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , 
     n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , 
     n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , 
     n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , 
     n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , 
     n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , 
     n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , 
     n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , 
     n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , 
     n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , 
     n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , 
     n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , 
     n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , 
     n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , 
     n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , 
     n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , 
     n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , 
     n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , 
     n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , 
     n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , 
     n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , 
     n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , 
     n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , 
     n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , 
     n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , 
     n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , 
     n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , 
     n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , 
     n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , 
     n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , 
     n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , 
     n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , 
     n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , 
     n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , 
     n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , 
     n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , 
     n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , 
     n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , 
     n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , 
     n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , 
     n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , 
     n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , 
     n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , 
     n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , 
     n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , 
     n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , 
     n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , 
     n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , 
     n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , 
     n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , 
     n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , 
     n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , 
     n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , 
     n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , 
     n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , 
     n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , 
     n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , 
     n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , 
     n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , 
     n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , 
     n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , 
     n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , 
     n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , 
     n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , 
     n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , 
     n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , 
     n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , 
     n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , 
     n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , 
     n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , 
     n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , 
     n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , 
     n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , 
     n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , 
     n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , 
     n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , 
     n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , 
     n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , 
     n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , 
     n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , 
     n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , 
     n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , 
     n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , 
     n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , 
     n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , 
     n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , 
     n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , 
     n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , 
     n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , 
     n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , 
     n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , 
     n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , 
     n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , 
     n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , 
     n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , 
     n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , 
     n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , 
     n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , 
     n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , 
     n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , 
     n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , 
     n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , 
     n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , 
     n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , 
     n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , 
     n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , 
     n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , 
     n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , 
     n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , 
     n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , 
     n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , 
     n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , 
     n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , 
     n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , 
     n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , 
     n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , 
     n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , 
     n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , 
     n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , 
     n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , 
     n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , 
     n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , 
     n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , 
     n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , 
     n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , 
     n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , 
     n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , 
     n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , 
     n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , 
     n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , 
     n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , 
     n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , 
     n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , 
     n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , 
     n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , 
     n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , 
     n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , 
     n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , 
     n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , 
     n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , 
     n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , 
     n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , 
     n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , 
     n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , 
     n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , 
     n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , 
     n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , 
     n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , 
     n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , 
     n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , 
     n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , 
     n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , 
     n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , 
     n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , 
     n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , 
     n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , 
     n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , 
     n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , 
     n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , 
     n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , 
     n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , 
     n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , 
     n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , 
     n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , 
     n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , 
     n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , 
     n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , 
     n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , 
     n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , 
     n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , 
     n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , 
     n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , 
     n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , 
     n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , 
     n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , 
     n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , 
     n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , 
     n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , 
     n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , 
     n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , 
     n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , 
     n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , 
     n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , 
     n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , 
     n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , 
     n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , 
     n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , 
     n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , 
     n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , 
     n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , 
     n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , 
     n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , 
     n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , 
     n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , 
     n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , 
     n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , 
     n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , 
     n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , 
     n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , 
     n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , 
     n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , 
     n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , 
     n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , 
     n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , 
     n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , 
     n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , 
     n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , 
     n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , 
     n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , 
     n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , 
     n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , 
     n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , 
     n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , 
     n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , 
     n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , 
     n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , 
     n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , 
     n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , 
     n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , 
     n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , 
     n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , 
     n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , 
     n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , 
     n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , 
     n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , 
     n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , 
     n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , 
     n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , 
     n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , 
     n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , 
     n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , 
     n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , 
     n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , 
     n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , 
     n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , 
     n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , 
     n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , 
     n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , 
     n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , 
     n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , 
     n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , 
     n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , 
     n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , 
     n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , 
     n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , 
     n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , 
     n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , 
     n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , 
     n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , 
     n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , 
     n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , 
     n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , 
     n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , 
     n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , 
     n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , 
     n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , 
     n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , 
     n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , 
     n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , 
     n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , 
     n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , 
     n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , 
     n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , 
     n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , 
     n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , 
     n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , 
     n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , 
     n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , 
     n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , 
     n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , 
     n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , 
     n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , 
     n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , 
     n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , 
     n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , 
     n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , 
     n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , 
     n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , 
     n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , 
     n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , 
     n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , 
     n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , 
     n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , 
     n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , 
     n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , 
     n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , 
     n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , 
     n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , 
     n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , 
     n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , 
     n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , 
     n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , 
     n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , 
     n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , 
     n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , 
     n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , 
     n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , 
     n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , 
     n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , 
     n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , 
     n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , 
     n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , 
     n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , 
     n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , 
     n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , 
     n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , 
     n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , 
     n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , 
     n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , 
     n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , 
     n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , 
     n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , 
     n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , 
     n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , 
     n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , 
     n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , 
     n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , 
     n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , 
     n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , 
     n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , 
     n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , 
     n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , 
     n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , 
     n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , 
     n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , 
     n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , 
     n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , 
     n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , 
     n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , 
     n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , 
     n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , 
     n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , 
     n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , 
     n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , 
     n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , 
     n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , 
     n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , 
     n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , 
     n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , 
     n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , 
     n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , 
     n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , 
     n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , 
     n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , 
     n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , 
     n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , 
     n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , 
     n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , 
     n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , 
     n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , 
     n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , 
     n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , 
     n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , 
     n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , 
     n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , 
     n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , 
     n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , 
     n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , 
     n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , 
     n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , 
     n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , 
     n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , 
     n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , 
     n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , 
     n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , 
     n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , 
     n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , 
     n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , 
     n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , 
     n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , 
     n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , 
     n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , 
     n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , 
     n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , 
     n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , 
     n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , 
     n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , 
     n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , 
     n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , 
     n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , 
     n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , 
     n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , 
     n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , 
     n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , 
     n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , 
     n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , 
     n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , 
     n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , 
     n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , 
     n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , 
     n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , 
     n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , 
     n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , 
     n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , 
     n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , 
     n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , 
     n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , 
     n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , 
     n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , 
     n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , 
     n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , 
     n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , 
     n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , 
     n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , 
     n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , 
     n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , 
     n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , 
     n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , 
     n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , 
     n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , 
     n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , 
     n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , 
     n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , 
     n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , 
     n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , 
     n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , 
     n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , 
     n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , 
     n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , 
     n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , 
     n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , 
     n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , 
     n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , 
     n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , 
     n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , 
     n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , 
     n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , 
     n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , 
     n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , 
     n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , 
     n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , 
     n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , 
     n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , 
     n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , 
     n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , 
     n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , 
     n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , 
     n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , 
     n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , 
     n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , 
     n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , 
     n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , 
     n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , 
     n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , 
     n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , 
     n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , 
     n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , 
     n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , 
     n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , 
     n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , 
     n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , 
     n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , 
     n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , 
     n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , 
     n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , 
     n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , 
     n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , 
     n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , 
     n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , 
     n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , 
     n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , 
     n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , 
     n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , 
     n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , 
     n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , 
     n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , 
     n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , 
     n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , 
     n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , 
     n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , 
     n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , 
     n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , 
     n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , 
     n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , 
     n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , 
     n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , 
     n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , 
     n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , 
     n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , 
     n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , 
     n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , 
     n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , 
     n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , 
     n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , 
     n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , 
     n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , 
     n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , 
     n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , 
     n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , 
     n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , 
     n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , 
     n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , 
     n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , 
     n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , 
     n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , 
     n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , 
     n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , 
     n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , 
     n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , 
     n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , 
     n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , 
     n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , 
     n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , 
     n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , 
     n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , 
     n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , 
     n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , 
     n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , 
     n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , 
     n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , 
     n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , 
     n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , 
     n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , 
     n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , 
     n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , 
     n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , 
     n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , 
     n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , 
     n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , 
     n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , 
     n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , 
     n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , 
     n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , 
     n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , 
     n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , 
     n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , 
     n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , 
     n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , 
     n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , 
     n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , 
     n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , 
     n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , 
     n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , 
     n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , 
     n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , 
     n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , 
     n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , 
     n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , 
     n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , 
     n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , 
     n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , 
     n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , 
     n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , 
     n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , 
     n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , 
     n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , 
     n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , 
     n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , 
     n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , 
     n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , 
     n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , 
     n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , 
     n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , 
     n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , 
     n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , 
     n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , 
     n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , 
     n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , 
     n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , 
     n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , 
     n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , 
     n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , 
     n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , 
     n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , 
     n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , 
     n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , 
     n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , 
     n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , 
     n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , 
     n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , 
     n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , 
     n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , 
     n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , 
     n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , 
     n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , 
     n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , 
     n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , 
     n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , 
     n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , 
     n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , 
     n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , 
     n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , 
     n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , 
     n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , 
     n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , 
     n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , 
     n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , 
     n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , 
     n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , 
     n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , 
     n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , 
     n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , 
     n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , 
     n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , 
     n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , 
     n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , 
     n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , 
     n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , 
     n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , 
     n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , 
     n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , 
     n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , 
     n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , 
     n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , 
     n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , 
     n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , 
     n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , 
     n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , 
     n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , 
     n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , 
     n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , 
     n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , 
     n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , 
     n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , 
     n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , 
     n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , 
     n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , 
     n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , 
     n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , 
     n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , 
     n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , 
     n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , 
     n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , 
     n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , 
     n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , 
     n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , 
     n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , 
     n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , 
     n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , 
     n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , 
     n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , 
     n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , 
     n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , 
     n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , 
     n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , 
     n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , 
     n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , 
     n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , 
     n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , 
     n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , 
     n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , 
     n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , 
     n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , 
     n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , 
     n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , 
     n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , 
     n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , 
     n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , 
     n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , 
     n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , 
     n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , 
     n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , 
     n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , 
     n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , 
     n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , 
     n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , 
     n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , 
     n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , 
     n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , 
     n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , 
     n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , 
     n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , 
     n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , 
     n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , 
     n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , 
     n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , 
     n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , 
     n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , 
     n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , 
     n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , 
     n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , 
     n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , 
     n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , 
     n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , 
     n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , 
     n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , 
     n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , 
     n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , 
     n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , 
     n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , 
     n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , 
     n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , 
     n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , 
     n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , 
     n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , 
     n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , 
     n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , 
     n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , 
     n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , 
     n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , 
     n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , 
     n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , 
     n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , 
     n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , 
     n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , 
     n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , 
     n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , 
     n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , 
     n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , 
     n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , 
     n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , 
     n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , 
     n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , 
     n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , 
     n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , 
     n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , 
     n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , 
     n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , 
     n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , 
     n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , 
     n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , 
     n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , 
     n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , 
     n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , 
     n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , 
     n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , 
     n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , 
     n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , 
     n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , 
     n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , 
     n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , 
     n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , 
     n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , 
     n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , 
     n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , 
     n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , 
     n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , 
     n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , 
     n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , 
     n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , 
     n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , 
     n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , 
     n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , 
     n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , 
     n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , 
     n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , 
     n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , 
     n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , 
     n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , 
     n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , 
     n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , 
     n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , 
     n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , 
     n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , 
     n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , 
     n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , 
     n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , 
     n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , 
     n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , 
     n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , 
     n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , 
     n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , 
     n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , 
     n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , 
     n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , 
     n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , 
     n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , 
     n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , 
     n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , 
     n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , 
     n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , 
     n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , 
     n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , 
     n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , 
     n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , 
     n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , 
     n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , 
     n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , 
     n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , 
     n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , 
     n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , 
     n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , 
     n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , 
     n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , 
     n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , 
     n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , 
     n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , 
     n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , 
     n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , 
     n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , 
     n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , 
     n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , 
     n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , 
     n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , 
     n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , 
     n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , 
     n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , 
     n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , 
     n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , 
     n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , 
     n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , 
     n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , 
     n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , 
     n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , 
     n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , 
     n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , 
     n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , 
     n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , 
     n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , 
     n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , 
     n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , 
     n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , 
     n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , 
     n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , 
     n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , 
     n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , 
     n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , 
     n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , 
     n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , 
     n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , 
     n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , 
     n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , 
     n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , 
     n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , 
     n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , 
     n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , 
     n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , 
     n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , 
     n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , 
     n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , 
     n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , 
     n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , 
     n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , 
     n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , 
     n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , 
     n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , 
     n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , 
     n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , 
     n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , 
     n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , 
     n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , 
     n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , 
     n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , 
     n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , 
     n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , 
     n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , 
     n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , 
     n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , 
     n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , 
     n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , 
     n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , 
     n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , 
     n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , 
     n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , 
     n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , 
     n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , 
     n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , 
     n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , 
     n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , 
     n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , 
     n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , 
     n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , 
     n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , 
     n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , 
     n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , 
     n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , 
     n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , 
     n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , 
     n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , 
     n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , 
     n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , 
     n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , 
     n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , 
     n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , 
     n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , 
     n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , 
     n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , 
     n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , 
     n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , 
     n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , 
     n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , 
     n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , 
     n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , 
     n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , 
     n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , 
     n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , 
     n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , 
     n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , 
     n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , 
     n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , 
     n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , 
     n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , 
     n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , 
     n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , 
     n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , 
     n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , 
     n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , 
     n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , 
     n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , 
     n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , 
     n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , 
     n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , 
     n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , 
     n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , 
     n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , 
     n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , 
     n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , 
     n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , 
     n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , 
     n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , 
     n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , 
     n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , 
     n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , 
     n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , 
     n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , 
     n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , 
     n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , 
     n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , 
     n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , 
     n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , 
     n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , 
     n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , 
     n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , 
     n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , 
     n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , 
     n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , 
     n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , 
     n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , 
     n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , 
     n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , 
     n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , 
     n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , 
     n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , 
     n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , 
     n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , 
     n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , 
     n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , 
     n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , 
     n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , 
     n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , 
     n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , 
     n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , 
     n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , 
     n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , 
     n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , 
     n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , 
     n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , 
     n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , 
     n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , 
     n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , 
     n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , 
     n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , 
     n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , 
     n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , 
     n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , 
     n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , 
     n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , 
     n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , 
     n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , 
     n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , 
     n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , 
     n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , 
     n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , 
     n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , 
     n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , 
     n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , 
     n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , 
     n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , 
     n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , 
     n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , 
     n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , 
     n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , 
     n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , 
     n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , 
     n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , 
     n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , 
     n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , 
     n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , 
     n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , 
     n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , 
     n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , 
     n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , 
     n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , 
     n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , 
     n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , 
     n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , 
     n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , 
     n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , 
     n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , 
     n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , 
     n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , 
     n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , 
     n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , 
     n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , 
     n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , 
     n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , 
     n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , 
     n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , 
     n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , 
     n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , 
     n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , 
     n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , 
     n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , 
     n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , 
     n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , 
     n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , 
     n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , 
     n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , 
     n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , 
     n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , 
     n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , 
     n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , 
     n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , 
     n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , 
     n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , 
     n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , 
     n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , 
     n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , 
     n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , 
     n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , 
     n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , 
     n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , 
     n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , 
     n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , 
     n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , 
     n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , 
     n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , 
     n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , 
     n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , 
     n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , 
     n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , 
     n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , 
     n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , 
     n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , 
     n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , 
     n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , 
     n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , 
     n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , 
     n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , 
     n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , 
     n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , 
     n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , 
     n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , 
     n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , 
     n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , 
     n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , 
     n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , 
     n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , 
     n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , 
     n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , 
     n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , 
     n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , 
     n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , 
     n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , 
     n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , 
     n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , 
     n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , 
     n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , 
     n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , 
     n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , 
     n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , 
     n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , 
     n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , 
     n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , 
     n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , 
     n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , 
     n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , 
     n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , 
     n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , 
     n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , 
     n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , 
     n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , 
     n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , 
     n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , 
     n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , 
     n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , 
     n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , 
     n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , 
     n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , 
     n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , 
     n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , 
     n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , 
     n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , 
     n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , 
     n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , 
     n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , 
     n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , 
     n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , 
     n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , 
     n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , 
     n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , 
     n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , 
     n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , 
     n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , 
     n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , 
     n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , 
     n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , 
     n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , 
     n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , 
     n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , 
     n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , 
     n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , 
     n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , 
     n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , 
     n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , 
     n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , 
     n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , 
     n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , 
     n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , 
     n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , 
     n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , 
     n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , 
     n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , 
     n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , 
     n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , 
     n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , 
     n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , 
     n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , 
     n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , 
     n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , 
     n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , 
     n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , 
     n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , 
     n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , 
     n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , 
     n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , 
     n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , 
     n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , 
     n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , 
     n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , 
     n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , 
     n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , 
     n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , 
     n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , 
     n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , 
     n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , 
     n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , 
     n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , 
     n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , 
     n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , 
     n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , 
     n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , 
     n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , 
     n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , 
     n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , 
     n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , 
     n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , 
     n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , 
     n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , 
     n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , 
     n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , 
     n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , 
     n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , 
     n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , 
     n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , 
     n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , 
     n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , 
     n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , 
     n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , 
     n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , 
     n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , 
     n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , 
     n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , 
     n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , 
     n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , 
     n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , 
     n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , 
     n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , 
     n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , 
     n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , 
     n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , 
     n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , 
     n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , 
     n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , 
     n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , 
     n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , 
     n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , 
     n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , 
     n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , 
     n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , 
     n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , 
     n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , 
     n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , 
     n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , 
     n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , 
     n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , 
     n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , 
     n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , 
     n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , 
     n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , 
     n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , 
     n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , 
     n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , 
     n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , 
     n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , 
     n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , 
     n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , 
     n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , 
     n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , 
     n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , 
     n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , 
     n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , 
     n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , 
     n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , 
     n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , 
     n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , 
     n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , 
     n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , 
     n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , 
     n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , 
     n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , 
     n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , 
     n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , 
     n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , 
     n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , 
     n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , 
     n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , 
     n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , 
     n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , 
     n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , 
     n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , 
     n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , 
     n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , 
     n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , 
     n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , 
     n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , 
     n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , 
     n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , 
     n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , 
     n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , 
     n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , 
     n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , 
     n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , 
     n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , 
     n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , 
     n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , 
     n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , 
     n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , 
     n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , 
     n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , 
     n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , 
     n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , 
     n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , 
     n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , 
     n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , 
     n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , 
     n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , 
     n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , 
     n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , 
     n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , 
     n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , 
     n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , 
     n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , 
     n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , 
     n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , 
     n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , 
     n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , 
     n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , 
     n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , 
     n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , 
     n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , 
     n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , 
     n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , 
     n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , 
     n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , 
     n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , 
     n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , 
     n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , 
     n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , 
     n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , 
     n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , 
     n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , 
     n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , 
     n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , 
     n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , 
     n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , 
     n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , 
     n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , 
     n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , 
     n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , 
     n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , 
     n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , 
     n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , 
     n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , 
     n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , 
     n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , 
     n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , 
     n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , 
     n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , 
     n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , 
     n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , 
     n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , 
     n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , 
     n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , 
     n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , 
     n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , 
     n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , 
     n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , 
     n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , 
     n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , 
     n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , 
     n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , 
     n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , 
     n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , 
     n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , 
     n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , 
     n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , 
     n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , 
     n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , 
     n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , 
     n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , 
     n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , 
     n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , 
     n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , 
     n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , 
     n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , 
     n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , 
     n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , 
     n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , 
     n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , 
     n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , 
     n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , 
     n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , 
     n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , 
     n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , 
     n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , 
     n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , 
     n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , 
     n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , 
     n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , 
     n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , 
     n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , 
     n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , 
     n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , 
     n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , 
     n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , 
     n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , 
     n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , 
     n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , 
     n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , 
     n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , 
     n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , 
     n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , 
     n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , 
     n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , 
     n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , 
     n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , 
     n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , 
     n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , 
     n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , 
     n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , 
     n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , 
     n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , 
     n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , 
     n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , 
     n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , 
     n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , 
     n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , 
     n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , 
     n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , 
     n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , 
     n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , 
     n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , 
     n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , 
     n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , 
     n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , 
     n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , 
     n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , 
     n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , 
     n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , 
     n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , 
     n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , 
     n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , 
     n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , 
     n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , 
     n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , 
     n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , 
     n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , 
     n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , 
     n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , 
     n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , 
     n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , 
     n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , 
     n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , 
     n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , 
     n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , 
     n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , 
     n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , 
     n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , 
     n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , 
     n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , 
     n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , 
     n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , 
     n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , 
     n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , 
     n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , 
     n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , 
     n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , 
     n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , 
     n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , 
     n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , 
     n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , 
     n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , 
     n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , 
     n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , 
     n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , 
     n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , 
     n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , 
     n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , 
     n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , 
     n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , 
     n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , 
     n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , 
     n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , 
     n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , 
     n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , 
     n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , 
     n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , 
     n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , 
     n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , 
     n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , 
     n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , 
     n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , 
     n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , 
     n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , 
     n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , 
     n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , 
     n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , 
     n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , 
     n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , 
     n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , 
     n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , 
     n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , 
     n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , 
     n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , 
     n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , 
     n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , 
     n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , 
     n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , 
     n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , 
     n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , 
     n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , 
     n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , 
     n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , 
     n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , 
     n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , 
     n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , 
     n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , 
     n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , 
     n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , 
     n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , 
     n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , 
     n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , 
     n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , 
     n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , 
     n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , 
     n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , 
     n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , 
     n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , 
     n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , 
     n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , 
     n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , 
     n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , 
     n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , 
     n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , 
     n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , 
     n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , 
     n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , 
     n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , 
     n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , 
     n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , 
     n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , 
     n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , 
     n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , 
     n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , 
     n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , 
     n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , 
     n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , 
     n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , 
     n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , 
     n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , 
     n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , 
     n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , 
     n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , 
     n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n51 , g50 );
buf ( n52 , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n62 , g61 );
buf ( n63 , g62 );
buf ( n64 , g63 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78 , g77 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n81 , g80 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n84 , g83 );
buf ( n85 , g84 );
buf ( n86 , g85 );
buf ( n87 , g86 );
buf ( n88 , g87 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n91 , g90 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n94 , g93 );
buf ( n95 , g94 );
buf ( n96 , g95 );
buf ( n97 , g96 );
buf ( n98 , g97 );
buf ( n99 , g98 );
buf ( n100 , g99 );
buf ( n101 , g100 );
buf ( n102 , g101 );
buf ( n103 , g102 );
buf ( n104 , g103 );
buf ( n105 , g104 );
buf ( n106 , g105 );
buf ( n107 , g106 );
buf ( n108 , g107 );
buf ( n109 , g108 );
buf ( n110 , g109 );
buf ( n111 , g110 );
buf ( n112 , g111 );
buf ( n113 , g112 );
buf ( n114 , g113 );
buf ( n115 , g114 );
buf ( n116 , g115 );
buf ( n117 , g116 );
buf ( n118 , g117 );
buf ( n119 , g118 );
buf ( n120 , g119 );
buf ( n121 , g120 );
buf ( n122 , g121 );
buf ( n123 , g122 );
buf ( n124 , g123 );
buf ( n125 , g124 );
buf ( n126 , g125 );
buf ( n127 , g126 );
buf ( n128 , g127 );
buf ( n129 , g128 );
buf ( n130 , g129 );
buf ( n131 , g130 );
buf ( n132 , g131 );
buf ( n133 , g132 );
buf ( n134 , g133 );
buf ( n135 , g134 );
buf ( n136 , g135 );
buf ( n137 , g136 );
buf ( n138 , g137 );
buf ( n139 , g138 );
buf ( n140 , g139 );
buf ( n141 , g140 );
buf ( n142 , g141 );
buf ( n143 , g142 );
buf ( n144 , g143 );
buf ( n145 , g144 );
buf ( n146 , g145 );
buf ( n147 , g146 );
buf ( n148 , g147 );
buf ( n149 , g148 );
buf ( n150 , g149 );
buf ( n151 , g150 );
buf ( n152 , g151 );
buf ( n153 , g152 );
buf ( n154 , g153 );
buf ( n155 , g154 );
buf ( n156 , g155 );
buf ( n157 , g156 );
buf ( n158 , g157 );
buf ( n159 , g158 );
buf ( n160 , g159 );
buf ( n161 , g160 );
buf ( n162 , g161 );
buf ( n163 , g162 );
buf ( n164 , g163 );
buf ( n165 , g164 );
buf ( n166 , g165 );
buf ( n167 , g166 );
buf ( n168 , g167 );
buf ( n169 , g168 );
buf ( n170 , g169 );
buf ( n171 , g170 );
buf ( n172 , g171 );
buf ( n173 , g172 );
buf ( n174 , g173 );
buf ( n175 , g174 );
buf ( n176 , g175 );
buf ( n177 , g176 );
buf ( n178 , g177 );
buf ( n179 , g178 );
buf ( n180 , g179 );
buf ( n181 , g180 );
buf ( n182 , g181 );
buf ( n183 , g182 );
buf ( n184 , g183 );
buf ( n185 , g184 );
buf ( n186 , g185 );
buf ( n187 , g186 );
buf ( n188 , g187 );
buf ( n189 , g188 );
buf ( n190 , g189 );
buf ( n191 , g190 );
buf ( n192 , g191 );
buf ( n193 , g192 );
buf ( n194 , g193 );
buf ( n195 , g194 );
buf ( n196 , g195 );
buf ( n197 , g196 );
buf ( n198 , g197 );
buf ( n199 , g198 );
buf ( n200 , g199 );
buf ( n201 , g200 );
buf ( n202 , g201 );
buf ( n203 , g202 );
buf ( n204 , g203 );
buf ( n205 , g204 );
buf ( n206 , g205 );
buf ( n207 , g206 );
buf ( n208 , g207 );
buf ( n209 , g208 );
buf ( n210 , g209 );
buf ( n211 , g210 );
buf ( n212 , g211 );
buf ( n213 , g212 );
buf ( n214 , g213 );
buf ( n215 , g214 );
buf ( n216 , g215 );
buf ( n217 , g216 );
buf ( n218 , g217 );
buf ( n219 , g218 );
buf ( n220 , g219 );
buf ( n221 , g220 );
buf ( n222 , g221 );
buf ( n223 , g222 );
buf ( n224 , g223 );
buf ( n225 , g224 );
buf ( n226 , g225 );
buf ( n227 , g226 );
buf ( n228 , g227 );
buf ( n229 , g228 );
buf ( n230 , g229 );
buf ( n231 , g230 );
buf ( n232 , g231 );
buf ( n233 , g232 );
buf ( n234 , g233 );
buf ( n235 , g234 );
buf ( n236 , g235 );
buf ( n237 , g236 );
buf ( n238 , g237 );
buf ( n239 , g238 );
buf ( n240 , g239 );
buf ( n241 , g240 );
buf ( n242 , g241 );
buf ( n243 , g242 );
buf ( n244 , g243 );
buf ( n245 , g244 );
buf ( n246 , g245 );
buf ( n247 , g246 );
buf ( n248 , g247 );
buf ( n249 , g248 );
buf ( n250 , g249 );
buf ( n251 , g250 );
buf ( n252 , g251 );
buf ( n253 , g252 );
buf ( n254 , g253 );
buf ( n255 , g254 );
buf ( n256 , g255 );
buf ( n257 , g256 );
buf ( n258 , g257 );
buf ( n259 , g258 );
buf ( n260 , g259 );
buf ( n261 , g260 );
buf ( n262 , g261 );
buf ( n263 , g262 );
buf ( n264 , g263 );
buf ( n265 , g264 );
buf ( n266 , g265 );
buf ( n267 , g266 );
buf ( n268 , g267 );
buf ( n269 , g268 );
buf ( n270 , g269 );
buf ( n271 , g270 );
buf ( n272 , g271 );
buf ( n273 , g272 );
buf ( n274 , g273 );
buf ( n275 , g274 );
buf ( n276 , g275 );
buf ( n277 , g276 );
buf ( n278 , g277 );
buf ( n279 , g278 );
buf ( n280 , g279 );
buf ( n281 , g280 );
buf ( n282 , g281 );
buf ( n283 , g282 );
buf ( n284 , g283 );
buf ( n285 , g284 );
buf ( n286 , g285 );
buf ( n287 , g286 );
buf ( n288 , g287 );
buf ( n289 , g288 );
buf ( n290 , g289 );
buf ( n291 , g290 );
buf ( n292 , g291 );
buf ( n293 , g292 );
buf ( n294 , g293 );
buf ( n295 , g294 );
buf ( n296 , g295 );
buf ( n297 , g296 );
buf ( n298 , g297 );
buf ( n299 , g298 );
buf ( n300 , g299 );
buf ( n301 , g300 );
buf ( n302 , g301 );
buf ( n303 , g302 );
buf ( n304 , g303 );
buf ( n305 , g304 );
buf ( n306 , g305 );
buf ( n307 , g306 );
buf ( n308 , g307 );
buf ( n309 , g308 );
buf ( n310 , g309 );
buf ( n311 , g310 );
buf ( n312 , g311 );
buf ( n313 , g312 );
buf ( n314 , g313 );
buf ( n315 , g314 );
buf ( n316 , g315 );
buf ( n317 , g316 );
buf ( n318 , g317 );
buf ( n319 , g318 );
buf ( n320 , g319 );
buf ( n321 , g320 );
buf ( n322 , g321 );
buf ( n323 , g322 );
buf ( n324 , g323 );
buf ( n325 , g324 );
buf ( n326 , g325 );
buf ( n327 , g326 );
buf ( n328 , g327 );
buf ( n329 , g328 );
buf ( n330 , g329 );
buf ( n331 , g330 );
buf ( n332 , g331 );
buf ( n333 , g332 );
buf ( n334 , g333 );
buf ( n335 , g334 );
buf ( n336 , g335 );
buf ( n337 , g336 );
buf ( n338 , g337 );
buf ( n339 , g338 );
buf ( n340 , g339 );
buf ( n341 , g340 );
buf ( n342 , g341 );
buf ( n343 , g342 );
buf ( n344 , g343 );
buf ( n345 , g344 );
buf ( n346 , g345 );
buf ( n347 , g346 );
buf ( n348 , g347 );
buf ( n349 , g348 );
buf ( n350 , g349 );
buf ( n351 , g350 );
buf ( n352 , g351 );
buf ( n353 , g352 );
buf ( n354 , g353 );
buf ( n355 , g354 );
buf ( n356 , g355 );
buf ( n357 , g356 );
buf ( n358 , g357 );
buf ( n359 , g358 );
buf ( n360 , g359 );
buf ( n361 , g360 );
buf ( n362 , g361 );
buf ( n363 , g362 );
buf ( n364 , g363 );
buf ( n365 , g364 );
buf ( n366 , g365 );
buf ( n367 , g366 );
buf ( n368 , g367 );
buf ( n369 , g368 );
buf ( n370 , g369 );
buf ( n371 , g370 );
buf ( n372 , g371 );
buf ( n373 , g372 );
buf ( n374 , g373 );
buf ( n375 , g374 );
buf ( n376 , g375 );
buf ( n377 , g376 );
buf ( n378 , g377 );
buf ( n379 , g378 );
buf ( n380 , g379 );
buf ( n381 , g380 );
buf ( n382 , g381 );
buf ( n383 , g382 );
buf ( n384 , g383 );
buf ( n385 , g384 );
buf ( n386 , g385 );
buf ( n387 , g386 );
buf ( n388 , g387 );
buf ( n389 , g388 );
buf ( n390 , g389 );
buf ( n391 , g390 );
buf ( n392 , g391 );
buf ( n393 , g392 );
buf ( n394 , g393 );
buf ( n395 , g394 );
buf ( n396 , g395 );
buf ( n397 , g396 );
buf ( n398 , g397 );
buf ( n399 , g398 );
buf ( n400 , g399 );
buf ( n401 , g400 );
buf ( n402 , g401 );
buf ( n403 , g402 );
buf ( n404 , g403 );
buf ( n405 , g404 );
buf ( n406 , g405 );
buf ( n407 , g406 );
buf ( n408 , g407 );
buf ( n409 , g408 );
buf ( n410 , g409 );
buf ( n411 , g410 );
buf ( n412 , g411 );
buf ( n413 , g412 );
buf ( n414 , g413 );
buf ( n415 , g414 );
buf ( n416 , g415 );
buf ( n417 , g416 );
buf ( n418 , g417 );
buf ( n419 , g418 );
buf ( n420 , g419 );
buf ( n421 , g420 );
buf ( n422 , g421 );
buf ( n423 , g422 );
buf ( n424 , g423 );
buf ( n425 , g424 );
buf ( n426 , g425 );
buf ( n427 , g426 );
buf ( n428 , g427 );
buf ( n429 , g428 );
buf ( n430 , g429 );
buf ( n431 , g430 );
buf ( n432 , g431 );
buf ( n433 , g432 );
buf ( n434 , g433 );
buf ( n435 , g434 );
buf ( n436 , g435 );
buf ( n437 , g436 );
buf ( n438 , g437 );
buf ( n439 , g438 );
buf ( n440 , g439 );
buf ( n441 , g440 );
buf ( n442 , g441 );
buf ( n443 , g442 );
buf ( n444 , g443 );
buf ( n445 , g444 );
buf ( n446 , g445 );
buf ( n447 , g446 );
buf ( n448 , g447 );
buf ( n449 , g448 );
buf ( n450 , g449 );
buf ( g450 , n451 );
buf ( g451 , n452 );
buf ( g452 , n453 );
buf ( g453 , n454 );
buf ( g454 , n455 );
buf ( g455 , n456 );
buf ( g456 , n457 );
buf ( g457 , n458 );
buf ( g458 , n459 );
buf ( g459 , n460 );
buf ( g460 , n461 );
buf ( g461 , n462 );
buf ( g462 , n463 );
buf ( g463 , n464 );
buf ( g464 , n465 );
buf ( g465 , n466 );
buf ( g466 , n467 );
buf ( g467 , n468 );
buf ( g468 , n469 );
buf ( g469 , n470 );
buf ( g470 , n471 );
buf ( g471 , n472 );
buf ( g472 , n473 );
buf ( g473 , n474 );
buf ( g474 , n475 );
buf ( g475 , n476 );
buf ( g476 , n477 );
buf ( g477 , n478 );
buf ( g478 , n479 );
buf ( g479 , n480 );
buf ( g480 , n481 );
buf ( g481 , n482 );
buf ( g482 , n483 );
buf ( g483 , n484 );
buf ( g484 , n485 );
buf ( g485 , n486 );
buf ( g486 , n487 );
buf ( g487 , n488 );
buf ( g488 , n489 );
buf ( g489 , n490 );
buf ( g490 , n491 );
buf ( g491 , n492 );
buf ( g492 , n493 );
buf ( g493 , n494 );
buf ( g494 , n495 );
buf ( g495 , n496 );
buf ( g496 , n497 );
buf ( g497 , n498 );
buf ( g498 , n499 );
buf ( g499 , n500 );
buf ( g500 , n501 );
buf ( g501 , n502 );
buf ( g502 , n503 );
buf ( g503 , n504 );
buf ( g504 , n505 );
buf ( g505 , n506 );
buf ( g506 , n507 );
buf ( g507 , n508 );
buf ( g508 , n509 );
buf ( g509 , n510 );
buf ( g510 , n511 );
buf ( g511 , n512 );
buf ( g512 , n513 );
buf ( g513 , n514 );
buf ( g514 , n515 );
buf ( g515 , n516 );
buf ( g516 , n517 );
buf ( g517 , n518 );
buf ( g518 , n519 );
buf ( g519 , n520 );
buf ( g520 , n521 );
buf ( g521 , n522 );
buf ( g522 , n523 );
buf ( g523 , n524 );
buf ( g524 , n525 );
buf ( g525 , n526 );
buf ( g526 , n527 );
buf ( g527 , n528 );
buf ( g528 , n529 );
buf ( g529 , n530 );
buf ( g530 , n531 );
buf ( g531 , n532 );
buf ( g532 , n533 );
buf ( g533 , n534 );
buf ( g534 , n535 );
buf ( g535 , n536 );
buf ( g536 , n537 );
buf ( g537 , n538 );
buf ( g538 , n539 );
buf ( g539 , n540 );
buf ( g540 , n541 );
buf ( g541 , n542 );
buf ( g542 , n543 );
buf ( g543 , n544 );
buf ( g544 , n545 );
buf ( g545 , n546 );
buf ( g546 , n547 );
buf ( g547 , n548 );
buf ( g548 , n549 );
buf ( g549 , n550 );
buf ( g550 , n551 );
buf ( g551 , n552 );
buf ( g552 , n553 );
buf ( g553 , n554 );
buf ( g554 , n555 );
buf ( g555 , n556 );
buf ( g556 , n557 );
buf ( g557 , n558 );
buf ( g558 , n559 );
buf ( g559 , n560 );
buf ( g560 , n561 );
buf ( g561 , n562 );
buf ( g562 , n563 );
buf ( g563 , n564 );
buf ( g564 , n565 );
buf ( g565 , n566 );
buf ( g566 , n567 );
buf ( g567 , n568 );
buf ( g568 , n569 );
buf ( g569 , n570 );
buf ( g570 , n571 );
buf ( g571 , n572 );
buf ( g572 , n573 );
buf ( g573 , n574 );
buf ( g574 , n575 );
buf ( g575 , n576 );
buf ( g576 , n577 );
buf ( g577 , n578 );
buf ( g578 , n579 );
buf ( g579 , n580 );
buf ( g580 , n581 );
buf ( g581 , n582 );
buf ( g582 , n583 );
buf ( g583 , n584 );
buf ( g584 , n585 );
buf ( g585 , n586 );
buf ( g586 , n587 );
buf ( g587 , n588 );
buf ( g588 , n589 );
buf ( g589 , n590 );
buf ( g590 , n591 );
buf ( g591 , n592 );
buf ( g592 , n593 );
buf ( g593 , n594 );
buf ( g594 , n595 );
buf ( g595 , n596 );
buf ( g596 , n597 );
buf ( g597 , n598 );
buf ( g598 , n599 );
buf ( g599 , n600 );
buf ( g600 , n601 );
buf ( g601 , n602 );
buf ( g602 , n603 );
buf ( g603 , n604 );
buf ( g604 , n605 );
buf ( g605 , n606 );
buf ( g606 , n607 );
buf ( g607 , n608 );
buf ( g608 , n609 );
buf ( g609 , n610 );
buf ( g610 , n611 );
buf ( g611 , n612 );
buf ( g612 , n613 );
buf ( g613 , n614 );
buf ( g614 , n615 );
buf ( g615 , n616 );
buf ( g616 , n617 );
buf ( g617 , n618 );
buf ( g618 , n619 );
buf ( g619 , n620 );
buf ( g620 , n621 );
buf ( g621 , n622 );
buf ( g622 , n623 );
buf ( g623 , n624 );
buf ( g624 , n625 );
buf ( g625 , n626 );
buf ( g626 , n627 );
buf ( g627 , n628 );
buf ( g628 , n629 );
buf ( g629 , n630 );
buf ( g630 , n631 );
buf ( g631 , n632 );
buf ( g632 , n633 );
buf ( g633 , n634 );
buf ( g634 , n635 );
buf ( g635 , n636 );
buf ( g636 , n637 );
buf ( g637 , n638 );
buf ( g638 , n639 );
buf ( g639 , n640 );
buf ( g640 , n641 );
buf ( g641 , n642 );
buf ( g642 , n643 );
buf ( g643 , n644 );
buf ( g644 , n645 );
buf ( g645 , n646 );
buf ( g646 , n647 );
buf ( g647 , n648 );
buf ( g648 , n649 );
buf ( g649 , n650 );
buf ( g650 , n651 );
buf ( g651 , n652 );
buf ( g652 , n653 );
buf ( g653 , n654 );
buf ( g654 , n655 );
buf ( g655 , n656 );
buf ( g656 , n657 );
buf ( g657 , n658 );
buf ( g658 , n659 );
buf ( g659 , n660 );
buf ( g660 , n661 );
buf ( g661 , n662 );
buf ( g662 , n663 );
buf ( g663 , n664 );
buf ( g664 , n665 );
buf ( g665 , n666 );
buf ( g666 , n667 );
buf ( g667 , n668 );
buf ( g668 , n669 );
buf ( g669 , n670 );
buf ( g670 , n671 );
buf ( g671 , n672 );
buf ( g672 , n673 );
buf ( g673 , n674 );
buf ( g674 , n675 );
buf ( g675 , n676 );
buf ( g676 , n677 );
buf ( g677 , n678 );
buf ( g678 , n679 );
buf ( g679 , n680 );
buf ( g680 , n681 );
buf ( g681 , n682 );
buf ( g682 , n683 );
buf ( g683 , n684 );
buf ( g684 , n685 );
buf ( g685 , n686 );
buf ( g686 , n687 );
buf ( g687 , n688 );
buf ( g688 , n689 );
buf ( g689 , n690 );
buf ( g690 , n691 );
buf ( g691 , n692 );
buf ( g692 , n693 );
buf ( g693 , n694 );
buf ( g694 , n695 );
buf ( g695 , n696 );
buf ( g696 , n697 );
buf ( g697 , n698 );
buf ( g698 , n699 );
buf ( g699 , n700 );
buf ( g700 , n701 );
buf ( g701 , n702 );
buf ( g702 , n703 );
buf ( g703 , n704 );
buf ( g704 , n705 );
buf ( g705 , n706 );
buf ( g706 , n707 );
buf ( g707 , n708 );
buf ( g708 , n709 );
buf ( g709 , n710 );
buf ( g710 , n711 );
buf ( g711 , n712 );
buf ( g712 , n713 );
buf ( g713 , n714 );
buf ( g714 , n715 );
buf ( g715 , n716 );
buf ( g716 , n717 );
buf ( g717 , n718 );
buf ( g718 , n719 );
buf ( g719 , n720 );
buf ( g720 , n721 );
buf ( g721 , n722 );
buf ( g722 , n723 );
buf ( g723 , n724 );
buf ( g724 , n725 );
buf ( g725 , n726 );
buf ( g726 , n727 );
buf ( g727 , n728 );
buf ( g728 , n729 );
buf ( g729 , n730 );
buf ( g730 , n731 );
buf ( g731 , n732 );
buf ( n451 , n19512 );
buf ( n452 , n19530 );
buf ( n453 , n13846 );
buf ( n454 , n20440 );
buf ( n455 , n20435 );
buf ( n456 , n7505 );
buf ( n457 , n9237 );
buf ( n458 , n19547 );
buf ( n459 , n20765 );
buf ( n460 , n20088 );
buf ( n461 , n20430 );
buf ( n462 , n18100 );
buf ( n463 , n19557 );
buf ( n464 , n16550 );
buf ( n465 , n18124 );
buf ( n466 , n20508 );
buf ( n467 , n19586 );
buf ( n468 , n20772 );
buf ( n469 , n20426 );
buf ( n470 , n19567 );
buf ( n471 , n19594 );
buf ( n472 , n19577 );
buf ( n473 , n14054 );
buf ( n474 , n14264 );
buf ( n475 , n20503 );
buf ( n476 , n19611 );
buf ( n477 , n13267 );
buf ( n478 , n9595 );
buf ( n479 , n11108 );
buf ( n480 , n20422 );
buf ( n481 , n20776 );
buf ( n482 , n20454 );
buf ( n483 , n20513 );
buf ( n484 , n20459 );
buf ( n485 , n20498 );
buf ( n486 , n20494 );
buf ( n487 , n18140 );
buf ( n488 , n19640 );
buf ( n489 , n12463 );
buf ( n490 , n14288 );
buf ( n491 , n20100 );
buf ( n492 , n14408 );
buf ( n493 , n18159 );
buf ( n494 , n8287 );
buf ( n495 , n19660 );
buf ( n496 , n14436 );
buf ( n497 , n8916 );
buf ( n498 , n20522 );
buf ( n499 , n20489 );
buf ( n500 , n20518 );
buf ( n501 , n20417 );
buf ( n502 , n20469 );
buf ( n503 , n20526 );
buf ( n504 , n20464 );
buf ( n505 , n20474 );
buf ( n506 , n20449 );
buf ( n507 , n20764 );
buf ( n508 , n20484 );
buf ( n509 , n20763 );
buf ( n510 , n20531 );
buf ( n511 , n20444 );
buf ( n512 , n20766 );
buf ( n513 , n20479 );
buf ( n514 , n20397 );
buf ( n515 , n20412 );
buf ( n516 , n20402 );
buf ( n517 , n20387 );
buf ( n518 , n18255 );
buf ( n519 , n18459 );
buf ( n520 , n9831 );
buf ( n521 , n18467 );
buf ( n522 , n10352 );
buf ( n523 , n18672 );
buf ( n524 , n20108 );
buf ( n525 , n14636 );
buf ( n526 , n19681 );
buf ( n527 , n19697 );
buf ( n528 , n19708 );
buf ( n529 , n20393 );
buf ( n530 , n15297 );
buf ( n531 , n18700 );
buf ( n532 , n2249 );
buf ( n533 , n20203 );
buf ( n534 , n3452 );
buf ( n535 , n18791 );
buf ( n536 , n18809 );
buf ( n537 , n18831 );
buf ( n538 , n19716 );
buf ( n539 , n20121 );
buf ( n540 , n20129 );
buf ( n541 , n18880 );
buf ( n542 , n19724 );
buf ( n543 , n18850 );
buf ( n544 , n19737 );
buf ( n545 , n11071 );
buf ( n546 , n18981 );
buf ( n547 , n19087 );
buf ( n548 , n20061 );
buf ( n549 , n20146 );
buf ( n550 , n11144 );
buf ( n551 , n15329 );
buf ( n552 , n11447 );
buf ( n553 , n12789 );
buf ( n554 , n19765 );
buf ( n555 , n15675 );
buf ( n556 , n20080 );
buf ( n557 , n16120 );
buf ( n558 , n16360 );
buf ( n559 , n19773 );
buf ( n560 , n19796 );
buf ( n561 , n13632 );
buf ( n562 , n11847 );
buf ( n563 , n12260 );
buf ( n564 , n19808 );
buf ( n565 , n4976 );
buf ( n566 , n19827 );
buf ( n567 , n20215 );
buf ( n568 , n19192 );
buf ( n569 , n18075 );
buf ( n570 , n19862 );
buf ( n571 , n19213 );
buf ( n572 , n19251 );
buf ( n573 , n19881 );
buf ( n574 , n19905 );
buf ( n575 , n19224 );
buf ( n576 , n16741 );
buf ( n577 , n16857 );
buf ( n578 , n16986 );
buf ( n579 , n20194 );
buf ( n580 , n11184 );
buf ( n581 , n5666 );
buf ( n582 , n19275 );
buf ( n583 , n17013 );
buf ( n584 , n20160 );
buf ( n585 , n19919 );
buf ( n586 , n13096 );
buf ( n587 , n19934 );
buf ( n588 , n17135 );
buf ( n589 , n19318 );
buf ( n590 , n13243 );
buf ( n591 , n19947 );
buf ( n592 , n17655 );
buf ( n593 , n20575 );
buf ( n594 , n19341 );
buf ( n595 , n19972 );
buf ( n596 , n17510 );
buf ( n597 , n19357 );
buf ( n598 , n17622 );
buf ( n599 , n19366 );
buf ( n600 , n19477 );
buf ( n601 , n20178 );
buf ( n602 , n20170 );
buf ( n603 , n6281 );
buf ( n604 , n20009 );
buf ( n605 , n20001 );
buf ( n606 , n20186 );
buf ( n607 , n20037 );
buf ( n608 , n19491 );
buf ( n609 , n17943 );
buf ( n610 , n17786 );
buf ( n611 , n17815 );
buf ( n612 , n17969 );
buf ( n613 , n13504 );
buf ( n614 , n16565 );
buf ( n615 , n13600 );
buf ( n616 , n106 );
buf ( n617 , n392 );
buf ( n618 , n20735 );
buf ( n619 , n392 );
buf ( n620 , n20691 );
buf ( n621 , n392 );
buf ( n622 , n20687 );
buf ( n623 , n392 );
buf ( n624 , n20551 );
buf ( n625 , n392 );
buf ( n626 , n20591 );
buf ( n627 , n392 );
buf ( n628 , n20663 );
buf ( n629 , n392 );
buf ( n630 , n20707 );
buf ( n631 , n392 );
buf ( n632 , n20651 );
buf ( n633 , n392 );
buf ( n634 , n20758 );
buf ( n635 , n392 );
buf ( n636 , n20599 );
buf ( n637 , n392 );
buf ( n638 , n20619 );
buf ( n639 , n392 );
buf ( n640 , n20559 );
buf ( n641 , n392 );
buf ( n642 , n20731 );
buf ( n643 , n392 );
buf ( n644 , n20579 );
buf ( n645 , n392 );
buf ( n646 , n20539 );
buf ( n647 , n392 );
buf ( n648 , n20679 );
buf ( n649 , n392 );
buf ( n650 , n20547 );
buf ( n651 , n392 );
buf ( n652 , n20567 );
buf ( n653 , n392 );
buf ( n654 , n20583 );
buf ( n655 , n392 );
buf ( n656 , n20711 );
buf ( n657 , n392 );
buf ( n658 , n20603 );
buf ( n659 , n392 );
buf ( n660 , n20543 );
buf ( n661 , n392 );
buf ( n662 , n20623 );
buf ( n663 , n392 );
buf ( n664 , n20659 );
buf ( n665 , n392 );
buf ( n666 , n20627 );
buf ( n667 , n392 );
buf ( n668 , n20719 );
buf ( n669 , n392 );
buf ( n670 , n20655 );
buf ( n671 , n392 );
buf ( n672 , n20753 );
buf ( n673 , n392 );
buf ( n674 , n20757 );
buf ( n675 , n392 );
buf ( n676 , n20715 );
buf ( n677 , n392 );
buf ( n678 , n20643 );
buf ( n679 , n392 );
buf ( n680 , n20667 );
buf ( n681 , n392 );
buf ( n682 , n20747 );
buf ( n683 , n392 );
buf ( n684 , n20675 );
buf ( n685 , n392 );
buf ( n686 , n20743 );
buf ( n687 , n392 );
buf ( n688 , n20615 );
buf ( n689 , n392 );
buf ( n690 , n20571 );
buf ( n691 , n392 );
buf ( n692 , n20587 );
buf ( n693 , n392 );
buf ( n694 , n20595 );
buf ( n695 , n392 );
buf ( n696 , n20631 );
buf ( n697 , n392 );
buf ( n698 , n20699 );
buf ( n699 , n392 );
buf ( n700 , n20749 );
buf ( n701 , n392 );
buf ( n702 , n20739 );
buf ( n703 , n392 );
buf ( n704 , n20555 );
buf ( n705 , n392 );
buf ( n706 , n20635 );
buf ( n707 , n392 );
buf ( n708 , n20639 );
buf ( n709 , n392 );
buf ( n710 , n20768 );
buf ( n711 , n392 );
buf ( n712 , n20647 );
buf ( n713 , n392 );
buf ( n714 , n20611 );
buf ( n715 , n392 );
buf ( n716 , n20607 );
buf ( n717 , n392 );
buf ( n718 , n20535 );
buf ( n719 , n392 );
buf ( n720 , n20695 );
buf ( n721 , n392 );
buf ( n722 , n20723 );
buf ( n723 , n392 );
buf ( n724 , n20683 );
buf ( n725 , n392 );
buf ( n726 , n20671 );
buf ( n727 , n392 );
buf ( n728 , n20727 );
buf ( n729 , n392 );
buf ( n730 , n20563 );
buf ( n731 , n392 );
buf ( n732 , n20703 );
not ( n735 , n164 );
nor ( n736 , n735 , n168 );
not ( n737 , n166 );
nand ( n738 , n736 , n737 );
not ( n739 , n164 );
nand ( n740 , n739 , n163 );
not ( n741 , n740 );
nand ( n742 , n741 , n165 );
nand ( n743 , n738 , n742 );
not ( n744 , n168 );
nand ( n745 , n744 , n163 );
not ( n746 , n745 );
nand ( n747 , n746 , n164 );
not ( n748 , n747 );
nand ( n749 , n167 , n169 );
or ( n750 , n743 , n748 , n749 );
not ( n751 , n164 );
nor ( n752 , n163 , n168 );
nand ( n753 , n751 , n752 );
not ( n754 , n167 );
nand ( n755 , n754 , n169 );
not ( n756 , n755 );
nand ( n757 , n753 , n756 );
nand ( n758 , n750 , n757 );
nand ( n759 , n163 , n164 );
not ( n760 , n759 );
nand ( n761 , n166 , n168 );
nand ( n762 , n760 , n761 );
not ( n763 , n762 );
nand ( n764 , n763 , n165 );
not ( n765 , n761 );
and ( n766 , n741 , n765 );
not ( n767 , n766 );
not ( n768 , n163 );
nand ( n769 , n768 , n168 );
not ( n770 , n769 );
nor ( n771 , n166 , n167 );
nand ( n772 , n770 , n771 );
and ( n773 , n764 , n767 , n772 );
nand ( n774 , n758 , n773 );
nor ( n775 , n165 , n166 );
nand ( n776 , n164 , n168 );
not ( n777 , n776 );
nand ( n778 , n775 , n777 );
not ( n779 , n169 );
and ( n780 , n778 , n779 );
nor ( n781 , n163 , n168 );
buf ( n782 , n781 );
buf ( n783 , n775 );
nand ( n784 , n782 , n783 );
buf ( n785 , n784 );
and ( n786 , n780 , n785 );
not ( n787 , n164 );
nor ( n788 , n787 , n163 );
not ( n789 , n788 );
nor ( n790 , n789 , n165 );
not ( n791 , n790 );
not ( n792 , n769 );
nand ( n793 , n792 , n164 );
nand ( n794 , n791 , n793 );
not ( n795 , n164 );
nand ( n796 , n795 , n166 );
not ( n797 , n796 );
nand ( n798 , n746 , n797 );
nand ( n799 , n798 , n167 );
or ( n800 , n794 , n799 );
nor ( n801 , n164 , n166 );
nand ( n802 , n163 , n168 );
not ( n803 , n802 );
nand ( n804 , n801 , n803 );
not ( n805 , n167 );
nand ( n806 , n804 , n805 );
nor ( n807 , n769 , n796 );
or ( n808 , n806 , n807 );
nand ( n809 , n800 , n808 );
nand ( n810 , n165 , n166 );
not ( n811 , n810 );
nand ( n812 , n811 , n163 );
nor ( n813 , n164 , n168 );
not ( n814 , n813 );
not ( n815 , n814 );
not ( n816 , n815 );
or ( n817 , n812 , n816 );
nand ( n818 , n786 , n809 , n817 );
and ( n819 , n774 , n818 );
not ( n820 , n166 );
nor ( n821 , n820 , n165 );
not ( n822 , n821 );
not ( n823 , n793 );
not ( n824 , n823 );
or ( n825 , n822 , n824 );
nand ( n826 , n825 , n170 );
not ( n827 , n826 );
not ( n828 , n746 );
nor ( n829 , n828 , n164 );
not ( n830 , n829 );
and ( n831 , n746 , n166 );
not ( n832 , n831 );
nand ( n833 , n830 , n832 );
not ( n834 , n164 );
nand ( n835 , n792 , n834 );
not ( n836 , n835 );
or ( n837 , n833 , n836 );
and ( n838 , n165 , n167 );
nand ( n839 , n837 , n838 );
not ( n840 , n165 );
nor ( n841 , n840 , n166 );
buf ( n842 , n841 );
nand ( n843 , n748 , n842 );
and ( n844 , n765 , n760 );
not ( n845 , n165 );
nand ( n846 , n845 , n163 );
not ( n847 , n846 );
and ( n848 , n847 , n801 );
nor ( n849 , n844 , n848 );
and ( n850 , n843 , n849 );
nor ( n851 , n850 , n167 );
not ( n852 , n851 );
nand ( n853 , n827 , n839 , n852 );
nor ( n854 , n819 , n853 );
not ( n855 , n164 );
nor ( n856 , n855 , n168 );
nand ( n857 , n847 , n856 );
not ( n858 , n857 );
not ( n859 , n164 );
nor ( n860 , n859 , n802 );
nand ( n861 , n860 , n811 );
nand ( n862 , n861 , n798 , n169 );
and ( n863 , n860 , n783 );
nor ( n864 , n862 , n863 );
not ( n865 , n864 );
or ( n866 , n858 , n865 );
nand ( n867 , n163 , n165 );
not ( n868 , n867 );
and ( n869 , n736 , n868 );
not ( n870 , n869 );
not ( n871 , n167 );
and ( n872 , n871 , n166 );
not ( n873 , n872 );
nor ( n874 , n870 , n873 );
not ( n875 , n801 );
not ( n876 , n165 );
nand ( n877 , n876 , n163 );
not ( n878 , n877 );
not ( n879 , n878 );
or ( n880 , n875 , n879 );
nand ( n881 , n880 , n779 );
nor ( n882 , n874 , n881 );
not ( n883 , n882 );
and ( n884 , n752 , n165 );
nand ( n885 , n884 , n834 );
not ( n886 , n885 );
or ( n887 , n883 , n886 );
nand ( n888 , n866 , n887 );
not ( n889 , n888 );
not ( n890 , n164 );
nand ( n891 , n890 , n168 );
not ( n892 , n891 );
nor ( n893 , n163 , n165 );
buf ( n894 , n893 );
nand ( n895 , n892 , n894 );
nor ( n896 , n895 , n166 );
nor ( n897 , n896 , n170 );
not ( n898 , n860 );
not ( n899 , n898 );
nand ( n900 , n760 , n165 );
not ( n901 , n165 );
nor ( n902 , n163 , n164 );
nand ( n903 , n901 , n902 );
nand ( n904 , n900 , n903 );
nand ( n905 , n904 , n166 );
not ( n906 , n905 );
or ( n907 , n899 , n906 );
not ( n908 , n167 );
nor ( n909 , n908 , n165 );
nand ( n910 , n907 , n909 );
nand ( n911 , n897 , n910 );
nand ( n912 , n842 , n760 );
not ( n913 , n168 );
nor ( n914 , n912 , n913 );
not ( n915 , n770 );
not ( n916 , n810 );
not ( n917 , n916 );
nor ( n918 , n915 , n917 );
nor ( n919 , n914 , n918 );
not ( n920 , n167 );
nand ( n921 , n919 , n920 );
nor ( n922 , n911 , n921 );
not ( n923 , n922 );
or ( n924 , n889 , n923 );
and ( n925 , n816 , n737 , n163 );
nor ( n926 , n925 , n884 );
not ( n927 , n926 );
not ( n928 , n882 );
or ( n929 , n927 , n928 );
and ( n930 , n841 , n168 );
not ( n931 , n930 );
not ( n932 , n164 );
nor ( n933 , n932 , n163 );
not ( n934 , n933 );
nor ( n935 , n931 , n934 );
not ( n936 , n903 );
nor ( n937 , n935 , n936 );
nand ( n938 , n864 , n937 );
nand ( n939 , n929 , n938 );
not ( n940 , n911 );
nand ( n941 , n939 , n940 , n167 );
nand ( n942 , n924 , n941 );
or ( n943 , n854 , n942 );
nand ( n944 , n878 , n765 );
nor ( n945 , n167 , n169 );
not ( n946 , n945 );
or ( n947 , n944 , n946 );
not ( n948 , n810 );
not ( n949 , n163 );
nand ( n950 , n948 , n892 , n949 );
nand ( n951 , n947 , n950 );
nand ( n952 , n166 , n167 );
not ( n953 , n952 );
not ( n954 , n953 );
not ( n955 , n168 );
nor ( n956 , n955 , n165 );
nand ( n957 , n741 , n956 );
not ( n958 , n957 );
not ( n959 , n958 );
or ( n960 , n954 , n959 );
nand ( n961 , n821 , n164 );
not ( n962 , n961 );
not ( n963 , n913 );
and ( n964 , n962 , n963 );
nor ( n965 , n964 , n766 );
or ( n966 , n965 , n749 );
nand ( n967 , n960 , n966 );
not ( n968 , n742 );
nand ( n969 , n968 , n953 );
nor ( n970 , n969 , n168 );
nor ( n971 , n951 , n967 , n970 );
nand ( n972 , n813 , n165 );
not ( n973 , n165 );
nand ( n974 , n973 , n168 );
nand ( n975 , n972 , n974 );
nand ( n976 , n975 , n846 );
nand ( n977 , n857 , n976 );
and ( n978 , n977 , n771 );
not ( n979 , n873 );
and ( n980 , n878 , n815 );
nand ( n981 , n979 , n980 );
not ( n982 , n870 );
nand ( n983 , n982 , n167 );
nand ( n984 , n981 , n983 );
or ( n985 , n978 , n984 );
nand ( n986 , n985 , n169 );
not ( n987 , n896 );
not ( n988 , n987 );
not ( n989 , n753 );
nand ( n990 , n989 , n842 );
not ( n991 , n990 );
or ( n992 , n988 , n991 );
not ( n993 , n169 );
nand ( n994 , n993 , n167 );
not ( n995 , n994 );
nand ( n996 , n992 , n995 );
and ( n997 , n971 , n986 , n996 );
nand ( n998 , n943 , n997 );
not ( n999 , n998 );
and ( n1000 , n811 , n788 , n168 );
not ( n1001 , n1000 );
not ( n1002 , n1001 );
not ( n1003 , n885 );
or ( n1004 , n1002 , n1003 );
nand ( n1005 , n1004 , n805 );
not ( n1006 , n1005 );
nand ( n1007 , n748 , n166 );
nand ( n1008 , n165 , n166 );
not ( n1009 , n1008 );
and ( n1010 , n1009 , n913 );
or ( n1011 , n807 , n1010 , n779 );
nand ( n1012 , n1011 , n749 );
nand ( n1013 , n930 , n741 );
not ( n1014 , n168 );
nor ( n1015 , n1014 , n164 );
and ( n1016 , n1015 , n165 );
not ( n1017 , n166 );
nand ( n1018 , n1017 , n167 );
not ( n1019 , n1018 );
nand ( n1020 , n1016 , n1019 );
and ( n1021 , n1007 , n1012 , n1013 , n1020 );
not ( n1022 , n1021 );
or ( n1023 , n1006 , n1022 );
nor ( n1024 , n1000 , n878 );
not ( n1025 , n1024 );
not ( n1026 , n885 );
or ( n1027 , n1025 , n1026 );
nand ( n1028 , n1027 , n920 );
not ( n1029 , n779 );
not ( n1030 , n753 );
or ( n1031 , n1029 , n1030 );
nand ( n1032 , n1031 , n946 );
not ( n1033 , n759 );
nand ( n1034 , n1033 , n166 );
not ( n1035 , n1034 );
not ( n1036 , n165 );
nand ( n1037 , n1035 , n1036 );
nand ( n1038 , n1028 , n1032 , n969 , n1037 );
nand ( n1039 , n1023 , n1038 );
nand ( n1040 , n884 , n164 );
nand ( n1041 , n936 , n913 );
not ( n1042 , n867 );
nand ( n1043 , n777 , n1042 );
nand ( n1044 , n1040 , n1041 , n1043 );
and ( n1045 , n1044 , n953 );
not ( n1046 , n898 );
not ( n1047 , n791 );
or ( n1048 , n1046 , n1047 );
nand ( n1049 , n1048 , n771 );
not ( n1050 , n170 );
nand ( n1051 , n1049 , n1050 );
nor ( n1052 , n1045 , n1051 );
nand ( n1053 , n1039 , n1052 );
not ( n1054 , n1053 );
not ( n1055 , n164 );
nand ( n1056 , n792 , n165 );
not ( n1057 , n1056 );
not ( n1058 , n1057 );
or ( n1059 , n1055 , n1058 );
nand ( n1060 , n1059 , n167 );
not ( n1061 , n1060 );
and ( n1062 , n775 , n163 );
and ( n1063 , n1062 , n168 );
not ( n1064 , n842 );
not ( n1065 , n856 );
nor ( n1066 , n1064 , n1065 );
nor ( n1067 , n1063 , n1066 );
nand ( n1068 , n1061 , n1067 );
nand ( n1069 , n1057 , n737 );
nand ( n1070 , n1069 , n805 );
and ( n1071 , n1068 , n1070 );
not ( n1072 , n165 );
nand ( n1073 , n1072 , n892 );
or ( n1074 , n1073 , n952 );
nand ( n1075 , n842 , n933 );
and ( n1076 , n1075 , n170 );
nand ( n1077 , n1074 , n1076 );
nor ( n1078 , n1071 , n1077 );
not ( n1079 , n961 );
nand ( n1080 , n1079 , n913 );
and ( n1081 , n1069 , n1080 );
not ( n1082 , n777 );
not ( n1083 , n877 );
or ( n1084 , n1082 , n1083 );
nand ( n1085 , n1084 , n1056 );
not ( n1086 , n972 );
or ( n1087 , n1085 , n1086 );
nand ( n1088 , n1087 , n805 );
nand ( n1089 , n1081 , n1088 );
not ( n1090 , n946 );
not ( n1091 , n881 );
or ( n1092 , n1090 , n1091 );
nand ( n1093 , n1092 , n772 );
or ( n1094 , n1089 , n1093 );
and ( n1095 , n782 , n1019 );
not ( n1096 , n771 );
not ( n1097 , n829 );
or ( n1098 , n1096 , n1097 );
nand ( n1099 , n1098 , n169 );
nor ( n1100 , n1095 , n1099 );
not ( n1101 , n953 );
not ( n1102 , n770 );
or ( n1103 , n1101 , n1102 );
nor ( n1104 , n810 , n949 );
nand ( n1105 , n1104 , n892 );
nand ( n1106 , n1103 , n1105 );
and ( n1107 , n975 , n167 );
nor ( n1108 , n1106 , n1107 );
nand ( n1109 , n1100 , n1108 );
nand ( n1110 , n1094 , n1109 );
nand ( n1111 , n1078 , n1110 );
not ( n1112 , n1111 );
or ( n1113 , n1054 , n1112 );
nand ( n1114 , n956 , n760 );
nand ( n1115 , n895 , n1114 );
nor ( n1116 , n847 , n1065 );
or ( n1117 , n1115 , n1116 );
nand ( n1118 , n1117 , n872 );
not ( n1119 , n957 );
nand ( n1120 , n933 , n765 );
not ( n1121 , n1120 );
or ( n1122 , n1119 , n1121 );
nand ( n1123 , n1122 , n167 );
and ( n1124 , n1123 , n169 );
nand ( n1125 , n1118 , n1124 );
nand ( n1126 , n975 , n163 );
nand ( n1127 , n856 , n894 );
and ( n1128 , n1126 , n1127 );
nor ( n1129 , n1128 , n1018 );
or ( n1130 , n1125 , n1129 );
not ( n1131 , n912 );
nor ( n1132 , n1131 , n169 );
not ( n1133 , n165 );
nand ( n1134 , n1133 , n741 );
not ( n1135 , n1134 );
nand ( n1136 , n1135 , n872 );
nand ( n1137 , n1132 , n1049 , n1136 );
nand ( n1138 , n1130 , n1137 );
nand ( n1139 , n782 , n797 );
buf ( n1140 , n842 );
nand ( n1141 , n1140 , n777 );
nand ( n1142 , n1105 , n1139 , n1141 );
and ( n1143 , n1142 , n995 );
not ( n1144 , n972 );
nand ( n1145 , n1144 , n166 );
and ( n1146 , n778 , n1145 );
nor ( n1147 , n1146 , n163 , n167 );
nor ( n1148 , n1143 , n1147 );
and ( n1149 , n1138 , n1148 );
nand ( n1150 , n1113 , n1149 );
not ( n1151 , n1150 );
and ( n1152 , n999 , n1151 );
not ( n1153 , n999 );
and ( n1154 , n1153 , n1150 );
nor ( n1155 , n1152 , n1154 );
not ( n1156 , n1155 );
not ( n1157 , n1156 );
nand ( n1158 , n1079 , n782 );
nand ( n1159 , n909 , n746 );
and ( n1160 , n990 , n1158 , n1159 );
nor ( n1161 , n976 , n989 );
or ( n1162 , n1161 , n779 );
nand ( n1163 , n1162 , n749 );
and ( n1164 , n1160 , n1163 );
nand ( n1165 , n944 , n1034 );
nand ( n1166 , n920 , n164 );
nor ( n1167 , n846 , n1166 );
nor ( n1168 , n1165 , n1167 );
not ( n1169 , n779 );
nand ( n1170 , n1010 , n949 );
not ( n1171 , n1170 );
or ( n1172 , n1169 , n1171 );
nand ( n1173 , n1172 , n994 );
and ( n1174 , n1168 , n1173 , n983 );
nor ( n1175 , n1164 , n1174 );
not ( n1176 , n167 );
nand ( n1177 , n989 , n783 );
nand ( n1178 , n1176 , n1177 );
not ( n1179 , n761 );
nand ( n1180 , n1179 , n894 );
nand ( n1181 , n1180 , n767 );
nor ( n1182 , n1178 , n1181 );
not ( n1183 , n783 );
not ( n1184 , n948 );
nand ( n1185 , n1183 , n1184 );
not ( n1186 , n1185 );
nor ( n1187 , n956 , n1042 );
nand ( n1188 , n1186 , n1187 );
not ( n1189 , n799 );
and ( n1190 , n1188 , n1189 , n1114 );
or ( n1191 , n1182 , n1190 );
nand ( n1192 , n1191 , n170 );
or ( n1193 , n1175 , n1192 );
nand ( n1194 , n823 , n167 );
nor ( n1195 , n918 , n779 );
nand ( n1196 , n1194 , n1195 );
and ( n1197 , n968 , n1019 );
or ( n1198 , n1196 , n1197 );
nand ( n1199 , n823 , n771 );
nand ( n1200 , n821 , n752 );
nand ( n1201 , n777 , n838 );
and ( n1202 , n1200 , n1201 );
nand ( n1203 , n1032 , n1199 , n1202 );
nand ( n1204 , n1198 , n1203 );
not ( n1205 , n821 );
not ( n1206 , n1205 );
not ( n1207 , n748 );
or ( n1208 , n1206 , n1207 );
not ( n1209 , n980 );
nand ( n1210 , n1208 , n1209 );
and ( n1211 , n1210 , n756 );
or ( n1212 , n920 , n163 , n1145 );
not ( n1213 , n1073 );
nand ( n1214 , n1213 , n1019 );
nand ( n1215 , n1212 , n1214 );
nor ( n1216 , n1211 , n1215 );
not ( n1217 , n894 );
not ( n1218 , n1217 );
not ( n1219 , n738 );
nand ( n1220 , n1218 , n1219 );
not ( n1221 , n1220 );
nor ( n1222 , n1013 , n167 );
nor ( n1223 , n1221 , n1222 , n170 );
nand ( n1224 , n1204 , n1216 , n1223 );
nand ( n1225 , n1193 , n1224 );
not ( n1226 , n779 );
nand ( n1227 , n831 , n1036 );
nor ( n1228 , n1227 , n164 );
not ( n1229 , n1228 );
nand ( n1230 , n913 , n953 , n933 );
nand ( n1231 , n1226 , n1229 , n1105 , n1230 );
not ( n1232 , n1178 );
not ( n1233 , n863 );
not ( n1234 , n782 );
nand ( n1235 , n1234 , n797 );
nand ( n1236 , n1233 , n1235 );
not ( n1237 , n1236 );
and ( n1238 , n1232 , n1237 );
not ( n1239 , n1069 );
nor ( n1240 , n1239 , n920 );
nor ( n1241 , n1238 , n1240 );
or ( n1242 , n1231 , n1241 );
and ( n1243 , n1220 , n1001 , n779 );
nand ( n1244 , n1120 , n167 );
not ( n1245 , n1244 );
nand ( n1246 , n1219 , n949 );
nand ( n1247 , n1245 , n1246 );
not ( n1248 , n1185 );
not ( n1249 , n829 );
or ( n1250 , n1248 , n1249 );
nand ( n1251 , n1250 , n1080 );
or ( n1252 , n1247 , n1251 );
not ( n1253 , n892 );
nand ( n1254 , n1217 , n761 );
not ( n1255 , n1254 );
not ( n1256 , n1255 );
or ( n1257 , n1253 , n1256 );
nor ( n1258 , n1034 , n974 );
nor ( n1259 , n1258 , n167 );
nand ( n1260 , n1257 , n1259 );
nand ( n1261 , n1252 , n1260 );
nand ( n1262 , n1243 , n1261 );
nand ( n1263 , n1242 , n1262 );
not ( n1264 , n871 );
not ( n1265 , n895 );
not ( n1266 , n1265 );
or ( n1267 , n1264 , n1266 );
nand ( n1268 , n1267 , n1201 );
nand ( n1269 , n1268 , n166 );
nand ( n1270 , n1225 , n1263 , n1269 );
not ( n1271 , n1270 );
not ( n1272 , n1271 );
not ( n1273 , n177 );
not ( n1274 , n174 );
nand ( n1275 , n1274 , n171 , n175 );
not ( n1276 , n172 );
nor ( n1277 , n1276 , n173 );
buf ( n1278 , n1277 );
or ( n1279 , n1275 , n1278 );
not ( n1280 , n176 );
nand ( n1281 , n1279 , n1280 );
not ( n1282 , n173 );
nand ( n1283 , n1282 , n171 );
nor ( n1284 , n1283 , n175 );
not ( n1285 , n174 );
and ( n1286 , n1284 , n1285 );
or ( n1287 , n1281 , n1286 );
nand ( n1288 , n174 , n175 );
nor ( n1289 , n1288 , n171 );
not ( n1290 , n1289 );
nand ( n1291 , n1290 , n176 );
nand ( n1292 , n1287 , n1291 );
not ( n1293 , n174 );
nor ( n1294 , n1293 , n171 );
nand ( n1295 , n1294 , n173 );
buf ( n1296 , n1295 );
not ( n1297 , n1296 );
not ( n1298 , n172 );
not ( n1299 , n1298 );
and ( n1300 , n1297 , n1299 );
not ( n1301 , n171 );
nor ( n1302 , n1301 , n175 );
nand ( n1303 , n1302 , n173 );
not ( n1304 , n1303 );
not ( n1305 , n176 );
nor ( n1306 , n1305 , n172 );
and ( n1307 , n1304 , n1306 );
nor ( n1308 , n1300 , n1307 );
nand ( n1309 , n1292 , n1308 );
not ( n1310 , n1309 );
or ( n1311 , n1273 , n1310 );
not ( n1312 , n173 );
nand ( n1313 , n1312 , n174 );
not ( n1314 , n1313 );
not ( n1315 , n175 );
nand ( n1316 , n1314 , n1315 );
not ( n1317 , n1316 );
nor ( n1318 , n171 , n174 );
not ( n1319 , n1318 );
not ( n1320 , n1319 );
nand ( n1321 , n172 , n173 );
not ( n1322 , n1321 );
nand ( n1323 , n1320 , n1322 );
not ( n1324 , n1323 );
or ( n1325 , n1317 , n1324 );
nand ( n1326 , n1325 , n176 );
not ( n1327 , n175 );
nor ( n1328 , n171 , n174 );
nand ( n1329 , n1327 , n1328 );
not ( n1330 , n1329 );
nor ( n1331 , n1330 , n1298 );
or ( n1332 , n1326 , n1331 );
not ( n1333 , n174 );
nor ( n1334 , n1333 , n175 );
nand ( n1335 , n1334 , n173 );
not ( n1336 , n1335 );
nand ( n1337 , n1336 , n171 );
nor ( n1338 , n172 , n176 );
not ( n1339 , n1338 );
or ( n1340 , n1337 , n1339 );
nand ( n1341 , n1332 , n1340 );
nor ( n1342 , n172 , n173 );
buf ( n1343 , n1342 );
not ( n1344 , n1343 );
not ( n1345 , n1344 );
not ( n1346 , n175 );
nor ( n1347 , n1346 , n174 , n171 );
buf ( n1348 , n1347 );
nand ( n1349 , n1345 , n1348 );
not ( n1350 , n178 );
nand ( n1351 , n1349 , n1350 );
nor ( n1352 , n1341 , n1351 );
nand ( n1353 , n1311 , n1352 );
nand ( n1354 , n173 , n176 );
not ( n1355 , n1354 );
not ( n1356 , n1294 );
not ( n1357 , n1356 );
nand ( n1358 , n1357 , n1338 );
not ( n1359 , n1358 );
or ( n1360 , n1355 , n1359 );
not ( n1361 , n1288 );
nand ( n1362 , n1360 , n1361 );
not ( n1363 , n1319 );
nand ( n1364 , n1363 , n1278 );
not ( n1365 , n1329 );
nand ( n1366 , n1365 , n176 );
and ( n1367 , n1362 , n1364 , n1366 );
nor ( n1368 , n1367 , n177 );
nor ( n1369 , n1353 , n1368 );
not ( n1370 , n177 );
not ( n1371 , n1370 );
not ( n1372 , n1323 );
or ( n1373 , n1371 , n1372 );
not ( n1374 , n177 );
nand ( n1375 , n1374 , n176 );
nand ( n1376 , n1373 , n1375 );
nand ( n1377 , n171 , n172 );
not ( n1378 , n1377 );
not ( n1379 , n1378 );
not ( n1380 , n1379 );
not ( n1381 , n173 );
nand ( n1382 , n1381 , n171 );
nor ( n1383 , n1382 , n176 );
not ( n1384 , n1383 );
not ( n1385 , n1384 );
or ( n1386 , n1380 , n1385 );
nand ( n1387 , n1314 , n1378 );
nand ( n1388 , n1387 , n1315 );
nand ( n1389 , n1386 , n1388 );
not ( n1390 , n1275 );
not ( n1391 , n1354 );
nand ( n1392 , n1390 , n1391 );
nand ( n1393 , n1376 , n1389 , n1392 );
not ( n1394 , n1280 );
not ( n1395 , n173 );
not ( n1396 , n174 );
nand ( n1397 , n1396 , n171 );
nor ( n1398 , n175 , n1397 );
not ( n1399 , n1398 );
or ( n1400 , n1395 , n1399 );
not ( n1401 , n171 );
nand ( n1402 , n1401 , n174 );
nor ( n1403 , n1402 , n173 );
not ( n1404 , n1403 );
nand ( n1405 , n1400 , n1404 );
not ( n1406 , n1405 );
or ( n1407 , n1394 , n1406 );
nor ( n1408 , n174 , n175 );
not ( n1409 , n1408 );
not ( n1410 , n1409 );
not ( n1411 , n172 );
nand ( n1412 , n1411 , n173 );
nor ( n1413 , n1412 , n171 );
nand ( n1414 , n1410 , n1413 );
not ( n1415 , n1397 );
not ( n1416 , n173 );
nand ( n1417 , n1416 , n176 );
not ( n1418 , n1417 );
nand ( n1419 , n1415 , n1418 );
nand ( n1420 , n1414 , n1419 );
nand ( n1421 , n1348 , n1278 );
nand ( n1422 , n1421 , n177 );
nor ( n1423 , n1420 , n1422 );
nand ( n1424 , n1407 , n1423 );
and ( n1425 , n1393 , n1424 );
nor ( n1426 , n1425 , n1350 );
or ( n1427 , n1369 , n1426 );
nand ( n1428 , n1289 , n1322 );
nand ( n1429 , n1428 , n1370 );
not ( n1430 , n1429 );
not ( n1431 , n1295 );
nand ( n1432 , n1431 , n1298 );
not ( n1433 , n1432 );
nand ( n1434 , n176 , n177 );
not ( n1435 , n1434 );
not ( n1436 , n1435 );
or ( n1437 , n1433 , n1436 );
nor ( n1438 , n172 , n173 );
not ( n1439 , n1438 );
nand ( n1440 , n171 , n174 );
nor ( n1441 , n1439 , n1440 );
nand ( n1442 , n1441 , n175 );
not ( n1443 , n172 );
nor ( n1444 , n1443 , n175 );
nand ( n1445 , n1319 , n1444 );
nor ( n1446 , n1370 , n176 );
nand ( n1447 , n1442 , n1445 , n1446 );
nand ( n1448 , n1328 , n1343 );
not ( n1449 , n1448 );
and ( n1450 , n1449 , n1315 );
or ( n1451 , n1447 , n1450 );
nand ( n1452 , n1437 , n1451 );
nor ( n1453 , n1397 , n175 );
nand ( n1454 , n1453 , n1278 );
not ( n1455 , n1335 );
nand ( n1456 , n1455 , n1378 );
nand ( n1457 , n1454 , n1456 );
nand ( n1458 , n172 , n176 );
not ( n1459 , n1458 );
and ( n1460 , n1348 , n1459 );
nor ( n1461 , n1457 , n1460 );
nand ( n1462 , n1452 , n1461 );
not ( n1463 , n1462 );
or ( n1464 , n1430 , n1463 );
not ( n1465 , n1313 );
nor ( n1466 , n171 , n175 );
not ( n1467 , n1466 );
not ( n1468 , n1467 );
nand ( n1469 , n1465 , n1468 );
not ( n1470 , n1469 );
not ( n1471 , n176 );
nand ( n1472 , n1471 , n172 );
not ( n1473 , n1472 );
and ( n1474 , n1470 , n1473 );
not ( n1475 , n173 );
nor ( n1476 , n1475 , n1288 );
and ( n1477 , n1476 , n1459 );
nor ( n1478 , n1474 , n1477 );
nand ( n1479 , n1464 , n1478 );
not ( n1480 , n1479 );
nand ( n1481 , n1427 , n1480 );
nand ( n1482 , n1277 , n175 );
not ( n1483 , n1482 );
nand ( n1484 , n171 , n174 );
not ( n1485 , n1484 );
nand ( n1486 , n1483 , n1485 );
nand ( n1487 , n1334 , n172 );
not ( n1488 , n173 );
nand ( n1489 , n1488 , n1466 );
nand ( n1490 , n1487 , n1489 );
not ( n1491 , n1490 );
not ( n1492 , n174 );
nor ( n1493 , n1492 , n175 );
nand ( n1494 , n1491 , n1493 );
nand ( n1495 , n1486 , n1494 , n1349 , n1280 );
not ( n1496 , n1298 );
not ( n1497 , n1319 );
or ( n1498 , n1496 , n1497 );
nand ( n1499 , n172 , n1402 );
nand ( n1500 , n1498 , n1499 );
not ( n1501 , n1500 );
and ( n1502 , n1501 , n175 );
nand ( n1503 , n172 , n173 );
not ( n1504 , n1503 );
nand ( n1505 , n1398 , n1504 );
not ( n1506 , n1505 );
nor ( n1507 , n1502 , n1506 );
nor ( n1508 , n1409 , n173 );
not ( n1509 , n171 );
nor ( n1510 , n1509 , n172 );
not ( n1511 , n1510 );
not ( n1512 , n1511 );
nand ( n1513 , n1508 , n1512 );
not ( n1514 , n1513 );
nor ( n1515 , n1482 , n174 );
nor ( n1516 , n1514 , n1515 , n1280 );
nand ( n1517 , n1507 , n1516 );
and ( n1518 , n1462 , n1495 , n1517 );
nor ( n1519 , n1481 , n1518 );
not ( n1520 , n1369 );
not ( n1521 , n1450 );
not ( n1522 , n175 );
nand ( n1523 , n1522 , n172 );
not ( n1524 , n1523 );
not ( n1525 , n1484 );
nand ( n1526 , n1524 , n1525 );
not ( n1527 , n1277 );
nor ( n1528 , n1527 , n1402 );
not ( n1529 , n1528 );
nand ( n1530 , n1521 , n1526 , n1529 , n1280 );
nand ( n1531 , n171 , n175 );
not ( n1532 , n1531 );
nand ( n1533 , n1314 , n1532 );
nand ( n1534 , n1533 , n176 );
not ( n1535 , n1534 );
nand ( n1536 , n1524 , n1415 );
not ( n1537 , n1527 );
and ( n1538 , n1285 , n1537 );
nor ( n1539 , n1538 , n1413 );
nand ( n1540 , n1535 , n1536 , n1539 );
nand ( n1541 , n1520 , n1530 , n1540 );
nand ( n1542 , n1519 , n1541 );
not ( n1543 , n1542 );
not ( n1544 , n1543 );
or ( n1545 , n1272 , n1544 );
nand ( n1546 , n1542 , n1270 );
nand ( n1547 , n1545 , n1546 );
not ( n1548 , n1547 );
or ( n1549 , n1157 , n1548 );
or ( n1550 , n1156 , n1547 );
nand ( n1551 , n1549 , n1550 );
not ( n1552 , n232 );
not ( n1553 , n153 );
not ( n1554 , n150 );
nor ( n1555 , n1554 , n146 );
nand ( n1556 , n1555 , n148 );
nor ( n1557 , n1556 , n151 );
or ( n1558 , n1557 , n152 );
not ( n1559 , n152 );
nand ( n1560 , n1559 , n149 );
nand ( n1561 , n1558 , n1560 );
not ( n1562 , n150 );
nor ( n1563 , n1562 , n148 );
buf ( n1564 , n1563 );
nand ( n1565 , n146 , n151 );
not ( n1566 , n1565 );
nand ( n1567 , n1564 , n1566 );
not ( n1568 , n150 );
nand ( n1569 , n147 , n151 );
nor ( n1570 , n1568 , n1569 );
not ( n1571 , n1570 );
not ( n1572 , n1569 );
buf ( n1573 , n1572 );
nor ( n1574 , n148 , n149 );
nand ( n1575 , n1573 , n1574 );
nand ( n1576 , n1561 , n1567 , n1571 , n1575 );
not ( n1577 , n1576 );
or ( n1578 , n1553 , n1577 );
nand ( n1579 , n149 , n153 );
not ( n1580 , n1579 );
not ( n1581 , n146 );
nand ( n1582 , n1581 , n151 );
not ( n1583 , n1582 );
not ( n1584 , n1583 );
nand ( n1585 , n147 , n148 );
nor ( n1586 , n1584 , n1585 );
nand ( n1587 , n1580 , n1586 );
nand ( n1588 , n1578 , n1587 );
nor ( n1589 , n146 , n151 );
and ( n1590 , n1589 , n147 );
nand ( n1591 , n1564 , n1590 );
and ( n1592 , n1591 , n152 );
nor ( n1593 , n148 , n151 );
and ( n1594 , n1593 , n146 );
not ( n1595 , n1594 );
nor ( n1596 , n146 , n147 );
nand ( n1597 , n1596 , n148 );
nand ( n1598 , n1595 , n1597 );
not ( n1599 , n147 );
and ( n1600 , n1589 , n1599 );
nor ( n1601 , n1600 , n149 );
nand ( n1602 , n1598 , n1601 );
not ( n1603 , n148 );
and ( n1604 , n1583 , n1603 , n149 );
not ( n1605 , n1604 );
not ( n1606 , n1597 );
nor ( n1607 , n150 , n151 );
nand ( n1608 , n1606 , n1607 );
and ( n1609 , n1605 , n1608 );
nand ( n1610 , n1592 , n1602 , n1609 );
and ( n1611 , n1588 , n1610 );
nor ( n1612 , n146 , n147 );
nand ( n1613 , n1603 , n1612 );
nor ( n1614 , n1613 , n151 );
not ( n1615 , n150 );
nand ( n1616 , n1614 , n1615 );
not ( n1617 , n149 );
nand ( n1618 , n1616 , n1617 );
not ( n1619 , n150 );
nor ( n1620 , n1619 , n147 );
nand ( n1621 , n1620 , n1566 );
nor ( n1622 , n1615 , n148 );
not ( n1623 , n151 );
nand ( n1624 , n1623 , n146 );
not ( n1625 , n1624 );
nand ( n1626 , n1622 , n1625 );
nand ( n1627 , n1621 , n1626 );
nor ( n1628 , n1618 , n1627 );
not ( n1629 , n148 );
nand ( n1630 , n1629 , n151 );
not ( n1631 , n1630 );
nand ( n1632 , n146 , n147 );
not ( n1633 , n1632 );
nand ( n1634 , n1631 , n1633 );
nand ( n1635 , n1634 , n149 );
not ( n1636 , n1635 );
nand ( n1637 , n1599 , n151 );
nand ( n1638 , n1637 , n148 );
not ( n1639 , n1555 );
not ( n1640 , n1639 );
and ( n1641 , n1638 , n1640 );
not ( n1642 , n151 );
not ( n1643 , n148 );
nor ( n1644 , n1643 , n150 );
not ( n1645 , n1644 );
not ( n1646 , n1645 );
and ( n1647 , n1642 , n1646 );
nor ( n1648 , n1641 , n1647 );
nand ( n1649 , n1636 , n1648 );
nand ( n1650 , n1649 , n153 );
or ( n1651 , n1628 , n1650 );
not ( n1652 , n147 );
nand ( n1653 , n1652 , n150 );
or ( n1654 , n1653 , n1624 );
not ( n1655 , n1654 );
not ( n1656 , n1574 );
not ( n1657 , n1656 );
and ( n1658 , n1655 , n1657 );
nand ( n1659 , n149 , n150 );
not ( n1660 , n1659 );
not ( n1661 , n148 );
nor ( n1662 , n1661 , n1632 );
and ( n1663 , n1660 , n1662 );
nor ( n1664 , n1658 , n1663 );
nand ( n1665 , n1651 , n1664 );
nor ( n1666 , n1611 , n1665 );
not ( n1667 , n151 );
nor ( n1668 , n1667 , n147 );
nand ( n1669 , n1668 , n148 );
not ( n1670 , n1669 );
nand ( n1671 , n1670 , n146 );
not ( n1672 , n1671 );
not ( n1673 , n149 );
and ( n1674 , n1672 , n1673 );
not ( n1675 , n147 );
nand ( n1676 , n1675 , n146 );
nor ( n1677 , n1676 , n148 );
or ( n1678 , n1557 , n1677 );
nand ( n1679 , n1678 , n149 );
not ( n1680 , n146 );
nand ( n1681 , n1680 , n147 );
not ( n1682 , n1681 );
buf ( n1683 , n1593 );
nand ( n1684 , n1682 , n1683 );
nand ( n1685 , n1679 , n1684 );
nor ( n1686 , n1674 , n1685 );
not ( n1687 , n1600 );
and ( n1688 , n1687 , n150 );
or ( n1689 , n1686 , n1688 );
nand ( n1690 , n1670 , n1615 );
not ( n1691 , n1690 );
not ( n1692 , n146 );
nor ( n1693 , n1692 , n151 );
and ( n1694 , n1693 , n147 );
buf ( n1695 , n1694 );
not ( n1696 , n1695 );
not ( n1697 , n1696 );
or ( n1698 , n1691 , n1697 );
and ( n1699 , n149 , n152 );
nand ( n1700 , n1698 , n1699 );
nand ( n1701 , n1612 , n151 );
not ( n1702 , n1701 );
nand ( n1703 , n1702 , n1603 );
not ( n1704 , n1703 );
nand ( n1705 , n1583 , n147 );
not ( n1706 , n1705 );
not ( n1707 , n1564 );
nand ( n1708 , n1706 , n1707 );
not ( n1709 , n1708 );
or ( n1710 , n1704 , n1709 );
not ( n1711 , n149 );
and ( n1712 , n1711 , n152 );
nand ( n1713 , n1710 , n1712 );
nand ( n1714 , n1693 , n148 );
not ( n1715 , n1714 );
nand ( n1716 , n1715 , n150 );
not ( n1717 , n1716 );
nand ( n1718 , n1717 , n152 );
and ( n1719 , n1700 , n1713 , n1718 );
nand ( n1720 , n1689 , n1719 );
nor ( n1721 , n149 , n150 );
and ( n1722 , n1625 , n1721 );
and ( n1723 , n148 , n149 );
or ( n1724 , n1722 , n1723 );
nand ( n1725 , n146 , n147 );
not ( n1726 , n1725 );
nand ( n1727 , n1724 , n1726 );
nand ( n1728 , n1600 , n149 );
not ( n1729 , n1589 );
not ( n1730 , n1729 );
nand ( n1731 , n1564 , n1730 );
and ( n1732 , n1727 , n1728 , n1731 );
nor ( n1733 , n1732 , n152 );
or ( n1734 , n1720 , n1733 );
not ( n1735 , n153 );
nand ( n1736 , n1734 , n1735 );
nor ( n1737 , n1653 , n1730 );
not ( n1738 , n1737 );
not ( n1739 , n1634 );
nand ( n1740 , n1739 , n1615 );
nand ( n1741 , n1738 , n1740 );
or ( n1742 , n1618 , n1741 );
nand ( n1743 , n1646 , n1625 );
not ( n1744 , n1743 );
or ( n1745 , n1744 , n1711 );
nand ( n1746 , n1742 , n1745 );
not ( n1747 , n1746 );
nand ( n1748 , n148 , n150 );
not ( n1749 , n1748 );
nand ( n1750 , n1749 , n151 );
nor ( n1751 , n1750 , n1676 );
not ( n1752 , n152 );
nand ( n1753 , n1590 , n1660 );
nor ( n1754 , n1637 , n148 );
nand ( n1755 , n1754 , n1640 );
nand ( n1756 , n1753 , n1755 );
nor ( n1757 , n1751 , n1752 , n1756 );
not ( n1758 , n1757 );
or ( n1759 , n1747 , n1758 );
nand ( n1760 , n1695 , n150 );
nand ( n1761 , n1564 , n1682 );
not ( n1762 , n1556 );
buf ( n1763 , n1668 );
nand ( n1764 , n1762 , n1763 );
not ( n1765 , n1613 );
not ( n1766 , n150 );
nand ( n1767 , n1766 , n151 );
not ( n1768 , n1767 );
nand ( n1769 , n1765 , n1768 );
nand ( n1770 , n1760 , n1761 , n1764 , n1769 );
nand ( n1771 , n1590 , n1615 );
nand ( n1772 , n1771 , n149 );
or ( n1773 , n1770 , n1772 );
and ( n1774 , n146 , n151 , n147 );
nand ( n1775 , n1774 , n1622 );
not ( n1776 , n1775 );
not ( n1777 , n1776 );
not ( n1778 , n1676 );
nand ( n1779 , n1778 , n1768 );
and ( n1780 , n1779 , n1617 );
nand ( n1781 , n1644 , n146 );
not ( n1782 , n1781 );
nor ( n1783 , n147 , n151 );
buf ( n1784 , n1783 );
nand ( n1785 , n1782 , n1784 );
not ( n1786 , n1729 );
nor ( n1787 , n148 , n150 );
nand ( n1788 , n1786 , n1787 );
nor ( n1789 , n1788 , n1599 );
not ( n1790 , n1789 );
nand ( n1791 , n1777 , n1780 , n1785 , n1790 );
nand ( n1792 , n1773 , n1791 );
not ( n1793 , n1748 );
nand ( n1794 , n1695 , n1793 );
not ( n1795 , n1794 );
nor ( n1796 , n1795 , n152 );
nand ( n1797 , n1792 , n1796 );
nand ( n1798 , n1759 , n1797 );
nand ( n1799 , n1666 , n1736 , n1798 );
not ( n1800 , n1799 );
not ( n1801 , n1800 );
or ( n1802 , n1552 , n1801 );
not ( n1803 , n1799 );
or ( n1804 , n232 , n1803 );
nand ( n1805 , n1802 , n1804 );
not ( n1806 , n1805 );
nand ( n1807 , n155 , n157 );
not ( n1808 , n1807 );
not ( n1809 , n1808 );
not ( n1810 , n156 );
nor ( n1811 , n1809 , n1810 );
nand ( n1812 , n1811 , n158 );
nor ( n1813 , n154 , n158 );
not ( n1814 , n156 );
nand ( n1815 , n1814 , n157 );
not ( n1816 , n1815 );
nand ( n1817 , n1813 , n1816 );
nand ( n1818 , n1812 , n1817 );
nand ( n1819 , n156 , n157 );
not ( n1820 , n1819 );
not ( n1821 , n1820 );
not ( n1822 , n158 );
nand ( n1823 , n1822 , n154 );
nor ( n1824 , n1821 , n1823 );
not ( n1825 , n155 );
and ( n1826 , n1824 , n1825 );
or ( n1827 , n1818 , n1826 );
not ( n1828 , n159 );
nand ( n1829 , n1827 , n1828 );
nand ( n1830 , n155 , n156 );
nor ( n1831 , n1830 , n157 );
not ( n1832 , n154 );
nand ( n1833 , n1832 , n158 );
not ( n1834 , n1833 );
nand ( n1835 , n1831 , n1834 );
and ( n1836 , n1835 , n161 );
nand ( n1837 , n1829 , n1836 );
not ( n1838 , n157 );
nand ( n1839 , n1838 , n155 );
not ( n1840 , n1839 );
not ( n1841 , n158 );
nand ( n1842 , n1840 , n1841 );
not ( n1843 , n1842 );
not ( n1844 , n159 );
nand ( n1845 , n1844 , n160 );
not ( n1846 , n1845 );
nand ( n1847 , n1843 , n1846 );
nand ( n1848 , n1840 , n1810 );
not ( n1849 , n157 );
nor ( n1850 , n1849 , n155 );
nand ( n1851 , n1850 , n158 );
nand ( n1852 , n1848 , n1851 );
not ( n1853 , n157 );
nor ( n1854 , n1853 , n155 );
nand ( n1855 , n1854 , n1810 );
not ( n1856 , n1855 );
or ( n1857 , n1852 , n1856 );
nand ( n1858 , n154 , n159 );
not ( n1859 , n1858 );
nand ( n1860 , n1857 , n1859 );
nand ( n1861 , n1847 , n1860 );
and ( n1862 , n1808 , n1810 );
nand ( n1863 , n1862 , n158 );
nor ( n1864 , n157 , n159 );
nor ( n1865 , n155 , n156 );
nand ( n1866 , n1864 , n1865 );
not ( n1867 , n1866 );
not ( n1868 , n160 );
nor ( n1869 , n1867 , n1868 );
nand ( n1870 , n1863 , n1869 );
nor ( n1871 , n1837 , n1861 , n1870 );
not ( n1872 , n1871 );
and ( n1873 , n1808 , n156 );
nand ( n1874 , n1873 , n1841 );
and ( n1875 , n1854 , n156 );
not ( n1876 , n1875 );
nand ( n1877 , n1874 , n1876 );
not ( n1878 , n1877 );
not ( n1879 , n1878 );
not ( n1880 , n1815 );
nor ( n1881 , n155 , n157 );
nand ( n1882 , n1881 , n156 );
not ( n1883 , n1882 );
nand ( n1884 , n1883 , n1841 );
not ( n1885 , n1884 );
or ( n1886 , n1880 , n1885 );
nand ( n1887 , n1886 , n159 );
not ( n1888 , n1887 );
or ( n1889 , n1879 , n1888 );
not ( n1890 , n154 );
and ( n1891 , n1876 , n1890 , n1884 );
nor ( n1892 , n154 , n159 );
nor ( n1893 , n1891 , n1892 );
nand ( n1894 , n1889 , n1893 );
not ( n1895 , n1894 );
or ( n1896 , n1872 , n1895 );
nand ( n1897 , n154 , n158 );
not ( n1898 , n1897 );
and ( n1899 , n1840 , n1898 );
nor ( n1900 , n1899 , n161 );
not ( n1901 , n1900 );
nand ( n1902 , n1824 , n155 );
not ( n1903 , n1902 );
or ( n1904 , n1901 , n1903 );
not ( n1905 , n161 );
nand ( n1906 , n1905 , n159 );
nand ( n1907 , n1904 , n1906 );
not ( n1908 , n1848 );
not ( n1909 , n1908 );
not ( n1910 , n1813 );
nor ( n1911 , n1909 , n1910 );
not ( n1912 , n155 );
nor ( n1913 , n1912 , n154 );
nand ( n1914 , n1913 , n1820 );
not ( n1915 , n1914 );
nand ( n1916 , n1915 , n159 );
nor ( n1917 , n156 , n157 );
nand ( n1918 , n1917 , n1890 );
not ( n1919 , n1918 );
nand ( n1920 , n158 , n159 );
not ( n1921 , n1920 );
nand ( n1922 , n1919 , n1921 );
nand ( n1923 , n1916 , n1922 );
nor ( n1924 , n1911 , n1923 );
nand ( n1925 , n1907 , n1924 );
not ( n1926 , n1925 );
nand ( n1927 , n1875 , n1892 );
nor ( n1928 , n154 , n158 );
nand ( n1929 , n155 , n156 );
not ( n1930 , n1929 );
and ( n1931 , n1928 , n1930 );
nand ( n1932 , n1931 , n157 );
nand ( n1933 , n1873 , n1898 );
nand ( n1934 , n1927 , n1932 , n1933 );
not ( n1935 , n1934 );
nand ( n1936 , n1856 , n158 );
not ( n1937 , n1823 );
not ( n1938 , n157 );
nand ( n1939 , n1938 , n156 );
not ( n1940 , n1939 );
nand ( n1941 , n1937 , n1940 );
nor ( n1942 , n1941 , n1825 );
nand ( n1943 , n1918 , n160 );
or ( n1944 , n1942 , n1943 );
nand ( n1945 , n1944 , n1845 );
nand ( n1946 , n1935 , n1936 , n1945 );
nand ( n1947 , n1875 , n154 );
not ( n1948 , n1947 );
not ( n1949 , n158 );
nor ( n1950 , n1949 , n159 );
nand ( n1951 , n1948 , n1950 );
or ( n1952 , n156 , n155 , n157 );
not ( n1953 , n1952 );
and ( n1954 , n1953 , n154 );
not ( n1955 , n159 );
nor ( n1956 , n1955 , n158 );
not ( n1957 , n1865 );
nand ( n1958 , n1956 , n1957 , n157 );
nor ( n1959 , n155 , n157 );
nand ( n1960 , n1959 , n1859 );
nand ( n1961 , n1817 , n1958 , n1960 , n1868 );
nor ( n1962 , n1954 , n1961 );
nand ( n1963 , n1951 , n1962 );
nand ( n1964 , n1946 , n1963 );
nand ( n1965 , n1926 , n1964 );
nand ( n1966 , n1896 , n1965 );
buf ( n1967 , n1831 );
not ( n1968 , n1967 );
nand ( n1969 , n1968 , n1936 );
not ( n1970 , n1969 );
nand ( n1971 , n1940 , n1890 );
nand ( n1972 , n1971 , n159 );
not ( n1973 , n1972 );
and ( n1974 , n1970 , n1973 );
nand ( n1975 , n1908 , n158 );
not ( n1976 , n1975 );
not ( n1977 , n1976 );
nand ( n1978 , n1862 , n1841 );
not ( n1979 , n159 );
and ( n1980 , n1977 , n1978 , n1979 );
nor ( n1981 , n1974 , n1980 );
nor ( n1982 , n1931 , n160 );
not ( n1983 , n154 );
nand ( n1984 , n1983 , n1881 );
not ( n1985 , n1984 );
nand ( n1986 , n1985 , n1841 );
nand ( n1987 , n1898 , n157 );
not ( n1988 , n1987 );
nand ( n1989 , n1988 , n1865 );
nand ( n1990 , n1982 , n1986 , n1989 , n1860 );
nor ( n1991 , n1981 , n1990 , n1837 );
or ( n1992 , n1966 , n1991 );
nand ( n1993 , n1954 , n1841 );
not ( n1994 , n1993 );
buf ( n1995 , n1911 );
not ( n1996 , n1995 );
not ( n1997 , n1996 );
or ( n1998 , n1994 , n1997 );
not ( n1999 , n160 );
nand ( n2000 , n1999 , n159 );
not ( n2001 , n2000 );
nand ( n2002 , n1998 , n2001 );
not ( n2003 , n159 );
not ( n2004 , n160 );
nand ( n2005 , n2003 , n2004 );
not ( n2006 , n2005 );
not ( n2007 , n2006 );
buf ( n2008 , n1808 );
and ( n2009 , n2008 , n158 );
not ( n2010 , n2009 );
or ( n2011 , n2007 , n2010 );
not ( n2012 , n1808 );
nor ( n2013 , n2012 , n156 , n1920 );
not ( n2014 , n2013 );
nand ( n2015 , n2011 , n2014 );
and ( n2016 , n2015 , n1890 );
not ( n2017 , n1909 );
nand ( n2018 , n2017 , n1898 );
and ( n2019 , n158 , n159 );
and ( n2020 , n2019 , n1816 , n154 );
nand ( n2021 , n2020 , n1825 );
nand ( n2022 , n2018 , n2021 );
nor ( n2023 , n2016 , n2022 );
nand ( n2024 , n2002 , n2023 );
not ( n2025 , n1936 );
nand ( n2026 , n2025 , n1892 );
not ( n2027 , n155 );
not ( n2028 , n154 );
nand ( n2029 , n2028 , n158 );
not ( n2030 , n2029 );
nand ( n2031 , n2030 , n156 );
not ( n2032 , n2031 );
not ( n2033 , n2032 );
or ( n2034 , n2027 , n2033 );
nand ( n2035 , n2034 , n1863 );
and ( n2036 , n2035 , n159 );
not ( n2037 , n1876 );
nand ( n2038 , n2037 , n1859 );
not ( n2039 , n1890 );
not ( n2040 , n1840 );
or ( n2041 , n2039 , n2040 );
nor ( n2042 , n155 , n156 );
nand ( n2043 , n2042 , n154 );
nand ( n2044 , n2041 , n2043 );
not ( n2045 , n156 );
nor ( n2046 , n2045 , n155 );
not ( n2047 , n2046 );
not ( n2048 , n154 );
nand ( n2049 , n2048 , n157 );
nor ( n2050 , n2047 , n2049 );
or ( n2051 , n2044 , n2050 );
nor ( n2052 , n158 , n159 );
nand ( n2053 , n2051 , n2052 );
nand ( n2054 , n2038 , n2053 );
nor ( n2055 , n2036 , n2054 );
and ( n2056 , n2026 , n2055 );
nor ( n2057 , n2056 , n1868 );
nor ( n2058 , n2024 , n2057 );
nand ( n2059 , n1992 , n2058 );
not ( n2060 , n2059 );
nor ( n2061 , n1851 , n1810 );
not ( n2062 , n156 );
nand ( n2063 , n2062 , n155 );
not ( n2064 , n2063 );
not ( n2065 , n158 );
nand ( n2066 , n2065 , n154 );
not ( n2067 , n2066 );
nand ( n2068 , n2064 , n2067 );
or ( n2069 , n2068 , n1864 );
nand ( n2070 , n2069 , n160 );
nor ( n2071 , n2061 , n2070 );
not ( n2072 , n2071 );
nor ( n2073 , n1897 , n155 );
not ( n2074 , n2073 );
not ( n2075 , n2074 );
not ( n2076 , n1975 );
or ( n2077 , n2075 , n2076 );
not ( n2078 , n159 );
nand ( n2079 , n2077 , n2078 );
not ( n2080 , n2079 );
or ( n2081 , n2072 , n2080 );
not ( n2082 , n2020 );
not ( n2083 , n154 );
nand ( n2084 , n2083 , n1979 );
not ( n2085 , n2084 );
not ( n2086 , n2031 );
or ( n2087 , n2085 , n2086 );
nand ( n2088 , n2087 , n157 );
not ( n2089 , n2004 );
not ( n2090 , n1952 );
or ( n2091 , n2089 , n2090 );
nand ( n2092 , n2091 , n2005 );
nand ( n2093 , n2082 , n2088 , n2092 );
nand ( n2094 , n2081 , n2093 );
not ( n2095 , n2094 );
not ( n2096 , n1921 );
nand ( n2097 , n1883 , n154 );
nand ( n2098 , n1811 , n154 );
nand ( n2099 , n2097 , n2098 );
not ( n2100 , n2099 );
or ( n2101 , n2096 , n2100 );
not ( n2102 , n1952 );
nand ( n2103 , n2102 , n158 );
not ( n2104 , n2103 );
not ( n2105 , n154 );
nand ( n2106 , n2105 , n159 );
not ( n2107 , n2106 );
nand ( n2108 , n2104 , n2107 );
nand ( n2109 , n2101 , n2108 );
not ( n2110 , n1971 );
not ( n2111 , n1811 );
not ( n2112 , n2111 );
or ( n2113 , n2110 , n2112 );
nand ( n2114 , n2113 , n2052 );
not ( n2115 , n2043 );
not ( n2116 , n154 );
nor ( n2117 , n2116 , n1929 );
nand ( n2118 , n2117 , n158 );
not ( n2119 , n2118 );
or ( n2120 , n2115 , n2119 );
nand ( n2121 , n2120 , n1864 );
nand ( n2122 , n2114 , n2121 , n1905 );
or ( n2123 , n2095 , n2109 , n2122 );
nor ( n2124 , n1830 , n157 );
and ( n2125 , n2124 , n154 );
nand ( n2126 , n1928 , n2008 );
not ( n2127 , n156 );
nor ( n2128 , n2127 , n155 );
nand ( n2129 , n2067 , n2128 );
nand ( n2130 , n2126 , n2129 );
or ( n2131 , n2125 , n2130 );
nand ( n2132 , n2131 , n159 );
and ( n2133 , n2064 , n1890 , n2019 );
nand ( n2134 , n1941 , n161 );
nor ( n2135 , n2133 , n2134 );
nand ( n2136 , n1840 , n154 );
not ( n2137 , n2136 );
nand ( n2138 , n2137 , n2052 );
nand ( n2139 , n2132 , n2135 , n2138 );
not ( n2140 , n2139 );
not ( n2141 , n2043 );
nor ( n2142 , n2141 , n1831 );
nor ( n2143 , n2117 , n2005 );
nand ( n2144 , n2142 , n2136 , n2143 );
nand ( n2145 , n1817 , n2001 );
and ( n2146 , n2144 , n2145 );
and ( n2147 , n2032 , n1825 );
nor ( n2148 , n1842 , n2107 );
nor ( n2149 , n2146 , n2147 , n2148 );
nand ( n2150 , n2140 , n2149 );
nand ( n2151 , n2123 , n2150 );
not ( n2152 , n1808 );
nor ( n2153 , n2152 , n156 );
and ( n2154 , n2153 , n154 );
nand ( n2155 , n2154 , n158 );
nand ( n2156 , n2155 , n160 );
not ( n2157 , n2052 );
not ( n2158 , n1856 );
or ( n2159 , n2157 , n2158 );
not ( n2160 , n1959 );
not ( n2161 , n158 );
and ( n2162 , n2160 , n2161 );
not ( n2163 , n1840 );
and ( n2164 , n2163 , n158 );
nor ( n2165 , n2162 , n2164 );
not ( n2166 , n1913 );
buf ( n2167 , n2166 );
nand ( n2168 , n2043 , n2167 );
or ( n2169 , n2165 , n2168 );
nand ( n2170 , n2169 , n159 );
nand ( n2171 , n2159 , n2170 );
or ( n2172 , n2156 , n2139 , n2171 );
not ( n2173 , n2172 );
or ( n2174 , n2151 , n2173 );
not ( n2175 , n2166 );
nor ( n2176 , n156 , n157 );
nand ( n2177 , n2175 , n2176 );
nand ( n2178 , n2177 , n1914 );
nand ( n2179 , n2128 , n154 );
nand ( n2180 , n1882 , n2179 );
or ( n2181 , n2178 , n2180 );
nand ( n2182 , n2181 , n1950 );
nand ( n2183 , n2182 , n160 );
not ( n2184 , n2183 );
not ( n2185 , n2126 );
nand ( n2186 , n2067 , n1816 );
nor ( n2187 , n2186 , n155 );
nor ( n2188 , n2185 , n2187 );
not ( n2189 , n1882 );
buf ( n2190 , n1813 );
nand ( n2191 , n2189 , n2190 );
and ( n2192 , n2124 , n158 );
not ( n2193 , n2192 );
nand ( n2194 , n2153 , n1890 );
nand ( n2195 , n2188 , n2191 , n2193 , n2194 );
not ( n2196 , n2195 );
and ( n2197 , n2184 , n2196 );
not ( n2198 , n1824 );
not ( n2199 , n2198 );
not ( n2200 , n2199 );
nand ( n2201 , n2200 , n2114 );
not ( n2202 , n1930 );
not ( n2203 , n2067 );
or ( n2204 , n2202 , n2203 );
nand ( n2205 , n2204 , n2001 );
nor ( n2206 , n2201 , n2104 , n2205 );
and ( n2207 , n2206 , n2155 );
nor ( n2208 , n2197 , n2207 );
nor ( n2209 , n2183 , n159 );
nand ( n2210 , n1834 , n1816 );
nand ( n2211 , n2210 , n2006 );
nor ( n2212 , n2201 , n2211 );
nor ( n2213 , n2209 , n2212 );
and ( n2214 , n2208 , n2213 );
nand ( n2215 , n2073 , n1864 );
not ( n2216 , n2215 );
not ( n2217 , n1858 );
nand ( n2218 , n1843 , n1828 );
not ( n2219 , n2218 );
or ( n2220 , n2217 , n2219 );
nand ( n2221 , n2220 , n1930 );
not ( n2222 , n2221 );
or ( n2223 , n2216 , n2222 );
nand ( n2224 , n2223 , n2168 );
not ( n2225 , n2224 );
nor ( n2226 , n2214 , n2225 );
nand ( n2227 , n2174 , n2226 );
buf ( n2228 , n2227 );
not ( n2229 , n2228 );
or ( n2230 , n2060 , n2229 );
not ( n2231 , n2059 );
not ( n2232 , n2227 );
nand ( n2233 , n2231 , n2232 );
nand ( n2234 , n2230 , n2233 );
not ( n2235 , n2234 );
not ( n2236 , n2235 );
or ( n2237 , n1806 , n2236 );
or ( n2238 , n1805 , n2235 );
nand ( n2239 , n2237 , n2238 );
not ( n2240 , n2239 );
and ( n2241 , n1551 , n2240 );
not ( n2242 , n1551 );
and ( n2243 , n2242 , n2239 );
nor ( n2244 , n2241 , n2243 );
or ( n2245 , n2244 , n1 );
not ( n2246 , n1 );
xnor ( n2247 , n232 , n233 );
or ( n2248 , n2246 , n2247 );
nand ( n2249 , n2245 , n2248 );
nand ( n2250 , n128 , n130 );
nand ( n2251 , n2250 , n131 );
not ( n2252 , n2251 );
not ( n2253 , n130 );
nand ( n2254 , n2253 , n129 );
not ( n2255 , n2254 );
not ( n2256 , n2255 );
not ( n2257 , n2256 );
or ( n2258 , n2252 , n2257 );
not ( n2259 , n128 );
nand ( n2260 , n2259 , n129 );
nand ( n2261 , n2258 , n2260 );
nand ( n2262 , n128 , n129 );
not ( n2263 , n2262 );
nand ( n2264 , n2263 , n131 );
nor ( n2265 , n133 , n134 );
and ( n2266 , n2261 , n2264 , n2265 );
not ( n2267 , n129 );
nand ( n2268 , n2267 , n130 );
not ( n2269 , n2268 );
not ( n2270 , n131 );
nand ( n2271 , n2269 , n2270 );
or ( n2272 , n2271 , n132 );
not ( n2273 , n134 );
nand ( n2274 , n2273 , n133 );
not ( n2275 , n2274 );
and ( n2276 , n2272 , n2275 );
nor ( n2277 , n2266 , n2276 );
not ( n2278 , n130 );
nand ( n2279 , n2278 , n128 );
not ( n2280 , n2279 );
nand ( n2281 , n2280 , n131 );
not ( n2282 , n2281 );
not ( n2283 , n132 );
nand ( n2284 , n2283 , n133 );
not ( n2285 , n2284 );
nand ( n2286 , n2282 , n2285 );
not ( n2287 , n2279 );
nor ( n2288 , n132 , n133 );
nand ( n2289 , n2287 , n2288 );
nand ( n2290 , n2286 , n2289 );
not ( n2291 , n131 );
nand ( n2292 , n2291 , n132 );
not ( n2293 , n2292 );
not ( n2294 , n2260 );
and ( n2295 , n2293 , n2294 );
or ( n2296 , n2277 , n2290 , n2295 );
nor ( n2297 , n2250 , n129 );
and ( n2298 , n2297 , n131 );
nand ( n2299 , n2298 , n132 );
not ( n2300 , n2299 );
not ( n2301 , n132 );
nor ( n2302 , n128 , n130 );
nand ( n2303 , n2301 , n2302 );
not ( n2304 , n2279 );
nand ( n2305 , n131 , n132 );
not ( n2306 , n2305 );
nand ( n2307 , n2304 , n2306 );
nand ( n2308 , n2303 , n2307 );
not ( n2309 , n131 );
nor ( n2310 , n128 , n129 );
buf ( n2311 , n2310 );
not ( n2312 , n2311 );
or ( n2313 , n2309 , n2312 );
not ( n2314 , n128 );
nor ( n2315 , n2314 , n131 );
not ( n2316 , n134 );
nor ( n2317 , n2315 , n2316 );
nand ( n2318 , n2313 , n2317 );
or ( n2319 , n2308 , n2318 );
not ( n2320 , n133 );
nand ( n2321 , n2320 , n134 );
nand ( n2322 , n2319 , n2321 );
not ( n2323 , n2268 );
not ( n2324 , n128 );
nand ( n2325 , n2323 , n2324 );
not ( n2326 , n2325 );
nor ( n2327 , n132 , n133 );
nand ( n2328 , n2326 , n2327 );
nand ( n2329 , n2322 , n2328 );
or ( n2330 , n2300 , n2329 );
nand ( n2331 , n2296 , n2330 );
nand ( n2332 , n2255 , n128 );
not ( n2333 , n2332 );
nand ( n2334 , n2333 , n131 );
not ( n2335 , n128 );
nor ( n2336 , n2335 , n129 );
nand ( n2337 , n2336 , n2270 );
not ( n2338 , n2337 );
nand ( n2339 , n2294 , n2301 );
not ( n2340 , n2339 );
or ( n2341 , n2338 , n2340 );
nor ( n2342 , n131 , n132 );
not ( n2343 , n2342 );
nand ( n2344 , n2341 , n2343 );
nand ( n2345 , n128 , n130 );
not ( n2346 , n2345 );
nand ( n2347 , n2342 , n2346 );
nand ( n2348 , n2334 , n2344 , n2347 );
and ( n2349 , n2348 , n133 );
not ( n2350 , n2327 );
not ( n2351 , n2282 );
or ( n2352 , n2350 , n2351 );
not ( n2353 , n2256 );
not ( n2354 , n132 );
nand ( n2355 , n2354 , n131 );
buf ( n2356 , n2355 );
not ( n2357 , n2356 );
and ( n2358 , n2353 , n2357 );
not ( n2359 , n135 );
nor ( n2360 , n2358 , n2359 );
nand ( n2361 , n2352 , n2360 );
nor ( n2362 , n2349 , n2361 );
nand ( n2363 , n2331 , n2362 );
not ( n2364 , n2363 );
not ( n2365 , n130 );
nand ( n2366 , n2365 , n2310 );
not ( n2367 , n2366 );
and ( n2368 , n2367 , n2270 );
and ( n2369 , n2302 , n129 );
nand ( n2370 , n2369 , n131 );
not ( n2371 , n130 );
nor ( n2372 , n2371 , n2262 );
nand ( n2373 , n2372 , n131 );
nand ( n2374 , n2370 , n2373 );
or ( n2375 , n2368 , n2374 );
nand ( n2376 , n132 , n133 );
not ( n2377 , n2376 );
nand ( n2378 , n2375 , n2377 );
not ( n2379 , n2262 );
nand ( n2380 , n2379 , n130 );
not ( n2381 , n2380 );
nand ( n2382 , n2255 , n2270 );
not ( n2383 , n2382 );
or ( n2384 , n2381 , n2383 );
nand ( n2385 , n2384 , n2288 );
and ( n2386 , n2385 , n2359 );
nand ( n2387 , n2378 , n2386 );
not ( n2388 , n2387 );
not ( n2389 , n130 );
nor ( n2390 , n2260 , n2389 );
nand ( n2391 , n2390 , n132 );
and ( n2392 , n2391 , n134 );
not ( n2393 , n2284 );
and ( n2394 , n2323 , n2301 );
nand ( n2395 , n2394 , n128 );
not ( n2396 , n2395 );
or ( n2397 , n2393 , n2396 );
nand ( n2398 , n2336 , n131 );
not ( n2399 , n2398 );
nand ( n2400 , n2397 , n2399 );
nand ( n2401 , n2392 , n2400 );
not ( n2402 , n131 );
nor ( n2403 , n2402 , n130 );
not ( n2404 , n2403 );
not ( n2405 , n2311 );
or ( n2406 , n2404 , n2405 );
nand ( n2407 , n131 , n132 );
not ( n2408 , n2407 );
nor ( n2409 , n2262 , n130 );
nand ( n2410 , n2408 , n2409 );
nand ( n2411 , n2406 , n2410 );
not ( n2412 , n2411 );
not ( n2413 , n129 );
nand ( n2414 , n2413 , n132 );
not ( n2415 , n2414 );
nand ( n2416 , n2287 , n2415 );
nor ( n2417 , n2305 , n128 );
not ( n2418 , n2417 );
nand ( n2419 , n2416 , n2418 );
not ( n2420 , n2419 );
and ( n2421 , n2412 , n2420 );
nor ( n2422 , n2421 , n133 );
or ( n2423 , n2401 , n2422 );
not ( n2424 , n133 );
not ( n2425 , n2424 );
not ( n2426 , n2411 );
or ( n2427 , n2425 , n2426 );
not ( n2428 , n2316 );
not ( n2429 , n2366 );
or ( n2430 , n2428 , n2429 );
not ( n2431 , n2265 );
nand ( n2432 , n2430 , n2431 );
nand ( n2433 , n2427 , n2432 );
nor ( n2434 , n131 , n133 );
not ( n2435 , n2434 );
not ( n2436 , n2435 );
nand ( n2437 , n2293 , n129 );
not ( n2438 , n2437 );
or ( n2439 , n2436 , n2438 );
nand ( n2440 , n2439 , n130 );
buf ( n2441 , n2323 );
nand ( n2442 , n2441 , n2377 , n131 );
nand ( n2443 , n2440 , n2442 );
or ( n2444 , n2433 , n2443 );
nand ( n2445 , n2423 , n2444 );
nand ( n2446 , n2388 , n2445 );
not ( n2447 , n2446 );
or ( n2448 , n2364 , n2447 );
and ( n2449 , n2310 , n132 );
not ( n2450 , n130 );
nand ( n2451 , n2449 , n2450 );
not ( n2452 , n2451 );
not ( n2453 , n2299 );
or ( n2454 , n2452 , n2453 );
nand ( n2455 , n2454 , n2275 );
not ( n2456 , n2385 );
buf ( n2457 , n2271 );
not ( n2458 , n2457 );
not ( n2459 , n133 );
nand ( n2460 , n2459 , n132 );
not ( n2461 , n2460 );
and ( n2462 , n2458 , n2461 );
nand ( n2463 , n129 , n130 );
nor ( n2464 , n2355 , n2463 );
nor ( n2465 , n2462 , n2464 );
not ( n2466 , n2465 );
or ( n2467 , n2456 , n2466 );
nand ( n2468 , n2467 , n2316 );
nor ( n2469 , n131 , n132 );
not ( n2470 , n2262 );
nand ( n2471 , n2469 , n2470 );
nand ( n2472 , n2311 , n2408 );
nand ( n2473 , n2471 , n2472 );
nor ( n2474 , n130 , n133 );
and ( n2475 , n2473 , n2474 );
nor ( n2476 , n2274 , n132 );
not ( n2477 , n2264 );
and ( n2478 , n2476 , n2477 );
nor ( n2479 , n2475 , n2478 );
and ( n2480 , n2468 , n2479 );
nand ( n2481 , n2455 , n2480 );
nor ( n2482 , n2301 , n2321 );
not ( n2483 , n2482 );
not ( n2484 , n2279 );
not ( n2485 , n129 );
nand ( n2486 , n2484 , n2485 );
nand ( n2487 , n2325 , n2486 , n2380 );
nand ( n2488 , n2487 , n2315 );
buf ( n2489 , n2369 );
nand ( n2490 , n2294 , n131 );
not ( n2491 , n2490 );
nor ( n2492 , n2489 , n2491 );
nand ( n2493 , n2488 , n2492 );
not ( n2494 , n2493 );
or ( n2495 , n2483 , n2494 );
or ( n2496 , n2325 , n2356 );
or ( n2497 , n2332 , n2301 );
not ( n2498 , n2250 );
and ( n2499 , n2498 , n2485 );
nand ( n2500 , n2499 , n2270 );
nand ( n2501 , n2496 , n2497 , n2500 , n2347 );
not ( n2502 , n2382 );
nand ( n2503 , n2502 , n2301 , n2324 );
not ( n2504 , n2503 );
or ( n2505 , n2501 , n2504 );
nand ( n2506 , n133 , n134 );
not ( n2507 , n2506 );
nand ( n2508 , n2505 , n2507 );
nand ( n2509 , n2495 , n2508 );
nor ( n2510 , n2481 , n2509 );
nand ( n2511 , n2448 , n2510 );
buf ( n2512 , n2511 );
not ( n2513 , n2512 );
not ( n2514 , n2513 );
not ( n2515 , n143 );
nor ( n2516 , n2515 , n139 );
not ( n2517 , n142 );
nand ( n2518 , n2516 , n2517 );
not ( n2519 , n140 );
nor ( n2520 , n2518 , n2519 );
not ( n2521 , n138 );
nand ( n2522 , n2520 , n2521 );
not ( n2523 , n138 );
nor ( n2524 , n2523 , n143 );
nor ( n2525 , n140 , n142 );
nand ( n2526 , n2524 , n2525 );
nor ( n2527 , n2526 , n139 );
not ( n2528 , n143 );
nor ( n2529 , n2528 , n138 );
not ( n2530 , n139 );
nor ( n2531 , n2530 , n140 );
nand ( n2532 , n2529 , n2531 );
nand ( n2533 , n139 , n143 );
not ( n2534 , n2533 );
nand ( n2535 , n2525 , n2534 );
nand ( n2536 , n2532 , n2535 );
nor ( n2537 , n2527 , n2536 );
not ( n2538 , n143 );
nand ( n2539 , n2538 , n138 , n139 );
not ( n2540 , n2539 );
nand ( n2541 , n2540 , n142 );
nand ( n2542 , n2522 , n2537 , n2541 );
nand ( n2543 , n2542 , n141 );
not ( n2544 , n2543 );
not ( n2545 , n138 );
nor ( n2546 , n2545 , n139 );
not ( n2547 , n2546 );
not ( n2548 , n140 );
nand ( n2549 , n2548 , n143 );
not ( n2550 , n2549 );
or ( n2551 , n2547 , n2550 );
not ( n2552 , n139 );
nor ( n2553 , n2552 , n138 );
buf ( n2554 , n2553 );
nor ( n2555 , n140 , n143 );
nand ( n2556 , n2554 , n2555 );
nand ( n2557 , n138 , n139 );
not ( n2558 , n2557 );
nand ( n2559 , n2550 , n2558 );
nand ( n2560 , n2551 , n2556 , n2559 );
not ( n2561 , n142 );
nor ( n2562 , n2561 , n141 );
and ( n2563 , n2560 , n2562 );
not ( n2564 , n144 );
nor ( n2565 , n2563 , n2564 );
not ( n2566 , n2565 );
or ( n2567 , n2544 , n2566 );
nor ( n2568 , n2549 , n141 );
not ( n2569 , n2568 );
not ( n2570 , n142 );
nor ( n2571 , n2570 , n138 );
not ( n2572 , n2571 );
nor ( n2573 , n2569 , n2572 );
not ( n2574 , n2573 );
not ( n2575 , n2533 );
nand ( n2576 , n2575 , n138 );
not ( n2577 , n2576 );
not ( n2578 , n140 );
nand ( n2579 , n2524 , n2578 );
buf ( n2580 , n2579 );
not ( n2581 , n2580 );
or ( n2582 , n2577 , n2581 );
nor ( n2583 , n141 , n142 );
not ( n2584 , n2583 );
not ( n2585 , n2584 );
nand ( n2586 , n2582 , n2585 );
not ( n2587 , n140 );
nor ( n2588 , n2587 , n142 );
nand ( n2589 , n138 , n143 );
not ( n2590 , n2589 );
nand ( n2591 , n2588 , n2590 );
and ( n2592 , n2591 , n2564 );
nand ( n2593 , n2574 , n2586 , n2592 );
nand ( n2594 , n2567 , n2593 );
not ( n2595 , n143 );
nand ( n2596 , n140 , n142 );
nor ( n2597 , n2595 , n2596 );
and ( n2598 , n2554 , n2597 );
nor ( n2599 , n139 , n143 );
not ( n2600 , n2599 );
nor ( n2601 , n2572 , n2600 );
not ( n2602 , n142 );
nand ( n2603 , n2602 , n140 );
not ( n2604 , n2558 );
nor ( n2605 , n2603 , n2604 );
or ( n2606 , n2598 , n2601 , n2605 );
not ( n2607 , n144 );
nand ( n2608 , n2607 , n141 );
not ( n2609 , n2608 );
nand ( n2610 , n2606 , n2609 );
nor ( n2611 , n2596 , n139 );
not ( n2612 , n2611 );
nor ( n2613 , n2612 , n138 );
nor ( n2614 , n140 , n142 );
nand ( n2615 , n2614 , n2558 );
not ( n2616 , n2615 );
or ( n2617 , n2613 , n2616 );
nor ( n2618 , n141 , n143 );
nand ( n2619 , n2617 , n2618 );
and ( n2620 , n2610 , n2619 );
and ( n2621 , n2594 , n2620 );
not ( n2622 , n2589 );
nand ( n2623 , n139 , n140 );
not ( n2624 , n2623 );
and ( n2625 , n2622 , n2624 );
nand ( n2626 , n2529 , n140 );
not ( n2627 , n2626 );
and ( n2628 , n2627 , n2564 );
nor ( n2629 , n2625 , n2628 );
nor ( n2630 , n139 , n143 );
and ( n2631 , n2630 , n138 );
nand ( n2632 , n2631 , n140 );
not ( n2633 , n140 );
nor ( n2634 , n138 , n139 );
nand ( n2635 , n2633 , n2634 );
not ( n2636 , n2635 );
nand ( n2637 , n2636 , n2595 );
and ( n2638 , n2629 , n2632 , n2637 );
and ( n2639 , n141 , n142 );
not ( n2640 , n2639 );
or ( n2641 , n2638 , n2640 );
not ( n2642 , n137 );
and ( n2643 , n2586 , n2642 );
nand ( n2644 , n2641 , n2643 );
not ( n2645 , n139 );
nor ( n2646 , n2645 , n143 );
not ( n2647 , n142 );
nor ( n2648 , n2647 , n138 );
nand ( n2649 , n2646 , n2648 );
nand ( n2650 , n2649 , n144 );
nand ( n2651 , n140 , n142 );
nor ( n2652 , n2651 , n139 );
or ( n2653 , n2650 , n2652 );
nand ( n2654 , n141 , n144 );
nand ( n2655 , n2653 , n2654 );
and ( n2656 , n2553 , n2588 );
not ( n2657 , n2618 );
and ( n2658 , n2656 , n2657 );
nand ( n2659 , n2590 , n142 );
nor ( n2660 , n2659 , n139 );
nor ( n2661 , n2658 , n2660 );
and ( n2662 , n2655 , n2661 );
not ( n2663 , n2564 );
not ( n2664 , n138 );
nand ( n2665 , n2664 , n2630 );
not ( n2666 , n2665 );
or ( n2667 , n2663 , n2666 );
nor ( n2668 , n141 , n144 );
not ( n2669 , n2668 );
nand ( n2670 , n2667 , n2669 );
not ( n2671 , n140 );
nand ( n2672 , n2671 , n142 );
not ( n2673 , n2672 );
nand ( n2674 , n2673 , n2590 );
and ( n2675 , n2670 , n2674 , n2569 );
or ( n2676 , n2662 , n2675 );
nor ( n2677 , n138 , n143 );
nand ( n2678 , n2677 , n140 );
nor ( n2679 , n2678 , n139 );
not ( n2680 , n2679 );
not ( n2681 , n2680 );
not ( n2682 , n2651 );
nand ( n2683 , n2540 , n2682 );
not ( n2684 , n2683 );
or ( n2685 , n2681 , n2684 );
not ( n2686 , n141 );
nand ( n2687 , n2685 , n2686 );
nand ( n2688 , n2676 , n2687 );
or ( n2689 , n2644 , n2688 );
not ( n2690 , n138 );
nor ( n2691 , n2690 , n139 );
not ( n2692 , n140 );
nand ( n2693 , n2692 , n142 );
and ( n2694 , n2691 , n2693 );
not ( n2695 , n2691 );
not ( n2696 , n141 );
nand ( n2697 , n2696 , n140 );
and ( n2698 , n2695 , n2697 );
nor ( n2699 , n2694 , n2698 );
not ( n2700 , n143 );
nor ( n2701 , n2700 , n138 );
nand ( n2702 , n2701 , n139 );
nand ( n2703 , n2699 , n2702 );
and ( n2704 , n2646 , n2583 );
not ( n2705 , n143 );
nand ( n2706 , n2705 , n139 );
nor ( n2707 , n2706 , n2603 );
nor ( n2708 , n2704 , n2707 );
not ( n2709 , n2564 );
not ( n2710 , n2539 );
or ( n2711 , n2709 , n2710 );
nand ( n2712 , n2711 , n2608 );
and ( n2713 , n2703 , n2708 , n2712 );
not ( n2714 , n2713 );
nand ( n2715 , n2701 , n2578 );
not ( n2716 , n2715 );
nand ( n2717 , n2716 , n2517 );
not ( n2718 , n2717 );
nand ( n2719 , n2546 , n2588 );
not ( n2720 , n2623 );
nand ( n2721 , n2524 , n2720 );
and ( n2722 , n2719 , n2721 , n2535 );
not ( n2723 , n2722 );
or ( n2724 , n2718 , n2723 );
nand ( n2725 , n2724 , n141 );
not ( n2726 , n2725 );
or ( n2727 , n2714 , n2726 );
nand ( n2728 , n2706 , n142 );
nand ( n2729 , n2600 , n2517 );
and ( n2730 , n2728 , n2729 );
nand ( n2731 , n2634 , n140 );
not ( n2732 , n140 );
nand ( n2733 , n2732 , n139 );
nand ( n2734 , n2731 , n2733 );
nor ( n2735 , n2730 , n2734 );
not ( n2736 , n2735 );
not ( n2737 , n2722 );
or ( n2738 , n2736 , n2737 );
nand ( n2739 , n2738 , n141 );
not ( n2740 , n2597 );
not ( n2741 , n2554 );
or ( n2742 , n2740 , n2741 );
nand ( n2743 , n2742 , n144 );
not ( n2744 , n143 );
nor ( n2745 , n2744 , n139 );
nand ( n2746 , n2745 , n2521 );
nor ( n2747 , n2746 , n2584 );
nor ( n2748 , n2743 , n2747 );
nand ( n2749 , n2739 , n2748 );
nand ( n2750 , n2727 , n2749 );
not ( n2751 , n141 );
nor ( n2752 , n2751 , n140 );
nand ( n2753 , n2554 , n2752 );
not ( n2754 , n2753 );
not ( n2755 , n2704 );
not ( n2756 , n2755 );
or ( n2757 , n2754 , n2756 );
buf ( n2758 , n2614 );
not ( n2759 , n2758 );
nand ( n2760 , n2757 , n2759 );
not ( n2761 , n2603 );
buf ( n2762 , n2524 );
nand ( n2763 , n2761 , n2762 );
and ( n2764 , n2760 , n2763 , n137 );
nand ( n2765 , n2750 , n2764 );
nand ( n2766 , n2689 , n2765 );
and ( n2767 , n2621 , n2766 );
not ( n2768 , n2767 );
and ( n2769 , n2514 , n2768 );
and ( n2770 , n2513 , n2767 );
nor ( n2771 , n2769 , n2770 );
and ( n2772 , n2771 , n236 );
not ( n2773 , n2771 );
not ( n2774 , n236 );
and ( n2775 , n2773 , n2774 );
nor ( n2776 , n2772 , n2775 );
nand ( n2777 , n123 , n124 );
nor ( n2778 , n2777 , n122 );
buf ( n2779 , n2778 );
nor ( n2780 , n120 , n121 );
not ( n2781 , n2780 );
not ( n2782 , n2781 );
nand ( n2783 , n2779 , n2782 );
not ( n2784 , n2783 );
not ( n2785 , n126 );
not ( n2786 , n2785 );
not ( n2787 , n124 );
nor ( n2788 , n2787 , n122 );
not ( n2789 , n121 );
nor ( n2790 , n2789 , n123 );
nand ( n2791 , n2788 , n2790 );
not ( n2792 , n2791 );
or ( n2793 , n2786 , n2792 );
not ( n2794 , n124 );
nand ( n2795 , n2794 , n123 );
nand ( n2796 , n2795 , n125 );
nand ( n2797 , n2796 , n2785 );
nand ( n2798 , n2793 , n2797 );
not ( n2799 , n2798 );
or ( n2800 , n2784 , n2799 );
not ( n2801 , n125 );
nand ( n2802 , n2801 , n123 );
not ( n2803 , n123 );
nand ( n2804 , n2803 , n124 );
nand ( n2805 , n2802 , n2804 );
not ( n2806 , n122 );
nand ( n2807 , n2806 , n123 );
not ( n2808 , n2807 );
or ( n2809 , n2805 , n2808 );
nor ( n2810 , n122 , n123 );
nand ( n2811 , n2810 , n125 );
nand ( n2812 , n2809 , n2811 );
not ( n2813 , n2812 );
nor ( n2814 , n123 , n124 );
buf ( n2815 , n2814 );
not ( n2816 , n125 );
nand ( n2817 , n2815 , n2816 );
or ( n2818 , n2817 , n121 );
nand ( n2819 , n2818 , n120 );
not ( n2820 , n2819 );
or ( n2821 , n2813 , n2820 );
not ( n2822 , n121 );
nand ( n2823 , n2822 , n125 );
not ( n2824 , n2823 );
not ( n2825 , n122 );
nand ( n2826 , n2825 , n124 );
nand ( n2827 , n2824 , n2826 );
not ( n2828 , n120 );
nor ( n2829 , n2827 , n2828 );
not ( n2830 , n123 );
nand ( n2831 , n2830 , n125 );
not ( n2832 , n2831 );
nand ( n2833 , n121 , n122 );
not ( n2834 , n2833 );
nand ( n2835 , n2832 , n2834 );
nand ( n2836 , n2835 , n126 );
nor ( n2837 , n2829 , n2836 );
nand ( n2838 , n2821 , n2837 );
nand ( n2839 , n2800 , n2838 );
not ( n2840 , n2839 );
not ( n2841 , n122 );
nor ( n2842 , n2841 , n125 , n123 );
not ( n2843 , n121 );
nand ( n2844 , n2842 , n2843 );
nand ( n2845 , n2808 , n125 );
not ( n2846 , n2845 );
not ( n2847 , n2843 );
and ( n2848 , n2846 , n2847 );
not ( n2849 , n125 );
nand ( n2850 , n2849 , n124 );
or ( n2851 , n121 , n123 );
nor ( n2852 , n2850 , n2851 );
nor ( n2853 , n2848 , n2852 );
not ( n2854 , n124 );
nand ( n2855 , n2842 , n2854 );
and ( n2856 , n2844 , n2853 , n2855 );
not ( n2857 , n120 );
or ( n2858 , n2856 , n2857 );
not ( n2859 , n126 );
nand ( n2860 , n2859 , n120 );
not ( n2861 , n2860 );
not ( n2862 , n2861 );
not ( n2863 , n124 );
nand ( n2864 , n2863 , n123 );
not ( n2865 , n2864 );
nand ( n2866 , n121 , n124 );
not ( n2867 , n2866 );
or ( n2868 , n2865 , n2867 );
nand ( n2869 , n2868 , n2802 );
not ( n2870 , n2869 );
or ( n2871 , n2862 , n2870 );
not ( n2872 , n2817 );
not ( n2873 , n2781 );
and ( n2874 , n2872 , n2873 );
not ( n2875 , n122 );
nor ( n2876 , n2875 , n124 );
not ( n2877 , n2876 );
not ( n2878 , n2824 );
or ( n2879 , n2877 , n2878 );
nand ( n2880 , n2879 , n127 );
nor ( n2881 , n2874 , n2880 );
nand ( n2882 , n2871 , n2881 );
not ( n2883 , n2882 );
nand ( n2884 , n2858 , n2883 );
or ( n2885 , n2840 , n2884 );
nor ( n2886 , n2828 , n121 );
not ( n2887 , n2886 );
nor ( n2888 , n2807 , n125 );
not ( n2889 , n2888 );
or ( n2890 , n2887 , n2889 );
nand ( n2891 , n2890 , n2785 );
not ( n2892 , n2834 );
buf ( n2893 , n2777 );
nor ( n2894 , n2892 , n2893 );
nor ( n2895 , n2891 , n2894 );
nor ( n2896 , n123 , n125 );
nand ( n2897 , n2896 , n121 );
not ( n2898 , n2897 );
not ( n2899 , n122 );
nand ( n2900 , n2899 , n121 );
not ( n2901 , n2900 );
nand ( n2902 , n2901 , n2815 );
not ( n2903 , n2902 );
or ( n2904 , n2898 , n2903 );
not ( n2905 , n120 );
nand ( n2906 , n2904 , n2905 );
nand ( n2907 , n2895 , n2906 );
not ( n2908 , n2804 );
nor ( n2909 , n121 , n122 );
nand ( n2910 , n2908 , n2909 );
not ( n2911 , n2910 );
nand ( n2912 , n2911 , n125 );
not ( n2913 , n2912 );
or ( n2914 , n2907 , n2913 );
not ( n2915 , n125 );
nand ( n2916 , n2915 , n124 );
nor ( n2917 , n2916 , n120 );
not ( n2918 , n2917 );
not ( n2919 , n2916 );
nand ( n2920 , n2919 , n2834 );
and ( n2921 , n2918 , n2920 , n126 );
nand ( n2922 , n121 , n125 );
not ( n2923 , n2922 );
not ( n2924 , n122 );
nand ( n2925 , n2795 , n2924 );
not ( n2926 , n2925 );
or ( n2927 , n2923 , n2926 );
nand ( n2928 , n2927 , n120 );
nand ( n2929 , n2921 , n2928 );
nand ( n2930 , n2914 , n2929 );
nand ( n2931 , n2908 , n122 );
not ( n2932 , n2931 );
not ( n2933 , n125 );
nand ( n2934 , n2933 , n2876 );
not ( n2935 , n2934 );
or ( n2936 , n2932 , n2935 );
nand ( n2937 , n2936 , n2782 );
not ( n2938 , n2796 );
nand ( n2939 , n120 , n121 );
not ( n2940 , n2939 );
nand ( n2941 , n2938 , n2940 );
not ( n2942 , n127 );
and ( n2943 , n2937 , n2941 , n2942 );
nand ( n2944 , n2930 , n2943 );
nand ( n2945 , n2885 , n2944 );
not ( n2946 , n2924 );
nand ( n2947 , n2946 , n2864 );
not ( n2948 , n2947 );
nand ( n2949 , n2948 , n2816 );
not ( n2950 , n2949 );
nand ( n2951 , n2779 , n125 );
not ( n2952 , n2951 );
or ( n2953 , n2950 , n2952 );
nand ( n2954 , n2953 , n2843 );
not ( n2955 , n2954 );
not ( n2956 , n2850 );
not ( n2957 , n2810 );
not ( n2958 , n2957 );
nand ( n2959 , n2956 , n2958 );
nand ( n2960 , n2815 , n2834 );
and ( n2961 , n2959 , n2960 );
not ( n2962 , n2961 );
or ( n2963 , n2955 , n2962 );
nand ( n2964 , n2963 , n2861 );
not ( n2965 , n2925 );
nand ( n2966 , n2965 , n121 );
buf ( n2967 , n2824 );
nand ( n2968 , n122 , n123 );
not ( n2969 , n2968 );
nand ( n2970 , n2967 , n2969 );
nand ( n2971 , n2966 , n2970 );
nand ( n2972 , n120 , n126 );
not ( n2973 , n2972 );
and ( n2974 , n2971 , n2973 );
not ( n2975 , n125 );
nand ( n2976 , n122 , n124 );
not ( n2977 , n2976 );
nand ( n2978 , n2975 , n2977 );
nor ( n2979 , n2978 , n121 );
not ( n2980 , n2979 );
not ( n2981 , n2980 );
not ( n2982 , n2937 );
or ( n2983 , n2981 , n2982 );
nand ( n2984 , n2983 , n126 );
not ( n2985 , n120 );
nand ( n2986 , n2985 , n121 );
not ( n2987 , n2986 );
nand ( n2988 , n2987 , n126 );
not ( n2989 , n2988 );
nand ( n2990 , n2826 , n125 );
not ( n2991 , n2990 );
and ( n2992 , n2989 , n2991 );
nor ( n2993 , n2986 , n126 );
and ( n2994 , n2948 , n2993 );
nor ( n2995 , n2992 , n2994 );
nand ( n2996 , n2984 , n2995 );
nor ( n2997 , n2974 , n2996 );
not ( n2998 , n120 );
not ( n2999 , n2897 );
nand ( n3000 , n2999 , n2876 );
not ( n3001 , n3000 );
nand ( n3002 , n2965 , n2816 );
not ( n3003 , n3002 );
or ( n3004 , n3001 , n3003 );
nand ( n3005 , n3004 , n2942 );
not ( n3006 , n2865 );
not ( n3007 , n2900 );
nand ( n3008 , n3006 , n3007 );
not ( n3009 , n3008 );
and ( n3010 , n2814 , n122 );
nand ( n3011 , n3010 , n2843 );
not ( n3012 , n3011 );
or ( n3013 , n3009 , n3012 );
nand ( n3014 , n3013 , n2816 );
nand ( n3015 , n3005 , n3014 );
nand ( n3016 , n2998 , n3015 );
nand ( n3017 , n2945 , n2964 , n2997 , n3016 );
not ( n3018 , n3017 );
not ( n3019 , n3018 );
buf ( n3020 , n3019 );
not ( n3021 , n3020 );
not ( n3022 , n3021 );
not ( n3023 , n114 );
nand ( n3024 , n3023 , n112 );
not ( n3025 , n3024 );
nor ( n3026 , n113 , n115 );
nand ( n3027 , n3025 , n3026 );
nand ( n3028 , n113 , n114 );
not ( n3029 , n3028 );
nand ( n3030 , n3029 , n115 );
and ( n3031 , n3027 , n3030 , n118 );
not ( n3032 , n3031 );
not ( n3033 , n114 );
nor ( n3034 , n3033 , n113 );
nor ( n3035 , n112 , n116 );
and ( n3036 , n3034 , n3035 );
not ( n3037 , n115 );
nand ( n3038 , n3036 , n3037 );
not ( n3039 , n3038 );
or ( n3040 , n3032 , n3039 );
not ( n3041 , n117 );
nand ( n3042 , n3041 , n118 );
nand ( n3043 , n3040 , n3042 );
not ( n3044 , n3043 );
nand ( n3045 , n115 , n116 );
nor ( n3046 , n3045 , n114 );
nand ( n3047 , n112 , n113 );
not ( n3048 , n3047 );
nand ( n3049 , n3046 , n3048 );
not ( n3050 , n115 );
nand ( n3051 , n3050 , n116 );
not ( n3052 , n3051 );
not ( n3053 , n113 );
nand ( n3054 , n3053 , n112 );
not ( n3055 , n3054 );
nand ( n3056 , n3052 , n3055 );
nand ( n3057 , n3049 , n3056 );
not ( n3058 , n114 );
nor ( n3059 , n3058 , n115 );
not ( n3060 , n3059 );
not ( n3061 , n112 );
nand ( n3062 , n3060 , n3061 );
nor ( n3063 , n116 , n117 );
not ( n3064 , n3063 );
nor ( n3065 , n3062 , n3064 );
nor ( n3066 , n3057 , n3065 );
not ( n3067 , n3066 );
or ( n3068 , n3044 , n3067 );
not ( n3069 , n113 );
nand ( n3070 , n3069 , n115 );
not ( n3071 , n116 );
or ( n3072 , n3070 , n3071 );
not ( n3073 , n113 );
nor ( n3074 , n3073 , n112 );
nand ( n3075 , n3074 , n114 );
nand ( n3076 , n3072 , n3075 , n117 );
not ( n3077 , n3076 );
not ( n3078 , n117 );
not ( n3079 , n114 );
nand ( n3080 , n3079 , n113 );
not ( n3081 , n3080 );
nand ( n3082 , n3081 , n112 );
not ( n3083 , n3082 );
not ( n3084 , n116 );
nand ( n3085 , n3083 , n3084 );
nand ( n3086 , n3078 , n3085 );
not ( n3087 , n3086 );
or ( n3088 , n3077 , n3087 );
not ( n3089 , n114 );
nor ( n3090 , n3089 , n112 );
not ( n3091 , n3090 );
not ( n3092 , n3091 );
not ( n3093 , n3092 );
not ( n3094 , n117 );
and ( n3095 , n3026 , n3094 );
not ( n3096 , n3095 );
or ( n3097 , n3093 , n3096 );
nand ( n3098 , n115 , n116 );
nor ( n3099 , n3098 , n117 );
buf ( n3100 , n3074 );
nand ( n3101 , n3099 , n3100 );
nand ( n3102 , n3097 , n3101 );
not ( n3103 , n115 );
nor ( n3104 , n3103 , n113 );
nand ( n3105 , n3104 , n3025 );
not ( n3106 , n118 );
nand ( n3107 , n3105 , n3106 );
nor ( n3108 , n3102 , n3107 );
nand ( n3109 , n3088 , n3108 );
nand ( n3110 , n3068 , n3109 );
not ( n3111 , n116 );
nand ( n3112 , n3111 , n115 );
not ( n3113 , n114 );
nor ( n3114 , n3112 , n3113 );
not ( n3115 , n3114 );
not ( n3116 , n3115 );
nand ( n3117 , n3116 , n3055 );
not ( n3118 , n3030 );
nand ( n3119 , n3118 , n116 );
nand ( n3120 , n3117 , n3119 );
not ( n3121 , n115 );
nand ( n3122 , n3121 , n3074 );
nor ( n3123 , n3122 , n114 );
not ( n3124 , n3123 );
not ( n3125 , n116 );
nor ( n3126 , n3125 , n112 );
nor ( n3127 , n113 , n114 );
and ( n3128 , n3126 , n3127 );
not ( n3129 , n3128 );
and ( n3130 , n117 , n119 );
nand ( n3131 , n3124 , n3129 , n3130 );
or ( n3132 , n3120 , n3131 );
buf ( n3133 , n3025 );
not ( n3134 , n3112 );
nand ( n3135 , n3133 , n3134 );
nand ( n3136 , n3059 , n3048 );
not ( n3137 , n119 );
nor ( n3138 , n3137 , n117 );
nand ( n3139 , n3135 , n3136 , n3138 );
nand ( n3140 , n3132 , n3139 );
nand ( n3141 , n3110 , n3140 );
not ( n3142 , n117 );
nand ( n3143 , n3141 , n3142 );
buf ( n3144 , n3081 );
not ( n3145 , n115 );
nand ( n3146 , n3145 , n3126 );
or ( n3147 , n3144 , n3146 );
buf ( n3148 , n3034 );
nand ( n3149 , n3148 , n3126 );
nand ( n3150 , n3147 , n3149 );
not ( n3151 , n3134 );
nor ( n3152 , n112 , n114 );
and ( n3153 , n3152 , n115 );
not ( n3154 , n3153 );
nor ( n3155 , n3151 , n3154 );
nor ( n3156 , n3150 , n3155 );
not ( n3157 , n113 );
nand ( n3158 , n112 , n114 );
nor ( n3159 , n3157 , n3158 );
buf ( n3160 , n3159 );
nand ( n3161 , n3160 , n3134 );
and ( n3162 , n3156 , n3161 );
or ( n3163 , n3143 , n3162 );
not ( n3164 , n117 );
not ( n3165 , n3164 );
not ( n3166 , n3123 );
or ( n3167 , n3165 , n3166 );
not ( n3168 , n116 );
nand ( n3169 , n3168 , n117 );
nand ( n3170 , n3167 , n3169 );
nand ( n3171 , n3055 , n115 );
nand ( n3172 , n3171 , n3122 );
nand ( n3173 , n3170 , n3172 );
not ( n3174 , n3098 );
and ( n3175 , n3159 , n3174 );
not ( n3176 , n3175 );
and ( n3177 , n3176 , n118 );
and ( n3178 , n3173 , n3177 );
not ( n3179 , n112 );
nand ( n3180 , n3179 , n114 );
not ( n3181 , n116 );
nand ( n3182 , n3181 , n115 );
nor ( n3183 , n3180 , n3182 );
not ( n3184 , n3183 );
nor ( n3185 , n3184 , n113 );
not ( n3186 , n3099 );
nor ( n3187 , n3186 , n113 );
nor ( n3188 , n3185 , n3187 );
not ( n3189 , n116 );
nand ( n3190 , n3189 , n3127 );
not ( n3191 , n3190 );
nand ( n3192 , n3191 , n3037 );
nor ( n3193 , n112 , n113 );
buf ( n3194 , n3193 );
nand ( n3195 , n3052 , n3194 );
and ( n3196 , n3192 , n3195 , n3136 , n3106 );
not ( n3197 , n3082 );
nand ( n3198 , n116 , n117 );
not ( n3199 , n3198 );
nand ( n3200 , n3197 , n3199 );
and ( n3201 , n3188 , n3196 , n3200 );
or ( n3202 , n3178 , n3201 );
not ( n3203 , n115 );
buf ( n3204 , n3152 );
nand ( n3205 , n3203 , n3204 );
not ( n3206 , n3205 );
not ( n3207 , n3091 );
not ( n3208 , n3070 );
nand ( n3209 , n3207 , n3208 );
not ( n3210 , n3209 );
or ( n3211 , n3206 , n3210 );
not ( n3212 , n3169 );
nand ( n3213 , n3211 , n3212 );
and ( n3214 , n3213 , n3137 );
nand ( n3215 , n3202 , n3214 );
nand ( n3216 , n3141 , n3215 );
nand ( n3217 , n3163 , n3216 );
not ( n3218 , n118 );
nand ( n3219 , n3144 , n3052 );
nor ( n3220 , n3219 , n3061 );
nor ( n3221 , n3220 , n117 );
not ( n3222 , n3221 );
or ( n3223 , n3218 , n3222 );
and ( n3224 , n3153 , n113 );
not ( n3225 , n3224 );
nand ( n3226 , n3081 , n3071 );
not ( n3227 , n3226 );
nor ( n3228 , n113 , n114 );
and ( n3229 , n3228 , n112 );
nand ( n3230 , n3229 , n116 );
not ( n3231 , n3230 );
or ( n3232 , n3227 , n3231 );
nand ( n3233 , n3232 , n3037 );
nand ( n3234 , n117 , n118 );
not ( n3235 , n3234 );
nand ( n3236 , n3225 , n3233 , n3235 );
nand ( n3237 , n3223 , n3236 );
not ( n3238 , n3158 );
nand ( n3239 , n3026 , n3238 );
buf ( n3240 , n3239 );
and ( n3241 , n3219 , n3240 , n117 );
not ( n3242 , n3241 );
nor ( n3243 , n3075 , n3037 );
nor ( n3244 , n3243 , n117 );
nand ( n3245 , n3244 , n3230 , n3105 );
and ( n3246 , n3242 , n3245 );
nor ( n3247 , n115 , n116 );
and ( n3248 , n112 , n114 );
and ( n3249 , n3247 , n3248 );
nor ( n3250 , n3249 , n118 );
not ( n3251 , n113 );
nand ( n3252 , n3046 , n3251 );
nand ( n3253 , n3250 , n3252 );
nor ( n3254 , n3246 , n3253 );
or ( n3255 , n3237 , n3254 );
and ( n3256 , n3118 , n3126 );
buf ( n3257 , n3035 );
nand ( n3258 , n3144 , n3257 );
not ( n3259 , n3258 );
or ( n3260 , n3256 , n3259 );
not ( n3261 , n3122 );
or ( n3262 , n3261 , n117 );
nand ( n3263 , n3260 , n3262 );
not ( n3264 , n3263 );
not ( n3265 , n116 );
nor ( n3266 , n3265 , n117 );
not ( n3267 , n3266 );
nor ( n3268 , n3267 , n3105 );
nor ( n3269 , n3264 , n3268 );
nand ( n3270 , n3255 , n3269 );
nor ( n3271 , n3217 , n3270 );
not ( n3272 , n3271 );
not ( n3273 , n137 );
not ( n3274 , n2702 );
nand ( n3275 , n3274 , n2758 );
not ( n3276 , n3275 );
nand ( n3277 , n2550 , n2546 );
nand ( n3278 , n3277 , n144 );
and ( n3279 , n2646 , n140 );
nor ( n3280 , n3278 , n3279 );
not ( n3281 , n3280 );
or ( n3282 , n3276 , n3281 );
not ( n3283 , n141 );
nand ( n3284 , n3283 , n144 );
nand ( n3285 , n3282 , n3284 );
not ( n3286 , n3285 );
not ( n3287 , n2583 );
nor ( n3288 , n3287 , n138 );
or ( n3289 , n3286 , n3288 );
or ( n3290 , n3284 , n2733 );
nand ( n3291 , n3289 , n3290 );
not ( n3292 , n3291 );
nand ( n3293 , n2652 , n2762 );
and ( n3294 , n3293 , n2674 );
not ( n3295 , n3294 );
or ( n3296 , n3292 , n3295 );
and ( n3297 , n2630 , n138 );
nand ( n3298 , n3297 , n2517 );
nand ( n3299 , n3298 , n2668 );
not ( n3300 , n3299 );
nand ( n3301 , n2691 , n140 );
or ( n3302 , n3301 , n2595 );
not ( n3303 , n2678 );
and ( n3304 , n3303 , n142 );
not ( n3305 , n2532 );
nor ( n3306 , n3304 , n3305 );
nand ( n3307 , n3302 , n3306 );
not ( n3308 , n3307 );
and ( n3309 , n3300 , n3308 );
nand ( n3310 , n2682 , n143 );
nand ( n3311 , n2677 , n139 );
and ( n3312 , n3310 , n3311 , n2609 );
and ( n3313 , n3302 , n3312 );
nor ( n3314 , n3309 , n3313 );
nand ( n3315 , n3296 , n3314 );
nand ( n3316 , n2590 , n2720 );
nor ( n3317 , n3316 , n142 );
not ( n3318 , n3317 );
nand ( n3319 , n2648 , n2516 );
nand ( n3320 , n3319 , n141 );
not ( n3321 , n3320 );
buf ( n3322 , n2646 );
nand ( n3323 , n3322 , n2682 );
nand ( n3324 , n3318 , n3321 , n3323 , n2637 );
not ( n3325 , n2719 );
not ( n3326 , n3325 );
nand ( n3327 , n2558 , n2555 );
nand ( n3328 , n3326 , n3327 , n2686 );
nand ( n3329 , n3324 , n3328 );
nand ( n3330 , n3315 , n3329 );
not ( n3331 , n3330 );
or ( n3332 , n3273 , n3331 );
buf ( n3333 , n2599 );
not ( n3334 , n3333 );
not ( n3335 , n3334 );
nand ( n3336 , n2673 , n3335 );
nand ( n3337 , n3336 , n2559 );
and ( n3338 , n3337 , n141 );
not ( n3339 , n2745 );
not ( n3340 , n3339 );
nand ( n3341 , n3340 , n2682 );
nand ( n3342 , n2615 , n3341 , n2564 );
nor ( n3343 , n3338 , n3342 );
not ( n3344 , n3343 );
nand ( n3345 , n3279 , n2521 );
not ( n3346 , n3345 );
not ( n3347 , n3302 );
or ( n3348 , n3346 , n3347 , n2660 );
nand ( n3349 , n3348 , n2686 );
not ( n3350 , n3349 );
or ( n3351 , n3344 , n3350 );
nand ( n3352 , n2758 , n3333 );
nand ( n3353 , n2680 , n3352 , n144 );
nor ( n3354 , n2674 , n139 );
or ( n3355 , n3353 , n3354 );
nand ( n3356 , n3355 , n3284 );
and ( n3357 , n3297 , n2673 );
nand ( n3358 , n3357 , n2686 );
nand ( n3359 , n3356 , n3358 );
nand ( n3360 , n3351 , n3359 );
nand ( n3361 , n2540 , n2761 );
not ( n3362 , n3361 );
nand ( n3363 , n3362 , n2686 );
not ( n3364 , n2600 );
nand ( n3365 , n2571 , n2686 );
nor ( n3366 , n3364 , n3365 );
not ( n3367 , n2534 );
nand ( n3368 , n3367 , n140 );
and ( n3369 , n3366 , n3368 );
not ( n3370 , n2731 );
and ( n3371 , n3370 , n2585 );
nor ( n3372 , n3369 , n3371 );
and ( n3373 , n3363 , n3372 );
nor ( n3374 , n3373 , n137 );
not ( n3375 , n2639 );
not ( n3376 , n3346 );
or ( n3377 , n3375 , n3376 );
not ( n3378 , n2665 );
not ( n3379 , n142 );
nand ( n3380 , n3379 , n141 );
not ( n3381 , n3380 );
nand ( n3382 , n3378 , n3381 );
not ( n3383 , n3382 );
nor ( n3384 , n138 , n139 );
nand ( n3385 , n2614 , n3384 );
not ( n3386 , n3385 );
nand ( n3387 , n3386 , n2595 );
not ( n3388 , n3387 );
nor ( n3389 , n3383 , n3388 );
nand ( n3390 , n3377 , n3389 );
nand ( n3391 , n3347 , n2562 );
not ( n3392 , n3391 );
nor ( n3393 , n3374 , n3390 , n3392 );
nand ( n3394 , n3360 , n3393 );
nand ( n3395 , n2631 , n2639 );
not ( n3396 , n2518 );
or ( n3397 , n3396 , n2571 );
nand ( n3398 , n3397 , n2550 );
nand ( n3399 , n3327 , n2564 );
nor ( n3400 , n3310 , n141 );
nor ( n3401 , n3399 , n3400 );
and ( n3402 , n3395 , n3398 , n3401 );
not ( n3403 , n3402 );
nand ( n3404 , n3274 , n140 );
not ( n3405 , n3404 );
nand ( n3406 , n3405 , n2517 );
not ( n3407 , n3406 );
or ( n3408 , n3403 , n3407 );
not ( n3409 , n140 );
nor ( n3410 , n138 , n143 );
nand ( n3411 , n3409 , n3410 );
not ( n3412 , n3411 );
nand ( n3413 , n2590 , n140 );
not ( n3414 , n3413 );
or ( n3415 , n3412 , n3414 );
nand ( n3416 , n3415 , n3381 );
and ( n3417 , n2636 , n2618 );
nor ( n3418 , n3417 , n2564 );
and ( n3419 , n2683 , n3416 , n3418 );
nor ( n3420 , n3419 , n137 );
nand ( n3421 , n3408 , n3420 );
not ( n3422 , n3385 );
not ( n3423 , n3406 );
or ( n3424 , n3422 , n3423 );
nand ( n3425 , n2642 , n141 );
not ( n3426 , n3425 );
nand ( n3427 , n3424 , n3426 );
nand ( n3428 , n3421 , n3427 );
nor ( n3429 , n3394 , n3428 );
nand ( n3430 , n3332 , n3429 );
not ( n3431 , n3430 );
and ( n3432 , n3272 , n3431 );
not ( n3433 , n3272 );
and ( n3434 , n3433 , n3430 );
nor ( n3435 , n3432 , n3434 );
not ( n3436 , n3435 );
not ( n3437 , n3436 );
or ( n3438 , n3022 , n3437 );
or ( n3439 , n3021 , n3436 );
nand ( n3440 , n3438 , n3439 );
not ( n3441 , n3440 );
and ( n3442 , n2776 , n3441 );
not ( n3443 , n2776 );
and ( n3444 , n3443 , n3440 );
nor ( n3445 , n3442 , n3444 );
or ( n3446 , n3445 , n1 );
and ( n3447 , n237 , n2774 );
not ( n3448 , n237 );
and ( n3449 , n3448 , n236 );
nor ( n3450 , n3447 , n3449 );
or ( n3451 , n2246 , n3450 );
nand ( n3452 , n3446 , n3451 );
nor ( n3453 , n205 , n206 );
nand ( n3454 , n3453 , n207 );
not ( n3455 , n3454 );
nand ( n3456 , n208 , n210 );
not ( n3457 , n3456 );
nand ( n3458 , n3455 , n3457 );
not ( n3459 , n210 );
nand ( n3460 , n206 , n207 );
nor ( n3461 , n3459 , n3460 );
not ( n3462 , n208 );
nand ( n3463 , n3461 , n3462 );
and ( n3464 , n3458 , n3463 );
not ( n3465 , n205 );
nand ( n3466 , n3465 , n206 );
not ( n3467 , n3466 );
not ( n3468 , n207 );
nand ( n3469 , n3467 , n3468 );
nor ( n3470 , n3469 , n208 );
not ( n3471 , n209 );
nor ( n3472 , n3470 , n3471 );
not ( n3473 , n205 );
nand ( n3474 , n3473 , n207 );
not ( n3475 , n3474 );
not ( n3476 , n210 );
nand ( n3477 , n3476 , n208 );
not ( n3478 , n3477 );
nand ( n3479 , n3475 , n3478 );
not ( n3480 , n3479 );
nand ( n3481 , n3480 , n206 );
and ( n3482 , n3464 , n3472 , n3481 );
and ( n3483 , n207 , n205 , n206 );
nand ( n3484 , n3483 , n208 );
not ( n3485 , n209 );
nand ( n3486 , n3484 , n3485 );
not ( n3487 , n3478 );
not ( n3488 , n206 );
nand ( n3489 , n3488 , n207 );
nor ( n3490 , n3487 , n3489 );
nor ( n3491 , n3486 , n3490 );
or ( n3492 , n3482 , n3491 );
nor ( n3493 , n206 , n208 );
not ( n3494 , n3493 );
not ( n3495 , n3494 );
not ( n3496 , n205 );
nor ( n3497 , n3496 , n207 );
not ( n3498 , n3497 );
not ( n3499 , n3498 );
or ( n3500 , n3495 , n3499 );
not ( n3501 , n209 );
nand ( n3502 , n3501 , n210 );
not ( n3503 , n3502 );
nand ( n3504 , n3500 , n3503 );
not ( n3505 , n208 );
nand ( n3506 , n3505 , n210 );
nor ( n3507 , n3506 , n205 );
not ( n3508 , n207 );
nand ( n3509 , n3508 , n206 );
not ( n3510 , n3509 );
nand ( n3511 , n3507 , n3510 );
not ( n3512 , n210 );
not ( n3513 , n206 );
nand ( n3514 , n3512 , n3513 , n207 , n205 );
and ( n3515 , n3504 , n3511 , n3514 , n212 );
nand ( n3516 , n3492 , n3515 );
not ( n3517 , n207 );
nor ( n3518 , n205 , n206 );
nand ( n3519 , n3517 , n3518 );
not ( n3520 , n3519 );
not ( n3521 , n210 );
nand ( n3522 , n3521 , n209 );
not ( n3523 , n3522 );
nand ( n3524 , n3520 , n3523 );
not ( n3525 , n211 );
and ( n3526 , n3524 , n3525 );
nand ( n3527 , n206 , n208 );
not ( n3528 , n3527 );
nand ( n3529 , n3528 , n3497 );
not ( n3530 , n3529 );
not ( n3531 , n205 );
nor ( n3532 , n3531 , n206 );
nand ( n3533 , n3532 , n208 );
not ( n3534 , n3533 );
nand ( n3535 , n3534 , n207 );
not ( n3536 , n3535 );
or ( n3537 , n3530 , n3536 );
nand ( n3538 , n3537 , n209 );
not ( n3539 , n207 );
not ( n3540 , n3466 );
or ( n3541 , n3539 , n3540 );
not ( n3542 , n210 );
nor ( n3543 , n3542 , n208 );
nand ( n3544 , n3541 , n3543 );
nor ( n3545 , n208 , n210 );
not ( n3546 , n3489 );
nand ( n3547 , n3545 , n3546 );
nand ( n3548 , n3544 , n3547 );
not ( n3549 , n3527 );
nor ( n3550 , n205 , n207 );
nand ( n3551 , n3549 , n3550 );
nor ( n3552 , n209 , n210 );
not ( n3553 , n3552 );
nor ( n3554 , n3551 , n3553 );
nor ( n3555 , n3548 , n3554 );
and ( n3556 , n3526 , n3538 , n3555 );
nand ( n3557 , n205 , n207 );
not ( n3558 , n3557 );
not ( n3559 , n3558 );
not ( n3560 , n3471 );
or ( n3561 , n3559 , n3560 );
not ( n3562 , n205 );
nor ( n3563 , n3562 , n207 );
not ( n3564 , n206 );
nand ( n3565 , n3563 , n3564 );
not ( n3566 , n3565 );
nand ( n3567 , n3566 , n208 );
nand ( n3568 , n3561 , n3567 );
not ( n3569 , n3485 );
not ( n3570 , n3520 );
or ( n3571 , n3569 , n3570 );
nand ( n3572 , n3571 , n211 );
nor ( n3573 , n3568 , n3572 );
nor ( n3574 , n3556 , n3573 );
or ( n3575 , n3516 , n3574 );
not ( n3576 , n205 );
not ( n3577 , n3461 );
or ( n3578 , n3576 , n3577 );
nand ( n3579 , n3578 , n3481 );
not ( n3580 , n3550 );
nor ( n3581 , n208 , n210 );
not ( n3582 , n3581 );
nor ( n3583 , n3580 , n3582 );
or ( n3584 , n3579 , n3583 );
nand ( n3585 , n3584 , n3485 );
not ( n3586 , n3456 );
not ( n3587 , n3586 );
not ( n3588 , n3587 );
buf ( n3589 , n3518 );
not ( n3590 , n3589 );
or ( n3591 , n3588 , n3590 );
nand ( n3592 , n3591 , n211 );
nand ( n3593 , n205 , n210 );
nor ( n3594 , n3527 , n3593 );
nor ( n3595 , n3592 , n3594 );
not ( n3596 , n206 );
nand ( n3597 , n3596 , n205 );
not ( n3598 , n3597 );
and ( n3599 , n207 , n209 );
nand ( n3600 , n3598 , n3599 , n210 );
nand ( n3601 , n3595 , n3600 );
not ( n3602 , n3553 );
and ( n3603 , n3510 , n3602 );
or ( n3604 , n3601 , n3603 );
not ( n3605 , n210 );
not ( n3606 , n3605 );
not ( n3607 , n207 );
nor ( n3608 , n3607 , n208 );
nand ( n3609 , n205 , n206 );
not ( n3610 , n3609 );
nand ( n3611 , n3608 , n3610 );
not ( n3612 , n3498 );
not ( n3613 , n3493 );
not ( n3614 , n3613 );
nand ( n3615 , n3612 , n3614 );
nand ( n3616 , n3611 , n3615 );
not ( n3617 , n3616 );
or ( n3618 , n3606 , n3617 );
not ( n3619 , n211 );
not ( n3620 , n3619 );
not ( n3621 , n3456 );
nand ( n3622 , n3621 , n3453 );
not ( n3623 , n3622 );
or ( n3624 , n3620 , n3623 );
nand ( n3625 , n3619 , n209 );
nand ( n3626 , n3624 , n3625 );
nand ( n3627 , n3618 , n3626 );
nand ( n3628 , n3604 , n3627 );
nand ( n3629 , n209 , n210 );
not ( n3630 , n3629 );
not ( n3631 , n3630 );
nand ( n3632 , n3475 , n3614 );
not ( n3633 , n3632 );
not ( n3634 , n3633 );
or ( n3635 , n3631 , n3634 );
not ( n3636 , n3625 );
buf ( n3637 , n3460 );
not ( n3638 , n3637 );
and ( n3639 , n3636 , n3638 , n3593 );
nor ( n3640 , n3639 , n212 );
nand ( n3641 , n3635 , n3640 );
nand ( n3642 , n3563 , n3462 );
nor ( n3643 , n3642 , n3629 );
nor ( n3644 , n3641 , n3643 );
nand ( n3645 , n3585 , n3628 , n3644 );
nand ( n3646 , n3575 , n3645 );
nand ( n3647 , n3545 , n3558 );
and ( n3648 , n3647 , n209 );
not ( n3649 , n3648 );
nand ( n3650 , n3470 , n3605 );
not ( n3651 , n3650 );
or ( n3652 , n3649 , n3651 );
not ( n3653 , n3565 );
not ( n3654 , n3653 );
nand ( n3655 , n3533 , n3654 );
not ( n3656 , n3655 );
nand ( n3657 , n3632 , n3485 );
not ( n3658 , n3657 );
and ( n3659 , n3656 , n3658 );
nor ( n3660 , n3659 , n3503 );
nand ( n3661 , n3652 , n3660 );
not ( n3662 , n3661 );
nor ( n3663 , n3503 , n211 );
not ( n3664 , n3663 );
not ( n3665 , n3494 );
nand ( n3666 , n3665 , n3558 );
nand ( n3667 , n3666 , n3619 );
nand ( n3668 , n3664 , n3667 );
not ( n3669 , n205 );
nand ( n3670 , n3669 , n3586 );
not ( n3671 , n3670 );
nand ( n3672 , n3671 , n3564 , n3599 );
and ( n3673 , n3668 , n3672 );
not ( n3674 , n3673 );
or ( n3675 , n3662 , n3674 );
not ( n3676 , n207 );
nand ( n3677 , n3676 , n210 );
not ( n3678 , n3677 );
nand ( n3679 , n3467 , n3678 );
not ( n3680 , n3679 );
nand ( n3681 , n3680 , n209 );
not ( n3682 , n208 );
nand ( n3683 , n206 , n207 );
nor ( n3684 , n3682 , n3683 );
not ( n3685 , n3684 );
not ( n3686 , n3685 );
nand ( n3687 , n3686 , n3602 );
and ( n3688 , n3681 , n3687 , n211 );
not ( n3689 , n3518 );
not ( n3690 , n3689 );
nand ( n3691 , n3690 , n3581 );
not ( n3692 , n3691 );
nand ( n3693 , n3692 , n3468 );
not ( n3694 , n3567 );
not ( n3695 , n210 );
nand ( n3696 , n3695 , n209 );
not ( n3697 , n3696 );
nand ( n3698 , n3694 , n3697 );
and ( n3699 , n3455 , n3543 );
not ( n3700 , n3699 );
nand ( n3701 , n3688 , n3693 , n3698 , n3700 );
nand ( n3702 , n3675 , n3701 );
not ( n3703 , n209 );
nor ( n3704 , n3514 , n3703 );
or ( n3705 , n3704 , n3594 );
nand ( n3706 , n208 , n209 );
nand ( n3707 , n3705 , n3706 );
nand ( n3708 , n3646 , n3702 , n3707 );
not ( n3709 , n3708 );
not ( n3710 , n184 );
nor ( n3711 , n181 , n182 );
buf ( n3712 , n3711 );
nand ( n3713 , n3710 , n3712 );
nand ( n3714 , n3713 , n185 );
not ( n3715 , n180 );
nand ( n3716 , n3714 , n3715 );
nand ( n3717 , n181 , n182 );
nor ( n3718 , n3717 , n180 );
nand ( n3719 , n3718 , n183 );
not ( n3720 , n181 );
nand ( n3721 , n3720 , n180 , n182 );
not ( n3722 , n3721 );
nand ( n3723 , n3722 , n183 );
and ( n3724 , n3716 , n3719 , n3723 );
not ( n3725 , n184 );
nand ( n3726 , n3725 , n183 );
not ( n3727 , n3726 );
not ( n3728 , n182 );
nand ( n3729 , n3728 , n181 );
not ( n3730 , n3729 );
nand ( n3731 , n3727 , n3730 );
not ( n3732 , n185 );
and ( n3733 , n3731 , n3732 );
or ( n3734 , n3724 , n3733 );
not ( n3735 , n3715 );
not ( n3736 , n183 );
nand ( n3737 , n3736 , n184 );
not ( n3738 , n3737 );
not ( n3739 , n3738 );
or ( n3740 , n3735 , n3739 );
nand ( n3741 , n3738 , n3730 );
nand ( n3742 , n3740 , n3741 );
not ( n3743 , n181 );
nand ( n3744 , n3743 , n180 );
not ( n3745 , n3744 );
nor ( n3746 , n183 , n184 );
buf ( n3747 , n3746 );
nand ( n3748 , n3745 , n3747 );
not ( n3749 , n186 );
nand ( n3750 , n3748 , n3749 );
nor ( n3751 , n3742 , n3750 );
nand ( n3752 , n3734 , n3751 );
not ( n3753 , n180 );
nor ( n3754 , n181 , n182 );
nand ( n3755 , n3753 , n3754 );
nand ( n3756 , n180 , n182 );
buf ( n3757 , n3756 );
nand ( n3758 , n3755 , n3757 , n186 );
nand ( n3759 , n185 , n186 );
nand ( n3760 , n3758 , n3759 );
not ( n3761 , n182 );
nor ( n3762 , n3761 , n181 );
not ( n3763 , n180 );
and ( n3764 , n3762 , n3763 );
nand ( n3765 , n3764 , n183 );
nand ( n3766 , n3760 , n3765 );
nand ( n3767 , n3752 , n3766 );
not ( n3768 , n3767 );
not ( n3769 , n3726 );
not ( n3770 , n180 );
nor ( n3771 , n3770 , n182 );
nand ( n3772 , n3769 , n3771 );
not ( n3773 , n181 );
nor ( n3774 , n3772 , n3773 );
not ( n3775 , n182 );
nand ( n3776 , n183 , n184 );
not ( n3777 , n3776 );
nand ( n3778 , n3775 , n3777 );
nor ( n3779 , n3744 , n3778 );
nor ( n3780 , n3774 , n3779 );
not ( n3781 , n3780 );
nand ( n3782 , n185 , n187 );
not ( n3783 , n3782 );
not ( n3784 , n184 );
nor ( n3785 , n3784 , n183 );
nand ( n3786 , n180 , n181 );
not ( n3787 , n3786 );
nand ( n3788 , n3785 , n3787 );
nand ( n3789 , n3783 , n3788 );
nor ( n3790 , n3729 , n183 );
and ( n3791 , n3790 , n3715 );
nor ( n3792 , n3789 , n3791 );
not ( n3793 , n3792 );
or ( n3794 , n3781 , n3793 );
not ( n3795 , n181 );
not ( n3796 , n3795 );
not ( n3797 , n3738 );
or ( n3798 , n3796 , n3797 );
nand ( n3799 , n3798 , n187 );
not ( n3800 , n3799 );
not ( n3801 , n184 );
nand ( n3802 , n3801 , n183 );
not ( n3803 , n3802 );
not ( n3804 , n181 );
nand ( n3805 , n3804 , n180 );
not ( n3806 , n3805 );
nand ( n3807 , n3803 , n3806 );
not ( n3808 , n182 );
nor ( n3809 , n3808 , n180 );
nand ( n3810 , n3809 , n184 );
not ( n3811 , n185 );
and ( n3812 , n3810 , n3811 );
not ( n3813 , n183 );
nor ( n3814 , n3813 , n3756 );
nand ( n3815 , n3814 , n181 );
nand ( n3816 , n3800 , n3807 , n3812 , n3815 );
nand ( n3817 , n3794 , n3816 );
not ( n3818 , n182 );
nand ( n3819 , n3818 , n181 , n3715 );
buf ( n3820 , n3819 );
not ( n3821 , n3738 );
nor ( n3822 , n3820 , n3821 );
or ( n3823 , n181 , n184 );
nor ( n3824 , n3757 , n3823 );
nor ( n3825 , n3822 , n3824 );
and ( n3826 , n3817 , n3825 );
not ( n3827 , n3826 );
or ( n3828 , n3768 , n3827 );
nor ( n3829 , n180 , n182 );
nand ( n3830 , n3829 , n3747 );
not ( n3831 , n3830 );
nand ( n3832 , n181 , n182 );
not ( n3833 , n3832 );
nand ( n3834 , n3833 , n184 );
not ( n3835 , n3834 );
not ( n3836 , n3715 );
and ( n3837 , n3835 , n3836 );
nor ( n3838 , n3837 , n3774 );
not ( n3839 , n3838 );
or ( n3840 , n3831 , n3839 );
nand ( n3841 , n3840 , n3811 );
nand ( n3842 , n3754 , n180 );
buf ( n3843 , n3842 );
not ( n3844 , n180 );
and ( n3845 , n3844 , n182 );
not ( n3846 , n3845 );
nand ( n3847 , n3843 , n3846 );
nand ( n3848 , n184 , n185 );
nor ( n3849 , n3848 , n183 );
and ( n3850 , n3847 , n3849 );
nor ( n3851 , n3850 , n187 );
and ( n3852 , n3841 , n3851 );
nor ( n3853 , n3715 , n3717 );
not ( n3854 , n184 );
nand ( n3855 , n3853 , n3854 );
nand ( n3856 , n3730 , n180 );
and ( n3857 , n3855 , n3856 , n3749 );
nor ( n3858 , n185 , n186 );
or ( n3859 , n3857 , n3858 );
nand ( n3860 , n183 , n184 );
not ( n3861 , n3860 );
nand ( n3862 , n3861 , n3712 );
not ( n3863 , n3862 );
nand ( n3864 , n3863 , n3732 );
nand ( n3865 , n3859 , n3864 );
not ( n3866 , n181 );
nand ( n3867 , n3866 , n182 );
nor ( n3868 , n3867 , n183 );
nand ( n3869 , n3868 , n3715 );
not ( n3870 , n3786 );
not ( n3871 , n182 );
nor ( n3872 , n3871 , n183 );
nand ( n3873 , n3870 , n3872 );
nand ( n3874 , n3869 , n3873 );
not ( n3875 , n3874 );
nor ( n3876 , n3875 , n184 );
or ( n3877 , n3865 , n3876 );
not ( n3878 , n3721 );
buf ( n3879 , n3878 );
not ( n3880 , n3848 );
nand ( n3881 , n3879 , n3880 );
and ( n3882 , n3777 , n3833 );
not ( n3883 , n3777 );
and ( n3884 , n3883 , n3712 );
nor ( n3885 , n3882 , n3884 );
not ( n3886 , n181 );
nor ( n3887 , n3886 , n180 );
nor ( n3888 , n184 , n185 );
nand ( n3889 , n3887 , n3888 );
nand ( n3890 , n3881 , n3885 , n3889 , n186 );
nand ( n3891 , n3877 , n3890 );
nand ( n3892 , n3852 , n3891 );
nand ( n3893 , n3828 , n3892 );
not ( n3894 , n181 );
nand ( n3895 , n3894 , n3746 );
not ( n3896 , n3895 );
not ( n3897 , n180 );
nor ( n3898 , n3897 , n182 );
nand ( n3899 , n3896 , n3898 );
nand ( n3900 , n3899 , n3732 );
nand ( n3901 , n3745 , n3872 );
nor ( n3902 , n3901 , n3854 );
nor ( n3903 , n3900 , n3902 );
not ( n3904 , n3895 );
nand ( n3905 , n3904 , n3845 );
not ( n3906 , n3905 );
not ( n3907 , n182 );
nor ( n3908 , n3907 , n181 );
nand ( n3909 , n3803 , n3908 );
not ( n3910 , n3909 );
nor ( n3911 , n3906 , n3910 );
and ( n3912 , n3903 , n3911 );
nand ( n3913 , n3791 , n3854 );
nand ( n3914 , n3913 , n185 );
not ( n3915 , n183 );
nand ( n3916 , n3915 , n3854 );
nor ( n3917 , n3757 , n3916 );
nor ( n3918 , n3914 , n3917 );
or ( n3919 , n3912 , n3918 );
not ( n3920 , n3842 );
nand ( n3921 , n3920 , n183 );
nand ( n3922 , n184 , n185 );
nor ( n3923 , n3921 , n3922 );
nor ( n3924 , n3923 , n186 );
nand ( n3925 , n3919 , n3924 );
not ( n3926 , n181 );
nand ( n3927 , n3727 , n3926 );
nor ( n3928 , n3927 , n3846 );
not ( n3929 , n3928 );
not ( n3930 , n3929 );
or ( n3931 , n3819 , n3854 );
not ( n3932 , n3931 );
or ( n3933 , n3930 , n3932 );
nand ( n3934 , n3933 , n185 );
nand ( n3935 , n3738 , n3898 );
not ( n3936 , n3935 );
not ( n3937 , n181 );
and ( n3938 , n3936 , n3937 );
nor ( n3939 , n3938 , n3749 );
not ( n3940 , n3755 );
nand ( n3941 , n3940 , n3747 );
not ( n3942 , n3726 );
nand ( n3943 , n3942 , n3787 );
or ( n3944 , n3943 , n185 );
nand ( n3945 , n3934 , n3939 , n3941 , n3944 );
nand ( n3946 , n3925 , n3945 );
not ( n3947 , n184 );
nand ( n3948 , n3947 , n185 );
not ( n3949 , n3948 );
or ( n3950 , n3949 , n3833 );
not ( n3951 , n3732 );
and ( n3952 , n184 , n181 , n183 );
not ( n3953 , n3952 );
or ( n3954 , n3951 , n3953 );
nand ( n3955 , n3954 , n3901 );
nand ( n3956 , n3950 , n3955 );
and ( n3957 , n3893 , n3946 , n3956 );
and ( n3958 , n3709 , n3957 );
not ( n3959 , n3709 );
not ( n3960 , n3957 );
and ( n3961 , n3959 , n3960 );
nor ( n3962 , n3958 , n3961 );
not ( n3963 , n3962 );
not ( n3964 , n197 );
nand ( n3965 , n3964 , n200 );
not ( n3966 , n3965 );
nand ( n3967 , n3966 , n198 );
not ( n3968 , n3967 );
not ( n3969 , n201 );
nand ( n3970 , n3969 , n199 );
buf ( n3971 , n3970 );
not ( n3972 , n3971 );
nand ( n3973 , n3968 , n3972 );
not ( n3974 , n198 );
nand ( n3975 , n197 , n200 );
nor ( n3976 , n3974 , n3975 );
not ( n3977 , n201 );
nor ( n3978 , n3977 , n199 );
and ( n3979 , n3976 , n3978 );
not ( n3980 , n3979 );
nand ( n3981 , n3973 , n3980 );
not ( n3982 , n3981 );
not ( n3983 , n3982 );
not ( n3984 , n3965 );
buf ( n3985 , n3984 );
not ( n3986 , n201 );
and ( n3987 , n3985 , n3986 );
not ( n3988 , n198 );
nand ( n3989 , n3988 , n197 );
not ( n3990 , n3989 );
nand ( n3991 , n199 , n201 );
not ( n3992 , n3991 );
nand ( n3993 , n3990 , n3992 );
not ( n3994 , n3993 );
nor ( n3995 , n197 , n198 );
not ( n3996 , n199 );
and ( n3997 , n3995 , n3996 );
nor ( n3998 , n3987 , n3994 , n3997 );
not ( n3999 , n3998 );
not ( n4000 , n200 );
nand ( n4001 , n4000 , n198 );
not ( n4002 , n4001 );
nand ( n4003 , n4002 , n197 );
not ( n4004 , n4003 );
nand ( n4005 , n4004 , n201 );
not ( n4006 , n199 );
nand ( n4007 , n4006 , n197 );
not ( n4008 , n200 );
nand ( n4009 , n4008 , n201 );
or ( n4010 , n4007 , n4009 );
nand ( n4011 , n4005 , n4010 );
not ( n4012 , n198 );
nand ( n4013 , n4012 , n201 );
not ( n4014 , n4013 );
nor ( n4015 , n197 , n200 );
buf ( n4016 , n4015 );
nand ( n4017 , n4014 , n4016 );
nand ( n4018 , n4017 , n203 );
nor ( n4019 , n4011 , n4018 );
not ( n4020 , n4019 );
or ( n4021 , n3999 , n4020 );
not ( n4022 , n199 );
nand ( n4023 , n4022 , n200 );
not ( n4024 , n4023 );
nor ( n4025 , n198 , n201 );
nand ( n4026 , n4024 , n4025 );
not ( n4027 , n197 );
nor ( n4028 , n4026 , n4027 );
not ( n4029 , n4028 );
nor ( n4030 , n3993 , n200 );
nor ( n4031 , n4030 , n3979 , n203 );
not ( n4032 , n200 );
nand ( n4033 , n4032 , n197 );
nor ( n4034 , n4033 , n3996 );
buf ( n4035 , n4034 );
not ( n4036 , n198 );
nand ( n4037 , n4035 , n4036 );
nand ( n4038 , n4029 , n4031 , n4037 );
nand ( n4039 , n4021 , n4038 );
not ( n4040 , n4039 );
or ( n4041 , n3983 , n4040 );
buf ( n4042 , n4019 );
buf ( n4043 , n4031 );
or ( n4044 , n4042 , n4043 );
nand ( n4045 , n4044 , n202 );
nand ( n4046 , n4041 , n4045 );
not ( n4047 , n200 );
nand ( n4048 , n3995 , n4047 );
not ( n4049 , n4048 );
not ( n4050 , n202 );
nor ( n4051 , n4050 , n201 );
nand ( n4052 , n4049 , n4051 );
nor ( n4053 , n199 , n201 );
and ( n4054 , n4015 , n4053 );
not ( n4055 , n4054 );
nor ( n4056 , n199 , n200 );
nand ( n4057 , n4051 , n4056 );
not ( n4058 , n204 );
and ( n4059 , n4052 , n4055 , n4057 , n4058 );
not ( n4060 , n4013 );
not ( n4061 , n3975 );
nand ( n4062 , n4060 , n4061 );
not ( n4063 , n4062 );
nand ( n4064 , n4004 , n3986 );
not ( n4065 , n4064 );
or ( n4066 , n4063 , n4065 );
not ( n4067 , n203 );
and ( n4068 , n4067 , n202 );
nand ( n4069 , n4066 , n4068 );
nand ( n4070 , n4061 , n198 );
nor ( n4071 , n4070 , n201 );
nand ( n4072 , n198 , n200 );
not ( n4073 , n4072 );
not ( n4074 , n4073 );
nor ( n4075 , n4074 , n3996 );
or ( n4076 , n4071 , n4075 );
nand ( n4077 , n202 , n203 );
not ( n4078 , n4077 );
nand ( n4079 , n4076 , n4078 );
not ( n4080 , n197 );
nand ( n4081 , n4080 , n198 );
nor ( n4082 , n4081 , n200 );
not ( n4083 , n4082 );
not ( n4084 , n4083 );
nand ( n4085 , n199 , n202 );
not ( n4086 , n4085 );
and ( n4087 , n4086 , n201 );
nand ( n4088 , n4084 , n4087 );
and ( n4089 , n4059 , n4069 , n4079 , n4088 );
nand ( n4090 , n4046 , n4089 );
not ( n4091 , n197 );
nor ( n4092 , n199 , n201 );
nand ( n4093 , n4091 , n4092 , n4073 );
not ( n4094 , n4093 );
and ( n4095 , n4061 , n201 );
not ( n4096 , n3992 );
nor ( n4097 , n198 , n200 );
nor ( n4098 , n4095 , n4096 , n4097 );
nor ( n4099 , n4094 , n4098 );
not ( n4100 , n3989 );
nor ( n4101 , n199 , n200 );
nand ( n4102 , n4100 , n4101 );
not ( n4103 , n4102 );
nor ( n4104 , n4103 , n203 );
not ( n4105 , n202 );
nand ( n4106 , n4105 , n201 );
not ( n4107 , n4106 );
nand ( n4108 , n3985 , n4107 );
nand ( n4109 , n4099 , n4104 , n4108 );
and ( n4110 , n199 , n3989 );
not ( n4111 , n199 );
not ( n4112 , n198 );
nand ( n4113 , n4112 , n200 );
not ( n4114 , n4113 );
not ( n4115 , n4114 );
and ( n4116 , n4111 , n4115 );
nor ( n4117 , n4110 , n4116 );
nor ( n4118 , n4117 , n4067 , n4095 );
not ( n4119 , n202 );
nand ( n4120 , n4119 , n203 );
not ( n4121 , n4120 );
or ( n4122 , n4118 , n4121 );
nand ( n4123 , n199 , n201 );
nand ( n4124 , n197 , n198 );
nor ( n4125 , n4123 , n4124 );
nand ( n4126 , n4125 , n200 );
not ( n4127 , n4023 );
nand ( n4128 , n3990 , n4127 );
and ( n4129 , n4126 , n4128 );
nand ( n4130 , n4122 , n4129 );
nand ( n4131 , n4109 , n4130 );
and ( n4132 , n4015 , n199 );
nand ( n4133 , n4132 , n198 );
not ( n4134 , n201 );
nor ( n4135 , n4134 , n197 );
nand ( n4136 , n4135 , n4073 );
nor ( n4137 , n4058 , n202 );
nand ( n4138 , n4133 , n4136 , n4102 , n4137 );
not ( n4139 , n4064 );
or ( n4140 , n4138 , n4139 );
nand ( n4141 , n4061 , n4025 );
nand ( n4142 , n4141 , n202 );
or ( n4143 , n4142 , n4058 );
nand ( n4144 , n4140 , n4143 );
and ( n4145 , n4082 , n3986 );
and ( n4146 , n4145 , n199 );
not ( n4147 , n198 );
not ( n4148 , n201 );
nand ( n4149 , n4147 , n4148 , n199 , n200 );
not ( n4150 , n4149 );
nand ( n4151 , n4150 , n197 );
not ( n4152 , n4151 );
nor ( n4153 , n4146 , n4152 );
nand ( n4154 , n4131 , n4144 , n4153 );
nand ( n4155 , n4090 , n4154 );
not ( n4156 , n3971 );
nand ( n4157 , n4049 , n4156 );
not ( n4158 , n4033 );
nand ( n4159 , n4060 , n4158 );
not ( n4160 , n202 );
and ( n4161 , n4159 , n4160 );
nand ( n4162 , n4157 , n4161 );
not ( n4163 , n4123 );
and ( n4164 , n4163 , n4027 );
not ( n4165 , n4002 );
not ( n4166 , n4165 );
nand ( n4167 , n4164 , n4166 );
not ( n4168 , n201 );
nand ( n4169 , n198 , n200 );
nor ( n4170 , n4168 , n4169 );
nand ( n4171 , n4170 , n3996 );
nand ( n4172 , n4167 , n4171 );
nor ( n4173 , n4162 , n4172 );
not ( n4174 , n202 );
nor ( n4175 , n198 , n197 );
nand ( n4176 , n4175 , n200 );
not ( n4177 , n4176 );
or ( n4178 , n4174 , n4177 );
nand ( n4179 , n201 , n202 );
nand ( n4180 , n4178 , n4179 );
nor ( n4181 , n3970 , n4169 );
nand ( n4182 , n4181 , n197 );
and ( n4183 , n4180 , n4182 , n4167 , n4055 );
or ( n4184 , n4173 , n4183 );
not ( n4185 , n4115 );
nand ( n4186 , n4164 , n4185 );
nand ( n4187 , n4184 , n4186 );
not ( n4188 , n4187 );
not ( n4189 , n4067 );
or ( n4190 , n4188 , n4189 );
nand ( n4191 , n3997 , n4047 );
not ( n4192 , n4124 );
nand ( n4193 , n4101 , n4192 );
and ( n4194 , n4017 , n4193 );
not ( n4195 , n4145 );
nand ( n4196 , n4191 , n4093 , n4194 , n4195 );
and ( n4197 , n4196 , n4121 );
not ( n4198 , n4128 );
nand ( n4199 , n4198 , n201 );
not ( n4200 , n4125 );
nand ( n4201 , n4151 , n4199 , n4200 );
and ( n4202 , n4201 , n4078 );
nor ( n4203 , n4197 , n4202 );
nand ( n4204 , n4190 , n4203 );
nor ( n4205 , n4191 , n4179 );
not ( n4206 , n4205 );
not ( n4207 , n4176 );
nand ( n4208 , n4207 , n4087 );
nand ( n4209 , n4206 , n4208 );
nor ( n4210 , n4204 , n4209 );
nand ( n4211 , n4155 , n4210 );
not ( n4212 , n3519 );
nand ( n4213 , n4212 , n208 );
and ( n4214 , n205 , n210 );
nand ( n4215 , n3546 , n4214 );
not ( n4216 , n4215 );
nand ( n4217 , n4216 , n208 );
nand ( n4218 , n4213 , n4217 );
and ( n4219 , n4218 , n3471 );
not ( n4220 , n3454 );
nand ( n4221 , n4220 , n208 );
not ( n4222 , n3484 );
nor ( n4223 , n205 , n207 );
not ( n4224 , n4223 );
nor ( n4225 , n4224 , n3613 );
nor ( n4226 , n4222 , n4225 );
and ( n4227 , n4221 , n4226 );
nor ( n4228 , n4227 , n3629 );
not ( n4229 , n3483 );
not ( n4230 , n4229 );
and ( n4231 , n3493 , n207 );
not ( n4232 , n4231 );
not ( n4233 , n4232 );
or ( n4234 , n4230 , n4233 );
nand ( n4235 , n4234 , n3552 );
not ( n4236 , n212 );
nand ( n4237 , n4235 , n4236 );
nor ( n4238 , n4219 , n4228 , n4237 );
not ( n4239 , n4238 );
not ( n4240 , n3669 );
nor ( n4241 , n4240 , n3683 );
nand ( n4242 , n4241 , n210 );
nand ( n4243 , n4242 , n211 );
not ( n4244 , n4243 );
not ( n4245 , n3670 );
not ( n4246 , n3597 );
nand ( n4247 , n4246 , n3678 );
not ( n4248 , n4247 );
or ( n4249 , n4245 , n4248 );
nand ( n4250 , n4249 , n3485 );
not ( n4251 , n3529 );
nand ( n4252 , n4251 , n3605 );
nand ( n4253 , n4244 , n3698 , n4250 , n4252 );
nand ( n4254 , n3519 , n3525 );
nand ( n4255 , n3510 , n208 );
nor ( n4256 , n4255 , n3605 );
nor ( n4257 , n4254 , n4256 );
nor ( n4258 , n209 , n211 );
or ( n4259 , n4257 , n4258 );
not ( n4260 , n3463 );
not ( n4261 , n206 );
nor ( n4262 , n4261 , n208 );
and ( n4263 , n4262 , n3485 );
nor ( n4264 , n4260 , n4263 );
nand ( n4265 , n4259 , n4264 );
nand ( n4266 , n4253 , n4265 );
not ( n4267 , n4266 );
or ( n4268 , n4239 , n4267 );
and ( n4269 , n210 , n3597 );
not ( n4270 , n210 );
and ( n4271 , n4270 , n3689 );
nor ( n4272 , n4269 , n4271 );
nand ( n4273 , n4223 , n208 );
not ( n4274 , n208 );
nand ( n4275 , n4274 , n205 );
nand ( n4276 , n4273 , n4275 );
nor ( n4277 , n4272 , n4276 );
not ( n4278 , n4277 );
nand ( n4279 , n3605 , n3608 , n3610 );
nand ( n4280 , n3532 , n207 , n208 );
and ( n4281 , n3479 , n4279 , n4280 );
not ( n4282 , n4281 );
or ( n4283 , n4278 , n4282 );
nand ( n4284 , n4283 , n209 );
not ( n4285 , n3469 );
not ( n4286 , n3533 );
or ( n4287 , n4285 , n4286 );
nand ( n4288 , n4287 , n3552 );
not ( n4289 , n4288 );
not ( n4290 , n210 );
not ( n4291 , n4251 );
or ( n4292 , n4290 , n4291 );
nand ( n4293 , n4292 , n211 );
nor ( n4294 , n4289 , n4293 );
nand ( n4295 , n4284 , n4294 );
and ( n4296 , n3510 , n3545 );
nor ( n4297 , n4296 , n3471 );
not ( n4298 , n4297 );
not ( n4299 , n4281 );
or ( n4300 , n4298 , n4299 );
nand ( n4301 , n3533 , n3484 , n4273 , n3485 );
nand ( n4302 , n4300 , n4301 );
nand ( n4303 , n3475 , n3543 );
not ( n4304 , n209 );
nand ( n4305 , n3564 , n3558 , n4304 );
not ( n4306 , n3597 );
nand ( n4307 , n4306 , n3552 );
nand ( n4308 , n4303 , n4305 , n4307 , n3525 );
and ( n4309 , n3534 , n3523 );
nor ( n4310 , n4308 , n4309 );
nand ( n4311 , n4302 , n4310 );
nand ( n4312 , n4295 , n4311 );
not ( n4313 , n3490 );
nand ( n4314 , n4313 , n212 );
nor ( n4315 , n3643 , n4314 );
nand ( n4316 , n4312 , n4315 );
nand ( n4317 , n4268 , n4316 );
not ( n4318 , n4262 );
and ( n4319 , n3475 , n4318 );
or ( n4320 , n3616 , n4319 );
nand ( n4321 , n4320 , n3503 );
and ( n4322 , n3633 , n3697 );
nor ( n4323 , n4322 , n3525 );
nand ( n4324 , n4321 , n4323 );
nor ( n4325 , n208 , n3509 );
and ( n4326 , n4325 , n205 );
or ( n4327 , n4326 , n4216 );
nand ( n4328 , n4327 , n209 );
nand ( n4329 , n4276 , n3697 , n206 );
nand ( n4330 , n4328 , n4329 );
nor ( n4331 , n4324 , n4330 );
not ( n4332 , n211 );
nand ( n4333 , n3558 , n208 );
nor ( n4334 , n4333 , n3522 );
not ( n4335 , n4334 );
not ( n4336 , n3529 );
nand ( n4337 , n4336 , n3630 );
not ( n4338 , n3460 );
nand ( n4339 , n3478 , n4338 );
buf ( n4340 , n4339 );
nand ( n4341 , n4332 , n4335 , n4337 , n4340 );
not ( n4342 , n209 );
not ( n4343 , n3589 );
or ( n4344 , n4342 , n4343 );
not ( n4345 , n4263 );
nand ( n4346 , n4344 , n4345 );
nand ( n4347 , n4346 , n3678 );
nand ( n4348 , n4235 , n4347 );
nor ( n4349 , n4341 , n4348 );
nor ( n4350 , n4331 , n4349 );
not ( n4351 , n3503 );
not ( n4352 , n4213 );
not ( n4353 , n4352 );
or ( n4354 , n4351 , n4353 );
not ( n4355 , n205 );
nor ( n4356 , n4355 , n210 );
and ( n4357 , n4231 , n4356 );
nand ( n4358 , n4357 , n3485 );
nand ( n4359 , n4354 , n4358 );
nor ( n4360 , n4350 , n4359 );
nand ( n4361 , n4317 , n4360 );
not ( n4362 , n4361 );
not ( n4363 , n4362 );
and ( n4364 , n4211 , n4363 );
not ( n4365 , n4211 );
not ( n4366 , n4362 );
not ( n4367 , n4366 );
and ( n4368 , n4365 , n4367 );
nor ( n4369 , n4364 , n4368 );
not ( n4370 , n4369 );
not ( n4371 , n4370 );
or ( n4372 , n3963 , n4371 );
not ( n4373 , n3962 );
nand ( n4374 , n4369 , n4373 );
nand ( n4375 , n4372 , n4374 );
not ( n4376 , n294 );
not ( n4377 , n4376 );
not ( n4378 , n192 );
nor ( n4379 , n4378 , n193 );
not ( n4380 , n4379 );
nor ( n4381 , n188 , n189 );
not ( n4382 , n190 );
and ( n4383 , n4381 , n4382 );
not ( n4384 , n4383 );
nor ( n4385 , n4384 , n191 );
nand ( n4386 , n4380 , n4385 );
not ( n4387 , n188 );
nand ( n4388 , n4387 , n189 , n192 );
nor ( n4389 , n4388 , n4382 );
not ( n4390 , n193 );
nand ( n4391 , n4389 , n4390 );
not ( n4392 , n4391 );
not ( n4393 , n191 );
nand ( n4394 , n4392 , n4393 );
not ( n4395 , n193 );
nor ( n4396 , n4395 , n192 );
and ( n4397 , n4396 , n4393 );
nand ( n4398 , n4397 , n4382 );
and ( n4399 , n4386 , n4394 , n4398 );
nor ( n4400 , n188 , n190 );
nand ( n4401 , n4400 , n4393 );
not ( n4402 , n4401 );
not ( n4403 , n189 );
nor ( n4404 , n4403 , n192 );
nand ( n4405 , n4402 , n4404 );
not ( n4406 , n192 );
nand ( n4407 , n188 , n190 );
not ( n4408 , n4407 );
nand ( n4409 , n4406 , n189 , n4408 );
not ( n4410 , n4409 );
not ( n4411 , n193 );
nand ( n4412 , n4411 , n191 );
not ( n4413 , n4412 );
nand ( n4414 , n4410 , n4413 );
not ( n4415 , n195 );
and ( n4416 , n4405 , n4414 , n4415 );
nand ( n4417 , n191 , n193 );
nor ( n4418 , n4388 , n4417 );
nand ( n4419 , n4418 , n4382 );
nand ( n4420 , n4399 , n4416 , n4419 );
not ( n4421 , n188 );
nor ( n4422 , n4421 , n190 );
buf ( n4423 , n4422 );
not ( n4424 , n4423 );
not ( n4425 , n4424 );
nand ( n4426 , n191 , n192 );
not ( n4427 , n4426 );
nand ( n4428 , n4425 , n4427 );
not ( n4429 , n4428 );
not ( n4430 , n189 );
nand ( n4431 , n4429 , n4430 );
nand ( n4432 , n188 , n189 );
or ( n4433 , n4432 , n190 );
not ( n4434 , n4433 );
not ( n4435 , n191 );
nand ( n4436 , n4435 , n193 );
not ( n4437 , n4436 );
nand ( n4438 , n4434 , n4437 );
nand ( n4439 , n4410 , n191 );
and ( n4440 , n4431 , n4438 , n4439 );
and ( n4441 , n4422 , n192 );
nand ( n4442 , n4441 , n4430 );
not ( n4443 , n189 );
nand ( n4444 , n4443 , n188 , n190 );
nor ( n4445 , n191 , n192 );
not ( n4446 , n4445 );
nor ( n4447 , n4444 , n4446 );
nor ( n4448 , n4447 , n194 );
nand ( n4449 , n4442 , n4448 );
not ( n4450 , n193 );
nor ( n4451 , n4450 , n194 );
not ( n4452 , n4451 );
and ( n4453 , n4449 , n4452 );
not ( n4454 , n4444 );
not ( n4455 , n4454 );
nor ( n4456 , n4455 , n4417 );
nor ( n4457 , n4453 , n4456 );
and ( n4458 , n4440 , n4457 );
not ( n4459 , n190 );
nor ( n4460 , n4459 , n188 );
not ( n4461 , n4460 );
not ( n4462 , n4461 );
nand ( n4463 , n4393 , n4462 );
not ( n4464 , n4463 );
not ( n4465 , n192 );
not ( n4466 , n4381 );
not ( n4467 , n4466 );
nand ( n4468 , n4465 , n4467 );
not ( n4469 , n4468 );
or ( n4470 , n4464 , n4469 );
nand ( n4471 , n4470 , n4390 );
nand ( n4472 , n188 , n191 );
not ( n4473 , n4472 );
nor ( n4474 , n190 , n192 );
nand ( n4475 , n4473 , n4474 );
not ( n4476 , n4472 );
not ( n4477 , n190 );
nand ( n4478 , n4477 , n189 );
not ( n4479 , n4478 );
nand ( n4480 , n4476 , n4479 );
nand ( n4481 , n4475 , n4480 );
not ( n4482 , n4481 );
nand ( n4483 , n4471 , n4482 , n194 );
not ( n4484 , n4413 );
not ( n4485 , n188 );
nor ( n4486 , n4485 , n189 );
nand ( n4487 , n4486 , n192 );
not ( n4488 , n4487 );
not ( n4489 , n4488 );
or ( n4490 , n4484 , n4489 );
buf ( n4491 , n4381 );
nand ( n4492 , n4491 , n191 );
nor ( n4493 , n4492 , n190 );
and ( n4494 , n192 , n193 );
nand ( n4495 , n189 , n190 );
not ( n4496 , n4495 );
and ( n4497 , n4494 , n4496 );
nor ( n4498 , n4493 , n4497 );
nand ( n4499 , n4490 , n4498 );
not ( n4500 , n4407 );
nand ( n4501 , n4500 , n189 );
not ( n4502 , n4501 );
buf ( n4503 , n4445 );
nand ( n4504 , n4502 , n4503 );
nor ( n4505 , n4504 , n4390 );
nor ( n4506 , n4483 , n4499 , n4505 );
nor ( n4507 , n4458 , n4506 );
or ( n4508 , n4420 , n4507 );
and ( n4509 , n4400 , n189 );
nand ( n4510 , n4509 , n192 );
not ( n4511 , n192 );
nand ( n4512 , n4511 , n188 );
not ( n4513 , n4512 );
nor ( n4514 , n189 , n190 );
nand ( n4515 , n4513 , n4514 );
not ( n4516 , n190 );
nand ( n4517 , n188 , n189 );
not ( n4518 , n4517 );
nand ( n4519 , n4516 , n4518 );
nand ( n4520 , n4510 , n4515 , n4519 );
and ( n4521 , n4460 , n191 );
nand ( n4522 , n4521 , n189 );
buf ( n4523 , n4522 );
not ( n4524 , n4523 );
or ( n4525 , n4520 , n4524 );
nand ( n4526 , n4525 , n4390 );
not ( n4527 , n4526 );
not ( n4528 , n4455 );
nor ( n4529 , n192 , n193 );
not ( n4530 , n4529 );
nand ( n4531 , n4528 , n4530 );
not ( n4532 , n4531 );
or ( n4533 , n4527 , n4532 );
not ( n4534 , n4515 );
nor ( n4535 , n4534 , n4393 );
nand ( n4536 , n4510 , n4523 , n4535 );
nand ( n4537 , n4533 , n4536 );
nand ( n4538 , n193 , n194 );
not ( n4539 , n4538 );
nand ( n4540 , n4539 , n191 );
not ( n4541 , n4408 );
or ( n4542 , n4540 , n4541 );
not ( n4543 , n4488 );
not ( n4544 , n189 );
nand ( n4545 , n4544 , n190 );
not ( n4546 , n4545 );
not ( n4547 , n192 );
nand ( n4548 , n4546 , n4547 );
nand ( n4549 , n4543 , n4548 );
nand ( n4550 , n4549 , n4539 );
not ( n4551 , n191 );
nand ( n4552 , n4551 , n192 );
not ( n4553 , n4552 );
not ( n4554 , n189 );
nor ( n4555 , n4554 , n188 );
nand ( n4556 , n4553 , n4555 );
not ( n4557 , n4556 );
not ( n4558 , n190 );
and ( n4559 , n4557 , n4558 );
nor ( n4560 , n4559 , n4415 );
nand ( n4561 , n4542 , n4550 , n4560 );
not ( n4562 , n194 );
nand ( n4563 , n4546 , n4513 );
nand ( n4564 , n4502 , n4427 );
nand ( n4565 , n4563 , n4564 );
not ( n4566 , n4565 );
or ( n4567 , n4562 , n4566 );
not ( n4568 , n4503 );
nand ( n4569 , n4462 , n189 );
nor ( n4570 , n4568 , n4569 );
nand ( n4571 , n4479 , n4427 );
nand ( n4572 , n4515 , n4571 );
not ( n4573 , n4521 );
nor ( n4574 , n4573 , n4396 );
or ( n4575 , n4570 , n4572 , n4574 );
not ( n4576 , n194 );
nand ( n4577 , n4575 , n4576 );
nand ( n4578 , n4567 , n4577 );
nor ( n4579 , n4561 , n4578 );
nand ( n4580 , n4537 , n4579 );
nand ( n4581 , n4508 , n4580 );
not ( n4582 , n192 );
nand ( n4583 , n4582 , n191 );
not ( n4584 , n4583 );
nand ( n4585 , n4383 , n4584 , n193 );
not ( n4586 , n4461 );
not ( n4587 , n189 );
nand ( n4588 , n4587 , n191 );
not ( n4589 , n4588 );
nand ( n4590 , n4586 , n4589 );
not ( n4591 , n4590 );
nand ( n4592 , n4591 , n4494 );
and ( n4593 , n4585 , n4592 );
and ( n4594 , n192 , n4496 );
not ( n4595 , n192 );
and ( n4596 , n4595 , n4514 );
or ( n4597 , n4594 , n4596 );
nand ( n4598 , n4555 , n4393 );
nor ( n4599 , n4597 , n4598 );
nand ( n4600 , n4491 , n4474 );
nand ( n4601 , n4479 , n4513 );
nand ( n4602 , n4600 , n4601 );
or ( n4603 , n4599 , n4493 , n4602 );
not ( n4604 , n194 );
nor ( n4605 , n4604 , n193 );
nand ( n4606 , n4603 , n4605 );
nor ( n4607 , n191 , n4444 );
nand ( n4608 , n4607 , n192 );
nor ( n4609 , n4608 , n4538 );
nand ( n4610 , n4518 , n192 );
and ( n4611 , n4563 , n4610 );
nor ( n4612 , n4611 , n4540 );
nor ( n4613 , n4609 , n4612 );
not ( n4614 , n4552 );
nand ( n4615 , n4502 , n4614 );
buf ( n4616 , n4400 );
and ( n4617 , n4445 , n4616 );
not ( n4618 , n4617 );
nand ( n4619 , n4615 , n4618 );
and ( n4620 , n4619 , n4451 );
and ( n4621 , n4451 , n4393 );
and ( n4622 , n4381 , n190 );
and ( n4623 , n4621 , n4622 );
nor ( n4624 , n4620 , n4623 );
and ( n4625 , n4593 , n4606 , n4613 , n4624 );
nand ( n4626 , n191 , n192 );
nor ( n4627 , n4626 , n188 );
nand ( n4628 , n4627 , n4546 );
not ( n4629 , n4552 );
not ( n4630 , n4629 );
not ( n4631 , n4630 );
nand ( n4632 , n4631 , n4383 );
not ( n4633 , n4632 );
nor ( n4634 , n4571 , n188 );
not ( n4635 , n4584 );
nor ( n4636 , n4635 , n4495 );
nor ( n4637 , n4634 , n4636 );
not ( n4638 , n4637 );
not ( n4639 , n4588 );
nand ( n4640 , n4423 , n4639 );
not ( n4641 , n4640 );
or ( n4642 , n4633 , n4638 , n4641 );
not ( n4643 , n4634 );
nand ( n4644 , n4643 , n193 );
nand ( n4645 , n4642 , n4644 );
nand ( n4646 , n4628 , n4645 );
nand ( n4647 , n4646 , n4576 );
and ( n4648 , n4581 , n4625 , n4647 );
not ( n4649 , n4648 );
not ( n4650 , n4649 );
not ( n4651 , n4650 );
or ( n4652 , n4377 , n4651 );
not ( n4653 , n4648 );
nand ( n4654 , n4653 , n294 );
nand ( n4655 , n4652 , n4654 );
not ( n4656 , n3732 );
nand ( n4657 , n3803 , n182 );
nor ( n4658 , n180 , n182 );
nand ( n4659 , n4658 , n183 );
nand ( n4660 , n4657 , n4659 );
nor ( n4661 , n3872 , n180 );
not ( n4662 , n4661 );
or ( n4663 , n4660 , n4662 );
not ( n4664 , n3730 );
or ( n4665 , n4664 , n184 );
nand ( n4666 , n4663 , n4665 );
not ( n4667 , n4666 );
or ( n4668 , n4656 , n4667 );
nand ( n4669 , n3787 , n183 );
not ( n4670 , n4669 );
not ( n4671 , n3855 );
or ( n4672 , n4670 , n4671 );
nand ( n4673 , n4672 , n185 );
and ( n4674 , n3940 , n184 );
nand ( n4675 , n3908 , n3738 );
nand ( n4676 , n4675 , n186 );
nor ( n4677 , n4674 , n4676 );
nand ( n4678 , n3878 , n184 );
and ( n4679 , n4673 , n4677 , n4678 );
nand ( n4680 , n4668 , n4679 );
nor ( n4681 , n3824 , n186 );
nor ( n4682 , n3832 , n180 );
nand ( n4683 , n4682 , n184 );
nand ( n4684 , n4681 , n4683 );
not ( n4685 , n3858 );
nand ( n4686 , n4684 , n4685 );
not ( n4687 , n3717 );
and ( n4688 , n4687 , n3785 );
nand ( n4689 , n4688 , n180 );
nand ( n4690 , n3764 , n3861 );
and ( n4691 , n4689 , n4690 );
nand ( n4692 , n4686 , n4691 );
nand ( n4693 , n4680 , n4692 );
not ( n4694 , n4693 );
nor ( n4695 , n3923 , n187 );
not ( n4696 , n3895 );
nand ( n4697 , n3940 , n3949 );
not ( n4698 , n4697 );
or ( n4699 , n4696 , n4698 );
nand ( n4700 , n3888 , n3908 );
nand ( n4701 , n4699 , n4700 );
nand ( n4702 , n4695 , n4701 );
not ( n4703 , n4689 );
not ( n4704 , n3774 );
not ( n4705 , n4704 );
or ( n4706 , n4703 , n4705 );
nand ( n4707 , n4706 , n3811 );
nor ( n4708 , n180 , n183 );
nand ( n4709 , n4687 , n4708 );
nor ( n4710 , n4709 , n184 );
not ( n4711 , n4710 );
not ( n4712 , n4711 );
not ( n4713 , n3765 );
or ( n4714 , n4712 , n4713 );
nand ( n4715 , n4714 , n3858 );
nand ( n4716 , n4707 , n4715 );
nor ( n4717 , n4702 , n4716 );
not ( n4718 , n4717 );
or ( n4719 , n4694 , n4718 );
not ( n4720 , n180 );
nand ( n4721 , n4720 , n181 );
nor ( n4722 , n4721 , n183 );
nand ( n4723 , n3809 , n183 );
not ( n4724 , n4723 );
not ( n4725 , n3834 );
or ( n4726 , n4722 , n4724 , n4725 );
not ( n4727 , n3759 );
nand ( n4728 , n4726 , n4727 );
not ( n4729 , n3802 );
not ( n4730 , n181 );
nor ( n4731 , n4730 , n4658 );
nand ( n4732 , n3949 , n4731 );
not ( n4733 , n4732 );
or ( n4734 , n4729 , n4733 );
not ( n4735 , n4682 );
nand ( n4736 , n4735 , n3843 );
nand ( n4737 , n4734 , n4736 );
and ( n4738 , n180 , n182 );
nand ( n4739 , n3952 , n4738 );
not ( n4740 , n4739 );
not ( n4741 , n4709 );
or ( n4742 , n4740 , n4741 );
nand ( n4743 , n4742 , n186 );
and ( n4744 , n4728 , n4737 , n4743 , n187 );
not ( n4745 , n181 );
nor ( n4746 , n4745 , n183 );
not ( n4747 , n4746 );
and ( n4748 , n3771 , n3854 );
not ( n4749 , n4748 );
or ( n4750 , n4747 , n4749 );
nand ( n4751 , n3730 , n3777 );
nand ( n4752 , n3806 , n3861 );
and ( n4753 , n4751 , n4752 );
nand ( n4754 , n4750 , n4753 );
nand ( n4755 , n3730 , n184 );
nor ( n4756 , n4755 , n185 );
or ( n4757 , n4754 , n4756 );
nand ( n4758 , n4757 , n3749 );
not ( n4759 , n3921 );
nor ( n4760 , n3786 , n3854 );
nand ( n4761 , n4760 , n3761 );
not ( n4762 , n4761 );
nor ( n4763 , n4762 , n3824 );
not ( n4764 , n4763 );
or ( n4765 , n4759 , n4764 );
nand ( n4766 , n4765 , n3811 );
not ( n4767 , n3869 );
nand ( n4768 , n4767 , n3759 );
and ( n4769 , n4758 , n4766 , n4768 );
nand ( n4770 , n4744 , n4769 );
nand ( n4771 , n4719 , n4770 );
not ( n4772 , n3759 );
nand ( n4773 , n4748 , n3773 );
not ( n4774 , n4773 );
not ( n4775 , n3803 );
or ( n4776 , n4774 , n4775 );
not ( n4777 , n4748 );
not ( n4778 , n3940 );
nand ( n4779 , n4777 , n4778 );
nand ( n4780 , n4776 , n4779 );
nand ( n4781 , n4780 , n3901 );
nand ( n4782 , n4781 , n186 );
not ( n4783 , n4782 );
or ( n4784 , n4772 , n4783 );
nor ( n4785 , n4741 , n3814 );
not ( n4786 , n4785 );
not ( n4787 , n185 );
nor ( n4788 , n180 , n181 );
buf ( n4789 , n4788 );
not ( n4790 , n4789 );
nand ( n4791 , n3738 , n3761 );
nor ( n4792 , n4790 , n4791 );
nor ( n4793 , n4787 , n4792 );
not ( n4794 , n4793 );
or ( n4795 , n4786 , n4794 );
nand ( n4796 , n4795 , n3948 );
not ( n4797 , n3719 );
nand ( n4798 , n4797 , n3854 );
nand ( n4799 , n4796 , n4798 );
nand ( n4800 , n4784 , n4799 );
not ( n4801 , n3854 );
not ( n4802 , n3820 );
not ( n4803 , n4802 );
not ( n4804 , n183 );
nand ( n4805 , n4804 , n3712 );
nand ( n4806 , n4803 , n3815 , n4805 );
not ( n4807 , n4806 );
or ( n4808 , n4801 , n4807 );
nand ( n4809 , n4808 , n4793 );
not ( n4810 , n3829 );
nor ( n4811 , n4810 , n3927 );
not ( n4812 , n4811 );
not ( n4813 , n3867 );
nand ( n4814 , n4813 , n184 );
nor ( n4815 , n4814 , n180 );
nor ( n4816 , n4815 , n185 );
buf ( n4817 , n3788 );
nand ( n4818 , n4812 , n4816 , n4817 );
and ( n4819 , n4809 , n4818 , n3749 );
nand ( n4820 , n183 , n185 );
or ( n4821 , n3931 , n4820 );
nand ( n4822 , n3952 , n3829 );
not ( n4823 , n4822 );
not ( n4824 , n3779 );
not ( n4825 , n4824 );
or ( n4826 , n4823 , n4825 );
nand ( n4827 , n4826 , n3749 );
nand ( n4828 , n4821 , n4827 );
nor ( n4829 , n4819 , n4828 );
nand ( n4830 , n4771 , n4800 , n4829 );
not ( n4831 , n4830 );
not ( n4832 , n4831 );
and ( n4833 , n3855 , n3748 );
nor ( n4834 , n4833 , n185 );
nand ( n4835 , n180 , n185 );
not ( n4836 , n4835 );
nand ( n4837 , n3803 , n4836 , n182 );
and ( n4838 , n3943 , n3749 );
not ( n4839 , n185 );
nand ( n4840 , n4839 , n184 );
not ( n4841 , n4840 );
nand ( n4842 , n4722 , n4841 );
nand ( n4843 , n4837 , n4838 , n4842 );
nor ( n4844 , n4834 , n4843 );
and ( n4845 , n3952 , n3845 );
or ( n4846 , n4845 , n4674 );
nand ( n4847 , n4846 , n185 );
and ( n4848 , n4844 , n4847 );
not ( n4849 , n3819 );
nand ( n4850 , n4849 , n183 );
not ( n4851 , n183 );
nand ( n4852 , n4851 , n3833 );
nand ( n4853 , n4850 , n4852 );
not ( n4854 , n3842 );
nand ( n4855 , n4854 , n3915 );
not ( n4856 , n4855 );
or ( n4857 , n4853 , n4856 );
nand ( n4858 , n4857 , n3949 );
nand ( n4859 , n4858 , n186 );
not ( n4860 , n3898 );
nor ( n4861 , n4746 , n4860 );
or ( n4862 , n3874 , n4861 );
nand ( n4863 , n4862 , n4841 );
not ( n4864 , n4709 );
not ( n4865 , n4678 );
or ( n4866 , n4864 , n4865 );
nand ( n4867 , n4866 , n185 );
nand ( n4868 , n4863 , n4867 );
nor ( n4869 , n4859 , n4868 );
nor ( n4870 , n4848 , n4869 );
not ( n4871 , n4659 );
nand ( n4872 , n4871 , n3795 );
nand ( n4873 , n3878 , n3861 );
and ( n4874 , n3855 , n4872 , n4873 , n3748 );
or ( n4875 , n185 , n187 );
or ( n4876 , n4874 , n4875 );
not ( n4877 , n3778 );
nand ( n4878 , n4877 , n4789 );
not ( n4879 , n4878 );
not ( n4880 , n3895 );
nand ( n4881 , n4880 , n4738 );
not ( n4882 , n4881 );
or ( n4883 , n4879 , n4882 );
nand ( n4884 , n4883 , n3811 );
nand ( n4885 , n4876 , n4884 );
nor ( n4886 , n4870 , n4885 );
nand ( n4887 , n4722 , n3949 );
nand ( n4888 , n3935 , n4887 , n3909 , n3749 );
not ( n4889 , n3878 );
or ( n4890 , n4889 , n185 );
not ( n4891 , n183 );
nor ( n4892 , n4891 , n185 );
nand ( n4893 , n4735 , n4860 , n4892 );
nand ( n4894 , n4890 , n4893 , n4700 );
or ( n4895 , n4888 , n4894 );
or ( n4896 , n3889 , n182 );
nor ( n4897 , n4845 , n3749 );
nand ( n4898 , n4896 , n4897 );
nand ( n4899 , n4895 , n4898 );
not ( n4900 , n4899 );
not ( n4901 , n4852 );
nand ( n4902 , n3771 , n183 );
not ( n4903 , n4902 );
or ( n4904 , n4901 , n4903 );
nand ( n4905 , n4904 , n3854 );
not ( n4906 , n4905 );
not ( n4907 , n3723 );
or ( n4908 , n4906 , n4907 );
nand ( n4909 , n4908 , n185 );
not ( n4910 , n187 );
not ( n4911 , n3909 );
or ( n4912 , n4910 , n4911 );
nand ( n4913 , n4912 , n3782 );
not ( n4914 , n3807 );
not ( n4915 , n183 );
nand ( n4916 , n4915 , n3845 );
nor ( n4917 , n4916 , n3848 );
nor ( n4918 , n4914 , n4917 );
not ( n4919 , n3872 );
nand ( n4920 , n3713 , n4919 );
not ( n4921 , n4814 );
or ( n4922 , n4920 , n4921 , n4871 );
nand ( n4923 , n4922 , n4727 );
and ( n4924 , n4909 , n4913 , n4918 , n4923 );
not ( n4925 , n4924 );
or ( n4926 , n4900 , n4925 );
not ( n4927 , n4723 );
not ( n4928 , n3948 );
and ( n4929 , n4927 , n4928 );
nand ( n4930 , n4761 , n186 );
nor ( n4931 , n4929 , n4930 );
or ( n4932 , n4815 , n4877 );
nand ( n4933 , n4932 , n3732 );
and ( n4934 , n4931 , n4798 , n4933 );
nand ( n4935 , n4817 , n3749 );
not ( n4936 , n185 );
nor ( n4937 , n4936 , n3755 );
nand ( n4938 , n3887 , n183 );
nor ( n4939 , n4938 , n3848 );
and ( n4940 , n4746 , n3732 );
nor ( n4941 , n4935 , n4937 , n4939 , n4940 );
or ( n4942 , n4934 , n4941 );
not ( n4943 , n183 );
nand ( n4944 , n4943 , n4788 );
not ( n4945 , n4944 );
nand ( n4946 , n4945 , n3761 );
nand ( n4947 , n3921 , n3815 , n4946 );
not ( n4948 , n3922 );
and ( n4949 , n4947 , n4948 );
nor ( n4950 , n4949 , n187 );
nand ( n4951 , n4942 , n4950 );
nand ( n4952 , n4926 , n4951 );
nand ( n4953 , n4886 , n4952 );
buf ( n4954 , n4953 );
not ( n4955 , n4954 );
not ( n4956 , n4955 );
or ( n4957 , n4832 , n4956 );
nand ( n4958 , n4954 , n4830 );
nand ( n4959 , n4957 , n4958 );
not ( n4960 , n4959 );
and ( n4961 , n4655 , n4960 );
not ( n4962 , n4655 );
and ( n4963 , n4962 , n4959 );
nor ( n4964 , n4961 , n4963 );
and ( n4965 , n4375 , n4964 );
not ( n4966 , n4375 );
not ( n4967 , n4964 );
and ( n4968 , n4966 , n4967 );
nor ( n4969 , n4965 , n4968 );
or ( n4970 , n4969 , n1 );
and ( n4971 , n295 , n4376 );
not ( n4972 , n295 );
and ( n4973 , n4972 , n294 );
nor ( n4974 , n4971 , n4973 );
or ( n4975 , n2246 , n4974 );
nand ( n4976 , n4970 , n4975 );
nand ( n4977 , n3898 , n181 , n183 );
not ( n4978 , n4977 );
nand ( n4979 , n4978 , n4841 );
not ( n4980 , n4820 );
and ( n4981 , n4980 , n3712 );
nor ( n4982 , n4721 , n3916 );
nor ( n4983 , n4981 , n4982 );
and ( n4984 , n4872 , n4983 );
and ( n4985 , n4979 , n4984 , n4732 );
nor ( n4986 , n4985 , n186 );
not ( n4987 , n4944 );
not ( n4988 , n3723 );
nand ( n4989 , n4988 , n3854 );
not ( n4990 , n4989 );
or ( n4991 , n4987 , n4990 );
nand ( n4992 , n4991 , n4727 );
not ( n4993 , n180 );
nor ( n4994 , n4993 , n3832 );
nand ( n4995 , n4994 , n3803 );
not ( n4996 , n4995 );
nor ( n4997 , n4814 , n3915 );
nor ( n4998 , n4997 , n185 );
not ( n4999 , n4998 );
or ( n5000 , n4996 , n4999 );
nand ( n5001 , n3873 , n185 );
not ( n5002 , n5001 );
not ( n5003 , n4944 );
nand ( n5004 , n5003 , n184 );
nand ( n5005 , n5002 , n5004 );
nand ( n5006 , n5000 , n5005 );
not ( n5007 , n187 );
and ( n5008 , n3905 , n5007 );
and ( n5009 , n4992 , n5006 , n5008 );
and ( n5010 , n4940 , n3898 );
nor ( n5011 , n5010 , n4740 );
not ( n5012 , n5011 );
not ( n5013 , n3931 );
nor ( n5014 , n3873 , n184 );
nor ( n5015 , n5013 , n5014 );
not ( n5016 , n5015 );
or ( n5017 , n5012 , n5016 );
nand ( n5018 , n5017 , n186 );
nand ( n5019 , n5009 , n5018 );
or ( n5020 , n4986 , n5019 );
not ( n5021 , n4982 );
buf ( n5022 , n3838 );
nand ( n5023 , n5021 , n5022 );
and ( n5024 , n5023 , n3732 );
nor ( n5025 , n3902 , n5007 );
not ( n5026 , n3764 );
nand ( n5027 , n5026 , n4755 );
or ( n5028 , n5027 , n4802 );
nand ( n5029 , n5028 , n4980 );
nand ( n5030 , n5025 , n5029 );
nor ( n5031 , n5024 , n5030 );
nand ( n5032 , n3856 , n4938 );
or ( n5033 , n5032 , n4748 , n3759 );
and ( n5034 , n3732 , n186 );
nand ( n5035 , n4778 , n5034 );
nand ( n5036 , n5033 , n5035 );
not ( n5037 , n5036 );
nand ( n5038 , n4683 , n3943 );
not ( n5039 , n4700 );
nor ( n5040 , n4978 , n5038 , n5039 );
not ( n5041 , n5040 );
or ( n5042 , n5037 , n5041 );
nor ( n5043 , n3805 , n183 );
nor ( n5044 , n5043 , n3878 , n3811 );
not ( n5045 , n5044 );
not ( n5046 , n3931 );
or ( n5047 , n5045 , n5046 );
nand ( n5048 , n3718 , n3854 );
nand ( n5049 , n4816 , n5048 );
nand ( n5050 , n5047 , n5049 );
nor ( n5051 , n3917 , n186 );
nand ( n5052 , n3747 , n3712 );
and ( n5053 , n5051 , n4822 , n5052 );
nand ( n5054 , n5050 , n5053 );
nand ( n5055 , n5042 , n5054 );
nand ( n5056 , n5031 , n5055 );
nand ( n5057 , n5020 , n5056 );
not ( n5058 , n4683 );
not ( n5059 , n4850 );
or ( n5060 , n5059 , n4741 );
nand ( n5061 , n5060 , n184 );
not ( n5062 , n5061 );
or ( n5063 , n5058 , n5062 );
nand ( n5064 , n5063 , n185 );
not ( n5065 , n5064 );
nand ( n5066 , n4978 , n185 );
not ( n5067 , n3821 );
and ( n5068 , n5067 , n4836 , n182 );
nor ( n5069 , n5068 , n3749 );
nand ( n5070 , n5066 , n5069 );
and ( n5071 , n4940 , n3829 , n184 );
not ( n5072 , n5071 );
nand ( n5073 , n3771 , n4746 );
not ( n5074 , n5073 );
or ( n5075 , n5074 , n4871 , n3868 );
nand ( n5076 , n5075 , n3888 );
nand ( n5077 , n5072 , n5076 );
nor ( n5078 , n5070 , n5077 );
not ( n5079 , n5078 );
or ( n5080 , n5065 , n5079 );
nand ( n5081 , n3749 , n185 );
nor ( n5082 , n4811 , n5081 );
and ( n5083 , n5082 , n5061 , n3905 );
nor ( n5084 , n4688 , n4685 );
nor ( n5085 , n5083 , n5084 );
nand ( n5086 , n5080 , n5085 );
and ( n5087 , n5057 , n5086 , n4690 );
not ( n5088 , n5087 );
and ( n5089 , n4163 , n4158 );
not ( n5090 , n5089 );
not ( n5091 , n5090 );
nor ( n5092 , n4004 , n4160 );
not ( n5093 , n5092 );
nand ( n5094 , n4016 , n3992 );
nor ( n5095 , n5094 , n198 );
nand ( n5096 , n3990 , n4053 );
nand ( n5097 , n4149 , n5096 );
nor ( n5098 , n5095 , n5097 );
not ( n5099 , n5098 );
or ( n5100 , n5093 , n5099 );
nor ( n5101 , n4176 , n199 );
not ( n5102 , n5101 );
buf ( n5103 , n3967 );
not ( n5104 , n5103 );
not ( n5105 , n3978 );
and ( n5106 , n5104 , n5105 );
nor ( n5107 , n5106 , n202 );
nand ( n5108 , n5102 , n5107 );
nand ( n5109 , n5100 , n5108 );
not ( n5110 , n5109 );
or ( n5111 , n5091 , n5110 );
nand ( n5112 , n5111 , n203 );
not ( n5113 , n199 );
not ( n5114 , n4124 );
not ( n5115 , n5114 );
or ( n5116 , n5113 , n5115 );
nand ( n5117 , n5116 , n5096 );
nor ( n5118 , n5117 , n4049 );
not ( n5119 , n5118 );
not ( n5120 , n5095 );
not ( n5121 , n5120 );
or ( n5122 , n5119 , n5121 );
nand ( n5123 , n5122 , n202 );
not ( n5124 , n5123 );
nor ( n5125 , n201 , n202 );
and ( n5126 , n4004 , n5125 );
nand ( n5127 , n4135 , n4056 );
not ( n5128 , n5127 );
nor ( n5129 , n5126 , n5128 );
not ( n5130 , n5129 );
or ( n5131 , n5124 , n5130 );
not ( n5132 , n203 );
nand ( n5133 , n5131 , n5132 );
not ( n5134 , n199 );
nand ( n5135 , n5134 , n4002 );
nor ( n5136 , n5135 , n201 );
nand ( n5137 , n5136 , n4027 );
not ( n5138 , n199 );
nor ( n5139 , n5138 , n4113 );
and ( n5140 , n5139 , n197 );
nand ( n5141 , n5140 , n5125 );
and ( n5142 , n5137 , n5141 );
nand ( n5143 , n5112 , n5133 , n5142 );
nand ( n5144 , n5143 , n4058 );
not ( n5145 , n5137 );
nor ( n5146 , n4026 , n197 );
not ( n5147 , n5146 );
nand ( n5148 , n5147 , n4186 );
nand ( n5149 , n4005 , n4068 );
nand ( n5150 , n3978 , n198 );
not ( n5151 , n5150 );
nand ( n5152 , n5151 , n4027 );
nand ( n5153 , n4195 , n5152 );
or ( n5154 , n5148 , n5149 , n5153 );
nand ( n5155 , n4004 , n3992 );
not ( n5156 , n4056 );
and ( n5157 , n5156 , n4025 , n197 );
nor ( n5158 , n202 , n203 );
not ( n5159 , n5158 );
nor ( n5160 , n5157 , n5159 );
nand ( n5161 , n5155 , n5160 , n3980 );
nand ( n5162 , n5154 , n5161 );
not ( n5163 , n5162 );
or ( n5164 , n5145 , n5163 );
nand ( n5165 , n5140 , n201 );
not ( n5166 , n5165 );
nor ( n5167 , n5166 , n5132 );
nand ( n5168 , n4156 , n4158 );
not ( n5169 , n5168 );
nand ( n5170 , n5169 , n202 );
not ( n5171 , n3984 );
nor ( n5172 , n5171 , n199 );
nand ( n5173 , n5172 , n4060 );
nor ( n5174 , n4083 , n4179 );
not ( n5175 , n5174 );
and ( n5176 , n5170 , n5173 , n5175 );
nand ( n5177 , n4049 , n4092 );
nand ( n5178 , n4053 , n5114 );
not ( n5179 , n200 );
nor ( n5180 , n5178 , n5179 );
not ( n5181 , n5180 );
not ( n5182 , n4015 );
nand ( n5183 , n5182 , n4060 );
nand ( n5184 , n5177 , n5181 , n5183 );
not ( n5185 , n202 );
nand ( n5186 , n5184 , n5185 );
nand ( n5187 , n5167 , n5176 , n5186 );
nand ( n5188 , n5164 , n5187 );
nand ( n5189 , n4127 , n4192 );
nand ( n5190 , n5189 , n202 );
not ( n5191 , n5190 );
not ( n5192 , n4114 );
nand ( n5193 , n5192 , n199 );
and ( n5194 , n5193 , n4135 );
and ( n5195 , n3972 , n4047 );
nor ( n5196 , n5194 , n5195 );
nand ( n5197 , n5191 , n5196 );
not ( n5198 , n5197 );
not ( n5199 , n4010 );
not ( n5200 , n5199 );
nand ( n5201 , n5200 , n5177 , n4062 , n5185 );
not ( n5202 , n5201 );
or ( n5203 , n5198 , n5202 );
not ( n5204 , n4170 );
not ( n5205 , n4107 );
not ( n5206 , n4132 );
or ( n5207 , n5205 , n5206 );
nand ( n5208 , n5207 , n5132 );
not ( n5209 , n5208 );
nand ( n5210 , n4127 , n4160 );
not ( n5211 , n5210 );
nand ( n5212 , n5211 , n198 );
nand ( n5213 , n4095 , n3996 );
nand ( n5214 , n5204 , n5209 , n5212 , n5213 );
not ( n5215 , n199 );
nor ( n5216 , n5215 , n197 );
nand ( n5217 , n4073 , n5216 );
nor ( n5218 , n5217 , n5185 );
or ( n5219 , n5214 , n5218 );
not ( n5220 , n5127 );
not ( n5221 , n4036 );
and ( n5222 , n5220 , n5221 );
nor ( n5223 , n5222 , n5132 );
not ( n5224 , n5172 );
not ( n5225 , n5224 );
not ( n5226 , n4007 );
not ( n5227 , n4176 );
or ( n5228 , n5226 , n5227 );
nand ( n5229 , n5228 , n4160 );
not ( n5230 , n5229 );
or ( n5231 , n5225 , n5230 );
nand ( n5232 , n5231 , n5210 );
not ( n5233 , n4157 );
not ( n5234 , n5233 );
nand ( n5235 , n5223 , n5232 , n5234 );
nand ( n5236 , n5219 , n5235 );
nand ( n5237 , n5203 , n5236 );
nand ( n5238 , n5237 , n204 );
not ( n5239 , n4160 );
not ( n5240 , n4102 );
or ( n5241 , n5239 , n5240 );
nand ( n5242 , n4200 , n4106 );
nand ( n5243 , n5241 , n5242 );
nand ( n5244 , n5144 , n5188 , n5238 , n5243 );
not ( n5245 , n5244 );
not ( n5246 , n5245 );
or ( n5247 , n5088 , n5246 );
not ( n5248 , n5087 );
nand ( n5249 , n5248 , n5244 );
nand ( n5250 , n5247 , n5249 );
nand ( n5251 , n4247 , n3485 );
nand ( n5252 , n3510 , n4356 );
not ( n5253 , n5252 );
or ( n5254 , n5251 , n5253 );
or ( n5255 , n3680 , n3471 );
nand ( n5256 , n5254 , n5255 );
not ( n5257 , n3691 );
nand ( n5258 , n4223 , n210 );
not ( n5259 , n5258 );
nand ( n5260 , n206 , n208 );
not ( n5261 , n5260 );
nand ( n5262 , n5259 , n5261 );
not ( n5263 , n3494 );
not ( n5264 , n3597 );
or ( n5265 , n5263 , n5264 );
nand ( n5266 , n5265 , n3599 );
nand ( n5267 , n5262 , n5266 );
nand ( n5268 , n3647 , n3525 );
nor ( n5269 , n5257 , n5267 , n5268 );
and ( n5270 , n5256 , n5269 );
not ( n5271 , n4241 );
not ( n5272 , n5271 );
not ( n5273 , n4255 );
or ( n5274 , n5272 , n5273 );
nand ( n5275 , n5274 , n209 );
nand ( n5276 , n3684 , n3593 );
nand ( n5277 , n3510 , n205 , n210 );
buf ( n5278 , n5277 );
nand ( n5279 , n3523 , n3475 );
and ( n5280 , n5275 , n5276 , n5278 , n5279 );
not ( n5281 , n4307 );
nor ( n5282 , n5281 , n3572 );
and ( n5283 , n5280 , n5282 );
nor ( n5284 , n5270 , n5283 );
not ( n5285 , n4296 );
not ( n5286 , n5285 );
or ( n5287 , n3579 , n5286 );
and ( n5288 , n209 , n212 );
not ( n5289 , n5288 );
nand ( n5290 , n5287 , n5289 );
nand ( n5291 , n3467 , n210 );
nand ( n5292 , n3469 , n5291 );
not ( n5293 , n3654 );
or ( n5294 , n5292 , n5293 );
not ( n5295 , n3706 );
nand ( n5296 , n5294 , n5295 );
not ( n5297 , n3593 );
nand ( n5298 , n4231 , n5297 );
and ( n5299 , n5298 , n212 );
nand ( n5300 , n5290 , n5296 , n5299 );
or ( n5301 , n5284 , n5300 );
and ( n5302 , n3684 , n3669 );
nand ( n5303 , n5302 , n3503 );
nand ( n5304 , n5303 , n4213 );
nand ( n5305 , n3690 , n5295 );
not ( n5306 , n206 );
nor ( n5307 , n5306 , n3550 );
nand ( n5308 , n3523 , n5307 );
nand ( n5309 , n5285 , n5305 , n5308 , n3525 );
or ( n5310 , n5304 , n5309 );
not ( n5311 , n5295 );
not ( n5312 , n3514 );
not ( n5313 , n5312 );
or ( n5314 , n5311 , n5313 );
nand ( n5315 , n4263 , n3475 );
nand ( n5316 , n5314 , n5315 );
not ( n5317 , n5316 );
nand ( n5318 , n3594 , n207 );
nand ( n5319 , n5318 , n211 );
not ( n5320 , n5319 );
not ( n5321 , n208 );
nor ( n5322 , n206 , n207 );
nand ( n5323 , n5321 , n5322 );
not ( n5324 , n5323 );
not ( n5325 , n3703 );
and ( n5326 , n5324 , n5325 );
nor ( n5327 , n5326 , n3680 );
not ( n5328 , n3611 );
nand ( n5329 , n5328 , n3605 );
nand ( n5330 , n5317 , n5320 , n5327 , n5329 );
nand ( n5331 , n5310 , n5330 );
not ( n5332 , n210 );
not ( n5333 , n3534 );
or ( n5334 , n5332 , n5333 );
not ( n5335 , n4339 );
nand ( n5336 , n5335 , n205 );
nand ( n5337 , n5334 , n5336 );
or ( n5338 , n5337 , n209 );
nand ( n5339 , n3611 , n209 );
nand ( n5340 , n5338 , n5339 );
not ( n5341 , n5323 );
not ( n5342 , n4356 );
nand ( n5343 , n5342 , n3629 );
and ( n5344 , n5341 , n5343 );
nor ( n5345 , n5344 , n212 );
nand ( n5346 , n5331 , n5340 , n5345 );
nand ( n5347 , n5301 , n5346 );
nand ( n5348 , n4241 , n5295 );
not ( n5349 , n5348 );
nor ( n5350 , n3679 , n209 );
nand ( n5351 , n5350 , n3462 );
not ( n5352 , n5351 );
or ( n5353 , n5349 , n5352 );
nand ( n5354 , n5353 , n211 );
not ( n5355 , n4246 );
nor ( n5356 , n5355 , n208 );
nor ( n5357 , n3474 , n4318 );
not ( n5358 , n4273 );
or ( n5359 , n5356 , n5357 , n5358 );
and ( n5360 , n3552 , n211 );
nand ( n5361 , n5359 , n5360 );
nand ( n5362 , n5354 , n5361 );
not ( n5363 , n3615 );
nand ( n5364 , n5363 , n3697 );
not ( n5365 , n5364 );
nand ( n5366 , n3478 , n4223 );
not ( n5367 , n5366 );
nand ( n5368 , n5367 , n3564 );
not ( n5369 , n5368 );
or ( n5370 , n5365 , n5369 );
nand ( n5371 , n5370 , n3636 );
not ( n5372 , n3543 );
not ( n5373 , n3558 );
or ( n5374 , n5372 , n5373 );
nand ( n5375 , n5374 , n5278 );
and ( n5376 , n209 , n211 );
and ( n5377 , n5375 , n5376 );
nor ( n5378 , n3593 , n211 );
not ( n5379 , n5378 );
not ( n5380 , n4263 );
or ( n5381 , n5379 , n5380 );
not ( n5382 , n5322 );
nor ( n5383 , n5382 , n3587 );
nand ( n5384 , n5383 , n205 );
nand ( n5385 , n5381 , n5384 );
nor ( n5386 , n5377 , n5385 );
not ( n5387 , n3551 );
or ( n5388 , n4326 , n5387 );
nand ( n5389 , n5388 , n3630 );
nand ( n5390 , n5371 , n5386 , n5389 );
nor ( n5391 , n5362 , n5390 );
nand ( n5392 , n5347 , n5391 );
not ( n5393 , n5392 );
not ( n5394 , n5393 );
not ( n5395 , n4361 );
not ( n5396 , n5395 );
or ( n5397 , n5394 , n5396 );
not ( n5398 , n5395 );
nand ( n5399 , n5398 , n5392 );
nand ( n5400 , n5397 , n5399 );
not ( n5401 , n5400 );
and ( n5402 , n5250 , n5401 );
not ( n5403 , n5250 );
and ( n5404 , n5403 , n5400 );
nor ( n5405 , n5402 , n5404 );
not ( n5406 , n3914 );
not ( n5407 , n5406 );
and ( n5408 , n4773 , n3935 , n4822 , n4678 );
not ( n5409 , n5408 );
or ( n5410 , n5407 , n5409 );
not ( n5411 , n3900 );
not ( n5412 , n3846 );
or ( n5413 , n4688 , n5412 );
nand ( n5414 , n5413 , n3810 , n4944 );
nand ( n5415 , n5411 , n5414 );
nand ( n5416 , n5410 , n5415 );
not ( n5417 , n5416 );
and ( n5418 , n4873 , n3749 );
not ( n5419 , n5418 );
or ( n5420 , n5417 , n5419 );
and ( n5421 , n3941 , n3810 );
not ( n5422 , n5421 );
not ( n5423 , n5015 );
or ( n5424 , n5422 , n5423 );
nand ( n5425 , n5424 , n3811 );
nand ( n5426 , n3910 , n185 );
not ( n5427 , n3822 );
or ( n5428 , n3843 , n3922 );
and ( n5429 , n5426 , n5427 , n4897 , n5428 );
nand ( n5430 , n5425 , n5429 );
nand ( n5431 , n5420 , n5430 );
not ( n5432 , n3868 );
nand ( n5433 , n5432 , n3811 );
or ( n5434 , n5059 , n5433 );
not ( n5435 , n3790 );
and ( n5436 , n5435 , n185 );
not ( n5437 , n5436 );
nand ( n5438 , n5434 , n5437 );
nand ( n5439 , n3939 , n5438 , n4812 );
nand ( n5440 , n4940 , n180 );
nor ( n5441 , n4760 , n186 );
not ( n5442 , n4688 );
and ( n5443 , n5440 , n3864 , n5441 , n5442 );
nand ( n5444 , n5066 , n5443 );
nand ( n5445 , n5439 , n5444 );
not ( n5446 , n5445 );
not ( n5447 , n4820 );
not ( n5448 , n4700 );
or ( n5449 , n5447 , n5448 );
nand ( n5450 , n5449 , n4738 );
not ( n5451 , n5450 );
and ( n5452 , n3738 , n3712 );
nor ( n5453 , n5452 , n4937 , n186 );
not ( n5454 , n5453 );
or ( n5455 , n5451 , n5454 );
not ( n5456 , n3821 );
not ( n5457 , n3856 );
not ( n5458 , n5457 );
or ( n5459 , n5456 , n5458 );
nand ( n5460 , n5459 , n5034 );
buf ( n5461 , n3791 );
nor ( n5462 , n5460 , n5461 );
nor ( n5463 , n4938 , n184 );
nor ( n5464 , n3879 , n5463 , n3759 );
or ( n5465 , n5462 , n5464 );
not ( n5466 , n4997 );
nand ( n5467 , n5465 , n5466 );
nand ( n5468 , n5455 , n5467 );
nand ( n5469 , n4797 , n3888 );
not ( n5470 , n3747 );
not ( n5471 , n5412 );
or ( n5472 , n5470 , n5471 );
nand ( n5473 , n5472 , n4878 );
nand ( n5474 , n5473 , n185 );
not ( n5475 , n3899 );
nor ( n5476 , n5475 , n187 );
and ( n5477 , n5469 , n5474 , n5476 );
nand ( n5478 , n5468 , n5477 );
nand ( n5479 , n5446 , n5478 );
not ( n5480 , n187 );
nand ( n5481 , n5002 , n4791 , n3927 , n4822 );
nand ( n5482 , n3941 , n4683 , n4675 , n3811 );
nand ( n5483 , n5481 , n5482 );
not ( n5484 , n5483 );
or ( n5485 , n5480 , n5484 );
nand ( n5486 , n5485 , n5478 );
and ( n5487 , n4767 , n4841 );
and ( n5488 , n3814 , n4948 );
nor ( n5489 , n5487 , n5488 );
nand ( n5490 , n5431 , n5479 , n5486 , n5489 );
not ( n5491 , n5490 );
not ( n5492 , n5491 );
not ( n5493 , n5492 );
not ( n5494 , n4519 );
nand ( n5495 , n5494 , n193 );
and ( n5496 , n4428 , n5495 , n194 );
nand ( n5497 , n4622 , n4547 );
not ( n5498 , n5497 );
nor ( n5499 , n4569 , n4584 );
or ( n5500 , n5498 , n5499 );
nand ( n5501 , n5500 , n4390 );
and ( n5502 , n4546 , n192 );
nand ( n5503 , n5502 , n4437 );
and ( n5504 , n5496 , n5501 , n5503 );
not ( n5505 , n4390 );
nand ( n5506 , n4423 , n4393 );
not ( n5507 , n5506 );
or ( n5508 , n5505 , n5507 );
nand ( n5509 , n5508 , n4518 );
or ( n5510 , n5509 , n4396 );
nand ( n5511 , n4584 , n4616 );
nand ( n5512 , n5510 , n5511 );
and ( n5513 , n4381 , n4382 );
not ( n5514 , n5513 );
not ( n5515 , n193 );
or ( n5516 , n5514 , n5515 );
nand ( n5517 , n5516 , n4604 );
nor ( n5518 , n5512 , n5517 );
nor ( n5519 , n5504 , n5518 );
nand ( n5520 , n4616 , n4494 );
not ( n5521 , n192 );
nand ( n5522 , n5521 , n4486 );
nand ( n5523 , n5520 , n5522 );
and ( n5524 , n5523 , n4401 , n193 );
not ( n5525 , n4555 );
nand ( n5526 , n188 , n191 );
and ( n5527 , n5525 , n5526 );
nand ( n5528 , n5524 , n5527 );
nor ( n5529 , n191 , n193 );
not ( n5530 , n5529 );
nor ( n5531 , n5530 , n4444 );
nand ( n5532 , n5531 , n192 );
nand ( n5533 , n4405 , n4415 , n5528 , n5532 );
nor ( n5534 , n5519 , n5533 );
not ( n5535 , n4504 );
not ( n5536 , n4446 );
nand ( n5537 , n5513 , n5536 );
not ( n5538 , n5537 );
or ( n5539 , n5535 , n5538 );
nand ( n5540 , n5539 , n4390 );
not ( n5541 , n188 );
nand ( n5542 , n4584 , n5541 );
not ( n5543 , n5542 );
nand ( n5544 , n5543 , n4546 );
not ( n5545 , n4616 );
nand ( n5546 , n4639 , n5545 , n4390 );
nand ( n5547 , n5544 , n5546 );
nand ( n5548 , n190 , n191 );
nor ( n5549 , n4487 , n5548 );
nor ( n5550 , n5549 , n4604 );
not ( n5551 , n5550 );
nor ( n5552 , n5547 , n5551 );
nand ( n5553 , n5540 , n5552 );
not ( n5554 , n4417 );
nand ( n5555 , n5554 , n4509 );
not ( n5556 , n4441 );
not ( n5557 , n5556 );
nand ( n5558 , n5557 , n4437 );
nand ( n5559 , n5555 , n5558 );
or ( n5560 , n5553 , n5559 );
not ( n5561 , n4628 );
not ( n5562 , n4480 );
nand ( n5563 , n4509 , n4393 );
not ( n5564 , n5563 );
nor ( n5565 , n5561 , n5562 , n4390 , n5564 );
nand ( n5566 , n4584 , n189 );
nor ( n5567 , n5566 , n188 );
nand ( n5568 , n4622 , n5536 );
not ( n5569 , n5568 );
nor ( n5570 , n5567 , n5569 );
and ( n5571 , n5565 , n5570 );
not ( n5572 , n4439 );
and ( n5573 , n4614 , n4486 );
nor ( n5574 , n5572 , n4607 , n5573 , n193 );
nor ( n5575 , n5571 , n5574 );
nand ( n5576 , n5560 , n5575 );
nand ( n5577 , n5534 , n5576 );
not ( n5578 , n5577 );
and ( n5579 , n4590 , n193 );
not ( n5580 , n5579 );
not ( n5581 , n5580 );
not ( n5582 , n190 );
nand ( n5583 , n5582 , n4629 );
and ( n5584 , n5542 , n4409 , n5583 );
nand ( n5585 , n5581 , n5584 );
nand ( n5586 , n4639 , n4408 );
and ( n5587 , n5586 , n4475 , n4390 );
nand ( n5588 , n5537 , n5587 );
and ( n5589 , n5585 , n5588 );
nor ( n5590 , n5589 , n4415 );
nand ( n5591 , n4509 , n4584 );
not ( n5592 , n5591 );
not ( n5593 , n5592 );
nand ( n5594 , n4423 , n4547 );
not ( n5595 , n4622 );
nand ( n5596 , n5594 , n5595 );
nand ( n5597 , n5596 , n4468 , n4390 );
nand ( n5598 , n4396 , n4462 );
nand ( n5599 , n5593 , n5597 , n5598 );
nand ( n5600 , n4632 , n194 );
or ( n5601 , n5599 , n5600 );
or ( n5602 , n4529 , n191 );
nand ( n5603 , n5602 , n4496 );
nor ( n5604 , n190 , n193 );
not ( n5605 , n5604 );
not ( n5606 , n4627 );
or ( n5607 , n5605 , n5606 );
nand ( n5608 , n5607 , n4576 );
and ( n5609 , n4584 , n4408 );
nor ( n5610 , n5608 , n5609 );
buf ( n5611 , n4389 );
nand ( n5612 , n5611 , n193 );
nand ( n5613 , n5603 , n5610 , n5612 );
nand ( n5614 , n5601 , n5613 );
nand ( n5615 , n5590 , n5614 );
not ( n5616 , n5615 );
nand ( n5617 , n5616 , n5576 );
not ( n5618 , n5617 );
or ( n5619 , n5578 , n5618 );
or ( n5620 , n5553 , n5559 );
not ( n5621 , n4405 );
not ( n5622 , n190 );
nand ( n5623 , n5622 , n192 );
nor ( n5624 , n4517 , n5623 );
nand ( n5625 , n5624 , n191 );
nand ( n5626 , n5625 , n4576 );
or ( n5627 , n5621 , n5626 );
nand ( n5628 , n5620 , n5627 );
not ( n5629 , n5628 );
not ( n5630 , n4529 );
not ( n5631 , n4641 );
or ( n5632 , n5630 , n5631 );
or ( n5633 , n4610 , n4417 );
nand ( n5634 , n5632 , n5633 );
nor ( n5635 , n5629 , n5634 );
nand ( n5636 , n5619 , n5635 );
not ( n5637 , n5636 );
or ( n5638 , n5493 , n5637 );
not ( n5639 , n5636 );
nand ( n5640 , n5639 , n5491 );
nand ( n5641 , n5638 , n5640 );
not ( n5642 , n324 );
not ( n5643 , n4955 );
or ( n5644 , n5642 , n5643 );
not ( n5645 , n4954 );
not ( n5646 , n5645 );
not ( n5647 , n324 );
nand ( n5648 , n5646 , n5647 );
nand ( n5649 , n5644 , n5648 );
not ( n5650 , n5649 );
and ( n5651 , n5641 , n5650 );
not ( n5652 , n5641 );
and ( n5653 , n5652 , n5649 );
nor ( n5654 , n5651 , n5653 );
and ( n5655 , n5405 , n5654 );
not ( n5656 , n5405 );
not ( n5657 , n5654 );
and ( n5658 , n5656 , n5657 );
nor ( n5659 , n5655 , n5658 );
or ( n5660 , n5659 , n1 );
and ( n5661 , n325 , n5647 );
not ( n5662 , n325 );
and ( n5663 , n5662 , n324 );
nor ( n5664 , n5661 , n5663 );
or ( n5665 , n2246 , n5664 );
nand ( n5666 , n5660 , n5665 );
and ( n5667 , n4171 , n5210 , n4067 );
nand ( n5668 , n4049 , n202 );
not ( n5669 , n5139 );
not ( n5670 , n5669 );
not ( n5671 , n4179 );
nand ( n5672 , n5670 , n5671 );
nand ( n5673 , n5667 , n5668 , n5672 );
not ( n5674 , n5673 );
not ( n5675 , n4037 );
nand ( n5676 , n5675 , n4051 );
nand ( n5677 , n4159 , n203 );
or ( n5678 , n4164 , n5677 );
nand ( n5679 , n5678 , n4077 );
nand ( n5680 , n5676 , n5679 , n4151 , n4136 );
not ( n5681 , n5680 );
or ( n5682 , n5674 , n5681 );
and ( n5683 , n4070 , n5135 );
not ( n5684 , n5125 );
nor ( n5685 , n5683 , n5684 );
nor ( n5686 , n4205 , n5685 );
nand ( n5687 , n4049 , n199 );
nand ( n5688 , n5687 , n4058 );
not ( n5689 , n5155 );
or ( n5690 , n5688 , n5689 );
nand ( n5691 , n4058 , n202 );
nand ( n5692 , n5690 , n5691 );
nand ( n5693 , n4133 , n4070 );
nand ( n5694 , n5693 , n4087 );
and ( n5695 , n5686 , n5692 , n5694 );
nand ( n5696 , n5682 , n5695 );
not ( n5697 , n5167 );
not ( n5698 , n197 );
nand ( n5699 , n4007 , n4009 );
nand ( n5700 , n5699 , n202 );
not ( n5701 , n5700 );
or ( n5702 , n5698 , n5701 );
nor ( n5703 , n197 , n198 );
nand ( n5704 , n5703 , n199 );
nand ( n5705 , n5704 , n4027 );
and ( n5706 , n4015 , n3986 );
or ( n5707 , n5705 , n5706 );
nand ( n5708 , n5707 , n202 );
nand ( n5709 , n4185 , n5125 );
nand ( n5710 , n5708 , n5709 );
nand ( n5711 , n5702 , n5710 );
not ( n5712 , n5711 );
or ( n5713 , n5697 , n5712 );
and ( n5714 , n5168 , n5152 );
not ( n5715 , n4068 );
not ( n5716 , n4026 );
or ( n5717 , n5715 , n5716 );
not ( n5718 , n4165 );
not ( n5719 , n5193 );
or ( n5720 , n5718 , n5719 );
nand ( n5721 , n5720 , n197 );
nand ( n5722 , n5721 , n5704 , n5158 );
nand ( n5723 , n5717 , n5722 );
nand ( n5724 , n4158 , n5125 );
nand ( n5725 , n5714 , n5723 , n5724 );
nand ( n5726 , n5713 , n5725 );
not ( n5727 , n198 );
not ( n5728 , n4034 );
or ( n5729 , n5727 , n5728 );
nand ( n5730 , n5729 , n202 );
not ( n5731 , n4081 );
nand ( n5732 , n4156 , n5731 );
nand ( n5733 , n4092 , n4061 );
nand ( n5734 , n5732 , n5733 , n204 );
or ( n5735 , n5730 , n5734 );
nand ( n5736 , n5168 , n4137 );
nand ( n5737 , n5735 , n5736 );
not ( n5738 , n3971 );
nand ( n5739 , n5738 , n4002 );
not ( n5740 , n5739 );
nand ( n5741 , n3996 , n3990 );
nor ( n5742 , n5741 , n4179 );
nor ( n5743 , n5740 , n5742 );
and ( n5744 , n5737 , n5743 );
nand ( n5745 , n5726 , n5744 );
nand ( n5746 , n5696 , n5745 );
nand ( n5747 , n4207 , n4156 );
and ( n5748 , n4128 , n5733 );
and ( n5749 , n5137 , n5747 , n4005 , n5748 );
or ( n5750 , n5749 , n4160 );
or ( n5751 , n4127 , n4081 );
nand ( n5752 , n5751 , n4102 , n5189 );
and ( n5753 , n5752 , n4107 );
nor ( n5754 , n5753 , n4067 );
nand ( n5755 , n5750 , n5754 );
not ( n5756 , n5685 );
not ( n5757 , n3972 );
not ( n5758 , n5757 );
not ( n5759 , n5114 );
not ( n5760 , n5759 );
and ( n5761 , n5758 , n5760 );
not ( n5762 , n4017 );
nor ( n5763 , n5761 , n5762 );
not ( n5764 , n5763 );
not ( n5765 , n5165 );
or ( n5766 , n5764 , n5765 );
nand ( n5767 , n5766 , n202 );
not ( n5768 , n4181 );
nand ( n5769 , n5768 , n4067 );
nor ( n5770 , n4106 , n4115 , n199 );
nor ( n5771 , n5769 , n5770 );
nand ( n5772 , n5756 , n5767 , n5771 );
and ( n5773 , n5755 , n5772 );
not ( n5774 , n5178 );
nand ( n5775 , n5774 , n5179 );
and ( n5776 , n5120 , n5775 );
nor ( n5777 , n5776 , n202 );
nor ( n5778 , n5773 , n5777 );
nand ( n5779 , n5746 , n5778 );
not ( n5780 , n5779 );
nand ( n5781 , n3997 , n3986 );
not ( n5782 , n5781 );
not ( n5783 , n4126 );
nor ( n5784 , n3981 , n5783 );
not ( n5785 , n5784 );
or ( n5786 , n5782 , n5785 );
nand ( n5787 , n5786 , n4160 );
not ( n5788 , n5103 );
not ( n5789 , n4071 );
not ( n5790 , n5789 );
or ( n5791 , n5788 , n5790 );
nand ( n5792 , n5791 , n4068 );
nor ( n5793 , n5127 , n4036 );
nand ( n5794 , n5793 , n202 );
not ( n5795 , n5742 );
and ( n5796 , n5792 , n5794 , n5795 , n4058 );
not ( n5797 , n4016 );
not ( n5798 , n3991 );
or ( n5799 , n5797 , n5798 );
nand ( n5800 , n5799 , n203 );
not ( n5801 , n5800 );
nand ( n5802 , n3992 , n4061 );
nand ( n5803 , n5801 , n5802 , n5709 );
and ( n5804 , n4004 , n5671 );
or ( n5805 , n5803 , n5804 );
not ( n5806 , n3986 );
nand ( n5807 , n5189 , n4102 );
not ( n5808 , n5807 );
or ( n5809 , n5806 , n5808 );
not ( n5810 , n5208 );
nand ( n5811 , n5809 , n5810 );
nand ( n5812 , n5805 , n5811 );
nand ( n5813 , n5787 , n5796 , n5812 );
not ( n5814 , n5813 );
not ( n5815 , n5140 );
not ( n5816 , n5815 );
not ( n5817 , n4036 );
not ( n5818 , n5706 );
or ( n5819 , n5817 , n5818 );
nand ( n5820 , n5819 , n5132 );
nor ( n5821 , n5730 , n5820 );
not ( n5822 , n5821 );
or ( n5823 , n5816 , n5822 );
nand ( n5824 , n5747 , n5158 );
nand ( n5825 , n5823 , n5824 );
not ( n5826 , n5136 );
nand ( n5827 , n3985 , n3978 );
not ( n5828 , n198 );
nand ( n5829 , n5828 , n3978 );
and ( n5830 , n5826 , n5827 , n5829 );
nand ( n5831 , n5825 , n5830 );
not ( n5832 , n5831 );
nand ( n5833 , n5759 , n203 );
or ( n5834 , n4049 , n5833 );
nand ( n5835 , n5834 , n4077 );
nand ( n5836 , n4037 , n5835 );
not ( n5837 , n5836 );
or ( n5838 , n5832 , n5837 );
nor ( n5839 , n4172 , n5101 );
and ( n5840 , n5839 , n3973 );
nor ( n5841 , n5840 , n5185 );
nand ( n5842 , n4064 , n204 );
not ( n5843 , n5842 );
not ( n5844 , n199 );
not ( n5845 , n3976 );
or ( n5846 , n5844 , n5845 );
nand ( n5847 , n5846 , n5739 );
nand ( n5848 , n5847 , n4160 );
not ( n5849 , n5156 );
not ( n5850 , n3989 );
or ( n5851 , n5849 , n5850 );
nand ( n5852 , n5851 , n4107 );
nand ( n5853 , n5843 , n5848 , n5173 , n5852 );
nor ( n5854 , n5841 , n5853 );
nand ( n5855 , n5838 , n5854 );
not ( n5856 , n5855 );
or ( n5857 , n5814 , n5856 );
not ( n5858 , n5146 );
nand ( n5859 , n5858 , n5178 );
and ( n5860 , n5859 , n202 );
nand ( n5861 , n5185 , n5114 );
nor ( n5862 , n4010 , n5861 );
not ( n5863 , n5862 );
nand ( n5864 , n5863 , n4067 );
nor ( n5865 , n5860 , n5864 );
not ( n5866 , n5137 );
nor ( n5867 , n5096 , n200 );
nor ( n5868 , n5867 , n5169 );
not ( n5869 , n5868 );
or ( n5870 , n5866 , n5869 );
nand ( n5871 , n5870 , n4160 );
nand ( n5872 , n5865 , n5871 , n4088 );
nor ( n5873 , n5793 , n5132 );
and ( n5874 , n5873 , n5177 );
nand ( n5875 , n3966 , n4060 );
and ( n5876 , n202 , n5875 );
not ( n5877 , n202 );
and ( n5878 , n5877 , n5768 );
or ( n5879 , n5876 , n5878 );
nand ( n5880 , n5676 , n5874 , n5879 );
and ( n5881 , n5872 , n5880 );
and ( n5882 , n202 , n4139 );
not ( n5883 , n202 );
not ( n5884 , n5802 );
and ( n5885 , n5883 , n5884 );
nor ( n5886 , n5882 , n5885 );
nor ( n5887 , n5886 , n4086 );
nor ( n5888 , n5881 , n5887 );
nand ( n5889 , n5857 , n5888 );
not ( n5890 , n5889 );
not ( n5891 , n5890 );
or ( n5892 , n5780 , n5891 );
not ( n5893 , n5779 );
nand ( n5894 , n5893 , n5889 );
nand ( n5895 , n5892 , n5894 );
not ( n5896 , n5895 );
not ( n5897 , n5288 );
not ( n5898 , n5252 );
or ( n5899 , n5897 , n5898 );
nand ( n5900 , n4221 , n4242 );
and ( n5901 , n3514 , n3471 );
and ( n5902 , n3615 , n212 );
nand ( n5903 , n5901 , n5902 );
or ( n5904 , n5900 , n5903 );
nand ( n5905 , n5899 , n5904 );
buf ( n5906 , n3479 );
not ( n5907 , n5906 );
nand ( n5908 , n5907 , n3564 );
and ( n5909 , n4252 , n5908 );
and ( n5910 , n5905 , n5909 );
not ( n5911 , n5910 );
nand ( n5912 , n3467 , n3462 );
and ( n5913 , n5912 , n4215 , n3670 );
not ( n5914 , n3468 );
nand ( n5915 , n4275 , n5260 );
not ( n5916 , n5915 );
or ( n5917 , n5914 , n5916 );
nand ( n5918 , n3506 , n207 );
nand ( n5919 , n5917 , n5918 );
not ( n5920 , n5919 );
nor ( n5921 , n5913 , n5920 );
and ( n5922 , n3619 , n3466 );
nor ( n5923 , n5922 , n3663 );
or ( n5924 , n5921 , n5923 , n5363 );
and ( n5925 , n4325 , n209 );
nor ( n5926 , n3629 , n3609 );
not ( n5927 , n3498 );
not ( n5928 , n5927 );
nor ( n5929 , n5928 , n3706 );
nor ( n5930 , n5925 , n5926 , n5929 );
not ( n5931 , n5319 );
not ( n5932 , n4326 );
nand ( n5933 , n5930 , n5931 , n5932 );
nand ( n5934 , n5924 , n5933 );
not ( n5935 , n5934 );
or ( n5936 , n5911 , n5935 );
nand ( n5937 , n3483 , n3543 );
and ( n5938 , n5384 , n5937 );
not ( n5939 , n4325 );
nor ( n5940 , n5939 , n5342 );
nor ( n5941 , n5940 , n3694 );
nand ( n5942 , n5938 , n5941 , n3481 , n4258 );
not ( n5943 , n3678 );
not ( n5944 , n3690 );
or ( n5945 , n5943 , n5944 );
nand ( n5946 , n5945 , n211 );
nand ( n5947 , n3665 , n5297 );
nand ( n5948 , n4215 , n5947 );
nor ( n5949 , n5946 , n5948 );
not ( n5950 , n208 );
nand ( n5951 , n5950 , n3550 );
and ( n5952 , n5937 , n5951 );
nand ( n5953 , n5927 , n208 );
not ( n5954 , n5953 );
or ( n5955 , n5954 , n3502 );
or ( n5956 , n3467 , n3553 );
nand ( n5957 , n5955 , n5956 );
nand ( n5958 , n5949 , n5952 , n5957 );
nand ( n5959 , n5942 , n5958 );
nand ( n5960 , n5949 , n5329 , n3685 , n209 );
nand ( n5961 , n5277 , n3514 );
not ( n5962 , n5961 );
nand ( n5963 , n5938 , n5962 , n3636 );
nand ( n5964 , n5960 , n5963 );
or ( n5965 , n5959 , n5964 );
and ( n5966 , n3697 , n3665 );
nand ( n5967 , n3691 , n4236 );
nor ( n5968 , n5966 , n5967 );
and ( n5969 , n5968 , n3524 , n3672 );
nand ( n5970 , n5965 , n5969 );
nand ( n5971 , n5936 , n5970 );
buf ( n5972 , n3478 );
not ( n5973 , n5972 );
and ( n5974 , n3520 , n5973 );
not ( n5975 , n3666 );
nor ( n5976 , n3474 , n5261 , n210 );
nor ( n5977 , n5974 , n5975 , n5976 );
not ( n5978 , n5977 );
not ( n5979 , n211 );
nor ( n5980 , n5979 , n209 );
not ( n5981 , n5980 );
not ( n5982 , n5981 );
and ( n5983 , n5978 , n5982 );
not ( n5984 , n4260 );
nand ( n5985 , n5984 , n5368 , n4247 );
and ( n5986 , n5985 , n4258 );
nor ( n5987 , n5983 , n5986 );
not ( n5988 , n3469 );
not ( n5989 , n3689 );
nand ( n5990 , n5989 , n3462 );
not ( n5991 , n5990 );
or ( n5992 , n5988 , n5991 );
nand ( n5993 , n5992 , n3605 );
nand ( n5994 , n5993 , n5336 );
nand ( n5995 , n5994 , n3636 );
not ( n5996 , n5262 );
not ( n5997 , n3458 );
or ( n5998 , n5996 , n5997 );
nand ( n5999 , n5998 , n3525 );
or ( n6000 , n4225 , n5387 );
nand ( n6001 , n6000 , n3630 );
and ( n6002 , n5995 , n5999 , n6001 );
not ( n6003 , n4333 );
not ( n6004 , n5932 );
or ( n6005 , n6003 , n6004 );
nand ( n6006 , n6005 , n210 );
not ( n6007 , n6006 );
not ( n6008 , n4252 );
or ( n6009 , n6007 , n6008 );
nand ( n6010 , n6009 , n5376 );
and ( n6011 , n5987 , n6002 , n6010 );
nand ( n6012 , n5971 , n6011 );
not ( n6013 , n6012 );
not ( n6014 , n4211 );
not ( n6015 , n6014 );
or ( n6016 , n6013 , n6015 );
not ( n6017 , n6012 );
nand ( n6018 , n4211 , n6017 );
nand ( n6019 , n6016 , n6018 );
not ( n6020 , n6019 );
or ( n6021 , n5896 , n6020 );
not ( n6022 , n6019 );
not ( n6023 , n5895 );
nand ( n6024 , n6022 , n6023 );
nand ( n6025 , n6021 , n6024 );
nand ( n6026 , n6025 , n2246 );
not ( n6027 , n4831 );
xor ( n6028 , n367 , n6027 );
nand ( n6029 , n4502 , n192 );
not ( n6030 , n6029 );
not ( n6031 , n4510 );
or ( n6032 , n6030 , n6031 );
nand ( n6033 , n6032 , n5554 );
not ( n6034 , n5625 );
nand ( n6035 , n5513 , n192 );
not ( n6036 , n6035 );
or ( n6037 , n6034 , n6036 );
not ( n6038 , n193 );
nand ( n6039 , n6037 , n6038 );
nand ( n6040 , n6033 , n6039 );
not ( n6041 , n4501 );
not ( n6042 , n192 );
nand ( n6043 , n6042 , n4479 );
not ( n6044 , n6043 );
or ( n6045 , n6041 , n6044 );
nor ( n6046 , n191 , n193 );
nand ( n6047 , n6045 , n6046 );
not ( n6048 , n6047 );
nor ( n6049 , n6048 , n195 );
nand ( n6050 , n4585 , n6049 );
nor ( n6051 , n6040 , n6050 );
nand ( n6052 , n4522 , n194 );
not ( n6053 , n4627 );
not ( n6054 , n6053 );
not ( n6055 , n4640 );
or ( n6056 , n6054 , n6055 );
not ( n6057 , n193 );
nand ( n6058 , n6056 , n6057 );
not ( n6059 , n5604 );
nand ( n6060 , n6059 , n5573 );
nand ( n6061 , n6058 , n6060 );
or ( n6062 , n6052 , n6061 );
not ( n6063 , n4530 );
not ( n6064 , n5566 );
or ( n6065 , n6063 , n6064 );
nand ( n6066 , n6065 , n190 );
nand ( n6067 , n5502 , n5554 );
nand ( n6068 , n6066 , n6067 );
or ( n6069 , n5517 , n6068 );
nand ( n6070 , n6062 , n6069 );
nand ( n6071 , n6051 , n6070 );
not ( n6072 , n6071 );
nand ( n6073 , n4546 , n5529 , n5541 );
not ( n6074 , n6073 );
not ( n6075 , n5550 );
or ( n6076 , n6074 , n6075 );
nor ( n6077 , n5567 , n194 );
nand ( n6078 , n4519 , n4547 );
nand ( n6079 , n4424 , n4466 , n4517 );
nand ( n6080 , n6078 , n6079 , n4390 );
not ( n6081 , n4396 );
not ( n6082 , n5506 );
nand ( n6083 , n6081 , n6082 );
not ( n6084 , n4548 );
nand ( n6085 , n6084 , n4437 );
nand ( n6086 , n6077 , n6080 , n6083 , n6085 );
nand ( n6087 , n6076 , n6086 );
not ( n6088 , n4513 );
not ( n6089 , n6088 );
not ( n6090 , n4556 );
or ( n6091 , n6089 , n6090 );
not ( n6092 , n4474 );
nand ( n6093 , n6092 , n5526 );
not ( n6094 , n6093 );
nand ( n6095 , n6091 , n6094 );
not ( n6096 , n5624 );
nand ( n6097 , n6095 , n6096 );
not ( n6098 , n6097 );
not ( n6099 , n193 );
or ( n6100 , n6098 , n6099 );
not ( n6101 , n5529 );
nor ( n6102 , n6101 , n5556 );
nor ( n6103 , n5522 , n4417 );
nand ( n6104 , n4629 , n4479 );
nand ( n6105 , n6104 , n195 );
nor ( n6106 , n6102 , n6103 , n6105 );
nand ( n6107 , n6100 , n6106 );
nand ( n6108 , n4491 , n192 );
nand ( n6109 , n6108 , n6088 );
or ( n6110 , n6109 , n4402 );
nand ( n6111 , n6110 , n4539 );
not ( n6112 , n4540 );
not ( n6113 , n4424 );
nand ( n6114 , n6112 , n6113 );
nand ( n6115 , n6111 , n6114 );
nor ( n6116 , n6107 , n6115 );
nand ( n6117 , n6087 , n6116 );
not ( n6118 , n6117 );
or ( n6119 , n6072 , n6118 );
not ( n6120 , n190 );
not ( n6121 , n6109 );
or ( n6122 , n6120 , n6121 );
not ( n6123 , n5545 );
nand ( n6124 , n6123 , n4404 );
nand ( n6125 , n6122 , n6124 );
nand ( n6126 , n6125 , n4393 );
and ( n6127 , n4563 , n4480 );
and ( n6128 , n6126 , n6127 );
nor ( n6129 , n6128 , n4538 );
not ( n6130 , n4413 );
nand ( n6131 , n4515 , n4409 );
not ( n6132 , n4509 );
nand ( n6133 , n6132 , n4388 );
nor ( n6134 , n6131 , n6133 );
or ( n6135 , n6134 , n4576 );
nand ( n6136 , n6135 , n6035 );
not ( n6137 , n6136 );
or ( n6138 , n6130 , n6137 );
or ( n6139 , n4548 , n4412 );
nand ( n6140 , n4614 , n4496 );
nand ( n6141 , n6139 , n6140 );
or ( n6142 , n6048 , n6141 );
nand ( n6143 , n6142 , n4604 );
nand ( n6144 , n6138 , n6143 );
or ( n6145 , n4493 , n5549 );
nand ( n6146 , n6145 , n4451 );
not ( n6147 , n4433 );
nor ( n6148 , n4446 , n193 );
nand ( n6149 , n6147 , n6148 );
not ( n6150 , n4610 );
nand ( n6151 , n6150 , n4621 );
nand ( n6152 , n6146 , n6149 , n6151 );
nor ( n6153 , n6129 , n6144 , n6152 );
nand ( n6154 , n6119 , n6153 );
not ( n6155 , n6154 );
not ( n6156 , n6155 );
not ( n6157 , n6156 );
not ( n6158 , n5580 );
and ( n6159 , n6158 , n194 );
and ( n6160 , n6140 , n4605 );
nor ( n6161 , n6159 , n6160 );
and ( n6162 , n5558 , n4618 );
nor ( n6163 , n6162 , n189 );
nor ( n6164 , n6161 , n6163 , n5592 );
not ( n6165 , n5566 );
nand ( n6166 , n6165 , n6113 );
not ( n6167 , n4404 );
nand ( n6168 , n6082 , n6167 );
nand ( n6169 , n6166 , n6168 );
or ( n6170 , n5621 , n6169 );
nand ( n6171 , n6170 , n4390 );
nand ( n6172 , n6171 , n4419 );
not ( n6173 , n4432 );
nand ( n6174 , n4445 , n6173 );
not ( n6175 , n6174 );
not ( n6176 , n5568 );
or ( n6177 , n6175 , n6176 );
nand ( n6178 , n6177 , n193 );
nand ( n6179 , n6178 , n4604 );
nor ( n6180 , n6172 , n6179 );
or ( n6181 , n6164 , n6180 );
not ( n6182 , n190 );
nor ( n6183 , n6182 , n4626 );
nand ( n6184 , n4390 , n6183 , n188 );
nand ( n6185 , n6181 , n6184 );
not ( n6186 , n6185 );
nor ( n6187 , n4444 , n4547 );
not ( n6188 , n6187 );
nand ( n6189 , n6188 , n6096 );
or ( n6190 , n4385 , n6189 );
nand ( n6191 , n6190 , n193 );
not ( n6192 , n4445 );
not ( n6193 , n4479 );
or ( n6194 , n6192 , n6193 );
nand ( n6195 , n6194 , n4576 );
not ( n6196 , n189 );
nand ( n6197 , n6196 , n4584 );
not ( n6198 , n6197 );
nor ( n6199 , n6195 , n6198 );
nand ( n6200 , n6191 , n6199 );
or ( n6201 , n5513 , n4518 , n4576 );
not ( n6202 , n6201 );
not ( n6203 , n4538 );
or ( n6204 , n6202 , n6203 );
nand ( n6205 , n6204 , n4442 );
nand ( n6206 , n6200 , n6205 );
not ( n6207 , n6206 );
not ( n6208 , n4556 );
nand ( n6209 , n6208 , n190 );
and ( n6210 , n4637 , n5497 , n6209 , n193 );
not ( n6211 , n4486 );
nand ( n6212 , n6211 , n6092 );
or ( n6213 , n6212 , n193 );
not ( n6214 , n6046 );
nand ( n6215 , n6213 , n6214 );
and ( n6216 , n6029 , n6215 , n6104 );
or ( n6217 , n6210 , n6216 );
nand ( n6218 , n5544 , n195 );
nor ( n6219 , n4433 , n191 );
nor ( n6220 , n6218 , n6219 );
nand ( n6221 , n6217 , n6220 );
not ( n6222 , n4521 );
not ( n6223 , n192 );
and ( n6224 , n6222 , n6223 );
and ( n6225 , n6073 , n192 );
nor ( n6226 , n6224 , n6225 );
and ( n6227 , n6205 , n6226 );
nor ( n6228 , n6221 , n6227 );
not ( n6229 , n6228 );
or ( n6230 , n6207 , n6229 );
not ( n6231 , n5608 );
not ( n6232 , n6231 );
or ( n6233 , n4392 , n6131 );
nand ( n6234 , n6233 , n4393 );
not ( n6235 , n6234 );
or ( n6236 , n6232 , n6235 );
not ( n6237 , n4545 );
not ( n6238 , n6214 );
and ( n6239 , n6237 , n6238 );
not ( n6240 , n4479 );
not ( n6241 , n5526 );
and ( n6242 , n6241 , n193 );
not ( n6243 , n6242 );
or ( n6244 , n6240 , n6243 );
not ( n6245 , n194 );
not ( n6246 , n4627 );
or ( n6247 , n6245 , n6246 );
nand ( n6248 , n5545 , n194 );
or ( n6249 , n6248 , n6183 );
nand ( n6250 , n6247 , n6249 );
nand ( n6251 , n6244 , n6250 );
nor ( n6252 , n6239 , n6251 );
nand ( n6253 , n4394 , n6252 );
nand ( n6254 , n6236 , n6253 );
nand ( n6255 , n6148 , n4467 );
nand ( n6256 , n4451 , n4496 , n5526 );
nand ( n6257 , n4496 , n6241 , n4390 );
nand ( n6258 , n6255 , n6256 , n6257 , n4415 );
not ( n6259 , n4397 );
not ( n6260 , n6147 );
or ( n6261 , n6259 , n6260 );
not ( n6262 , n6103 );
nand ( n6263 , n6261 , n6262 );
nor ( n6264 , n6124 , n4417 );
nor ( n6265 , n6258 , n6263 , n6264 );
nand ( n6266 , n6254 , n6265 );
nand ( n6267 , n6230 , n6266 );
nand ( n6268 , n6186 , n6267 );
not ( n6269 , n6268 );
and ( n6270 , n6157 , n6269 );
not ( n6271 , n6154 );
not ( n6272 , n6271 );
and ( n6273 , n6272 , n6268 );
nor ( n6274 , n6270 , n6273 );
xnor ( n6275 , n6028 , n6274 );
or ( n6276 , n6026 , n6275 );
xnor ( n6277 , n367 , n368 );
or ( n6278 , n6277 , n2246 );
not ( n6279 , n6025 );
nand ( n6280 , n6279 , n6275 , n2246 );
nand ( n6281 , n6276 , n6278 , n6280 );
not ( n6282 , n21 );
nand ( n6283 , n6282 , n20 );
not ( n6284 , n6283 );
nand ( n6285 , n6284 , n22 );
not ( n6286 , n6285 );
not ( n6287 , n24 );
nand ( n6288 , n6286 , n6287 );
not ( n6289 , n24 );
nor ( n6290 , n6289 , n20 );
and ( n6291 , n6290 , n21 , n22 );
not ( n6292 , n6291 );
nand ( n6293 , n6288 , n6292 );
nand ( n6294 , n21 , n24 );
not ( n6295 , n6294 );
not ( n6296 , n20 );
nand ( n6297 , n6295 , n23 , n6296 );
buf ( n6298 , n6297 );
not ( n6299 , n25 );
nand ( n6300 , n6298 , n6299 );
or ( n6301 , n6293 , n6300 );
not ( n6302 , n22 );
nand ( n6303 , n6302 , n21 );
not ( n6304 , n6303 );
nand ( n6305 , n20 , n24 );
not ( n6306 , n6305 );
nand ( n6307 , n6304 , n6306 );
nand ( n6308 , n6307 , n25 );
nand ( n6309 , n6301 , n6308 );
nor ( n6310 , n20 , n21 );
not ( n6311 , n6310 );
nor ( n6312 , n6311 , n22 );
buf ( n6313 , n6312 );
nand ( n6314 , n23 , n25 );
not ( n6315 , n6314 );
and ( n6316 , n6313 , n6315 );
not ( n6317 , n6305 );
nor ( n6318 , n22 , n23 );
nand ( n6319 , n6317 , n6318 );
not ( n6320 , n26 );
and ( n6321 , n6319 , n6320 );
not ( n6322 , n6321 );
not ( n6323 , n20 );
nand ( n6324 , n6323 , n21 );
not ( n6325 , n6324 );
not ( n6326 , n6325 );
not ( n6327 , n6326 );
nand ( n6328 , n22 , n23 );
not ( n6329 , n6328 );
buf ( n6330 , n6329 );
nand ( n6331 , n6327 , n6330 );
not ( n6332 , n6331 );
nor ( n6333 , n6316 , n6322 , n6332 );
nand ( n6334 , n6309 , n6333 );
not ( n6335 , n6334 );
nor ( n6336 , n20 , n21 );
and ( n6337 , n6336 , n6287 );
nand ( n6338 , n6337 , n22 );
nand ( n6339 , n25 , n26 );
not ( n6340 , n6339 );
not ( n6341 , n6310 );
not ( n6342 , n6341 );
not ( n6343 , n23 );
nand ( n6344 , n6342 , n6343 );
not ( n6345 , n6344 );
not ( n6346 , n6297 );
or ( n6347 , n6345 , n6346 );
not ( n6348 , n22 );
nand ( n6349 , n6347 , n6348 );
and ( n6350 , n6338 , n6340 , n6349 );
not ( n6351 , n23 );
nor ( n6352 , n6351 , n22 );
nand ( n6353 , n6352 , n24 );
not ( n6354 , n6353 );
nand ( n6355 , n6354 , n6342 );
not ( n6356 , n25 );
nand ( n6357 , n6355 , n6356 );
not ( n6358 , n6357 );
and ( n6359 , n26 , n6358 );
nor ( n6360 , n6350 , n6359 );
not ( n6361 , n6360 );
or ( n6362 , n6335 , n6361 );
nand ( n6363 , n6329 , n21 );
not ( n6364 , n6363 );
nand ( n6365 , n6364 , n6356 );
not ( n6366 , n24 );
nor ( n6367 , n6366 , n20 );
not ( n6368 , n6367 );
nor ( n6369 , n6365 , n6368 );
not ( n6370 , n6369 );
not ( n6371 , n23 );
nor ( n6372 , n6371 , n24 );
nand ( n6373 , n6284 , n6372 );
not ( n6374 , n6373 );
nand ( n6375 , n22 , n25 );
not ( n6376 , n6375 );
and ( n6377 , n6374 , n6376 );
and ( n6378 , n6310 , n6318 );
nand ( n6379 , n6378 , n6287 );
not ( n6380 , n6379 );
nor ( n6381 , n6377 , n6380 );
buf ( n6382 , n6337 );
not ( n6383 , n25 );
nor ( n6384 , n6383 , n23 );
and ( n6385 , n6382 , n6384 );
not ( n6386 , n6385 );
and ( n6387 , n6370 , n6381 , n6386 );
nand ( n6388 , n6362 , n6387 );
not ( n6389 , n6388 );
not ( n6390 , n20 );
not ( n6391 , n21 );
nor ( n6392 , n6391 , n24 );
nand ( n6393 , n6390 , n6392 );
not ( n6394 , n6393 );
and ( n6395 , n6394 , n6315 );
not ( n6396 , n6395 );
nand ( n6397 , n6396 , n19 );
not ( n6398 , n6397 );
nand ( n6399 , n6367 , n6304 );
not ( n6400 , n6399 );
nand ( n6401 , n20 , n21 );
not ( n6402 , n6401 );
nor ( n6403 , n23 , n24 );
nand ( n6404 , n6402 , n6403 );
nor ( n6405 , n6404 , n22 );
or ( n6406 , n6400 , n6286 , n6405 );
nand ( n6407 , n6406 , n6340 );
not ( n6408 , n25 );
nor ( n6409 , n6408 , n24 );
and ( n6410 , n6284 , n6409 );
nor ( n6411 , n6363 , n6299 );
not ( n6412 , n6403 );
not ( n6413 , n20 );
nor ( n6414 , n6413 , n22 );
nor ( n6415 , n6412 , n6414 , n25 );
or ( n6416 , n6410 , n6411 , n6415 );
or ( n6417 , n25 , n26 );
and ( n6418 , n6417 , n6339 );
nand ( n6419 , n6416 , n6418 );
nand ( n6420 , n6312 , n6287 );
buf ( n6421 , n6420 );
not ( n6422 , n6421 );
not ( n6423 , n23 );
nand ( n6424 , n6423 , n22 );
not ( n6425 , n6424 );
nand ( n6426 , n6425 , n20 );
not ( n6427 , n6426 );
and ( n6428 , n21 , n24 );
nand ( n6429 , n6427 , n6428 );
not ( n6430 , n21 );
and ( n6431 , n6329 , n6430 );
nand ( n6432 , n6431 , n20 );
nand ( n6433 , n6429 , n6432 );
not ( n6434 , n6433 );
not ( n6435 , n6434 );
or ( n6436 , n6422 , n6435 );
nand ( n6437 , n6436 , n25 );
nand ( n6438 , n6398 , n6407 , n6419 , n6437 );
and ( n6439 , n6336 , n24 );
buf ( n6440 , n6439 );
nand ( n6441 , n6440 , n6343 );
nor ( n6442 , n21 , n22 );
buf ( n6443 , n6442 );
nand ( n6444 , n6443 , n6306 );
buf ( n6445 , n6444 );
nand ( n6446 , n6441 , n6445 , n6320 );
not ( n6447 , n26 );
nand ( n6448 , n6447 , n25 );
nand ( n6449 , n6446 , n6448 );
nor ( n6450 , n21 , n24 );
nand ( n6451 , n6450 , n22 );
not ( n6452 , n6451 );
not ( n6453 , n25 );
nand ( n6454 , n6453 , n23 );
not ( n6455 , n6454 );
and ( n6456 , n6452 , n6455 );
not ( n6457 , n6303 );
and ( n6458 , n6457 , n6299 );
buf ( n6459 , n6458 );
not ( n6460 , n20 );
nor ( n6461 , n6460 , n24 );
buf ( n6462 , n6461 );
and ( n6463 , n6459 , n6462 );
nor ( n6464 , n6456 , n6463 );
nand ( n6465 , n6449 , n6464 , n6292 );
buf ( n6466 , n6424 );
not ( n6467 , n6466 );
nand ( n6468 , n6467 , n6367 );
nand ( n6469 , n6445 , n26 , n6468 );
buf ( n6470 , n6339 );
nand ( n6471 , n6469 , n6470 );
not ( n6472 , n23 );
nor ( n6473 , n6472 , n6294 );
nand ( n6474 , n6473 , n6348 );
buf ( n6475 , n6474 );
not ( n6476 , n20 );
nand ( n6477 , n6476 , n6329 );
not ( n6478 , n6477 );
not ( n6479 , n24 );
nor ( n6480 , n6479 , n21 );
not ( n6481 , n6480 );
not ( n6482 , n6481 );
nand ( n6483 , n6478 , n6482 );
nand ( n6484 , n6471 , n6475 , n6483 );
and ( n6485 , n6465 , n6484 );
or ( n6486 , n6438 , n6485 );
not ( n6487 , n6421 );
nand ( n6488 , n6487 , n6470 );
nand ( n6489 , n6428 , n22 );
not ( n6490 , n22 );
nand ( n6491 , n6490 , n6450 );
nand ( n6492 , n6489 , n6491 );
not ( n6493 , n6384 );
not ( n6494 , n6493 );
nand ( n6495 , n6492 , n6494 );
nand ( n6496 , n6329 , n6306 );
nor ( n6497 , n6496 , n21 );
not ( n6498 , n6497 );
nand ( n6499 , n6488 , n6495 , n6498 , n26 );
not ( n6500 , n6499 );
nand ( n6501 , n6440 , n6315 );
nand ( n6502 , n6501 , n6320 );
not ( n6503 , n6502 );
not ( n6504 , n6445 );
not ( n6505 , n20 );
nand ( n6506 , n6505 , n21 , n6343 );
nor ( n6507 , n6506 , n22 );
nor ( n6508 , n6504 , n6507 );
not ( n6509 , n23 );
nor ( n6510 , n6509 , n22 );
or ( n6511 , n6427 , n6510 );
not ( n6512 , n21 );
nor ( n6513 , n6512 , n24 );
nand ( n6514 , n6511 , n6513 );
nand ( n6515 , n6503 , n6508 , n6365 , n6514 );
not ( n6516 , n6515 );
or ( n6517 , n6500 , n6516 );
nand ( n6518 , n6284 , n24 );
not ( n6519 , n6518 );
nand ( n6520 , n6519 , n22 );
nor ( n6521 , n23 , n25 );
not ( n6522 , n6521 );
nor ( n6523 , n6520 , n6522 );
not ( n6524 , n23 );
nor ( n6525 , n6524 , n24 );
not ( n6526 , n6525 );
nor ( n6527 , n6342 , n6526 );
nand ( n6528 , n20 , n21 );
not ( n6529 , n6528 );
not ( n6530 , n6529 );
nand ( n6531 , n6530 , n22 );
buf ( n6532 , n6531 );
and ( n6533 , n6527 , n6532 );
nor ( n6534 , n20 , n24 );
buf ( n6535 , n6534 );
and ( n6536 , n6467 , n6535 );
nor ( n6537 , n6533 , n6536 );
or ( n6538 , n6537 , n25 );
not ( n6539 , n19 );
nand ( n6540 , n6538 , n6539 );
and ( n6541 , n6348 , n6534 );
not ( n6542 , n6541 );
buf ( n6543 , n6528 );
not ( n6544 , n24 );
nand ( n6545 , n6544 , n22 );
nor ( n6546 , n6543 , n6545 );
not ( n6547 , n6546 );
and ( n6548 , n6542 , n6547 );
nor ( n6549 , n6548 , n6493 );
nor ( n6550 , n6523 , n6540 , n6549 );
nand ( n6551 , n6517 , n6550 );
nand ( n6552 , n6486 , n6551 );
nand ( n6553 , n6389 , n6552 );
buf ( n6554 , n6553 );
not ( n6555 , n6554 );
not ( n6556 , n6555 );
not ( n6557 , n6339 );
nand ( n6558 , n6373 , n6477 , n26 );
not ( n6559 , n6558 );
or ( n6560 , n6557 , n6559 );
not ( n6561 , n6529 );
nor ( n6562 , n6561 , n6545 );
nand ( n6563 , n6562 , n6343 );
nand ( n6564 , n6560 , n6563 );
not ( n6565 , n6564 );
and ( n6566 , n6461 , n22 );
nand ( n6567 , n6566 , n6384 );
and ( n6568 , n6567 , n6297 );
and ( n6569 , n6565 , n6568 );
nor ( n6570 , n6458 , n26 );
not ( n6571 , n6341 );
not ( n6572 , n6363 );
or ( n6573 , n6571 , n6572 );
nand ( n6574 , n6573 , n6409 );
and ( n6575 , n6474 , n6570 , n6574 );
nor ( n6576 , n6569 , n6575 );
not ( n6577 , n6401 );
nand ( n6578 , n6577 , n24 );
nand ( n6579 , n6348 , n6480 );
nand ( n6580 , n6578 , n6579 );
nand ( n6581 , n6580 , n6343 );
nor ( n6582 , n6497 , n19 );
and ( n6583 , n6581 , n6582 , n6338 );
and ( n6584 , n6539 , n25 );
or ( n6585 , n6583 , n6584 );
nor ( n6586 , n6578 , n6348 );
not ( n6587 , n6586 );
nand ( n6588 , n6439 , n22 );
nand ( n6589 , n6587 , n6588 , n6420 );
nand ( n6590 , n6589 , n6315 );
nand ( n6591 , n6585 , n6590 );
or ( n6592 , n6576 , n6591 );
not ( n6593 , n22 );
nand ( n6594 , n6593 , n6529 );
not ( n6595 , n6594 );
nand ( n6596 , n6290 , n22 );
not ( n6597 , n6596 );
or ( n6598 , n6595 , n6597 );
nand ( n6599 , n6598 , n6343 );
nand ( n6600 , n6599 , n6447 );
nor ( n6601 , n6518 , n6348 );
nor ( n6602 , n6600 , n6601 );
not ( n6603 , n6401 );
nand ( n6604 , n6603 , n6352 );
nand ( n6605 , n6604 , n25 );
nor ( n6606 , n22 , n23 );
nand ( n6607 , n6284 , n6606 );
not ( n6608 , n6607 );
nor ( n6609 , n6605 , n6608 );
not ( n6610 , n6329 );
not ( n6611 , n6461 );
or ( n6612 , n6610 , n6611 );
nand ( n6613 , n6325 , n6343 );
nand ( n6614 , n6612 , n6613 );
and ( n6615 , n6614 , n6513 );
or ( n6616 , n6609 , n6615 );
nand ( n6617 , n6616 , n6417 );
or ( n6618 , n6602 , n6617 );
not ( n6619 , n6461 );
nor ( n6620 , n6619 , n22 );
nand ( n6621 , n6620 , n6315 );
and ( n6622 , n6284 , n6521 );
nand ( n6623 , n6622 , n22 );
not ( n6624 , n6466 );
not ( n6625 , n6481 );
nand ( n6626 , n6624 , n6625 );
and ( n6627 , n6621 , n6623 , n6626 , n19 );
nand ( n6628 , n6618 , n6627 );
nand ( n6629 , n6592 , n6628 );
not ( n6630 , n6363 );
nand ( n6631 , n6630 , n6462 );
nand ( n6632 , n6631 , n25 );
not ( n6633 , n6305 );
nand ( n6634 , n6633 , n22 );
or ( n6635 , n6634 , n23 );
not ( n6636 , n6341 );
nand ( n6637 , n6636 , n6525 );
nand ( n6638 , n6635 , n6637 );
or ( n6639 , n6632 , n6638 );
nand ( n6640 , n6519 , n6606 );
not ( n6641 , n6450 );
nor ( n6642 , n6641 , n6477 );
nor ( n6643 , n6642 , n25 );
nand ( n6644 , n6640 , n6643 );
nand ( n6645 , n6639 , n6644 , n6470 );
nand ( n6646 , n6629 , n6645 );
not ( n6647 , n6646 );
nand ( n6648 , n6459 , n6525 );
not ( n6649 , n6466 );
nand ( n6650 , n6649 , n6428 );
not ( n6651 , n6522 );
nand ( n6652 , n6651 , n6580 );
and ( n6653 , n6648 , n6650 , n6652 , n6447 );
not ( n6654 , n6653 );
and ( n6655 , n6457 , n6403 );
not ( n6656 , n6655 );
not ( n6657 , n6656 );
not ( n6658 , n6356 );
and ( n6659 , n6657 , n6658 );
nand ( n6660 , n6624 , n6284 );
not ( n6661 , n6660 );
nor ( n6662 , n6659 , n6661 );
nand ( n6663 , n6444 , n6634 );
nor ( n6664 , n6531 , n6367 );
or ( n6665 , n6663 , n6664 );
nand ( n6666 , n6665 , n6356 );
nand ( n6667 , n6354 , n6296 );
nand ( n6668 , n6662 , n6666 , n6667 );
buf ( n6669 , n6622 );
or ( n6670 , n6668 , n6669 );
nand ( n6671 , n6670 , n19 );
not ( n6672 , n6671 );
or ( n6673 , n6654 , n6672 );
nand ( n6674 , n6414 , n6450 );
nand ( n6675 , n6307 , n6674 );
buf ( n6676 , n6457 );
nor ( n6677 , n6676 , n6368 );
or ( n6678 , n6675 , n6677 );
not ( n6679 , n6454 );
nand ( n6680 , n6678 , n6679 );
nand ( n6681 , n6680 , n26 );
not ( n6682 , n6681 );
not ( n6683 , n6466 );
not ( n6684 , n6393 );
and ( n6685 , n6683 , n6684 );
not ( n6686 , n6307 );
and ( n6687 , n6686 , n6343 );
nor ( n6688 , n6685 , n6687 );
nand ( n6689 , n6439 , n6606 );
not ( n6690 , n6689 );
nor ( n6691 , n6518 , n6343 );
nor ( n6692 , n6690 , n6691 );
nand ( n6693 , n6414 , n6392 );
nand ( n6694 , n6688 , n6692 , n6693 );
nand ( n6695 , n6694 , n25 );
nand ( n6696 , n6682 , n6695 );
nand ( n6697 , n6673 , n6696 );
nand ( n6698 , n6647 , n6697 );
not ( n6699 , n6698 );
not ( n6700 , n6699 );
not ( n6701 , n28 );
nand ( n6702 , n6701 , n29 );
not ( n6703 , n6702 );
not ( n6704 , n30 );
nand ( n6705 , n6703 , n6704 );
not ( n6706 , n27 );
nor ( n6707 , n6705 , n6706 );
not ( n6708 , n28 );
not ( n6709 , n29 );
nor ( n6710 , n6709 , n27 );
not ( n6711 , n6710 );
or ( n6712 , n6708 , n6711 );
not ( n6713 , n30 );
nor ( n6714 , n6713 , n28 );
nor ( n6715 , n27 , n29 );
nand ( n6716 , n6714 , n6715 );
nand ( n6717 , n6712 , n6716 );
or ( n6718 , n6707 , n6717 );
not ( n6719 , n31 );
nand ( n6720 , n6718 , n6719 );
not ( n6721 , n29 );
nand ( n6722 , n6721 , n30 , n28 );
not ( n6723 , n6722 );
nand ( n6724 , n6723 , n31 );
not ( n6725 , n30 );
nand ( n6726 , n6725 , n28 );
not ( n6727 , n6726 );
not ( n6728 , n29 );
nor ( n6729 , n6728 , n27 );
nand ( n6730 , n6727 , n6729 );
and ( n6731 , n6724 , n6730 );
nand ( n6732 , n6720 , n6731 );
and ( n6733 , n6732 , n32 );
not ( n6734 , n28 );
nor ( n6735 , n6734 , n27 );
nor ( n6736 , n29 , n30 );
nand ( n6737 , n6735 , n6736 );
nand ( n6738 , n28 , n30 );
not ( n6739 , n6738 );
nand ( n6740 , n6729 , n6739 );
nand ( n6741 , n6737 , n6740 );
not ( n6742 , n6741 );
not ( n6743 , n30 );
nor ( n6744 , n6743 , n28 );
not ( n6745 , n6744 );
nor ( n6746 , n6745 , n6710 );
not ( n6747 , n6746 );
and ( n6748 , n6742 , n6747 );
not ( n6749 , n32 );
nand ( n6750 , n6749 , n31 );
nor ( n6751 , n6748 , n6750 );
or ( n6752 , n6733 , n6751 );
nand ( n6753 , n6752 , n33 );
not ( n6754 , n30 );
not ( n6755 , n27 );
nor ( n6756 , n6755 , n31 );
and ( n6757 , n6756 , n28 );
not ( n6758 , n6757 );
or ( n6759 , n6754 , n6758 );
nor ( n6760 , n28 , n29 );
buf ( n6761 , n6760 );
not ( n6762 , n30 );
nand ( n6763 , n6762 , n31 );
not ( n6764 , n6763 );
nand ( n6765 , n6761 , n6764 );
nand ( n6766 , n6759 , n6765 );
nand ( n6767 , n27 , n31 );
not ( n6768 , n6767 );
nand ( n6769 , n6768 , n29 );
nor ( n6770 , n6769 , n6726 );
or ( n6771 , n6766 , n6770 );
not ( n6772 , n33 );
and ( n6773 , n6772 , n32 );
nand ( n6774 , n6771 , n6773 );
nor ( n6775 , n27 , n29 );
nand ( n6776 , n6739 , n6775 );
nor ( n6777 , n6776 , n31 );
not ( n6778 , n28 );
and ( n6779 , n6768 , n6778 );
and ( n6780 , n6779 , n6736 );
or ( n6781 , n6777 , n6780 );
not ( n6782 , n32 );
nand ( n6783 , n6781 , n6782 );
not ( n6784 , n27 );
not ( n6785 , n30 );
nor ( n6786 , n6785 , n29 );
nand ( n6787 , n6784 , n6786 );
not ( n6788 , n6787 );
nand ( n6789 , n28 , n29 );
not ( n6790 , n6789 );
nand ( n6791 , n6790 , n30 );
not ( n6792 , n6791 );
or ( n6793 , n6788 , n6792 );
nor ( n6794 , n31 , n32 );
nand ( n6795 , n6793 , n6794 );
not ( n6796 , n6795 );
not ( n6797 , n29 );
nor ( n6798 , n6797 , n30 , n27 );
not ( n6799 , n6750 );
and ( n6800 , n6798 , n6799 );
nand ( n6801 , n29 , n30 );
not ( n6802 , n6801 );
and ( n6803 , n6756 , n6802 );
nor ( n6804 , n6800 , n6803 );
not ( n6805 , n6804 );
or ( n6806 , n6796 , n6805 );
not ( n6807 , n33 );
nand ( n6808 , n6806 , n6807 );
and ( n6809 , n6774 , n6783 , n6808 );
nand ( n6810 , n6753 , n6809 );
not ( n6811 , n6810 );
not ( n6812 , n34 );
and ( n6813 , n6795 , n6812 );
nor ( n6814 , n28 , n29 );
nand ( n6815 , n30 , n6814 );
not ( n6816 , n6815 );
nand ( n6817 , n6816 , n27 );
not ( n6818 , n28 );
nand ( n6819 , n6818 , n6715 );
nor ( n6820 , n6819 , n30 );
not ( n6821 , n6820 );
nand ( n6822 , n6817 , n6821 );
not ( n6823 , n6791 );
nand ( n6824 , n6823 , n27 );
not ( n6825 , n6824 );
or ( n6826 , n6822 , n6825 );
nand ( n6827 , n31 , n32 );
not ( n6828 , n6827 );
nand ( n6829 , n6826 , n6828 );
nand ( n6830 , n6813 , n6829 );
not ( n6831 , n27 );
nor ( n6832 , n6831 , n30 );
nand ( n6833 , n6761 , n6832 );
not ( n6834 , n6722 );
nand ( n6835 , n27 , n31 );
buf ( n6836 , n6835 );
not ( n6837 , n6836 );
nand ( n6838 , n6834 , n6837 );
and ( n6839 , n6833 , n6838 );
nor ( n6840 , n6839 , n32 );
nor ( n6841 , n6830 , n6840 );
not ( n6842 , n6841 );
not ( n6843 , n29 );
nor ( n6844 , n6843 , n30 );
nand ( n6845 , n6757 , n6844 );
not ( n6846 , n6702 );
and ( n6847 , n30 , n31 );
nand ( n6848 , n6846 , n6847 );
buf ( n6849 , n6848 );
nand ( n6850 , n6845 , n6849 );
not ( n6851 , n6763 );
not ( n6852 , n6851 );
not ( n6853 , n29 );
nand ( n6854 , n6853 , n28 );
not ( n6855 , n6854 );
not ( n6856 , n6855 );
or ( n6857 , n6852 , n6856 );
nand ( n6858 , n6857 , n6782 );
not ( n6859 , n6858 );
not ( n6860 , n6835 );
nand ( n6861 , n6778 , n6860 );
nand ( n6862 , n6861 , n33 );
not ( n6863 , n6862 );
and ( n6864 , n6859 , n6863 );
not ( n6865 , n6756 );
not ( n6866 , n6865 );
nand ( n6867 , n6727 , n6866 );
nand ( n6868 , n32 , n33 );
not ( n6869 , n6868 );
and ( n6870 , n6867 , n6869 );
nor ( n6871 , n6864 , n6870 );
or ( n6872 , n6850 , n6871 );
nand ( n6873 , n6802 , n31 );
nor ( n6874 , n6873 , n27 );
not ( n6875 , n6874 );
not ( n6876 , n31 );
not ( n6877 , n30 );
nand ( n6878 , n6877 , n29 );
nor ( n6879 , n6876 , n6878 );
and ( n6880 , n27 , n32 );
nand ( n6881 , n6879 , n6880 );
not ( n6882 , n32 );
and ( n6883 , n6729 , n6882 );
not ( n6884 , n6883 );
nand ( n6885 , n6875 , n6881 , n6884 , n6807 );
and ( n6886 , n6761 , n6704 );
nand ( n6887 , n6886 , n32 );
not ( n6888 , n6887 );
or ( n6889 , n6885 , n6888 );
nand ( n6890 , n6872 , n6889 );
not ( n6891 , n6890 );
or ( n6892 , n6842 , n6891 );
nand ( n6893 , n6745 , n27 );
nor ( n6894 , n6789 , n30 );
nor ( n6895 , n6893 , n6894 );
not ( n6896 , n6895 );
not ( n6897 , n6865 );
nand ( n6898 , n6897 , n6855 );
nand ( n6899 , n6898 , n32 );
not ( n6900 , n6899 );
or ( n6901 , n6896 , n6900 );
not ( n6902 , n6858 );
buf ( n6903 , n6855 );
nand ( n6904 , n6902 , n6903 );
nand ( n6905 , n6901 , n6904 );
not ( n6906 , n31 );
nor ( n6907 , n6906 , n27 );
nand ( n6908 , n6907 , n30 );
nor ( n6909 , n6908 , n28 );
not ( n6910 , n6909 );
not ( n6911 , n32 );
nor ( n6912 , n6911 , n31 );
nand ( n6913 , n6798 , n6912 );
nand ( n6914 , n6910 , n6913 , n6807 );
nor ( n6915 , n6905 , n6914 );
not ( n6916 , n31 );
not ( n6917 , n6855 );
or ( n6918 , n6916 , n6917 );
not ( n6919 , n6814 );
nor ( n6920 , n6919 , n31 );
not ( n6921 , n6920 );
nand ( n6922 , n6918 , n6921 );
nor ( n6923 , n28 , n30 );
nand ( n6924 , n6923 , n27 );
not ( n6925 , n6735 );
nand ( n6926 , n6924 , n6925 );
or ( n6927 , n6922 , n6926 );
nand ( n6928 , n6927 , n32 );
not ( n6929 , n6928 );
not ( n6930 , n6794 );
not ( n6931 , n6705 );
not ( n6932 , n6931 );
or ( n6933 , n6930 , n6932 );
nand ( n6934 , n6933 , n33 );
nor ( n6935 , n6929 , n6934 , n6770 );
or ( n6936 , n6915 , n6935 );
nor ( n6937 , n27 , n31 );
not ( n6938 , n6789 );
nand ( n6939 , n6937 , n6938 );
nand ( n6940 , n6735 , n6764 );
and ( n6941 , n32 , n34 );
and ( n6942 , n6939 , n6940 , n6941 );
not ( n6943 , n6722 );
nand ( n6944 , n6943 , n27 );
not ( n6945 , n31 );
nand ( n6946 , n6945 , n6714 );
not ( n6947 , n6946 );
nand ( n6948 , n6947 , n27 );
nand ( n6949 , n6942 , n6944 , n6948 );
nand ( n6950 , n6898 , n6782 , n34 );
and ( n6951 , n6949 , n6950 );
not ( n6952 , n6786 );
nor ( n6953 , n6865 , n6952 );
nor ( n6954 , n6951 , n6953 );
nand ( n6955 , n6936 , n6954 );
nand ( n6956 , n6892 , n6955 );
nand ( n6957 , n6811 , n6956 );
not ( n6958 , n6957 );
not ( n6959 , n6958 );
or ( n6960 , n6700 , n6959 );
nand ( n6961 , n6957 , n6698 );
nand ( n6962 , n6960 , n6961 );
not ( n6963 , n6962 );
not ( n6964 , n6963 );
or ( n6965 , n6556 , n6964 );
or ( n6966 , n6963 , n6555 );
nand ( n6967 , n6965 , n6966 );
not ( n6968 , n14 );
nor ( n6969 , n6968 , n12 );
nand ( n6970 , n11 , n15 );
not ( n6971 , n6970 );
and ( n6972 , n6969 , n6971 );
nand ( n6973 , n6972 , n16 );
nand ( n6974 , n14 , n15 );
not ( n6975 , n6974 );
nor ( n6976 , n12 , n13 );
nand ( n6977 , n6975 , n6976 );
not ( n6978 , n17 );
and ( n6979 , n6977 , n6978 );
not ( n6980 , n13 );
nor ( n6981 , n6980 , n14 );
nand ( n6982 , n11 , n12 );
not ( n6983 , n6982 );
buf ( n6984 , n6983 );
nand ( n6985 , n6981 , n6984 );
and ( n6986 , n6973 , n6979 , n6985 );
not ( n6987 , n14 );
nand ( n6988 , n6987 , n11 );
not ( n6989 , n6988 );
nand ( n6990 , n12 , n15 );
not ( n6991 , n6990 );
and ( n6992 , n6989 , n6991 );
not ( n6993 , n13 );
nor ( n6994 , n6993 , n14 );
nand ( n6995 , n6994 , n6971 );
not ( n6996 , n6995 );
not ( n6997 , n11 );
nand ( n6998 , n6997 , n12 );
not ( n6999 , n6998 );
not ( n7000 , n15 );
nand ( n7001 , n7000 , n14 );
not ( n7002 , n7001 );
nand ( n7003 , n6999 , n7002 );
not ( n7004 , n7003 );
or ( n7005 , n6992 , n6996 , n7004 );
not ( n7006 , n16 );
nand ( n7007 , n7005 , n7006 );
nand ( n7008 , n13 , n16 );
not ( n7009 , n7008 );
not ( n7010 , n12 );
nor ( n7011 , n11 , n14 );
not ( n7012 , n7011 );
not ( n7013 , n7012 );
nand ( n7014 , n7010 , n7013 );
not ( n7015 , n7014 );
nand ( n7016 , n7009 , n7015 );
nand ( n7017 , n6986 , n7007 , n7016 );
nor ( n7018 , n14 , n15 );
nand ( n7019 , n6999 , n7018 );
not ( n7020 , n7019 );
not ( n7021 , n6995 );
not ( n7022 , n13 );
nand ( n7023 , n7022 , n7011 );
not ( n7024 , n7023 );
or ( n7025 , n7021 , n7024 );
not ( n7026 , n12 );
nand ( n7027 , n7025 , n7026 );
not ( n7028 , n7027 );
or ( n7029 , n7020 , n7028 );
nand ( n7030 , n7029 , n16 );
not ( n7031 , n15 );
nor ( n7032 , n7031 , n11 );
nand ( n7033 , n7026 , n7032 );
not ( n7034 , n7033 );
not ( n7035 , n14 );
nand ( n7036 , n7034 , n7035 );
not ( n7037 , n16 );
nand ( n7038 , n7037 , n13 );
nor ( n7039 , n7036 , n7038 );
nor ( n7040 , n7039 , n6978 );
nand ( n7041 , n7030 , n7040 );
nand ( n7042 , n7017 , n7041 );
nor ( n7043 , n11 , n14 );
not ( n7044 , n15 );
and ( n7045 , n7043 , n7044 );
nor ( n7046 , n12 , n13 );
nand ( n7047 , n7045 , n7046 );
not ( n7048 , n7038 );
nand ( n7049 , n6992 , n7048 );
not ( n7050 , n16 );
nor ( n7051 , n7050 , n13 );
buf ( n7052 , n7051 );
nand ( n7053 , n7045 , n7052 );
not ( n7054 , n11 );
nand ( n7055 , n7054 , n14 );
not ( n7056 , n7055 );
not ( n7057 , n15 );
nand ( n7058 , n7057 , n13 );
not ( n7059 , n7058 );
nand ( n7060 , n7056 , n7059 );
not ( n7061 , n7060 );
nand ( n7062 , n12 , n16 );
not ( n7063 , n7062 );
nand ( n7064 , n7061 , n7063 );
and ( n7065 , n7047 , n7049 , n7053 , n7064 );
nand ( n7066 , n11 , n14 );
and ( n7067 , n7066 , n12 );
not ( n7068 , n7067 );
not ( n7069 , n7068 );
nor ( n7070 , n7058 , n7013 );
not ( n7071 , n7070 );
or ( n7072 , n7069 , n7071 );
not ( n7073 , n7018 );
not ( n7074 , n7073 );
nand ( n7075 , n7056 , n15 );
buf ( n7076 , n7075 );
not ( n7077 , n7076 );
or ( n7078 , n7074 , n7077 );
not ( n7079 , n13 );
nand ( n7080 , n7079 , n12 );
not ( n7081 , n7080 );
nand ( n7082 , n7078 , n7081 );
nand ( n7083 , n7072 , n7082 );
nor ( n7084 , n10 , n16 );
nand ( n7085 , n7083 , n7084 );
and ( n7086 , n7042 , n7065 , n7085 );
nand ( n7087 , n12 , n13 );
not ( n7088 , n7087 );
and ( n7089 , n7032 , n7035 , n7088 );
not ( n7090 , n13 );
nor ( n7091 , n7090 , n12 );
and ( n7092 , n7091 , n6971 );
nor ( n7093 , n7089 , n7092 );
not ( n7094 , n6969 );
nand ( n7095 , n7094 , n7044 );
not ( n7096 , n7095 );
nor ( n7097 , n13 , n16 );
not ( n7098 , n7097 );
not ( n7099 , n7098 );
nand ( n7100 , n7096 , n7099 );
nand ( n7101 , n7093 , n7100 , n17 );
not ( n7102 , n13 );
nand ( n7103 , n7102 , n14 );
not ( n7104 , n7103 );
not ( n7105 , n15 );
nand ( n7106 , n7105 , n11 );
not ( n7107 , n7106 );
nand ( n7108 , n7104 , n7107 );
nor ( n7109 , n7108 , n12 );
nand ( n7110 , n7056 , n12 );
not ( n7111 , n7110 );
nor ( n7112 , n7109 , n7111 );
and ( n7113 , n6989 , n7026 );
nand ( n7114 , n7113 , n15 );
and ( n7115 , n7112 , n7114 );
not ( n7116 , n16 );
nor ( n7117 , n7115 , n7116 );
or ( n7118 , n7101 , n7117 );
not ( n7119 , n6992 );
nand ( n7120 , n7059 , n6999 );
not ( n7121 , n7120 );
not ( n7122 , n11 );
nor ( n7123 , n7122 , n12 );
nand ( n7124 , n7123 , n7002 );
not ( n7125 , n7124 );
or ( n7126 , n7121 , n7125 );
not ( n7127 , n16 );
nand ( n7128 , n7126 , n7127 );
nand ( n7129 , n7119 , n7128 );
not ( n7130 , n7129 );
not ( n7131 , n17 );
and ( n7132 , n7131 , n16 );
not ( n7133 , n7132 );
nand ( n7134 , n7056 , n7044 );
not ( n7135 , n7134 );
not ( n7136 , n11 );
nor ( n7137 , n7136 , n7087 );
nor ( n7138 , n7135 , n7137 );
not ( n7139 , n7138 );
or ( n7140 , n7133 , n7139 );
and ( n7141 , n7043 , n15 );
not ( n7142 , n13 );
nand ( n7143 , n7141 , n7142 );
nor ( n7144 , n16 , n17 );
nand ( n7145 , n7143 , n7144 );
nand ( n7146 , n7140 , n7145 );
nand ( n7147 , n7130 , n7146 );
nand ( n7148 , n7118 , n7147 );
not ( n7149 , n7148 );
not ( n7150 , n7059 );
not ( n7151 , n6989 );
or ( n7152 , n7150 , n7151 );
nand ( n7153 , n7152 , n16 );
not ( n7154 , n15 );
nor ( n7155 , n7154 , n7066 );
nand ( n7156 , n7155 , n7081 );
nand ( n7157 , n13 , n14 );
not ( n7158 , n7157 );
nand ( n7159 , n7158 , n6999 );
buf ( n7160 , n7159 );
nand ( n7161 , n7156 , n7160 );
not ( n7162 , n7012 );
nor ( n7163 , n12 , n15 );
nand ( n7164 , n7162 , n7163 );
not ( n7165 , n7164 );
or ( n7166 , n7153 , n7161 , n7165 );
not ( n7167 , n6974 );
nor ( n7168 , n11 , n12 );
nand ( n7169 , n7167 , n7168 );
not ( n7170 , n16 );
nand ( n7171 , n7169 , n7170 );
not ( n7172 , n7171 );
not ( n7173 , n14 );
nand ( n7174 , n7173 , n15 );
nor ( n7175 , n13 , n7174 );
nand ( n7176 , n7175 , n12 );
nand ( n7177 , n7172 , n7176 );
nand ( n7178 , n7166 , n7177 );
not ( n7179 , n7178 );
or ( n7180 , n7149 , n7179 );
nand ( n7181 , n7180 , n10 );
not ( n7182 , n7052 );
not ( n7183 , n7182 );
not ( n7184 , n16 );
nand ( n7185 , n7045 , n7184 );
not ( n7186 , n7185 );
or ( n7187 , n7183 , n7186 );
nand ( n7188 , n11 , n15 );
not ( n7189 , n7188 );
nand ( n7190 , n7189 , n12 );
not ( n7191 , n11 );
nor ( n7192 , n12 , n15 );
nand ( n7193 , n7191 , n7192 );
nand ( n7194 , n7190 , n7193 );
nand ( n7195 , n7187 , n7194 );
not ( n7196 , n7159 );
nand ( n7197 , n7196 , n15 );
nand ( n7198 , n7195 , n7197 );
not ( n7199 , n7198 );
not ( n7200 , n17 );
or ( n7201 , n7199 , n7200 );
nor ( n7202 , n7095 , n7067 );
nand ( n7203 , n7202 , n7052 );
nand ( n7204 , n7201 , n7203 );
nand ( n7205 , n6989 , n7026 );
nand ( n7206 , n7002 , n6983 );
nand ( n7207 , n7205 , n7206 );
nand ( n7208 , n7207 , n7142 );
not ( n7209 , n7107 );
not ( n7210 , n13 );
nor ( n7211 , n7210 , n12 );
not ( n7212 , n7211 );
or ( n7213 , n7209 , n7212 );
nand ( n7214 , n7213 , n7169 );
not ( n7215 , n6984 );
nor ( n7216 , n7038 , n7215 );
nor ( n7217 , n7214 , n7216 );
nand ( n7218 , n7141 , n7009 );
and ( n7219 , n7208 , n7217 , n7218 );
nor ( n7220 , n7219 , n17 );
or ( n7221 , n7204 , n7220 );
not ( n7222 , n10 );
nand ( n7223 , n7221 , n7222 );
and ( n7224 , n7086 , n7181 , n7223 );
buf ( n7225 , n7224 );
not ( n7226 , n7225 );
not ( n7227 , n9 );
not ( n7228 , n6 );
nand ( n7229 , n7228 , n2 );
not ( n7230 , n7229 );
nor ( n7231 , n3 , n4 );
buf ( n7232 , n7231 );
nand ( n7233 , n7230 , n7232 );
not ( n7234 , n7233 );
not ( n7235 , n2 );
nand ( n7236 , n7235 , n5 );
not ( n7237 , n7236 );
nand ( n7238 , n7237 , n4 );
not ( n7239 , n7238 );
not ( n7240 , n3 );
nand ( n7241 , n7239 , n7240 );
not ( n7242 , n7241 );
or ( n7243 , n7234 , n7242 );
nand ( n7244 , n7243 , n7 );
not ( n7245 , n7244 );
not ( n7246 , n3 );
nor ( n7247 , n7246 , n4 );
nand ( n7248 , n7247 , n6 );
not ( n7249 , n7248 );
not ( n7250 , n7249 );
not ( n7251 , n5 );
not ( n7252 , n7251 );
or ( n7253 , n7250 , n7252 );
not ( n7254 , n6 );
nand ( n7255 , n7254 , n3 );
nand ( n7256 , n7237 , n7255 );
nor ( n7257 , n5 , n6 );
nand ( n7258 , n7257 , n4 );
nand ( n7259 , n7256 , n7258 );
nand ( n7260 , n5 , n6 );
not ( n7261 , n7260 );
nand ( n7262 , n7261 , n4 );
nand ( n7263 , n7238 , n7262 );
or ( n7264 , n7259 , n7263 );
not ( n7265 , n7 );
nand ( n7266 , n7264 , n7265 );
nand ( n7267 , n7253 , n7266 );
not ( n7268 , n7267 );
not ( n7269 , n7268 );
or ( n7270 , n7245 , n7269 );
not ( n7271 , n8 );
nand ( n7272 , n7270 , n7271 );
nor ( n7273 , n7241 , n7 );
not ( n7274 , n3 );
nand ( n7275 , n7274 , n4 );
not ( n7276 , n7275 );
not ( n7277 , n2 );
nand ( n7278 , n7277 , n6 );
not ( n7279 , n7278 );
nand ( n7280 , n7276 , n7279 );
not ( n7281 , n7280 );
not ( n7282 , n4 );
not ( n7283 , n6 );
nand ( n7284 , n7283 , n5 );
not ( n7285 , n7284 );
nand ( n7286 , n7282 , n7285 );
nand ( n7287 , n3 , n7 );
nor ( n7288 , n7286 , n7287 );
nor ( n7289 , n7273 , n7281 , n7288 );
nor ( n7290 , n3 , n7 );
nand ( n7291 , n7290 , n7230 , n7251 );
not ( n7292 , n7291 );
nand ( n7293 , n2 , n3 );
not ( n7294 , n7293 );
nand ( n7295 , n7294 , n4 );
not ( n7296 , n7295 );
nand ( n7297 , n7296 , n7285 );
not ( n7298 , n7297 );
or ( n7299 , n7292 , n7298 );
nand ( n7300 , n7299 , n8 );
nand ( n7301 , n7272 , n7289 , n7300 );
not ( n7302 , n7301 );
or ( n7303 , n7227 , n7302 );
not ( n7304 , n7240 );
not ( n7305 , n7262 );
not ( n7306 , n7305 );
or ( n7307 , n7304 , n7306 );
or ( n7308 , n2 , n5 );
not ( n7309 , n7308 );
not ( n7310 , n7255 );
nand ( n7311 , n7309 , n7310 );
nand ( n7312 , n7307 , n7311 );
not ( n7313 , n7297 );
or ( n7314 , n7312 , n7313 );
not ( n7315 , n8 );
and ( n7316 , n7315 , n7 );
nand ( n7317 , n7314 , n7316 );
not ( n7318 , n4 );
nor ( n7319 , n7318 , n3 );
nand ( n7320 , n2 , n6 );
not ( n7321 , n7320 );
nand ( n7322 , n7319 , n7321 );
not ( n7323 , n7322 );
nor ( n7324 , n2 , n4 );
nand ( n7325 , n7324 , n6 );
not ( n7326 , n7325 );
nand ( n7327 , n2 , n5 );
not ( n7328 , n7327 );
nand ( n7329 , n7328 , n6 );
not ( n7330 , n7329 );
or ( n7331 , n7326 , n7330 );
nand ( n7332 , n7331 , n7290 );
not ( n7333 , n7332 );
or ( n7334 , n7323 , n7333 );
nand ( n7335 , n7334 , n7271 );
nor ( n7336 , n2 , n5 );
not ( n7337 , n4 );
and ( n7338 , n7336 , n7337 );
nor ( n7339 , n7338 , n7 );
not ( n7340 , n2 );
not ( n7341 , n7260 );
nand ( n7342 , n7340 , n7231 , n7341 );
nand ( n7343 , n7342 , n7311 );
nand ( n7344 , n7339 , n7343 );
not ( n7345 , n4 );
nand ( n7346 , n7345 , n7230 );
not ( n7347 , n7346 );
not ( n7348 , n3 );
nor ( n7349 , n7348 , n7 );
and ( n7350 , n7349 , n7271 );
nand ( n7351 , n7347 , n7350 );
and ( n7352 , n7335 , n7344 , n7351 );
not ( n7353 , n2 );
nand ( n7354 , n7353 , n5 , n6 );
not ( n7355 , n7354 );
nand ( n7356 , n3 , n4 );
not ( n7357 , n7356 );
nand ( n7358 , n7355 , n7357 );
not ( n7359 , n7358 );
not ( n7360 , n6 );
nor ( n7361 , n2 , n5 );
nand ( n7362 , n7360 , n7361 );
not ( n7363 , n7362 );
nand ( n7364 , n7363 , n4 );
not ( n7365 , n7364 );
or ( n7366 , n7359 , n7365 );
nand ( n7367 , n7366 , n7265 );
not ( n7368 , n7367 );
nand ( n7369 , n7247 , n7321 );
not ( n7370 , n7 );
not ( n7371 , n2 );
nor ( n7372 , n7371 , n4 );
nand ( n7373 , n7370 , n7372 );
nand ( n7374 , n7369 , n7373 );
nand ( n7375 , n7230 , n4 );
nor ( n7376 , n7375 , n7287 );
or ( n7377 , n7374 , n7376 );
nand ( n7378 , n7377 , n7271 );
not ( n7379 , n7378 );
or ( n7380 , n7368 , n7379 );
not ( n7381 , n9 );
nand ( n7382 , n7380 , n7381 );
and ( n7383 , n7317 , n7352 , n7382 );
nand ( n7384 , n7303 , n7383 );
or ( n7385 , n7356 , n5 );
not ( n7386 , n7385 );
not ( n7387 , n3 );
nor ( n7388 , n7387 , n6 );
nand ( n7389 , n7237 , n7388 );
not ( n7390 , n7389 );
or ( n7391 , n7386 , n7390 );
nand ( n7392 , n7391 , n7265 );
not ( n7393 , n6 );
nor ( n7394 , n7393 , n5 );
not ( n7395 , n7293 );
nand ( n7396 , n7394 , n7395 );
nand ( n7397 , n7392 , n7396 );
not ( n7398 , n6 );
nand ( n7399 , n7398 , n2 , n5 , n4 );
nor ( n7400 , n7399 , n3 );
nand ( n7401 , n7285 , n4 );
not ( n7402 , n3 );
nand ( n7403 , n7402 , n7 );
nor ( n7404 , n7401 , n7403 );
or ( n7405 , n7397 , n7400 , n7404 );
nand ( n7406 , n7405 , n7381 );
not ( n7407 , n7406 );
not ( n7408 , n7372 );
not ( n7409 , n5 );
nand ( n7410 , n7409 , n6 );
not ( n7411 , n7410 );
nand ( n7412 , n7408 , n7411 );
not ( n7413 , n7412 );
not ( n7414 , n5 );
nor ( n7415 , n7414 , n4 );
nor ( n7416 , n2 , n6 );
nand ( n7417 , n7415 , n7416 );
nand ( n7418 , n7415 , n7321 );
nand ( n7419 , n7417 , n7418 );
not ( n7420 , n7419 );
not ( n7421 , n7420 );
or ( n7422 , n7413 , n7421 );
nand ( n7423 , n7422 , n7349 );
nand ( n7424 , n7372 , n7285 );
not ( n7425 , n7424 );
nand ( n7426 , n7355 , n3 );
not ( n7427 , n7426 );
or ( n7428 , n7425 , n7427 );
nand ( n7429 , n7428 , n7 );
not ( n7430 , n2 );
nand ( n7431 , n7337 , n5 );
nand ( n7432 , n7258 , n7431 );
not ( n7433 , n7432 );
or ( n7434 , n7430 , n7433 );
nor ( n7435 , n2 , n4 );
nand ( n7436 , n7411 , n7435 );
nand ( n7437 , n7434 , n7436 );
not ( n7438 , n7403 );
nand ( n7439 , n7437 , n7438 );
nand ( n7440 , n7423 , n7429 , n7439 );
or ( n7441 , n7407 , n7440 );
nand ( n7442 , n7441 , n8 );
not ( n7443 , n6 );
nor ( n7444 , n7443 , n2 , n5 );
nand ( n7445 , n7444 , n4 );
not ( n7446 , n7329 );
not ( n7447 , n7446 );
nand ( n7448 , n7445 , n7447 );
nor ( n7449 , n7265 , n7356 );
nand ( n7450 , n7448 , n7449 );
not ( n7451 , n7316 );
not ( n7452 , n7362 );
not ( n7453 , n7452 );
or ( n7454 , n7451 , n7453 );
nand ( n7455 , n7454 , n7332 );
not ( n7456 , n7455 );
not ( n7457 , n7287 );
not ( n7458 , n2 );
not ( n7459 , n4 );
nand ( n7460 , n7459 , n7257 );
not ( n7461 , n7460 );
nand ( n7462 , n7457 , n7458 , n7461 );
and ( n7463 , n7450 , n7456 , n7462 );
nor ( n7464 , n7463 , n9 );
not ( n7465 , n7237 );
and ( n7466 , n3 , n7465 );
not ( n7467 , n3 );
and ( n7468 , n7467 , n7308 );
nor ( n7469 , n7466 , n7468 );
or ( n7470 , n7469 , n7432 );
nand ( n7471 , n7470 , n8 );
nand ( n7472 , n7355 , n4 );
nand ( n7473 , n7231 , n2 );
not ( n7474 , n7473 );
not ( n7475 , n7251 );
and ( n7476 , n7474 , n7475 );
and ( n7477 , n7319 , n7394 );
nor ( n7478 , n7476 , n7477 );
and ( n7479 , n7471 , n7472 , n7478 );
nor ( n7480 , n7479 , n7265 , n7381 );
nor ( n7481 , n7464 , n7480 );
nand ( n7482 , n7442 , n7481 );
nor ( n7483 , n7384 , n7482 );
not ( n7484 , n7483 );
buf ( n7485 , n7484 );
not ( n7486 , n7485 );
not ( n7487 , n7486 );
not ( n7488 , n41 );
and ( n7489 , n7487 , n7488 );
not ( n7490 , n7485 );
and ( n7491 , n7490 , n41 );
nor ( n7492 , n7489 , n7491 );
not ( n7493 , n7492 );
or ( n7494 , n7226 , n7493 );
or ( n7495 , n7492 , n7225 );
nand ( n7496 , n7494 , n7495 );
and ( n7497 , n6967 , n7496 );
not ( n7498 , n6967 );
not ( n7499 , n7496 );
and ( n7500 , n7498 , n7499 );
nor ( n7501 , n7497 , n7500 );
or ( n7502 , n7501 , n1 );
xnor ( n7503 , n41 , n42 );
or ( n7504 , n2246 , n7503 );
nand ( n7505 , n7502 , n7504 );
nor ( n7506 , n6985 , n15 );
not ( n7507 , n7506 );
not ( n7508 , n7157 );
not ( n7509 , n15 );
nor ( n7510 , n7509 , n11 );
nand ( n7511 , n7508 , n7510 );
buf ( n7512 , n7174 );
not ( n7513 , n7512 );
nand ( n7514 , n7211 , n7513 );
nand ( n7515 , n7511 , n7514 );
not ( n7516 , n7515 );
nand ( n7517 , n6976 , n11 );
nor ( n7518 , n7517 , n7073 );
nor ( n7519 , n7518 , n7170 );
nand ( n7520 , n7507 , n7516 , n7519 , n7143 );
not ( n7521 , n11 );
nand ( n7522 , n7081 , n7521 );
not ( n7523 , n15 );
nand ( n7524 , n7523 , n14 );
nor ( n7525 , n7522 , n7524 );
not ( n7526 , n7525 );
nand ( n7527 , n13 , n15 );
nor ( n7528 , n7527 , n12 );
not ( n7529 , n7066 );
nand ( n7530 , n7528 , n7529 );
nand ( n7531 , n7184 , n7530 );
not ( n7532 , n7531 );
nand ( n7533 , n7526 , n7532 , n7108 );
nand ( n7534 , n7520 , n7533 );
not ( n7535 , n7534 );
not ( n7536 , n7143 );
nand ( n7537 , n7536 , n7026 );
not ( n7538 , n7197 );
nor ( n7539 , n7538 , n17 );
and ( n7540 , n7537 , n7539 );
not ( n7541 , n7540 );
or ( n7542 , n7535 , n7541 );
nand ( n7543 , n6972 , n7142 );
not ( n7544 , n16 );
nand ( n7545 , n7544 , n17 );
nor ( n7546 , n7070 , n7545 );
nand ( n7547 , n7543 , n7546 );
not ( n7548 , n7047 );
or ( n7549 , n7547 , n7548 );
nand ( n7550 , n7056 , n7081 );
not ( n7551 , n7550 );
and ( n7552 , n16 , n17 );
not ( n7553 , n7552 );
or ( n7554 , n7551 , n7553 );
nand ( n7555 , n7549 , n7554 );
not ( n7556 , n7218 );
not ( n7557 , n7059 );
nor ( n7558 , n7557 , n7205 );
not ( n7559 , n7524 );
and ( n7560 , n7137 , n7559 );
nor ( n7561 , n7556 , n7558 , n7560 );
nand ( n7562 , n7555 , n7561 );
nand ( n7563 , n7542 , n7562 );
not ( n7564 , n10 );
nand ( n7565 , n7045 , n7081 );
nand ( n7566 , n7565 , n17 );
nor ( n7567 , n14 , n15 );
and ( n7568 , n6983 , n7567 );
and ( n7569 , n7170 , n7568 );
not ( n7570 , n7170 );
and ( n7571 , n7570 , n7113 );
nor ( n7572 , n7569 , n7571 );
not ( n7573 , n6981 );
nor ( n7574 , n7573 , n7033 );
not ( n7575 , n7056 );
or ( n7576 , n12 , n16 );
nor ( n7577 , n7575 , n7576 );
nor ( n7578 , n7574 , n7577 );
nand ( n7579 , n7572 , n7578 );
or ( n7580 , n7566 , n7579 );
not ( n7581 , n16 );
not ( n7582 , n6992 );
or ( n7583 , n7581 , n7582 );
not ( n7584 , n7211 );
not ( n7585 , n7529 );
or ( n7586 , n7584 , n7585 );
nand ( n7587 , n7586 , n7131 );
nand ( n7588 , n6999 , n6994 );
nor ( n7589 , n7588 , n16 );
nor ( n7590 , n7587 , n7589 );
nand ( n7591 , n7583 , n7590 );
and ( n7592 , n7142 , n7576 );
buf ( n7593 , n7188 );
nor ( n7594 , n7592 , n7593 );
or ( n7595 , n7591 , n7594 );
nand ( n7596 , n7580 , n7595 );
not ( n7597 , n7596 );
or ( n7598 , n7564 , n7597 );
nand ( n7599 , n7163 , n14 );
not ( n7600 , n7599 );
not ( n7601 , n7588 );
or ( n7602 , n7600 , n7601 );
nand ( n7603 , n7602 , n16 );
not ( n7604 , n15 );
nand ( n7605 , n7604 , n12 );
and ( n7606 , n7605 , n7103 );
nor ( n7607 , n7603 , n7606 );
nor ( n7608 , n7607 , n10 );
nand ( n7609 , n7107 , n7097 );
not ( n7610 , n7609 );
nand ( n7611 , n7610 , n12 , n14 );
and ( n7612 , n7537 , n7608 , n7611 );
nand ( n7613 , n7160 , n17 );
not ( n7614 , n16 );
nand ( n7615 , n6989 , n7614 );
not ( n7616 , n7528 );
nand ( n7617 , n7616 , n7605 );
nor ( n7618 , n7615 , n7617 );
nor ( n7619 , n7613 , n7618 );
not ( n7620 , n7075 );
nand ( n7621 , n7620 , n16 );
nand ( n7622 , n7619 , n7621 );
nand ( n7623 , n7051 , n11 );
nor ( n7624 , n7623 , n7605 );
or ( n7625 , n7622 , n7624 );
not ( n7626 , n17 );
not ( n7627 , n7626 );
not ( n7628 , n7045 );
not ( n7629 , n7628 );
or ( n7630 , n7627 , n7629 );
not ( n7631 , n7144 );
nand ( n7632 , n7630 , n7631 );
nand ( n7633 , n7104 , n7510 );
nor ( n7634 , n7633 , n16 );
and ( n7635 , n6981 , n7168 );
nand ( n7636 , n14 , n15 );
nor ( n7637 , n7636 , n7062 );
nor ( n7638 , n7634 , n7635 , n7637 );
nand ( n7639 , n7632 , n7638 );
nand ( n7640 , n7625 , n7639 );
nand ( n7641 , n7612 , n7640 );
nand ( n7642 , n7598 , n7641 );
not ( n7643 , n7522 );
not ( n7644 , n6981 );
nor ( n7645 , n7644 , n12 );
nor ( n7646 , n6972 , n7643 , n7645 );
not ( n7647 , n7153 );
and ( n7648 , n7646 , n7647 );
not ( n7649 , n7157 );
nand ( n7650 , n7649 , n7168 );
nand ( n7651 , n7649 , n7107 );
and ( n7652 , n7650 , n7651 , n7170 );
and ( n7653 , n7047 , n7652 );
nor ( n7654 , n7648 , n7653 );
nand ( n7655 , n7641 , n7654 );
not ( n7656 , n7637 );
not ( n7657 , n7575 );
nand ( n7658 , n7657 , n7192 );
nand ( n7659 , n7656 , n7658 );
not ( n7660 , n7088 );
nand ( n7661 , n7038 , n7660 );
nand ( n7662 , n7659 , n7661 );
nand ( n7663 , n7563 , n7642 , n7655 , n7662 );
not ( n7664 , n7663 );
not ( n7665 , n7664 );
not ( n7666 , n78 );
and ( n7667 , n7665 , n7666 );
not ( n7668 , n7663 );
and ( n7669 , n7668 , n78 );
nor ( n7670 , n7667 , n7669 );
nand ( n7671 , n7362 , n7265 );
buf ( n7672 , n7258 );
nand ( n7673 , n7435 , n5 );
and ( n7674 , n7672 , n7673 );
or ( n7675 , n7671 , n7674 );
not ( n7676 , n5 );
nand ( n7677 , n7676 , n2 );
not ( n7678 , n7677 );
nand ( n7679 , n7678 , n7337 );
not ( n7680 , n7679 );
and ( n7681 , n7680 , n7 );
nor ( n7682 , n5 , n6 );
nand ( n7683 , n7319 , n7458 , n7682 );
not ( n7684 , n7683 );
nor ( n7685 , n7681 , n7684 , n7315 );
not ( n7686 , n7248 );
nand ( n7687 , n7686 , n7336 );
nand ( n7688 , n7675 , n7685 , n7687 );
not ( n7689 , n7688 );
not ( n7690 , n7373 );
or ( n7691 , n7690 , n7395 );
nand ( n7692 , n7691 , n6 );
not ( n7693 , n7692 );
nand ( n7694 , n7394 , n2 );
not ( n7695 , n7694 );
buf ( n7696 , n7695 );
nand ( n7697 , n4 , n7 );
not ( n7698 , n7697 );
and ( n7699 , n7696 , n7698 );
nand ( n7700 , n7309 , n7357 );
nor ( n7701 , n7700 , n7 );
not ( n7702 , n7395 );
nor ( n7703 , n7431 , n7702 );
or ( n7704 , n7703 , n8 );
nor ( n7705 , n7699 , n7701 , n7704 );
not ( n7706 , n7705 );
or ( n7707 , n7693 , n7706 );
not ( n7708 , n7375 );
not ( n7709 , n7236 );
buf ( n7710 , n7709 );
not ( n7711 , n7710 );
not ( n7712 , n7711 );
or ( n7713 , n7708 , n7712 );
not ( n7714 , n6 );
nand ( n7715 , n7237 , n7714 );
and ( n7716 , n7715 , n7295 , n7 );
nand ( n7717 , n7713 , n7716 );
nand ( n7718 , n7710 , n7357 );
nand ( n7719 , n7717 , n7718 , n8 );
nand ( n7720 , n7680 , n7714 );
not ( n7721 , n3 );
nor ( n7722 , n7721 , n4 );
not ( n7723 , n7722 );
nand ( n7724 , n7723 , n7695 );
and ( n7725 , n7720 , n7724 );
nor ( n7726 , n7725 , n7 );
or ( n7727 , n7719 , n7726 );
nand ( n7728 , n7362 , n7262 , n7316 );
not ( n7729 , n7728 );
nand ( n7730 , n7709 , n7240 );
not ( n7731 , n7730 );
nand ( n7732 , n7731 , n6 );
nor ( n7733 , n7 , n8 );
nand ( n7734 , n7732 , n7733 );
not ( n7735 , n7734 );
or ( n7736 , n7729 , n7735 );
nand ( n7737 , n7336 , n7722 );
nand ( n7738 , n7736 , n7737 );
nand ( n7739 , n7727 , n7738 );
not ( n7740 , n7265 );
not ( n7741 , n7400 );
or ( n7742 , n7740 , n7741 );
nor ( n7743 , n7325 , n3 );
nand ( n7744 , n7743 , n7251 );
nand ( n7745 , n7742 , n7744 );
and ( n7746 , n7362 , n3 );
not ( n7747 , n7286 );
not ( n7748 , n7700 );
or ( n7749 , n7747 , n7748 );
nand ( n7750 , n7749 , n7 );
nor ( n7751 , n7746 , n7750 );
nor ( n7752 , n7745 , n7751 , n9 );
nand ( n7753 , n7739 , n7752 );
nand ( n7754 , n7707 , n7753 );
not ( n7755 , n7754 );
not ( n7756 , n7755 );
or ( n7757 , n7689 , n7756 );
not ( n7758 , n6 );
and ( n7759 , n7231 , n7361 );
nand ( n7760 , n7758 , n7759 );
not ( n7761 , n3 );
nor ( n7762 , n7761 , n4 );
nand ( n7763 , n7710 , n7762 );
nand ( n7764 , n7760 , n7763 , n7265 );
nand ( n7765 , n7310 , n7328 );
not ( n7766 , n7765 );
or ( n7767 , n7764 , n7766 );
nand ( n7768 , n7418 , n7 );
not ( n7769 , n7768 );
not ( n7770 , n7275 );
not ( n7771 , n2 );
and ( n7772 , n7770 , n7771 );
and ( n7773 , n7762 , n7251 );
nor ( n7774 , n7772 , n7773 );
nand ( n7775 , n7769 , n7774 );
nand ( n7776 , n7767 , n7775 );
not ( n7777 , n6 );
nand ( n7778 , n7777 , n7678 );
not ( n7779 , n7778 );
and ( n7780 , n7779 , n7457 );
nor ( n7781 , n7780 , n7381 );
nand ( n7782 , n7776 , n7781 );
not ( n7783 , n7782 );
not ( n7784 , n7753 );
or ( n7785 , n7783 , n7784 );
nor ( n7786 , n7431 , n2 , n6 );
and ( n7787 , n7786 , n7349 );
and ( n7788 , n7305 , n7457 );
nor ( n7789 , n7787 , n7788 );
nand ( n7790 , n7785 , n7789 );
not ( n7791 , n7444 );
not ( n7792 , n7791 );
nand ( n7793 , n7792 , n7240 );
buf ( n7794 , n7232 );
nand ( n7795 , n7779 , n7794 );
nand ( n7796 , n7793 , n7 , n7795 );
nand ( n7797 , n7249 , n7251 );
nand ( n7798 , n7296 , n7682 );
nand ( n7799 , n7426 , n7797 , n7798 , n7315 );
or ( n7800 , n7796 , n7799 );
buf ( n7801 , n7389 );
nand ( n7802 , n7328 , n3 );
not ( n7803 , n4 );
nand ( n7804 , n7803 , n7416 );
not ( n7805 , n7804 );
not ( n7806 , n7805 );
and ( n7807 , n7801 , n7802 , n7806 );
nand ( n7808 , n7807 , n7285 );
not ( n7809 , n7248 );
nand ( n7810 , n7809 , n7328 );
buf ( n7811 , n7733 );
nand ( n7812 , n7808 , n7810 , n7811 );
nand ( n7813 , n7800 , n7812 );
buf ( n7814 , n7358 );
and ( n7815 , n7814 , n7744 );
and ( n7816 , n7813 , n7815 );
nand ( n7817 , n7773 , n7230 );
not ( n7818 , n7730 );
nand ( n7819 , n7818 , n7698 );
and ( n7820 , n7817 , n7819 , n7297 );
not ( n7821 , n7310 );
nor ( n7822 , n7821 , n7336 );
not ( n7823 , n7822 );
nor ( n7824 , n7320 , n3 );
buf ( n7825 , n7415 );
nand ( n7826 , n7824 , n7825 );
nand ( n7827 , n7823 , n7760 , n7826 , n8 );
nand ( n7828 , n7 , n8 );
nand ( n7829 , n7827 , n7828 );
nand ( n7830 , n7444 , n7457 );
and ( n7831 , n7820 , n7829 , n7830 );
nor ( n7832 , n7816 , n7831 );
nor ( n7833 , n7790 , n7832 );
nand ( n7834 , n7757 , n7833 );
not ( n7835 , n7834 );
not ( n7836 , n7835 );
nand ( n7837 , n6820 , n6719 );
nand ( n7838 , n7837 , n6882 );
not ( n7839 , n6740 );
not ( n7840 , n7839 );
not ( n7841 , n6719 );
or ( n7842 , n7840 , n7841 );
not ( n7843 , n6851 );
nor ( n7844 , n7843 , n6761 );
not ( n7845 , n7844 );
nand ( n7846 , n7842 , n7845 );
or ( n7847 , n7838 , n7846 );
not ( n7848 , n6702 );
nand ( n7849 , n7848 , n6706 );
not ( n7850 , n6764 );
nor ( n7851 , n7849 , n7850 );
or ( n7852 , n7851 , n6899 );
nand ( n7853 , n7847 , n7852 );
nor ( n7854 , n6815 , n6827 );
nor ( n7855 , n7854 , n6770 , n6807 );
nand ( n7856 , n7853 , n7855 );
not ( n7857 , n7856 );
not ( n7858 , n6724 );
nor ( n7859 , n7858 , n6782 );
not ( n7860 , n7859 );
nor ( n7861 , n27 , n28 , n30 , n31 );
and ( n7862 , n7861 , n29 );
and ( n7863 , n6920 , n30 );
not ( n7864 , n6923 );
nor ( n7865 , n6769 , n7864 );
nor ( n7866 , n6909 , n7862 , n7863 , n7865 );
not ( n7867 , n7866 );
or ( n7868 , n7860 , n7867 );
not ( n7869 , n31 );
nor ( n7870 , n7869 , n27 );
nand ( n7871 , n6823 , n7870 );
nand ( n7872 , n6894 , n6719 );
nand ( n7873 , n7871 , n7872 , n6867 , n6782 );
nand ( n7874 , n7868 , n7873 );
nand ( n7875 , n6838 , n6807 );
not ( n7876 , n30 );
nor ( n7877 , n7876 , n27 , n31 );
not ( n7878 , n7877 );
nor ( n7879 , n7878 , n28 , n29 );
nor ( n7880 , n7875 , n7879 );
nand ( n7881 , n7874 , n7880 );
not ( n7882 , n7881 );
or ( n7883 , n7857 , n7882 );
not ( n7884 , n6854 );
nand ( n7885 , n7884 , n6907 );
not ( n7886 , n7885 );
nand ( n7887 , n7886 , n6704 );
not ( n7888 , n7887 );
and ( n7889 , n7888 , n6782 );
nand ( n7890 , n6739 , n27 );
not ( n7891 , n7890 );
and ( n7892 , n7891 , n6828 );
nor ( n7893 , n7889 , n7892 );
nand ( n7894 , n7883 , n7893 );
not ( n7895 , n7894 );
not ( n7896 , n6866 );
not ( n7897 , n6844 );
or ( n7898 , n7896 , n7897 );
nand ( n7899 , n6722 , n32 );
not ( n7900 , n7899 );
nand ( n7901 , n7898 , n7900 );
not ( n7902 , n7901 );
and ( n7903 , n7848 , n6706 );
nand ( n7904 , n7903 , n6704 );
nand ( n7905 , n6744 , n29 );
not ( n7906 , n7905 );
not ( n7907 , n6907 );
and ( n7908 , n7906 , n7907 );
nor ( n7909 , n7908 , n32 );
nand ( n7910 , n7904 , n7909 );
not ( n7911 , n7910 );
or ( n7912 , n7902 , n7911 );
not ( n7913 , n6855 );
nor ( n7914 , n7913 , n6836 );
buf ( n7915 , n7914 );
not ( n7916 , n7915 );
nand ( n7917 , n7912 , n7916 );
not ( n7918 , n7917 );
not ( n7919 , n33 );
or ( n7920 , n7918 , n7919 );
nand ( n7921 , n6727 , n6706 );
not ( n7922 , n7921 );
nand ( n7923 , n6761 , n6837 );
not ( n7924 , n7923 );
or ( n7925 , n7922 , n7924 );
nand ( n7926 , n7925 , n32 );
not ( n7927 , n7926 );
nor ( n7928 , n6886 , n6719 );
not ( n7929 , n7928 );
and ( n7930 , n7927 , n7929 );
nor ( n7931 , n7879 , n34 );
nand ( n7932 , n6894 , n27 );
not ( n7933 , n7932 );
nand ( n7934 , n7933 , n6794 );
nand ( n7935 , n7931 , n7934 );
nor ( n7936 , n7930 , n7935 );
nand ( n7937 , n7920 , n7936 );
nand ( n7938 , n6761 , n7870 );
nand ( n7939 , n6887 , n7938 );
not ( n7940 , n7939 );
nand ( n7941 , n27 , n32 );
nand ( n7942 , n6855 , n6794 );
and ( n7943 , n7941 , n7942 );
buf ( n7944 , n6738 );
nor ( n7945 , n7943 , n7944 );
not ( n7946 , n7945 );
and ( n7947 , n7940 , n7946 );
nor ( n7948 , n7947 , n33 );
or ( n7949 , n7937 , n7948 );
nand ( n7950 , n6761 , n6704 );
not ( n7951 , n7950 );
not ( n7952 , n29 );
nand ( n7953 , n6735 , n7952 );
nand ( n7954 , n7953 , n6924 );
not ( n7955 , n7954 );
or ( n7956 , n7951 , n7955 );
nand ( n7957 , n7956 , n33 );
nand ( n7958 , n7957 , n6868 );
not ( n7959 , n7958 );
not ( n7960 , n6716 );
nand ( n7961 , n7960 , n31 );
not ( n7962 , n7961 );
nor ( n7963 , n7849 , n6882 );
nor ( n7964 , n6833 , n31 );
nor ( n7965 , n7962 , n7963 , n7964 );
not ( n7966 , n7965 );
or ( n7967 , n7959 , n7966 );
not ( n7968 , n6772 );
not ( n7969 , n7923 );
or ( n7970 , n7968 , n7969 );
not ( n7971 , n6773 );
nand ( n7972 , n7970 , n7971 );
and ( n7973 , n6883 , n30 );
nand ( n7974 , n7870 , n6938 );
nand ( n7975 , n7974 , n6873 );
nor ( n7976 , n7973 , n7975 );
nand ( n7977 , n7906 , n6880 );
nand ( n7978 , n7972 , n7976 , n7977 );
nand ( n7979 , n7967 , n7978 );
nand ( n7980 , n7979 , n34 );
nand ( n7981 , n7949 , n7980 );
or ( n7982 , n7937 , n7948 );
not ( n7983 , n7838 );
and ( n7984 , n6851 , n6938 );
not ( n7985 , n7984 );
and ( n7986 , n7885 , n7985 );
and ( n7987 , n7983 , n7986 );
nand ( n7988 , n6740 , n32 );
not ( n7989 , n6778 );
not ( n7990 , n7870 );
or ( n7991 , n7989 , n7990 );
nor ( n7992 , n6865 , n29 );
not ( n7993 , n7992 );
nand ( n7994 , n7991 , n7993 );
not ( n7995 , n6702 );
nand ( n7996 , n7995 , n6764 );
not ( n7997 , n7996 );
nor ( n7998 , n7988 , n7994 , n7997 );
nor ( n7999 , n7987 , n7998 );
nand ( n8000 , n7982 , n7999 );
nand ( n8001 , n7895 , n7981 , n8000 );
not ( n8002 , n8001 );
not ( n8003 , n8002 );
or ( n8004 , n7836 , n8003 );
nand ( n8005 , n8001 , n7834 );
nand ( n8006 , n8004 , n8005 );
xor ( n8007 , n7670 , n8006 );
not ( n8008 , n24 );
nor ( n8009 , n8008 , n23 );
not ( n8010 , n8009 );
not ( n8011 , n6285 );
not ( n8012 , n8011 );
or ( n8013 , n8010 , n8012 );
nand ( n8014 , n8013 , n6491 );
nand ( n8015 , n8014 , n25 );
not ( n8016 , n8015 );
not ( n8017 , n6307 );
nand ( n8018 , n8017 , n6343 );
nand ( n8019 , n8018 , n26 );
and ( n8020 , n6586 , n23 );
nor ( n8021 , n8016 , n8019 , n8020 );
not ( n8022 , n6526 );
nand ( n8023 , n6458 , n24 );
not ( n8024 , n8023 );
or ( n8025 , n8022 , n8024 );
nand ( n8026 , n8025 , n6327 );
and ( n8027 , n8021 , n8026 );
not ( n8028 , n6338 );
not ( n8029 , n6535 );
nand ( n8030 , n8029 , n6384 , n21 );
not ( n8031 , n6375 );
nand ( n8032 , n8031 , n6342 );
nand ( n8033 , n8030 , n8032 , n6656 , n6447 );
nor ( n8034 , n8028 , n6369 , n8033 );
nor ( n8035 , n8027 , n8034 );
and ( n8036 , n6291 , n25 );
and ( n8037 , n6442 , n20 );
and ( n8038 , n6534 , n22 );
nor ( n8039 , n8037 , n8038 );
and ( n8040 , n8039 , n6399 );
nor ( n8041 , n8040 , n6522 );
nor ( n8042 , n8036 , n8041 );
not ( n8043 , n8042 );
not ( n8044 , n6326 );
nand ( n8045 , n8044 , n23 );
not ( n8046 , n8045 );
nand ( n8047 , n8046 , n6348 , n6287 , n6299 );
not ( n8048 , n8047 );
or ( n8049 , n8043 , n8048 );
nand ( n8050 , n8049 , n26 );
not ( n8051 , n8050 );
nand ( n8052 , n6608 , n6287 );
not ( n8053 , n6491 );
nand ( n8054 , n8053 , n6315 );
and ( n8055 , n8052 , n8054 , n6539 );
or ( n8056 , n6433 , n25 );
nand ( n8057 , n8056 , n6308 );
nand ( n8058 , n8055 , n8057 );
nor ( n8059 , n8035 , n8051 , n8058 );
not ( n8060 , n6528 );
nand ( n8061 , n8060 , n23 );
not ( n8062 , n8061 );
not ( n8063 , n6287 );
and ( n8064 , n8062 , n8063 );
nand ( n8065 , n6325 , n24 );
nor ( n8066 , n8065 , n6466 );
nor ( n8067 , n8064 , n8066 );
nand ( n8068 , n8067 , n6656 );
not ( n8069 , n8068 );
nor ( n8070 , n6382 , n25 );
and ( n8071 , n8069 , n8070 );
nand ( n8072 , n6367 , n6343 );
nand ( n8073 , n6513 , n22 );
and ( n8074 , n8072 , n25 , n8065 , n8073 );
nor ( n8075 , n8071 , n8074 );
nand ( n8076 , n6529 , n6525 );
and ( n8077 , n8076 , n26 );
not ( n8078 , n6669 );
nand ( n8079 , n6292 , n6650 , n8077 , n8078 );
or ( n8080 , n8075 , n8079 );
not ( n8081 , n6299 );
not ( n8082 , n8068 );
or ( n8083 , n8081 , n8082 );
nand ( n8084 , n6373 , n6356 );
not ( n8085 , n8084 );
not ( n8086 , n6404 );
not ( n8087 , n8086 );
and ( n8088 , n8085 , n8087 );
nand ( n8089 , n6579 , n25 );
nor ( n8090 , n6519 , n8089 );
nor ( n8091 , n8088 , n8090 );
not ( n8092 , n6378 );
nand ( n8093 , n6478 , n6513 );
nand ( n8094 , n6321 , n8092 , n8093 );
nor ( n8095 , n8091 , n8094 , n6395 );
nand ( n8096 , n8083 , n8095 );
and ( n8097 , n8080 , n8096 );
nand ( n8098 , n6284 , n6354 );
nand ( n8099 , n8098 , n19 );
nand ( n8100 , n6287 , n6284 );
and ( n8101 , n8045 , n6393 , n8100 );
nor ( n8102 , n8101 , n6375 );
nor ( n8103 , n8099 , n8102 );
nand ( n8104 , n8050 , n8103 );
nor ( n8105 , n8097 , n8104 );
or ( n8106 , n8059 , n8105 );
not ( n8107 , n6337 );
not ( n8108 , n8107 );
nand ( n8109 , n8108 , n6649 );
nand ( n8110 , n8052 , n8109 , n6320 , n6454 );
nand ( n8111 , n6354 , n20 );
and ( n8112 , n8111 , n8077 );
not ( n8113 , n6594 );
nand ( n8114 , n8113 , n6679 , n6447 );
and ( n8115 , n8114 , n6299 );
nor ( n8116 , n8112 , n8115 );
and ( n8117 , n8110 , n8116 );
not ( n8118 , n6693 );
nand ( n8119 , n6394 , n22 );
not ( n8120 , n8119 );
or ( n8121 , n8118 , n8120 );
nand ( n8122 , n8121 , n6315 );
nand ( n8123 , n6431 , n6462 );
nand ( n8124 , n8122 , n8123 );
nor ( n8125 , n8117 , n8124 );
nand ( n8126 , n8106 , n8125 );
not ( n8127 , n8126 );
and ( n8128 , n8127 , n6698 );
not ( n8129 , n8127 );
not ( n8130 , n6698 );
and ( n8131 , n8129 , n8130 );
nor ( n8132 , n8128 , n8131 );
not ( n8133 , n8132 );
not ( n8134 , n6869 );
nand ( n8135 , n6844 , n27 );
and ( n8136 , n6946 , n7905 , n8135 );
not ( n8137 , n8136 );
or ( n8138 , n8134 , n8137 );
not ( n8139 , n32 );
nand ( n8140 , n8139 , n33 );
not ( n8141 , n8140 );
nand ( n8142 , n7950 , n8141 );
nand ( n8143 , n8138 , n8142 );
and ( n8144 , n27 , n30 );
nand ( n8145 , n6703 , n8144 );
not ( n8146 , n8145 );
not ( n8147 , n8146 );
not ( n8148 , n6803 );
and ( n8149 , n7985 , n8147 , n8148 , n7942 );
nand ( n8150 , n8143 , n8149 );
not ( n8151 , n8150 );
nand ( n8152 , n7996 , n6787 );
nor ( n8153 , n8152 , n7899 );
not ( n8154 , n7872 );
nor ( n8155 , n6858 , n8154 );
or ( n8156 , n8153 , n8155 );
not ( n8157 , n7865 );
or ( n8158 , n27 , n31 );
nor ( n8159 , n8158 , n7944 );
nor ( n8160 , n8159 , n33 );
and ( n8161 , n6760 , n6937 );
not ( n8162 , n8161 );
and ( n8163 , n8157 , n8160 , n8162 );
nand ( n8164 , n8156 , n8163 );
not ( n8165 , n8164 );
or ( n8166 , n8151 , n8165 );
not ( n8167 , n6854 );
nand ( n8168 , n8167 , n6704 );
or ( n8169 , n8168 , n6706 );
not ( n8170 , n8169 );
nand ( n8171 , n6848 , n6705 );
or ( n8172 , n8170 , n8171 );
nand ( n8173 , n8172 , n6880 );
not ( n8174 , n6855 );
not ( n8175 , n6908 );
not ( n8176 , n8175 );
or ( n8177 , n8174 , n8176 );
nand ( n8178 , n8177 , n34 );
not ( n8179 , n8178 );
and ( n8180 , n8173 , n8179 );
nand ( n8181 , n8166 , n8180 );
not ( n8182 , n8145 );
nand ( n8183 , n8182 , n6719 );
nand ( n8184 , n6823 , n6837 );
and ( n8185 , n8183 , n8184 , n7871 );
not ( n8186 , n8185 );
buf ( n8187 , n6937 );
nand ( n8188 , n8187 , n6844 );
not ( n8189 , n8188 );
or ( n8190 , n8186 , n8189 );
nand ( n8191 , n8190 , n6882 );
not ( n8192 , n8191 );
or ( n8193 , n8181 , n8192 );
not ( n8194 , n27 );
nand ( n8195 , n8194 , n6736 );
not ( n8196 , n8195 );
nor ( n8197 , n8196 , n6868 );
not ( n8198 , n8197 );
buf ( n8199 , n6786 );
nand ( n8200 , n6757 , n8199 );
not ( n8201 , n8200 );
or ( n8202 , n8198 , n8201 );
not ( n8203 , n6745 );
nand ( n8204 , n6710 , n8203 );
nand ( n8205 , n8204 , n8141 );
nand ( n8206 , n8202 , n8205 );
not ( n8207 , n8206 );
nand ( n8208 , n7839 , n6719 );
and ( n8209 , n8208 , n8184 , n7996 );
not ( n8210 , n8209 );
or ( n8211 , n8207 , n8210 );
nand ( n8212 , n6761 , n6880 );
and ( n8213 , n8188 , n8212 , n6807 );
not ( n8214 , n6833 );
and ( n8215 , n7864 , n6912 , n29 );
nor ( n8216 , n8214 , n8215 );
not ( n8217 , n6750 );
nand ( n8218 , n8146 , n8217 );
nand ( n8219 , n8213 , n8216 , n8218 );
nand ( n8220 , n8211 , n8219 );
nand ( n8221 , n6757 , n6802 );
not ( n8222 , n8221 );
or ( n8223 , n8222 , n7915 , n32 );
not ( n8224 , n6775 );
not ( n8225 , n6764 );
or ( n8226 , n8224 , n8225 );
not ( n8227 , n7988 );
nand ( n8228 , n8226 , n8227 );
nand ( n8229 , n8223 , n8228 );
nor ( n8230 , n8168 , n31 );
nand ( n8231 , n8230 , n6706 );
not ( n8232 , n8231 );
nor ( n8233 , n8232 , n34 );
nand ( n8234 , n8220 , n8229 , n8233 );
nand ( n8235 , n8193 , n8234 );
nand ( n8236 , n8231 , n6773 );
or ( n8237 , n8236 , n7964 );
not ( n8238 , n28 );
not ( n8239 , n8175 );
or ( n8240 , n8238 , n8239 );
nor ( n8241 , n7984 , n6807 );
nand ( n8242 , n8240 , n8241 );
nand ( n8243 , n8237 , n8242 );
not ( n8244 , n8243 );
nand ( n8245 , n6879 , n6926 );
not ( n8246 , n8245 );
or ( n8247 , n8244 , n8246 );
and ( n8248 , n7974 , n6782 );
nor ( n8249 , n8248 , n8141 );
nand ( n8250 , n8247 , n8249 );
not ( n8251 , n7904 );
nand ( n8252 , n8251 , n8217 );
not ( n8253 , n8204 );
or ( n8254 , n8253 , n7954 );
not ( n8255 , n6794 );
not ( n8256 , n8255 );
nand ( n8257 , n8254 , n8256 );
nand ( n8258 , n8252 , n8257 , n7977 );
and ( n8259 , n8258 , n33 );
and ( n8260 , n7914 , n6704 );
nor ( n8261 , n8259 , n8260 );
and ( n8262 , n8250 , n8261 );
nand ( n8263 , n8235 , n8262 );
buf ( n8264 , n8263 );
not ( n8265 , n8264 );
nand ( n8266 , n6811 , n6956 );
not ( n8267 , n8266 );
not ( n8268 , n8267 );
not ( n8269 , n8268 );
or ( n8270 , n8265 , n8269 );
not ( n8271 , n8264 );
not ( n8272 , n6957 );
nand ( n8273 , n8271 , n8272 );
nand ( n8274 , n8270 , n8273 );
not ( n8275 , n8274 );
or ( n8276 , n8133 , n8275 );
or ( n8277 , n8132 , n8274 );
nand ( n8278 , n8276 , n8277 );
and ( n8279 , n8007 , n8278 );
not ( n8280 , n8007 );
not ( n8281 , n8278 );
and ( n8282 , n8280 , n8281 );
nor ( n8283 , n8279 , n8282 );
or ( n8284 , n8283 , n1 );
xnor ( n8285 , n78 , n92 );
or ( n8286 , n2246 , n8285 );
nand ( n8287 , n8284 , n8286 );
not ( n8288 , n8267 );
buf ( n8289 , n6707 );
and ( n8290 , n8289 , n8256 );
not ( n8291 , n30 );
not ( n8292 , n7995 );
not ( n8293 , n8292 );
or ( n8294 , n8291 , n8293 );
nand ( n8295 , n8294 , n7870 );
not ( n8296 , n6952 );
and ( n8297 , n8296 , n8187 );
nor ( n8298 , n8297 , n33 );
nand ( n8299 , n8295 , n8298 );
nor ( n8300 , n8290 , n8299 );
not ( n8301 , n8300 );
not ( n8302 , n6921 );
nand ( n8303 , n8302 , n6704 );
nand ( n8304 , n8303 , n7932 );
not ( n8305 , n6944 );
or ( n8306 , n8304 , n8305 );
nand ( n8307 , n8306 , n32 );
not ( n8308 , n8307 );
or ( n8309 , n8301 , n8308 );
nand ( n8310 , n33 , n7944 );
or ( n8311 , n6886 , n8310 );
nand ( n8312 , n8311 , n6868 );
nand ( n8313 , n8312 , n8169 );
nand ( n8314 , n8309 , n8313 );
nand ( n8315 , n6943 , n6719 );
not ( n8316 , n7851 );
or ( n8317 , n6727 , n6775 );
nand ( n8318 , n8317 , n8217 );
and ( n8319 , n8315 , n8316 , n8318 );
nand ( n8320 , n8314 , n8319 );
nand ( n8321 , n6779 , n8199 );
and ( n8322 , n7904 , n6875 , n8321 , n6941 );
not ( n8323 , n8183 );
not ( n8324 , n8323 );
and ( n8325 , n8322 , n8324 );
not ( n8326 , n32 );
nand ( n8327 , n8326 , n34 );
nor ( n8328 , n6825 , n6953 , n8327 );
nor ( n8329 , n8325 , n8328 );
or ( n8330 , n8320 , n8329 );
not ( n8331 , n32 );
not ( n8332 , n7858 );
or ( n8333 , n8331 , n8332 );
not ( n8334 , n6934 );
nand ( n8335 , n8333 , n8334 );
not ( n8336 , n6882 );
not ( n8337 , n8154 );
or ( n8338 , n8336 , n8337 );
not ( n8339 , n6769 );
not ( n8340 , n6761 );
not ( n8341 , n8340 );
or ( n8342 , n8339 , n8341 );
nand ( n8343 , n8342 , n6861 );
nand ( n8344 , n8338 , n8343 );
nor ( n8345 , n8335 , n8344 );
not ( n8346 , n7905 );
nand ( n8347 , n6823 , n6719 );
not ( n8348 , n8347 );
or ( n8349 , n8346 , n8348 );
nand ( n8350 , n8349 , n32 );
nand ( n8351 , n6741 , n6719 );
and ( n8352 , n8350 , n7972 , n8351 );
or ( n8353 , n8345 , n8352 );
not ( n8354 , n6940 );
not ( n8355 , n7961 );
or ( n8356 , n8354 , n8355 );
nand ( n8357 , n8356 , n32 );
and ( n8358 , n8357 , n6812 );
nand ( n8359 , n8353 , n8358 );
not ( n8360 , n7861 );
not ( n8361 , n8360 );
not ( n8362 , n8185 );
or ( n8363 , n8361 , n8362 );
nand ( n8364 , n8363 , n6782 );
not ( n8365 , n8364 );
or ( n8366 , n8359 , n8365 );
nand ( n8367 , n8330 , n8366 );
and ( n8368 , n6764 , n6778 );
nor ( n8369 , n8368 , n6782 );
nand ( n8370 , n8369 , n6779 , n7952 );
not ( n8371 , n8370 );
not ( n8372 , n6776 );
nand ( n8373 , n8372 , n8217 );
not ( n8374 , n8373 );
nor ( n8375 , n8371 , n8374 );
not ( n8376 , n8375 );
buf ( n8377 , n8230 );
not ( n8378 , n8377 );
not ( n8379 , n7879 );
nand ( n8380 , n8378 , n8379 );
nand ( n8381 , n6898 , n6782 );
or ( n8382 , n8380 , n8381 , n33 );
or ( n8383 , n7862 , n7971 , n8159 );
nand ( n8384 , n8382 , n8383 );
not ( n8385 , n8384 );
or ( n8386 , n8376 , n8385 );
nand ( n8387 , n8377 , n6880 );
or ( n8388 , n7997 , n6868 );
or ( n8389 , n6803 , n8140 );
nand ( n8390 , n8388 , n8389 );
nand ( n8391 , n8387 , n7961 , n7837 , n8390 );
nand ( n8392 , n8386 , n8391 );
not ( n8393 , n6912 );
or ( n8394 , n6787 , n8393 );
nor ( n8395 , n6769 , n32 );
not ( n8396 , n8395 );
nand ( n8397 , n8394 , n8396 );
nand ( n8398 , n8397 , n28 );
and ( n8399 , n8392 , n8398 );
nand ( n8400 , n8367 , n8399 );
not ( n8401 , n8400 );
not ( n8402 , n8401 );
or ( n8403 , n8288 , n8402 );
buf ( n8404 , n8266 );
nand ( n8405 , n8400 , n8404 );
nand ( n8406 , n8403 , n8405 );
not ( n8407 , n8406 );
not ( n8408 , n8130 );
not ( n8409 , n6340 );
and ( n8410 , n6427 , n6450 );
not ( n8411 , n8410 );
or ( n8412 , n8409 , n8411 );
not ( n8413 , n6640 );
nand ( n8414 , n8413 , n25 );
nand ( n8415 , n8412 , n8414 );
not ( n8416 , n20 );
not ( n8417 , n6365 );
not ( n8418 , n8417 );
or ( n8419 , n8416 , n8418 );
not ( n8420 , n26 );
nor ( n8421 , n8420 , n6489 );
nand ( n8422 , n8421 , n6521 );
nand ( n8423 , n8419 , n8422 );
nor ( n8424 , n8415 , n8423 );
buf ( n8425 , n6689 );
not ( n8426 , n8425 );
and ( n8427 , n8052 , n8098 , n6660 , n6299 );
not ( n8428 , n8427 );
or ( n8429 , n8426 , n8428 );
nand ( n8430 , n6483 , n25 );
not ( n8431 , n8430 );
and ( n8432 , n6655 , n6296 );
not ( n8433 , n8432 );
and ( n8434 , n8431 , n8433 , n6319 );
nor ( n8435 , n8434 , n26 );
nand ( n8436 , n8429 , n8435 );
not ( n8437 , n6355 );
or ( n8438 , n8437 , n6380 , n6395 );
nand ( n8439 , n8438 , n26 );
and ( n8440 , n8424 , n8436 , n8439 );
not ( n8441 , n26 );
not ( n8442 , n6305 );
not ( n8443 , n8107 );
or ( n8444 , n8442 , n8443 );
nand ( n8445 , n8444 , n6339 );
and ( n8446 , n6288 , n8445 );
not ( n8447 , n8446 );
or ( n8448 , n8441 , n8447 );
not ( n8449 , n6547 );
not ( n8450 , n6520 );
or ( n8451 , n8449 , n8450 );
nand ( n8452 , n8451 , n25 );
not ( n8453 , n6409 );
not ( n8454 , n6344 );
not ( n8455 , n8454 );
or ( n8456 , n8453 , n8455 );
not ( n8457 , n24 );
not ( n8458 , n6326 );
or ( n8459 , n8457 , n8458 );
nand ( n8460 , n8459 , n6510 );
nand ( n8461 , n6606 , n6625 );
and ( n8462 , n8460 , n8461 , n6320 );
nand ( n8463 , n8456 , n8462 );
nor ( n8464 , n8119 , n6522 );
nor ( n8465 , n8463 , n8464 );
nand ( n8466 , n8452 , n8465 );
nand ( n8467 , n8448 , n8466 );
not ( n8468 , n8467 );
nand ( n8469 , n6519 , n6343 );
not ( n8470 , n6510 );
nor ( n8471 , n8470 , n20 );
nand ( n8472 , n8471 , n6513 );
or ( n8473 , n6462 , n6443 );
nand ( n8474 , n8473 , n6679 );
and ( n8475 , n8469 , n8472 , n8474 , n19 );
nand ( n8476 , n6676 , n6535 );
nand ( n8477 , n6474 , n8476 );
buf ( n8478 , n8066 );
or ( n8479 , n8477 , n8430 , n8478 );
not ( n8480 , n6587 );
not ( n8481 , n6626 );
or ( n8482 , n8480 , n8481 , n25 );
nand ( n8483 , n8479 , n8482 );
nand ( n8484 , n8475 , n8483 );
or ( n8485 , n8468 , n8484 );
nand ( n8486 , n6502 , n6348 );
nand ( n8487 , n6342 , n6356 , n6330 );
not ( n8488 , n8487 );
nor ( n8489 , n8488 , n19 );
not ( n8490 , n6448 );
buf ( n8491 , n6578 );
or ( n8492 , n8491 , n23 );
nand ( n8493 , n8492 , n8065 );
nand ( n8494 , n8490 , n8493 );
nand ( n8495 , n6541 , n6521 );
nand ( n8496 , n8486 , n8489 , n8494 , n8495 );
and ( n8497 , n6343 , n6675 );
and ( n8498 , n6344 , n26 );
nor ( n8499 , n8497 , n8498 );
not ( n8500 , n8067 );
nand ( n8501 , n8500 , n6299 );
nand ( n8502 , n8499 , n8501 , n6621 );
or ( n8503 , n8496 , n8502 );
nand ( n8504 , n8485 , n8503 );
nand ( n8505 , n8440 , n8504 );
not ( n8506 , n8505 );
not ( n8507 , n8506 );
or ( n8508 , n8408 , n8507 );
nand ( n8509 , n6698 , n8505 );
nand ( n8510 , n8508 , n8509 );
not ( n8511 , n8510 );
or ( n8512 , n8407 , n8511 );
or ( n8513 , n8510 , n8406 );
nand ( n8514 , n8512 , n8513 );
not ( n8515 , n69 );
nand ( n8516 , n7658 , n6995 );
not ( n8517 , n7633 );
not ( n8518 , n8517 );
not ( n8519 , n6999 );
nor ( n8520 , n8519 , n7512 );
not ( n8521 , n8520 );
nand ( n8522 , n8518 , n8521 );
or ( n8523 , n8516 , n8522 );
not ( n8524 , n7023 );
or ( n8525 , n8524 , n7170 );
nand ( n8526 , n8523 , n8525 );
not ( n8527 , n7108 );
and ( n8528 , n8527 , n7576 );
nor ( n8529 , n8528 , n7222 );
and ( n8530 , n8526 , n8529 );
not ( n8531 , n8530 );
not ( n8532 , n7649 );
not ( n8533 , n7192 );
nand ( n8534 , n8532 , n8533 );
nand ( n8535 , n8534 , n11 );
not ( n8536 , n7605 );
nand ( n8537 , n8536 , n14 );
and ( n8538 , n8535 , n8537 );
nor ( n8539 , n8538 , n7170 );
nand ( n8540 , n7649 , n7189 );
nor ( n8541 , n8540 , n7026 );
not ( n8542 , n8541 );
nand ( n8543 , n8542 , n7124 );
or ( n8544 , n8539 , n8543 , n7131 );
not ( n8545 , n7088 );
not ( n8546 , n7510 );
nor ( n8547 , n8545 , n8546 );
or ( n8548 , n8547 , n6989 );
nand ( n8549 , n8548 , n7661 );
not ( n8550 , n7517 );
buf ( n8551 , n7513 );
nand ( n8552 , n8550 , n8551 );
nand ( n8553 , n8549 , n8552 , n7658 , n7131 );
nand ( n8554 , n8544 , n8553 );
not ( n8555 , n8554 );
or ( n8556 , n8531 , n8555 );
nand ( n8557 , n7111 , n7059 );
not ( n8558 , n8557 );
nor ( n8559 , n7621 , n13 );
not ( n8560 , n7531 );
not ( n8561 , n7649 );
not ( n8562 , n7107 );
or ( n8563 , n8561 , n8562 );
nand ( n8564 , n8563 , n7530 );
not ( n8565 , n8564 );
or ( n8566 , n8560 , n8565 );
nand ( n8567 , n7003 , n6978 );
or ( n8568 , n7109 , n8567 );
not ( n8569 , n7132 );
nand ( n8570 , n8568 , n8569 );
nand ( n8571 , n8566 , n8570 );
nor ( n8572 , n8558 , n8559 , n8571 );
not ( n8573 , n7190 );
not ( n8574 , n7543 );
or ( n8575 , n8573 , n8574 );
nand ( n8576 , n8575 , n16 );
nand ( n8577 , n7096 , n7614 , n8534 );
nor ( n8578 , n7575 , n7142 );
nand ( n8579 , n8578 , n7605 );
nand ( n8580 , n8577 , n8579 );
nor ( n8581 , n7615 , n13 );
nor ( n8582 , n8580 , n8581 );
nand ( n8583 , n8576 , n8582 );
nand ( n8584 , n7045 , n13 );
nand ( n8585 , n8584 , n17 );
nor ( n8586 , n8583 , n8585 );
or ( n8587 , n8572 , n8586 );
nor ( n8588 , n7649 , n7168 );
nand ( n8589 , n8588 , n7628 );
nand ( n8590 , n8589 , n7531 , n7008 );
nor ( n8591 , n7615 , n6990 );
or ( n8592 , n8591 , n7015 );
nand ( n8593 , n8592 , n7142 );
nor ( n8594 , n8521 , n7008 );
nor ( n8595 , n8594 , n10 );
and ( n8596 , n8590 , n8593 , n8595 );
nand ( n8597 , n8587 , n8596 );
nand ( n8598 , n8556 , n8597 );
not ( n8599 , n17 );
not ( n8600 , n7206 );
nand ( n8601 , n8600 , n7142 );
not ( n8602 , n8601 );
or ( n8603 , n8599 , n8602 );
nand ( n8604 , n6989 , n7044 );
not ( n8605 , n7636 );
nand ( n8606 , n8605 , n6984 );
nand ( n8607 , n8604 , n8606 );
or ( n8608 , n8607 , n7015 );
nand ( n8609 , n8608 , n7142 );
nor ( n8610 , n7089 , n17 );
nand ( n8611 , n8609 , n8610 );
nand ( n8612 , n8603 , n8611 );
not ( n8613 , n8610 );
or ( n8614 , n7026 , n7636 );
nand ( n8615 , n8614 , n7124 );
and ( n8616 , n8613 , n8615 , n13 );
nor ( n8617 , n8616 , n7170 );
not ( n8618 , n8584 );
nand ( n8619 , n8618 , n7026 );
nand ( n8620 , n8612 , n8617 , n8619 );
nand ( n8621 , n7093 , n7565 , n7060 , n7144 );
not ( n8622 , n7215 );
not ( n8623 , n7175 );
or ( n8624 , n8622 , n8623 );
nand ( n8625 , n8624 , n7164 );
or ( n8626 , n8585 , n8625 , n7171 );
nand ( n8627 , n8620 , n8621 , n8626 );
nand ( n8628 , n8626 , n7506 );
nand ( n8629 , n8598 , n8627 , n8628 );
not ( n8630 , n8629 );
not ( n8631 , n8630 );
or ( n8632 , n8515 , n8631 );
buf ( n8633 , n8629 );
not ( n8634 , n69 );
nand ( n8635 , n8633 , n8634 );
nand ( n8636 , n8632 , n8635 );
not ( n8637 , n6775 );
not ( n8638 , n8637 );
not ( n8639 , n7950 );
or ( n8640 , n8638 , n8639 );
nand ( n8641 , n8640 , n6912 );
nand ( n8642 , n8641 , n8162 , n6812 );
nor ( n8643 , n8371 , n8642 );
not ( n8644 , n8643 );
not ( n8645 , n7871 );
nand ( n8646 , n7995 , n6719 );
and ( n8647 , n6727 , n6860 );
nor ( n8648 , n8647 , n32 );
or ( n8649 , n27 , n28 , n30 );
and ( n8650 , n8646 , n8648 , n7885 , n8649 );
not ( n8651 , n8650 );
or ( n8652 , n8645 , n8651 );
nand ( n8653 , n7885 , n32 );
not ( n8654 , n8653 );
nand ( n8655 , n6802 , n27 );
nand ( n8656 , n8654 , n8347 , n8655 );
nand ( n8657 , n8652 , n8656 );
nand ( n8658 , n6765 , n33 );
nor ( n8659 , n7858 , n8658 );
nand ( n8660 , n8657 , n8659 );
not ( n8661 , n6939 );
nand ( n8662 , n8661 , n6704 );
nand ( n8663 , n8169 , n8662 , n6882 );
or ( n8664 , n8663 , n8323 );
nand ( n8665 , n8315 , n32 );
nand ( n8666 , n8664 , n8665 );
nand ( n8667 , n7984 , n32 );
nand ( n8668 , n8667 , n6807 );
nor ( n8669 , n8260 , n8668 );
nand ( n8670 , n8666 , n8669 , n7871 );
nand ( n8671 , n8660 , n8670 );
not ( n8672 , n8671 );
or ( n8673 , n8644 , n8672 );
nand ( n8674 , n8184 , n6730 );
nand ( n8675 , n8674 , n33 );
not ( n8676 , n8675 );
and ( n8677 , n6849 , n6817 , n8315 , n6868 );
not ( n8678 , n8677 );
or ( n8679 , n8676 , n8678 );
and ( n8680 , n6727 , n27 );
nor ( n8681 , n8680 , n6782 );
not ( n8682 , n6798 );
nand ( n8683 , n6938 , n31 );
and ( n8684 , n8681 , n8682 , n8683 );
nor ( n8685 , n8684 , n6773 );
nand ( n8686 , n8679 , n8685 );
not ( n8687 , n8199 );
not ( n8688 , n6837 );
or ( n8689 , n8687 , n8688 );
nand ( n8690 , n8187 , n6802 );
not ( n8691 , n8690 );
nand ( n8692 , n6750 , n6836 );
or ( n8693 , n8691 , n8692 );
buf ( n8694 , n6846 );
nand ( n8695 , n8693 , n8694 );
nand ( n8696 , n8689 , n8695 );
and ( n8697 , n8696 , n6807 );
not ( n8698 , n6737 );
and ( n8699 , n8698 , n6868 );
not ( n8700 , n8203 );
not ( n8701 , n7992 );
or ( n8702 , n8700 , n8701 );
nand ( n8703 , n8702 , n34 );
nor ( n8704 , n8699 , n8703 );
not ( n8705 , n6882 );
not ( n8706 , n6757 );
not ( n8707 , n8706 );
or ( n8708 , n8705 , n8707 );
nand ( n8709 , n8708 , n8154 );
nand ( n8710 , n8704 , n8709 );
nor ( n8711 , n8697 , n8710 );
nand ( n8712 , n8686 , n8711 );
nand ( n8713 , n8673 , n8712 );
not ( n8714 , n6845 );
not ( n8715 , n8714 );
not ( n8716 , n7890 );
not ( n8717 , n6730 );
or ( n8718 , n8716 , n8717 );
nand ( n8719 , n8718 , n31 );
nand ( n8720 , n8719 , n6869 );
not ( n8721 , n8720 );
and ( n8722 , n8715 , n8721 );
not ( n8723 , n6704 );
not ( n8724 , n8646 );
not ( n8725 , n8724 );
or ( n8726 , n8723 , n8725 );
nor ( n8727 , n8161 , n33 );
nand ( n8728 , n8726 , n8727 );
nor ( n8729 , n8728 , n8222 );
nor ( n8730 , n8722 , n8729 );
nor ( n8731 , n6765 , n27 );
not ( n8732 , n8731 );
nand ( n8733 , n8732 , n8157 );
or ( n8734 , n8730 , n8733 );
not ( n8735 , n6947 );
nand ( n8736 , n8655 , n8195 , n33 );
not ( n8737 , n8736 );
not ( n8738 , n8737 );
or ( n8739 , n8735 , n8738 );
and ( n8740 , n6765 , n6776 , n6782 );
not ( n8741 , n8740 );
not ( n8742 , n6821 );
or ( n8743 , n8741 , n8742 );
or ( n8744 , n32 , n33 );
nand ( n8745 , n8743 , n8744 );
nand ( n8746 , n8739 , n8745 );
nand ( n8747 , n8734 , n8746 );
not ( n8748 , n7964 );
nand ( n8749 , n6903 , n6764 );
nand ( n8750 , n8748 , n6875 , n8749 );
not ( n8751 , n8744 );
and ( n8752 , n8750 , n8751 );
and ( n8753 , n8157 , n8321 );
nor ( n8754 , n8753 , n33 );
nor ( n8755 , n8752 , n8754 );
and ( n8756 , n8747 , n8755 );
nand ( n8757 , n8713 , n8756 );
not ( n8758 , n8757 );
not ( n8759 , n8758 );
nand ( n8760 , n7426 , n7763 );
not ( n8761 , n4 );
nor ( n8762 , n8761 , n7320 );
not ( n8763 , n8762 );
not ( n8764 , n8763 );
not ( n8765 , n7826 );
or ( n8766 , n8764 , n8765 );
nand ( n8767 , n8766 , n7 );
nand ( n8768 , n8767 , n7311 );
nor ( n8769 , n8760 , n8768 );
and ( n8770 , n7319 , n5 );
not ( n8771 , n8770 );
nand ( n8772 , n8771 , n7672 );
not ( n8773 , n7431 );
nor ( n8774 , n8773 , n6 );
not ( n8775 , n8774 );
or ( n8776 , n8772 , n8775 );
nand ( n8777 , n7678 , n7240 );
nand ( n8778 , n8776 , n8777 );
not ( n8779 , n7810 );
or ( n8780 , n8778 , n8779 );
nand ( n8781 , n8780 , n7265 );
and ( n8782 , n8769 , n8781 );
nor ( n8783 , n8782 , n7271 );
not ( n8784 , n7810 );
not ( n8785 , n7239 );
not ( n8786 , n7310 );
nor ( n8787 , n8785 , n8786 );
not ( n8788 , n8787 );
not ( n8789 , n8788 );
or ( n8790 , n8784 , n8789 );
nand ( n8791 , n8790 , n7271 );
nand ( n8792 , n7444 , n7457 , n4 );
and ( n8793 , n7766 , n7316 );
not ( n8794 , n7759 );
nand ( n8795 , n8794 , n7381 );
nor ( n8796 , n8793 , n8795 );
and ( n8797 , n8791 , n8792 , n8796 );
not ( n8798 , n7438 );
not ( n8799 , n7315 );
not ( n8800 , n7355 );
or ( n8801 , n8799 , n8800 );
nor ( n8802 , n7452 , n7435 );
nand ( n8803 , n8801 , n8802 );
not ( n8804 , n8803 );
or ( n8805 , n8798 , n8804 );
not ( n8806 , n7715 );
nand ( n8807 , n8806 , n4 );
not ( n8808 , n7473 );
nand ( n8809 , n8808 , n7285 );
nand ( n8810 , n8807 , n8809 );
nor ( n8811 , n7694 , n7275 );
buf ( n8812 , n8811 );
or ( n8813 , n8810 , n8812 );
nand ( n8814 , n8813 , n7811 );
nand ( n8815 , n8805 , n8814 );
not ( n8816 , n8815 );
nand ( n8817 , n8797 , n8816 );
or ( n8818 , n8783 , n8817 );
and ( n8819 , n7 , n9 );
not ( n8820 , n8819 );
nor ( n8821 , n7327 , n6 );
nand ( n8822 , n8821 , n7240 );
not ( n8823 , n8822 );
or ( n8824 , n8820 , n8823 );
not ( n8825 , n7732 );
nor ( n8826 , n8825 , n7381 );
nand ( n8827 , n7396 , n7265 );
nor ( n8828 , n8827 , n7786 );
nand ( n8829 , n8826 , n7445 , n8828 );
nand ( n8830 , n8824 , n8829 );
nand ( n8831 , n7296 , n7251 );
nand ( n8832 , n7814 , n8831 );
nand ( n8833 , n8808 , n7411 );
nor ( n8834 , n7385 , n7278 );
not ( n8835 , n8834 );
nand ( n8836 , n8833 , n7417 , n8835 );
or ( n8837 , n8832 , n8836 );
nand ( n8838 , n8837 , n7271 );
nand ( n8839 , n7296 , n7341 );
nand ( n8840 , n8839 , n7424 );
and ( n8841 , n8840 , n8 );
and ( n8842 , n7346 , n7401 , n7802 );
or ( n8843 , n8842 , n7828 );
not ( n8844 , n8821 );
not ( n8845 , n8844 );
not ( n8846 , n7791 );
or ( n8847 , n8845 , n8846 );
nand ( n8848 , n8847 , n7276 );
nand ( n8849 , n8843 , n8848 );
and ( n8850 , n7350 , n7678 );
nor ( n8851 , n8841 , n8849 , n8850 );
nand ( n8852 , n8830 , n8838 , n8851 );
nand ( n8853 , n8818 , n8852 );
nand ( n8854 , n7801 , n7369 );
or ( n8855 , n7684 , n8854 );
nand ( n8856 , n8855 , n7733 );
not ( n8857 , n7262 );
not ( n8858 , n7424 );
or ( n8859 , n8857 , n8858 );
nand ( n8860 , n8859 , n3 );
not ( n8861 , n8860 );
or ( n8862 , n7400 , n8861 );
not ( n8863 , n7828 );
nand ( n8864 , n8862 , n8863 );
not ( n8865 , n8835 );
not ( n8866 , n7798 );
or ( n8867 , n8865 , n8866 );
nand ( n8868 , n8867 , n7315 );
and ( n8869 , n8856 , n8864 , n8868 );
not ( n8870 , n7714 );
not ( n8871 , n8777 );
not ( n8872 , n8871 );
or ( n8873 , n8870 , n8872 );
nand ( n8874 , n8873 , n8794 );
nand ( n8875 , n7446 , n7276 );
not ( n8876 , n8875 );
or ( n8877 , n8874 , n8876 );
nand ( n8878 , n8877 , n7316 );
not ( n8879 , n7462 );
nand ( n8880 , n7678 , n7310 );
nor ( n8881 , n8880 , n7697 );
nor ( n8882 , n8879 , n8881 );
and ( n8883 , n8878 , n8882 );
nand ( n8884 , n7452 , n7275 );
nand ( n8885 , n7341 , n7435 );
nand ( n8886 , n8884 , n8833 , n8885 );
not ( n8887 , n7793 );
or ( n8888 , n8886 , n8887 );
or ( n8889 , n7315 , n7 );
not ( n8890 , n8889 );
nand ( n8891 , n8888 , n8890 );
and ( n8892 , n8869 , n8883 , n8891 );
nand ( n8893 , n8853 , n8892 );
not ( n8894 , n8893 );
not ( n8895 , n8894 );
or ( n8896 , n8759 , n8895 );
buf ( n8897 , n8893 );
nand ( n8898 , n8897 , n8757 );
nand ( n8899 , n8896 , n8898 );
not ( n8900 , n8899 );
and ( n8901 , n8636 , n8900 );
not ( n8902 , n8636 );
and ( n8903 , n8902 , n8899 );
nor ( n8904 , n8901 , n8903 );
and ( n8905 , n8514 , n8904 );
not ( n8906 , n8514 );
not ( n8907 , n8904 );
and ( n8908 , n8906 , n8907 );
nor ( n8909 , n8905 , n8908 );
or ( n8910 , n8909 , n1 );
and ( n8911 , n97 , n8634 );
not ( n8912 , n97 );
and ( n8913 , n8912 , n69 );
nor ( n8914 , n8911 , n8913 );
or ( n8915 , n2246 , n8914 );
nand ( n8916 , n8910 , n8915 );
buf ( n8917 , n6698 );
not ( n8918 , n8917 );
not ( n8919 , n8918 );
nand ( n8920 , n8168 , n6769 , n32 );
not ( n8921 , n8920 );
not ( n8922 , n7863 );
nand ( n8923 , n8922 , n6782 );
not ( n8924 , n8923 );
or ( n8925 , n8921 , n8924 );
not ( n8926 , n6727 );
not ( n8927 , n6883 );
or ( n8928 , n8926 , n8927 );
nand ( n8929 , n6736 , n27 );
not ( n8930 , n8929 );
nand ( n8931 , n8930 , n6799 );
nand ( n8932 , n8928 , n8931 );
buf ( n8933 , n8146 );
nor ( n8934 , n8932 , n8933 );
nand ( n8935 , n8925 , n8934 );
not ( n8936 , n8935 );
not ( n8937 , n6807 );
or ( n8938 , n8936 , n8937 );
nand ( n8939 , n6704 , n6925 , n6794 );
nand ( n8940 , n6875 , n8321 , n8939 );
and ( n8941 , n8940 , n33 );
nand ( n8942 , n6855 , n27 );
and ( n8943 , n8662 , n8942 , n8204 );
nor ( n8944 , n8943 , n6868 );
nor ( n8945 , n8941 , n8944 );
nand ( n8946 , n8938 , n8945 );
and ( n8947 , n6821 , n7996 , n6941 );
and ( n8948 , n8221 , n8947 , n7916 );
not ( n8949 , n6948 );
not ( n8950 , n8327 );
nand ( n8951 , n8950 , n6776 );
nor ( n8952 , n8949 , n8951 );
nor ( n8953 , n8948 , n8952 );
or ( n8954 , n8946 , n8953 );
not ( n8955 , n27 );
not ( n8956 , n6789 );
or ( n8957 , n8955 , n8956 );
nand ( n8958 , n8957 , n7844 );
nand ( n8959 , n6866 , n6923 );
nand ( n8960 , n8200 , n8958 , n8959 );
and ( n8961 , n8960 , n6782 );
nor ( n8962 , n8961 , n34 );
not ( n8963 , n7854 );
not ( n8964 , n6879 );
not ( n8965 , n8964 );
not ( n8966 , n8646 );
or ( n8967 , n8965 , n8966 );
nand ( n8968 , n8967 , n6706 );
nand ( n8969 , n8963 , n8968 );
nor ( n8970 , n8395 , n8372 , n33 );
nand ( n8971 , n6845 , n8970 );
or ( n8972 , n8969 , n8971 );
and ( n8973 , n6820 , n6782 );
not ( n8974 , n6838 );
nor ( n8975 , n8973 , n8974 );
not ( n8976 , n33 );
not ( n8977 , n8393 );
or ( n8978 , n8976 , n8977 );
nand ( n8979 , n8978 , n8736 );
nand ( n8980 , n8975 , n8979 );
nand ( n8981 , n8972 , n8980 );
not ( n8982 , n8360 );
not ( n8983 , n6845 );
or ( n8984 , n8982 , n8983 );
nand ( n8985 , n8984 , n32 );
nand ( n8986 , n8962 , n8981 , n8985 );
nand ( n8987 , n8954 , n8986 );
nand ( n8988 , n8169 , n6849 , n6782 );
or ( n8989 , n8988 , n8933 );
not ( n8990 , n7938 );
or ( n8991 , n7988 , n8990 );
nand ( n8992 , n8989 , n8991 );
nand ( n8993 , n8694 , n6837 );
not ( n8994 , n8993 );
nor ( n8995 , n8994 , n8159 );
and ( n8996 , n8992 , n8995 );
nor ( n8997 , n8996 , n33 );
not ( n8998 , n7961 );
not ( n8999 , n8140 );
and ( n9000 , n8998 , n8999 );
not ( n9001 , n8218 );
nor ( n9002 , n9000 , n9001 );
not ( n9003 , n8303 );
not ( n9004 , n8260 );
not ( n9005 , n9004 );
or ( n9006 , n9003 , n9005 );
nand ( n9007 , n9006 , n7838 );
not ( n9008 , n6778 );
not ( n9009 , n6874 );
or ( n9010 , n9008 , n9009 );
nand ( n9011 , n9010 , n8162 );
or ( n9012 , n9011 , n8214 );
nand ( n9013 , n9012 , n6869 );
nand ( n9014 , n9002 , n9007 , n9013 );
nor ( n9015 , n8997 , n9014 );
nand ( n9016 , n8987 , n9015 );
not ( n9017 , n9016 );
not ( n9018 , n9017 );
not ( n9019 , n8827 );
nand ( n9020 , n9019 , n8807 );
not ( n9021 , n7694 );
nand ( n9022 , n9021 , n4 );
not ( n9023 , n9022 );
or ( n9024 , n9020 , n9023 );
nand ( n9025 , n7769 , n7737 );
nand ( n9026 , n9024 , n9025 );
nand ( n9027 , n7231 , n7341 );
and ( n9028 , n8831 , n9027 );
nand ( n9029 , n9026 , n9028 );
not ( n9030 , n9029 );
not ( n9031 , n7400 );
not ( n9032 , n8786 );
not ( n9033 , n8777 );
or ( n9034 , n9032 , n9033 );
nand ( n9035 , n9034 , n7372 );
and ( n9036 , n9031 , n9035 , n7830 , n8885 );
and ( n9037 , n9030 , n9036 );
nor ( n9038 , n9037 , n8 );
nand ( n9039 , n7822 , n7337 );
nand ( n9040 , n7276 , n7682 );
and ( n9041 , n9040 , n7265 );
and ( n9042 , n9039 , n9041 , n7765 );
not ( n9043 , n9042 );
not ( n9044 , n7472 );
nand ( n9045 , n9044 , n7240 );
not ( n9046 , n9045 );
or ( n9047 , n9043 , n9046 );
nand ( n9048 , n7461 , n7240 );
nand ( n9049 , n9031 , n9048 , n7 );
nand ( n9050 , n9047 , n9049 );
nor ( n9051 , n8762 , n7805 );
nor ( n9052 , n9051 , n7457 );
not ( n9053 , n9052 );
not ( n9054 , n7671 );
or ( n9055 , n9053 , n9054 );
nand ( n9056 , n9055 , n7814 );
not ( n9057 , n9056 );
not ( n9058 , n8 );
or ( n9059 , n9057 , n9058 );
and ( n9060 , n7296 , n7733 );
nor ( n9061 , n9060 , n9 );
nand ( n9062 , n9059 , n9061 );
not ( n9063 , n9062 );
nand ( n9064 , n9050 , n9063 );
or ( n9065 , n9038 , n9064 );
not ( n9066 , n7271 );
not ( n9067 , n7716 );
or ( n9068 , n9066 , n9067 );
nand ( n9069 , n7444 , n7240 );
nand ( n9070 , n9069 , n7733 );
nand ( n9071 , n9068 , n9070 );
nand ( n9072 , n7357 , n7416 );
not ( n9073 , n9072 );
not ( n9074 , n7424 );
or ( n9075 , n9073 , n9074 );
nand ( n9076 , n9075 , n7265 );
not ( n9077 , n9076 );
nor ( n9078 , n9077 , n9023 );
nand ( n9079 , n9071 , n9078 );
nor ( n9080 , n9079 , n9029 );
buf ( n9081 , n8785 );
nand ( n9082 , n9081 , n8809 );
and ( n9083 , n7695 , n7337 );
or ( n9084 , n9082 , n9083 );
nand ( n9085 , n9084 , n7 );
nand ( n9086 , n8774 , n7290 );
and ( n9087 , n7369 , n8 , n9086 , n8835 );
and ( n9088 , n9085 , n9087 );
or ( n9089 , n9080 , n9088 );
nand ( n9090 , n8875 , n7718 );
not ( n9091 , n9090 );
and ( n9092 , n7435 , n7682 );
not ( n9093 , n9092 );
and ( n9094 , n8880 , n9093 , n8819 );
nand ( n9095 , n9091 , n9094 );
not ( n9096 , n7477 );
nor ( n9097 , n7381 , n7 );
nand ( n9098 , n9096 , n8885 , n9097 );
nand ( n9099 , n9095 , n9098 );
nand ( n9100 , n9089 , n9099 );
nand ( n9101 , n9065 , n9100 );
not ( n9102 , n9021 );
not ( n9103 , n9102 );
and ( n9104 , n9103 , n7722 );
nor ( n9105 , n9104 , n7759 );
nand ( n9106 , n9105 , n7364 );
nand ( n9107 , n9106 , n8863 );
nand ( n9108 , n7452 , n7438 );
and ( n9109 , n9107 , n9108 , n7760 );
not ( n9110 , n7265 );
not ( n9111 , n7687 );
or ( n9112 , n9110 , n9111 );
not ( n9113 , n8788 );
or ( n9114 , n9113 , n8890 );
nand ( n9115 , n9112 , n9114 );
nand ( n9116 , n9023 , n7349 );
and ( n9117 , n9109 , n9115 , n9116 );
nand ( n9118 , n9101 , n9117 );
not ( n9119 , n9118 );
not ( n9120 , n9119 );
or ( n9121 , n9018 , n9120 );
nand ( n9122 , n9118 , n9016 );
nand ( n9123 , n9121 , n9122 );
not ( n9124 , n9123 );
not ( n9125 , n9124 );
or ( n9126 , n8919 , n9125 );
nand ( n9127 , n8917 , n9123 );
nand ( n9128 , n9126 , n9127 );
not ( n9129 , n7075 );
not ( n9130 , n7046 );
not ( n9131 , n9130 );
and ( n9132 , n9129 , n9131 );
and ( n9133 , n7076 , n9130 );
nor ( n9134 , n9132 , n9133 );
and ( n9135 , n9134 , n7116 );
nor ( n9136 , n9135 , n7132 );
not ( n9137 , n9136 );
nand ( n9138 , n7123 , n7104 );
nand ( n9139 , n7124 , n9138 , n7511 , n16 );
and ( n9140 , n7568 , n7142 );
nor ( n9141 , n9139 , n9140 );
nand ( n9142 , n9141 , n7537 );
not ( n9143 , n9142 );
or ( n9144 , n9137 , n9143 );
nor ( n9145 , n7080 , n7636 );
nor ( n9146 , n7560 , n9145 );
nand ( n9147 , n8584 , n9146 );
and ( n9148 , n9147 , n7132 );
not ( n9149 , n6999 );
nand ( n9150 , n9149 , n6988 , n7097 , n15 );
nand ( n9151 , n7081 , n6971 );
nand ( n9152 , n9150 , n9151 );
and ( n9153 , n9152 , n7131 );
nor ( n9154 , n9148 , n9153 );
nand ( n9155 , n9144 , n9154 );
not ( n9156 , n9155 );
and ( n9157 , n7123 , n7170 );
nor ( n9158 , n7092 , n9157 );
nand ( n9159 , n7632 , n9158 );
not ( n9160 , n9159 );
nand ( n9161 , n7063 , n13 );
nor ( n9162 , n9161 , n7106 );
not ( n9163 , n9162 );
and ( n9164 , n9160 , n9163 );
and ( n9165 , n6995 , n17 );
not ( n9166 , n14 );
nand ( n9167 , n9166 , n7088 );
not ( n9168 , n9167 );
not ( n9169 , n7060 );
or ( n9170 , n9168 , n9169 );
nand ( n9171 , n9170 , n7006 );
nand ( n9172 , n7004 , n7052 );
and ( n9173 , n9165 , n9171 , n9172 , n8601 );
nor ( n9174 , n9164 , n9173 );
nand ( n9175 , n7197 , n7019 );
and ( n9176 , n9175 , n7006 );
nor ( n9177 , n9176 , n8594 );
nand ( n9178 , n8606 , n7164 );
nand ( n9179 , n7009 , n9178 );
nand ( n9180 , n9177 , n9150 , n9179 , n7222 );
or ( n9181 , n9174 , n9180 );
nand ( n9182 , n7512 , n12 );
not ( n9183 , n9182 );
nand ( n9184 , n7058 , n7056 );
not ( n9185 , n9184 );
or ( n9186 , n9183 , n9185 );
nand ( n9187 , n7550 , n16 );
nand ( n9188 , n9186 , n9187 );
nor ( n9189 , n7202 , n9188 );
nand ( n9190 , n7514 , n6978 );
and ( n9191 , n7051 , n7192 , n11 );
or ( n9192 , n9189 , n9190 , n9191 );
not ( n9193 , n8604 );
not ( n9194 , n7110 );
or ( n9195 , n9193 , n9194 );
nand ( n9196 , n9195 , n7099 );
nor ( n9197 , n7560 , n6978 );
nand ( n9198 , n9196 , n9197 );
nand ( n9199 , n9192 , n9198 );
not ( n9200 , n8578 );
nand ( n9201 , n7018 , n12 );
nand ( n9202 , n9200 , n7023 , n9201 , n7094 );
and ( n9203 , n9202 , n7552 );
and ( n9204 , n7176 , n9138 );
nor ( n9205 , n9204 , n7116 );
and ( n9206 , n7091 , n16 );
nand ( n9207 , n9206 , n7559 );
nor ( n9208 , n7184 , n6974 );
nand ( n9209 , n9208 , n6999 );
nand ( n9210 , n7081 , n7510 );
nand ( n9211 , n9207 , n9209 , n9210 , n10 );
nor ( n9212 , n9203 , n9205 , n9211 );
nand ( n9213 , n9199 , n9212 );
nand ( n9214 , n9181 , n9213 );
nand ( n9215 , n9156 , n9214 );
not ( n9216 , n9215 );
not ( n9217 , n9216 );
not ( n9218 , n7484 );
not ( n9219 , n9218 );
or ( n9220 , n9217 , n9219 );
not ( n9221 , n9215 );
or ( n9222 , n9221 , n9218 );
nand ( n9223 , n9220 , n9222 );
not ( n9224 , n9223 );
and ( n9225 , n43 , n9224 );
not ( n9226 , n43 );
and ( n9227 , n9226 , n9223 );
nor ( n9228 , n9225 , n9227 );
not ( n9229 , n9228 );
and ( n9230 , n9128 , n9229 );
not ( n9231 , n9128 );
and ( n9232 , n9231 , n9228 );
nor ( n9233 , n9230 , n9232 );
or ( n9234 , n9233 , n1 );
xnor ( n9235 , n43 , n44 );
or ( n9236 , n2246 , n9235 );
nand ( n9237 , n9234 , n9236 );
not ( n9238 , n73 );
not ( n9239 , n8630 );
or ( n9240 , n9238 , n9239 );
not ( n9241 , n73 );
nand ( n9242 , n9241 , n8629 );
nand ( n9243 , n9240 , n9242 );
not ( n9244 , n9216 );
not ( n9245 , n7543 );
nand ( n9246 , n7135 , n7046 );
nor ( n9247 , n7589 , n17 );
and ( n9248 , n9246 , n9247 );
not ( n9249 , n9248 );
or ( n9250 , n9245 , n9249 );
not ( n9251 , n7215 );
not ( n9252 , n7621 );
or ( n9253 , n9251 , n9252 );
not ( n9254 , n8532 );
nand ( n9255 , n9253 , n9254 );
nand ( n9256 , n7660 , n7013 );
and ( n9257 , n7609 , n9256 , n17 );
nand ( n9258 , n9255 , n9257 );
nand ( n9259 , n9250 , n9258 );
not ( n9260 , n9259 );
not ( n9261 , n7593 );
and ( n9262 , n8532 , n7132 , n9261 );
not ( n9263 , n7141 );
nand ( n9264 , n9263 , n7524 );
and ( n9265 , n9206 , n9264 );
nor ( n9266 , n9262 , n9265 );
not ( n9267 , n9266 );
or ( n9268 , n9260 , n9267 );
nand ( n9269 , n9268 , n7222 );
not ( n9270 , n7574 );
and ( n9271 , n7047 , n9270 );
not ( n9272 , n9271 );
or ( n9273 , n7525 , n7153 );
nand ( n9274 , n7184 , n9151 );
nand ( n9275 , n9273 , n9274 );
not ( n9276 , n9275 );
or ( n9277 , n9272 , n9276 );
nand ( n9278 , n9277 , n17 );
nor ( n9279 , n7621 , n9130 );
nor ( n9280 , n7035 , n7038 , n7215 );
nor ( n9281 , n9279 , n9280 );
not ( n9282 , n7018 );
not ( n9283 , n7046 );
or ( n9284 , n9282 , n9283 );
not ( n9285 , n8532 );
not ( n9286 , n7188 );
and ( n9287 , n9285 , n9286 );
and ( n9288 , n7175 , n6983 );
nor ( n9289 , n9287 , n9288 );
nand ( n9290 , n9284 , n9289 );
nand ( n9291 , n9290 , n7084 );
and ( n9292 , n9278 , n9281 , n9291 );
not ( n9293 , n7116 );
not ( n9294 , n9140 );
or ( n9295 , n9293 , n9294 );
not ( n9296 , n7211 );
nand ( n9297 , n15 , n6988 );
not ( n9298 , n9297 );
or ( n9299 , n9296 , n9298 );
not ( n9300 , n17 );
nand ( n9301 , n9299 , n9300 );
nor ( n9302 , n7033 , n13 );
nor ( n9303 , n9301 , n9302 );
nand ( n9304 , n9295 , n9303 );
not ( n9305 , n7044 );
not ( n9306 , n8524 );
or ( n9307 , n9305 , n9306 );
nand ( n9308 , n9307 , n7206 );
not ( n9309 , n9308 );
not ( n9310 , n16 );
or ( n9311 , n9309 , n9310 );
buf ( n9312 , n9209 );
nand ( n9313 , n9311 , n9312 );
or ( n9314 , n9304 , n9313 );
not ( n9315 , n7185 );
or ( n9316 , n7636 , n16 );
nand ( n9317 , n9316 , n7003 , n17 );
or ( n9318 , n9315 , n9317 );
nand ( n9319 , n9314 , n9318 );
nand ( n9320 , n7123 , n7567 );
nand ( n9321 , n9320 , n16 );
nor ( n9322 , n9288 , n9321 );
not ( n9323 , n9322 );
not ( n9324 , n7093 );
or ( n9325 , n9323 , n9324 );
not ( n9326 , n16 );
nand ( n9327 , n9326 , n7524 );
or ( n9328 , n9327 , n7168 );
nand ( n9329 , n9328 , n7098 );
nand ( n9330 , n9329 , n9210 , n8606 );
nand ( n9331 , n9325 , n9330 );
nor ( n9332 , n7558 , n8517 );
nand ( n9333 , n9331 , n9332 );
not ( n9334 , n9333 );
nand ( n9335 , n9319 , n9334 );
nand ( n9336 , n9335 , n10 );
not ( n9337 , n8594 );
not ( n9338 , n9337 );
nor ( n9339 , n7103 , n11 );
and ( n9340 , n9339 , n7033 );
nor ( n9341 , n7511 , n12 );
nor ( n9342 , n9340 , n9341 , n16 );
not ( n9343 , n9342 );
not ( n9344 , n7537 );
or ( n9345 , n9343 , n9344 );
nand ( n9346 , n7519 , n6977 );
nand ( n9347 , n9345 , n9346 );
not ( n9348 , n9347 );
or ( n9349 , n9338 , n9348 );
nand ( n9350 , n9349 , n6978 );
nand ( n9351 , n9269 , n9292 , n9336 , n9350 );
not ( n9352 , n9351 );
not ( n9353 , n9352 );
or ( n9354 , n9244 , n9353 );
not ( n9355 , n9221 );
nand ( n9356 , n9351 , n9355 );
nand ( n9357 , n9354 , n9356 );
xnor ( n9358 , n9243 , n9357 );
not ( n9359 , n9218 );
not ( n9360 , n7733 );
not ( n9361 , n7714 );
not ( n9362 , n7818 );
or ( n9363 , n9361 , n9362 );
nand ( n9364 , n9363 , n7241 );
nand ( n9365 , n7722 , n7355 );
not ( n9366 , n9365 );
not ( n9367 , n7744 );
nor ( n9368 , n9360 , n9364 , n9366 , n9367 );
and ( n9369 , n7795 , n7 , n9027 , n7315 );
or ( n9370 , n9368 , n9369 );
nand ( n9371 , n9370 , n8792 );
and ( n9372 , n7290 , n7230 );
and ( n9373 , n7295 , n5 );
nand ( n9374 , n7385 , n7677 );
nor ( n9375 , n9373 , n9374 );
nor ( n9376 , n9372 , n9375 );
not ( n9377 , n9376 );
not ( n9378 , n8880 );
not ( n9379 , n7426 );
or ( n9380 , n9378 , n9379 );
nand ( n9381 , n9380 , n7 );
not ( n9382 , n9381 );
or ( n9383 , n9377 , n9382 );
not ( n9384 , n7781 );
nand ( n9385 , n9383 , n9384 );
or ( n9386 , n7819 , n6 );
not ( n9387 , n8 );
not ( n9388 , n7322 );
or ( n9389 , n9387 , n9388 );
nand ( n9390 , n9389 , n7828 );
nand ( n9391 , n9386 , n9390 );
nand ( n9392 , n7687 , n7760 );
nor ( n9393 , n9391 , n9392 );
nand ( n9394 , n9385 , n9393 );
nand ( n9395 , n9371 , n9394 );
not ( n9396 , n7824 );
nand ( n9397 , n9102 , n9396 );
and ( n9398 , n9397 , n7316 );
and ( n9399 , n7286 , n7436 );
nor ( n9400 , n9399 , n7287 );
nor ( n9401 , n9398 , n9400 , n9 );
not ( n9402 , n9401 );
and ( n9403 , n7420 , n7460 );
nor ( n9404 , n9403 , n3 );
not ( n9405 , n3 );
not ( n9406 , n7446 );
or ( n9407 , n9405 , n9406 );
nand ( n9408 , n9021 , n7276 );
nand ( n9409 , n9407 , n9408 );
or ( n9410 , n9404 , n9409 );
not ( n9411 , n7240 );
not ( n9412 , n7419 );
or ( n9413 , n9411 , n9412 );
nand ( n9414 , n9413 , n7 );
nand ( n9415 , n9410 , n9414 );
not ( n9416 , n7701 );
nand ( n9417 , n9415 , n9416 );
not ( n9418 , n9409 );
nand ( n9419 , n9048 , n8 );
not ( n9420 , n9419 );
and ( n9421 , n9418 , n9420 );
nor ( n9422 , n9421 , n8863 );
nand ( n9423 , n9417 , n9422 );
not ( n9424 , n9423 );
or ( n9425 , n9402 , n9424 );
not ( n9426 , n7291 );
not ( n9427 , n8844 );
not ( n9428 , n7354 );
or ( n9429 , n9427 , n9428 );
nand ( n9430 , n9429 , n7 );
not ( n9431 , n9430 );
or ( n9432 , n9426 , n9431 );
nand ( n9433 , n9432 , n4 );
not ( n9434 , n7743 );
not ( n9435 , n6 );
not ( n9436 , n7677 );
or ( n9437 , n9435 , n9436 );
nand ( n9438 , n9437 , n7722 );
and ( n9439 , n9434 , n9438 , n7315 );
nand ( n9440 , n9433 , n9108 , n9439 );
nor ( n9441 , n7315 , n7341 );
not ( n9442 , n9441 );
not ( n9443 , n7362 );
or ( n9444 , n9442 , n9443 );
nand ( n9445 , n9444 , n7828 );
nand ( n9446 , n8807 , n9445 );
nand ( n9447 , n9440 , n9446 );
not ( n9448 , n7265 );
not ( n9449 , n4 );
not ( n9450 , n7446 );
or ( n9451 , n9449 , n9450 );
nand ( n9452 , n9451 , n7280 );
not ( n9453 , n9452 );
or ( n9454 , n9448 , n9453 );
nand ( n9455 , n9454 , n8826 );
not ( n9456 , n7349 );
not ( n9457 , n7435 );
nand ( n9458 , n9457 , n7284 );
not ( n9459 , n9458 );
or ( n9460 , n9456 , n9459 );
nand ( n9461 , n9460 , n7817 );
nor ( n9462 , n9455 , n9461 );
nor ( n9463 , n8811 , n8834 );
not ( n9464 , n9463 );
nand ( n9465 , n7720 , n7369 );
or ( n9466 , n9464 , n9465 );
nand ( n9467 , n9466 , n7 );
nand ( n9468 , n9447 , n9462 , n9467 );
nand ( n9469 , n9425 , n9468 );
and ( n9470 , n7296 , n7265 , n5 );
not ( n9471 , n7342 );
and ( n9472 , n9471 , n7 );
nor ( n9473 , n9470 , n9472 );
and ( n9474 , n9395 , n9469 , n9473 );
not ( n9475 , n9474 );
or ( n9476 , n9359 , n9475 );
or ( n9477 , n7490 , n9474 );
nand ( n9478 , n9476 , n9477 );
or ( n9479 , n6614 , n6541 , n6447 );
nand ( n9480 , n9479 , n6470 );
nand ( n9481 , n6637 , n9480 );
nand ( n9482 , n6519 , n23 );
nand ( n9483 , n8037 , n23 );
nand ( n9484 , n9482 , n9483 );
or ( n9485 , n9481 , n9484 );
nor ( n9486 , n6405 , n26 );
not ( n9487 , n9486 );
not ( n9488 , n6288 );
or ( n9489 , n9487 , n9488 );
nand ( n9490 , n9489 , n6448 );
not ( n9491 , n8491 );
nand ( n9492 , n9491 , n6510 );
and ( n9493 , n9492 , n8123 );
nand ( n9494 , n9490 , n9493 );
nand ( n9495 , n9485 , n9494 );
nor ( n9496 , n6378 , n19 );
nand ( n9497 , n9495 , n9496 );
not ( n9498 , n6382 );
not ( n9499 , n6443 );
nand ( n9500 , n9499 , n6447 );
not ( n9501 , n9500 );
and ( n9502 , n9498 , n9501 );
not ( n9503 , n8421 );
and ( n9504 , n9503 , n23 );
nor ( n9505 , n9502 , n9504 );
not ( n9506 , n8076 );
not ( n9507 , n9506 );
nand ( n9508 , n9507 , n8469 );
or ( n9509 , n9505 , n9508 );
nor ( n9510 , n6443 , n6447 );
and ( n9511 , n6489 , n9510 );
not ( n9512 , n6382 );
nand ( n9513 , n9511 , n9512 , n8491 );
nand ( n9514 , n9509 , n9513 );
and ( n9515 , n9514 , n8431 );
not ( n9516 , n9492 );
nor ( n9517 , n9516 , n8478 , n25 );
nor ( n9518 , n9515 , n9517 );
or ( n9519 , n9497 , n9518 );
and ( n9520 , n8469 , n6298 , n6588 , n6674 );
or ( n9521 , n9520 , n25 );
nor ( n9522 , n6468 , n21 );
not ( n9523 , n6563 );
nor ( n9524 , n6404 , n6299 );
nor ( n9525 , n9522 , n9523 , n9524 , n6539 );
nand ( n9526 , n9521 , n9525 );
not ( n9527 , n8020 );
nand ( n9528 , n9527 , n26 );
not ( n9529 , n9528 );
not ( n9530 , n8061 );
or ( n9531 , n6566 , n9530 );
nand ( n9532 , n9531 , n25 );
nand ( n9533 , n6676 , n6409 );
and ( n9534 , n9532 , n9533 , n6693 );
and ( n9535 , n9529 , n9534 );
or ( n9536 , n6507 , n6431 );
and ( n9537 , n9536 , n24 );
nand ( n9538 , n8046 , n6356 );
nand ( n9539 , n9538 , n6331 , n6674 , n6320 );
nor ( n9540 , n9537 , n9539 );
nor ( n9541 , n9535 , n9540 );
or ( n9542 , n9526 , n9541 );
nand ( n9543 , n9519 , n9542 );
and ( n9544 , n8113 , n6525 );
not ( n9545 , n6496 );
nor ( n9546 , n9544 , n9523 , n9545 );
or ( n9547 , n9546 , n6299 );
nor ( n9548 , n9512 , n6467 );
not ( n9549 , n6489 );
not ( n9550 , n8072 );
not ( n9551 , n9550 );
or ( n9552 , n9549 , n9551 );
nand ( n9553 , n9552 , n6445 );
or ( n9554 , n9548 , n9553 );
nand ( n9555 , n9554 , n6299 );
nand ( n9556 , n9547 , n9555 , n26 );
not ( n9557 , n8084 );
and ( n9558 , n9557 , n8109 , n6475 );
not ( n9559 , n6429 );
nor ( n9560 , n9559 , n6356 );
not ( n9561 , n9560 );
not ( n9562 , n6287 );
not ( n9563 , n6506 );
not ( n9564 , n9563 );
or ( n9565 , n9562 , n9564 );
nand ( n9566 , n9565 , n8092 );
nor ( n9567 , n9561 , n9566 );
or ( n9568 , n9558 , n9567 );
and ( n9569 , n8093 , n6483 , n6447 );
nand ( n9570 , n9568 , n9569 );
and ( n9571 , n9556 , n9570 );
and ( n9572 , n6421 , n8119 );
nor ( n9573 , n9572 , n6314 );
nor ( n9574 , n9571 , n9573 );
nand ( n9575 , n9543 , n9574 );
or ( n9576 , n8757 , n9575 );
nand ( n9577 , n9575 , n8757 );
nand ( n9578 , n9576 , n9577 );
not ( n9579 , n9578 );
and ( n9580 , n9478 , n9579 );
not ( n9581 , n9478 );
and ( n9582 , n9581 , n9578 );
nor ( n9583 , n9580 , n9582 );
and ( n9584 , n9358 , n9583 );
not ( n9585 , n9358 );
not ( n9586 , n9583 );
and ( n9587 , n9585 , n9586 );
nor ( n9588 , n9584 , n9587 );
or ( n9589 , n9588 , n1 );
and ( n9590 , n74 , n9241 );
not ( n9591 , n74 );
and ( n9592 , n9591 , n73 );
nor ( n9593 , n9590 , n9592 );
or ( n9594 , n2246 , n9593 );
nand ( n9595 , n9589 , n9594 );
not ( n9596 , n5745 );
not ( n9597 , n5696 );
or ( n9598 , n9596 , n9597 );
nand ( n9599 , n9598 , n5778 );
nand ( n9600 , n5912 , n3529 );
and ( n9601 , n3605 , n9600 );
not ( n9602 , n3605 );
and ( n9603 , n9602 , n5261 );
nor ( n9604 , n9601 , n9603 );
not ( n9605 , n9604 );
not ( n9606 , n208 );
not ( n9607 , n5961 );
or ( n9608 , n9606 , n9607 );
not ( n9609 , n5366 );
not ( n9610 , n208 );
nand ( n9611 , n9610 , n3678 );
nor ( n9612 , n9611 , n3589 );
nor ( n9613 , n9609 , n9612 );
nand ( n9614 , n9608 , n9613 );
not ( n9615 , n9614 );
not ( n9616 , n9615 );
or ( n9617 , n9605 , n9616 );
not ( n9618 , n9600 );
and ( n9619 , n9618 , n3697 );
and ( n9620 , n5939 , n3630 );
nor ( n9621 , n9619 , n9620 );
nand ( n9622 , n9617 , n9621 );
nand ( n9623 , n3455 , n3630 );
not ( n9624 , n3667 );
and ( n9625 , n9623 , n9624 );
nand ( n9626 , n9622 , n9625 );
not ( n9627 , n4225 );
nand ( n9628 , n9627 , n211 );
nor ( n9629 , n9614 , n9628 );
or ( n9630 , n9629 , n5376 );
nand ( n9631 , n3685 , n5323 );
nand ( n9632 , n9631 , n3697 );
and ( n9633 , n9632 , n4217 );
nand ( n9634 , n9630 , n9633 );
nand ( n9635 , n9626 , n9634 );
not ( n9636 , n4251 );
nand ( n9637 , n9636 , n5951 );
and ( n9638 , n9637 , n3697 );
nor ( n9639 , n9638 , n212 );
nand ( n9640 , n9635 , n9639 );
not ( n9641 , n3471 );
and ( n9642 , n3455 , n3605 );
not ( n9643 , n9642 );
or ( n9644 , n9641 , n9643 );
not ( n9645 , n5302 );
nand ( n9646 , n3653 , n209 );
nand ( n9647 , n3630 , n5261 );
and ( n9648 , n9645 , n9646 , n9647 );
nand ( n9649 , n9644 , n9648 );
not ( n9650 , n5383 );
not ( n9651 , n9650 );
not ( n9652 , n4326 );
not ( n9653 , n9652 );
or ( n9654 , n9651 , n9653 );
not ( n9655 , n209 );
nand ( n9656 , n9654 , n9655 );
not ( n9657 , n9656 );
or ( n9658 , n9649 , n9657 );
nand ( n9659 , n9658 , n3619 );
not ( n9660 , n3464 );
not ( n9661 , n3619 );
and ( n9662 , n9660 , n9661 );
not ( n9663 , n5357 );
nand ( n9664 , n3533 , n9663 );
nor ( n9665 , n5940 , n9664 );
not ( n9666 , n5376 );
or ( n9667 , n9665 , n9666 );
nand ( n9668 , n5360 , n3468 , n4275 );
nand ( n9669 , n9667 , n9668 );
nor ( n9670 , n9662 , n9669 );
and ( n9671 , n3679 , n9627 , n5288 );
not ( n9672 , n9671 );
not ( n9673 , n5337 );
not ( n9674 , n9673 );
or ( n9675 , n9672 , n9674 );
nand ( n9676 , n5906 , n3471 );
not ( n9677 , n9676 );
nor ( n9678 , n5975 , n4236 );
nand ( n9679 , n9677 , n9678 );
nand ( n9680 , n9675 , n9679 );
nand ( n9681 , n9659 , n9670 , n9680 );
nand ( n9682 , n9640 , n9681 );
nand ( n9683 , n5989 , n3605 );
not ( n9684 , n9683 );
not ( n9685 , n4242 );
or ( n9686 , n9684 , n9685 );
nand ( n9687 , n9686 , n3462 );
nand ( n9688 , n4213 , n5384 , n9687 );
not ( n9689 , n9688 );
not ( n9690 , n209 );
or ( n9691 , n9689 , n9690 );
nand ( n9692 , n9691 , n211 );
not ( n9693 , n5384 );
nand ( n9694 , n5989 , n3543 );
and ( n9695 , n9694 , n3611 , n3636 );
not ( n9696 , n9695 );
or ( n9697 , n9693 , n9696 );
nand ( n9698 , n4241 , n3582 );
not ( n9699 , n209 );
nand ( n9700 , n3567 , n9698 , n9699 );
nand ( n9701 , n9697 , n9700 );
nand ( n9702 , n3671 , n206 );
nand ( n9703 , n9701 , n9702 , n3647 );
and ( n9704 , n9692 , n9703 );
nand ( n9705 , n3699 , n5980 );
nand ( n9706 , n9705 , n3693 , n5303 , n3524 );
nor ( n9707 , n9704 , n9706 );
nand ( n9708 , n9682 , n9707 );
not ( n9709 , n9708 );
not ( n9710 , n9709 );
not ( n9711 , n3812 );
not ( n9712 , n3931 );
or ( n9713 , n9711 , n9712 );
nand ( n9714 , n4892 , n3832 );
nand ( n9715 , n9713 , n9714 );
not ( n9716 , n9715 );
not ( n9717 , n4989 );
and ( n9718 , n3803 , n3829 );
nor ( n9719 , n9717 , n9718 );
not ( n9720 , n9719 );
or ( n9721 , n9716 , n9720 );
nand ( n9722 , n4798 , n3830 , n185 );
nand ( n9723 , n9721 , n9722 );
not ( n9724 , n9723 );
not ( n9725 , n4722 );
not ( n9726 , n3854 );
and ( n9727 , n9725 , n9726 );
not ( n9728 , n4797 );
not ( n9729 , n5435 );
nor ( n9730 , n9729 , n184 );
and ( n9731 , n9728 , n9730 );
nor ( n9732 , n9727 , n9731 );
not ( n9733 , n3955 );
nand ( n9734 , n9733 , n5428 , n3749 );
or ( n9735 , n9732 , n9734 );
nor ( n9736 , n3755 , n185 );
or ( n9737 , n9736 , n3949 );
nand ( n9738 , n4669 , n4944 );
nand ( n9739 , n9737 , n9738 );
nand ( n9740 , n9739 , n4873 , n186 );
nand ( n9741 , n9735 , n9740 );
not ( n9742 , n9741 );
or ( n9743 , n9724 , n9742 );
nand ( n9744 , n9743 , n5007 );
nand ( n9745 , n3861 , n4789 );
and ( n9746 , n4709 , n9745 );
not ( n9747 , n9746 );
not ( n9748 , n4773 );
or ( n9749 , n9747 , n9748 );
nand ( n9750 , n9749 , n3811 );
or ( n9751 , n3764 , n3952 );
nand ( n9752 , n9751 , n185 );
and ( n9753 , n4977 , n9752 , n3749 );
nand ( n9754 , n9750 , n9753 );
nand ( n9755 , n4824 , n186 );
nand ( n9756 , n4661 , n3888 );
nand ( n9757 , n4817 , n9756 );
nor ( n9758 , n9755 , n9757 );
or ( n9759 , n9758 , n5007 );
not ( n9760 , n183 );
not ( n9761 , n3908 );
or ( n9762 , n9760 , n9761 );
nand ( n9763 , n9762 , n5073 );
nor ( n9764 , n9763 , n4710 );
or ( n9765 , n9764 , n3782 );
nand ( n9766 , n9759 , n9765 );
and ( n9767 , n9754 , n9766 );
and ( n9768 , n3772 , n3901 , n3811 );
nor ( n9769 , n9768 , n5007 );
not ( n9770 , n9769 );
not ( n9771 , n5013 );
nand ( n9772 , n4995 , n185 );
not ( n9773 , n9772 );
nand ( n9774 , n9771 , n5466 , n4946 , n9773 );
not ( n9775 , n9774 );
or ( n9776 , n9770 , n9775 );
and ( n9777 , n4979 , n4697 , n3941 );
nand ( n9778 , n9776 , n9777 );
nor ( n9779 , n9767 , n9778 );
not ( n9780 , n4761 );
nor ( n9781 , n4978 , n185 );
not ( n9782 , n9781 );
or ( n9783 , n9780 , n9782 );
or ( n9784 , n4805 , n3922 );
nand ( n9785 , n9784 , n5002 );
nand ( n9786 , n9783 , n9785 );
not ( n9787 , n3922 );
or ( n9788 , n5001 , n9787 );
not ( n9789 , n3765 );
nand ( n9790 , n9788 , n9789 );
buf ( n9791 , n4751 );
and ( n9792 , n9790 , n5051 , n9791 );
nand ( n9793 , n9786 , n9792 );
or ( n9794 , n3765 , n3922 );
nand ( n9795 , n4856 , n4841 );
nand ( n9796 , n9794 , n9795 );
nand ( n9797 , n9793 , n9796 );
not ( n9798 , n3741 );
nand ( n9799 , n9798 , n180 );
and ( n9800 , n5052 , n186 );
and ( n9801 , n9799 , n4872 , n9800 );
nor ( n9802 , n9801 , n5034 );
nand ( n9803 , n9793 , n9802 );
nand ( n9804 , n9744 , n9779 , n9797 , n9803 );
not ( n9805 , n9804 );
not ( n9806 , n9805 );
or ( n9807 , n9710 , n9806 );
not ( n9808 , n9709 );
nand ( n9809 , n9804 , n9808 );
nand ( n9810 , n9807 , n9809 );
xor ( n9811 , n9599 , n9810 );
not ( n9812 , n196 );
not ( n9813 , n9812 );
not ( n9814 , n4954 );
not ( n9815 , n9814 );
not ( n9816 , n6155 );
or ( n9817 , n9815 , n9816 );
nand ( n9818 , n4954 , n6154 );
nand ( n9819 , n9817 , n9818 );
not ( n9820 , n9819 );
or ( n9821 , n9813 , n9820 );
or ( n9822 , n9819 , n9812 );
nand ( n9823 , n9821 , n9822 );
xnor ( n9824 , n9811 , n9823 );
or ( n9825 , n9824 , n1 );
and ( n9826 , n213 , n9812 );
not ( n9827 , n213 );
and ( n9828 , n9827 , n196 );
nor ( n9829 , n9826 , n9828 );
or ( n9830 , n2246 , n9829 );
nand ( n9831 , n9825 , n9830 );
not ( n9832 , n124 );
not ( n9833 , n2970 );
not ( n9834 , n9833 );
or ( n9835 , n9832 , n9834 );
nand ( n9836 , n2919 , n121 );
nand ( n9837 , n9836 , n2897 );
nand ( n9838 , n9837 , n122 );
nand ( n9839 , n9835 , n9838 );
buf ( n9840 , n2909 );
nand ( n9841 , n2938 , n9840 );
nand ( n9842 , n9841 , n2785 );
not ( n9843 , n9842 );
and ( n9844 , n123 , n124 );
not ( n9845 , n9844 );
not ( n9846 , n9845 );
nand ( n9847 , n9846 , n121 );
nor ( n9848 , n9847 , n2816 );
not ( n9849 , n9848 );
nand ( n9850 , n9843 , n9849 );
or ( n9851 , n9839 , n9850 );
not ( n9852 , n2845 );
not ( n9853 , n9837 );
not ( n9854 , n9853 );
or ( n9855 , n9852 , n9854 );
nand ( n9856 , n9855 , n120 );
nand ( n9857 , n2832 , n2977 );
nor ( n9858 , n9857 , n121 );
nor ( n9859 , n9858 , n2785 );
nor ( n9860 , n122 , n124 );
nor ( n9861 , n9860 , n2908 );
nand ( n9862 , n2968 , n121 );
not ( n9863 , n9862 );
and ( n9864 , n9861 , n9863 );
nand ( n9865 , n2815 , n2780 );
not ( n9866 , n9865 );
nand ( n9867 , n9866 , n122 );
not ( n9868 , n9867 );
nor ( n9869 , n9864 , n9868 );
nand ( n9870 , n9856 , n9859 , n9869 );
nand ( n9871 , n9851 , n9870 );
not ( n9872 , n9871 );
not ( n9873 , n2788 );
not ( n9874 , n9873 );
nand ( n9875 , n2832 , n9874 );
not ( n9876 , n9875 );
nand ( n9877 , n9876 , n2828 );
not ( n9878 , n2835 );
nand ( n9879 , n9878 , n2854 );
and ( n9880 , n9877 , n9879 , n127 );
not ( n9881 , n2834 );
not ( n9882 , n2816 );
or ( n9883 , n9881 , n9882 );
nor ( n9884 , n122 , n124 );
not ( n9885 , n9884 );
nor ( n9886 , n9885 , n125 );
not ( n9887 , n9886 );
nand ( n9888 , n9883 , n9887 );
not ( n9889 , n2811 );
or ( n9890 , n9888 , n9889 );
nand ( n9891 , n9890 , n2785 );
not ( n9892 , n9891 );
nand ( n9893 , n121 , n125 );
not ( n9894 , n9893 );
nand ( n9895 , n2815 , n9894 );
and ( n9896 , n9895 , n2960 );
not ( n9897 , n9896 );
not ( n9898 , n2934 );
nor ( n9899 , n9897 , n9898 );
not ( n9900 , n9899 );
or ( n9901 , n9892 , n9900 );
nand ( n9902 , n9901 , n2857 );
nor ( n9903 , n124 , n125 );
and ( n9904 , n2810 , n9903 );
not ( n9905 , n9857 );
or ( n9906 , n9904 , n9905 );
buf ( n9907 , n2886 );
nand ( n9908 , n9906 , n9907 );
and ( n9909 , n9880 , n9902 , n9908 );
not ( n9910 , n9909 );
or ( n9911 , n9872 , n9910 );
buf ( n9912 , n2815 );
not ( n9913 , n9912 );
not ( n9914 , n2967 );
or ( n9915 , n9913 , n9914 );
nand ( n9916 , n9915 , n2844 );
not ( n9917 , n9847 );
or ( n9918 , n9916 , n9917 );
not ( n9919 , n120 );
nand ( n9920 , n9918 , n9919 );
not ( n9921 , n2911 );
and ( n9922 , n2920 , n9921 );
and ( n9923 , n9920 , n9922 );
nand ( n9924 , n2977 , n121 );
and ( n9925 , n2855 , n9924 );
not ( n9926 , n9925 );
or ( n9927 , n9926 , n126 );
nor ( n9928 , n120 , n126 );
not ( n9929 , n9928 );
nand ( n9930 , n9927 , n9929 );
and ( n9931 , n9923 , n9930 , n2966 );
nand ( n9932 , n3007 , n2832 );
not ( n9933 , n9932 );
not ( n9934 , n2857 );
and ( n9935 , n9933 , n9934 );
not ( n9936 , n9874 );
nand ( n9937 , n2824 , n123 );
not ( n9938 , n9937 );
not ( n9939 , n9938 );
or ( n9940 , n9936 , n9939 );
and ( n9941 , n2909 , n120 );
nand ( n9942 , n3006 , n9941 );
nand ( n9943 , n9940 , n9942 );
nor ( n9944 , n9935 , n9943 );
and ( n9945 , n9944 , n9859 );
or ( n9946 , n9931 , n9945 );
nand ( n9947 , n9860 , n125 );
nand ( n9948 , n9947 , n2978 );
and ( n9949 , n9948 , n2940 );
and ( n9950 , n120 , n125 );
buf ( n9951 , n9950 );
nand ( n9952 , n3006 , n9951 );
nand ( n9953 , n9952 , n2942 );
nor ( n9954 , n9949 , n9953 );
not ( n9955 , n2958 );
not ( n9956 , n2917 );
or ( n9957 , n9955 , n9956 );
nand ( n9958 , n9886 , n2987 );
nand ( n9959 , n9957 , n9958 );
nand ( n9960 , n124 , n125 );
nor ( n9961 , n2968 , n9960 );
not ( n9962 , n9961 );
not ( n9963 , n9962 );
nor ( n9964 , n9959 , n9963 );
nand ( n9965 , n2965 , n125 );
and ( n9966 , n9954 , n9964 , n9965 );
nand ( n9967 , n9946 , n9966 );
nand ( n9968 , n9911 , n9967 );
not ( n9969 , n2785 );
not ( n9970 , n2966 );
or ( n9971 , n9969 , n9970 );
nand ( n9972 , n9971 , n2797 );
not ( n9973 , n9963 );
not ( n9974 , n9973 );
not ( n9975 , n120 );
and ( n9976 , n9974 , n9975 );
not ( n9977 , n9907 );
nor ( n9978 , n9977 , n2855 );
nor ( n9979 , n9976 , n9978 );
nand ( n9980 , n9972 , n9979 );
nand ( n9981 , n2864 , n2824 );
and ( n9982 , n9981 , n126 );
and ( n9983 , n2940 , n2842 );
not ( n9984 , n3000 );
nor ( n9985 , n9983 , n9984 );
not ( n9986 , n2978 );
buf ( n9987 , n2780 );
nand ( n9988 , n9986 , n9987 );
nand ( n9989 , n9982 , n9985 , n9877 , n9988 );
and ( n9990 , n9980 , n9989 );
or ( n9991 , n9921 , n120 );
buf ( n9992 , n9838 );
nand ( n9993 , n9991 , n9992 );
nor ( n9994 , n9990 , n9993 );
nand ( n9995 , n9968 , n9994 );
not ( n9996 , n9995 );
not ( n9997 , n9996 );
nand ( n9998 , n3160 , n116 );
not ( n9999 , n9998 );
nand ( n10000 , n9999 , n3037 );
and ( n10001 , n10000 , n119 );
not ( n10002 , n3209 );
nor ( n10003 , n3047 , n115 );
buf ( n10004 , n10003 );
nor ( n10005 , n10002 , n10004 );
not ( n10006 , n10005 );
nand ( n10007 , n113 , n114 );
not ( n10008 , n10007 );
nand ( n10009 , n10008 , n3052 );
and ( n10010 , n9998 , n10009 );
not ( n10011 , n10010 );
or ( n10012 , n10006 , n10011 );
nand ( n10013 , n10012 , n3164 );
nor ( n10014 , n10007 , n115 );
nand ( n10015 , n10014 , n3257 );
not ( n10016 , n10015 );
not ( n10017 , n3117 );
or ( n10018 , n10016 , n10017 );
nand ( n10019 , n10018 , n117 );
buf ( n10020 , n3070 );
not ( n10021 , n10020 );
or ( n10022 , n3062 , n10021 );
nand ( n10023 , n3052 , n112 );
nand ( n10024 , n10022 , n10023 );
not ( n10025 , n3042 );
nand ( n10026 , n10024 , n10025 );
and ( n10027 , n10019 , n10026 );
nand ( n10028 , n10001 , n10013 , n10027 );
nand ( n10029 , n9998 , n3117 );
not ( n10030 , n3045 );
nand ( n10031 , n3144 , n10030 );
buf ( n10032 , n3180 );
nor ( n10033 , n10032 , n115 );
not ( n10034 , n10033 );
not ( n10035 , n118 );
nand ( n10036 , n10035 , n117 );
not ( n10037 , n10036 );
and ( n10038 , n10031 , n10034 , n10037 );
nand ( n10039 , n3248 , n113 );
nor ( n10040 , n117 , n118 );
and ( n10041 , n10039 , n3129 , n10040 );
nor ( n10042 , n10038 , n10041 );
nor ( n10043 , n10029 , n10042 );
not ( n10044 , n10043 );
and ( n10045 , n3104 , n3238 );
not ( n10046 , n10045 );
not ( n10047 , n10046 );
nand ( n10048 , n3127 , n116 );
nand ( n10049 , n3075 , n10048 );
not ( n10050 , n112 );
nand ( n10051 , n10050 , n3228 );
not ( n10052 , n10051 );
or ( n10053 , n10049 , n10052 );
nand ( n10054 , n115 , n117 );
not ( n10055 , n10054 );
nand ( n10056 , n10053 , n10055 );
not ( n10057 , n10056 );
or ( n10058 , n10047 , n10057 );
nand ( n10059 , n10058 , n3212 );
not ( n10060 , n10059 );
nand ( n10061 , n3144 , n3247 );
not ( n10062 , n116 );
nor ( n10063 , n10062 , n10054 );
not ( n10064 , n3025 );
not ( n10065 , n10064 );
nand ( n10066 , n10063 , n10065 );
and ( n10067 , n10061 , n10066 );
not ( n10068 , n10067 );
or ( n10069 , n10060 , n10068 );
nand ( n10070 , n10069 , n3106 );
not ( n10071 , n10070 );
or ( n10072 , n10044 , n10071 );
nor ( n10073 , n3105 , n116 );
not ( n10074 , n10073 );
nand ( n10075 , n3204 , n113 );
not ( n10076 , n10075 );
nand ( n10077 , n10076 , n3134 );
nor ( n10078 , n10048 , n115 );
nor ( n10079 , n10078 , n3106 );
nand ( n10080 , n10074 , n10077 , n10079 , n3049 );
nand ( n10081 , n10072 , n10080 );
not ( n10082 , n10081 );
or ( n10083 , n10028 , n10082 );
nand ( n10084 , n3160 , n115 );
not ( n10085 , n10084 );
not ( n10086 , n10085 );
and ( n10087 , n3054 , n117 );
nor ( n10088 , n10087 , n3212 );
not ( n10089 , n10088 );
and ( n10090 , n10086 , n10089 );
not ( n10091 , n10007 );
and ( n10092 , n3247 , n10091 );
nor ( n10093 , n10092 , n117 );
nand ( n10094 , n10030 , n3055 );
and ( n10095 , n10093 , n3135 , n10094 , n10048 );
nor ( n10096 , n10090 , n10095 );
not ( n10097 , n3081 );
not ( n10098 , n112 );
nand ( n10099 , n10098 , n116 );
nor ( n10100 , n10097 , n10099 );
nor ( n10101 , n10100 , n10035 );
and ( n10102 , n3160 , n3247 );
not ( n10103 , n10102 );
not ( n10104 , n3036 );
nand ( n10105 , n10101 , n10103 , n10104 , n3027 );
or ( n10106 , n10096 , n10105 );
not ( n10107 , n10040 );
not ( n10108 , n10020 );
or ( n10109 , n10107 , n10108 );
nand ( n10110 , n3251 , n3037 );
nand ( n10111 , n10110 , n3204 );
not ( n10112 , n10111 );
nand ( n10113 , n3204 , n116 );
not ( n10114 , n10113 );
or ( n10115 , n10112 , n10114 );
not ( n10116 , n10030 );
nand ( n10117 , n10115 , n10116 );
nand ( n10118 , n10117 , n10035 );
nand ( n10119 , n10109 , n10118 );
not ( n10120 , n3239 );
nand ( n10121 , n10120 , n3071 );
nand ( n10122 , n10119 , n10121 );
nand ( n10123 , n10106 , n10122 );
not ( n10124 , n3144 );
nor ( n10125 , n10124 , n115 );
not ( n10126 , n10125 );
nand ( n10127 , n10126 , n10094 );
and ( n10128 , n3051 , n3115 );
not ( n10129 , n3100 );
nor ( n10130 , n10128 , n10129 );
or ( n10131 , n10127 , n10130 );
nand ( n10132 , n10131 , n117 );
not ( n10133 , n3105 );
and ( n10134 , n10133 , n3094 );
nand ( n10135 , n3124 , n3137 );
nor ( n10136 , n10134 , n10135 );
not ( n10137 , n3102 );
and ( n10138 , n10132 , n10136 , n10137 );
nand ( n10139 , n10070 , n10123 , n10138 );
nand ( n10140 , n10083 , n10139 );
not ( n10141 , n10104 );
not ( n10142 , n3220 );
not ( n10143 , n10142 );
or ( n10144 , n10141 , n10143 );
not ( n10145 , n117 );
nand ( n10146 , n10144 , n10145 );
not ( n10147 , n3200 );
nand ( n10148 , n10147 , n115 );
not ( n10149 , n3161 );
not ( n10150 , n3234 );
and ( n10151 , n10149 , n10150 );
not ( n10152 , n10025 );
not ( n10153 , n10133 );
or ( n10154 , n10152 , n10153 );
not ( n10155 , n10124 );
not ( n10156 , n3146 );
nand ( n10157 , n10155 , n10156 , n118 );
nand ( n10158 , n10154 , n10157 );
nor ( n10159 , n10151 , n10158 );
nor ( n10160 , n3054 , n116 );
not ( n10161 , n10160 );
or ( n10162 , n10161 , n115 );
nand ( n10163 , n10162 , n3209 );
or ( n10164 , n10163 , n3175 );
nand ( n10165 , n10164 , n10040 );
and ( n10166 , n10146 , n10148 , n10159 , n10165 );
nand ( n10167 , n10140 , n10166 );
not ( n10168 , n10167 );
not ( n10169 , n10168 );
or ( n10170 , n9997 , n10169 );
nand ( n10171 , n10167 , n9995 );
nand ( n10172 , n10170 , n10171 );
not ( n10173 , n128 );
nand ( n10174 , n10173 , n130 );
not ( n10175 , n10174 );
nand ( n10176 , n10175 , n2415 );
and ( n10177 , n10176 , n133 );
buf ( n10178 , n2307 );
nand ( n10179 , n2357 , n2372 );
nand ( n10180 , n10178 , n10179 );
not ( n10181 , n10180 );
not ( n10182 , n2368 );
and ( n10183 , n10177 , n10181 , n10182 );
nor ( n10184 , n2490 , n2389 );
buf ( n10185 , n10184 );
not ( n10186 , n10185 );
not ( n10187 , n2486 );
not ( n10188 , n10187 );
not ( n10189 , n130 );
nor ( n10190 , n10189 , n2305 );
not ( n10191 , n10190 );
and ( n10192 , n10186 , n10188 , n10191 );
and ( n10193 , n10183 , n10192 );
and ( n10194 , n2369 , n2301 );
not ( n10195 , n10194 );
nand ( n10196 , n10195 , n2424 );
not ( n10197 , n2434 );
not ( n10198 , n2499 );
or ( n10199 , n10197 , n10198 );
nor ( n10200 , n129 , n130 );
nand ( n10201 , n10200 , n131 );
not ( n10202 , n10201 );
nand ( n10203 , n10202 , n2461 );
nand ( n10204 , n10199 , n10203 );
or ( n10205 , n10196 , n10185 , n10204 );
nand ( n10206 , n10205 , n2316 );
nor ( n10207 , n10193 , n10206 );
nand ( n10208 , n2357 , n2294 );
not ( n10209 , n2256 );
nand ( n10210 , n10209 , n2315 );
and ( n10211 , n10208 , n10210 , n2424 );
or ( n10212 , n10183 , n10211 );
buf ( n10213 , n2390 );
nand ( n10214 , n10213 , n2270 );
not ( n10215 , n10214 );
and ( n10216 , n2297 , n2469 );
nor ( n10217 , n10216 , n2282 );
not ( n10218 , n10217 );
or ( n10219 , n10215 , n10218 );
nand ( n10220 , n10219 , n2507 );
not ( n10221 , n131 );
not ( n10222 , n132 );
nor ( n10223 , n10222 , n2463 );
nand ( n10224 , n10221 , n10223 );
not ( n10225 , n10224 );
nand ( n10226 , n2255 , n2417 );
not ( n10227 , n10226 );
or ( n10228 , n10225 , n10227 );
nand ( n10229 , n10228 , n134 );
and ( n10230 , n2317 , n2327 , n2485 );
nor ( n10231 , n10230 , n2359 );
and ( n10232 , n10220 , n10229 , n10231 );
nand ( n10233 , n10212 , n10232 );
or ( n10234 , n10207 , n10233 );
not ( n10235 , n2284 );
not ( n10236 , n10235 );
not ( n10237 , n10200 );
not ( n10238 , n10237 );
nand ( n10239 , n10238 , n2270 );
not ( n10240 , n2463 );
nand ( n10241 , n10240 , n131 );
nand ( n10242 , n10239 , n10241 );
not ( n10243 , n10242 );
or ( n10244 , n10236 , n10243 );
nand ( n10245 , n10244 , n2410 );
nand ( n10246 , n10245 , n134 );
nand ( n10247 , n2333 , n2357 );
not ( n10248 , n10247 );
and ( n10249 , n10248 , n2424 );
buf ( n10250 , n2302 );
nor ( n10251 , n10250 , n2414 , n133 );
nand ( n10252 , n10251 , n2251 );
nor ( n10253 , n2356 , n133 );
buf ( n10254 , n2311 );
nand ( n10255 , n10253 , n10254 );
nand ( n10256 , n10252 , n10255 , n2359 );
nor ( n10257 , n10249 , n10256 );
not ( n10258 , n2321 );
nand ( n10259 , n2368 , n10258 );
not ( n10260 , n131 );
nand ( n10261 , n10260 , n2311 );
not ( n10262 , n10261 );
not ( n10263 , n2298 );
not ( n10264 , n10263 );
or ( n10265 , n10262 , n10264 );
nand ( n10266 , n10265 , n10235 );
nand ( n10267 , n10246 , n10257 , n10259 , n10266 );
nand ( n10268 , n10234 , n10267 );
not ( n10269 , n2359 );
not ( n10270 , n2293 );
not ( n10271 , n2326 );
or ( n10272 , n10270 , n10271 );
nand ( n10273 , n2489 , n2377 );
nand ( n10274 , n10272 , n10273 );
not ( n10275 , n10274 );
nand ( n10276 , n2356 , n2292 );
nand ( n10277 , n10276 , n2499 );
or ( n10278 , n10174 , n132 );
not ( n10279 , n10278 );
not ( n10280 , n2332 );
or ( n10281 , n10279 , n10280 );
nand ( n10282 , n10281 , n2270 );
nand ( n10283 , n10190 , n2424 );
nand ( n10284 , n10275 , n10277 , n10282 , n10283 );
not ( n10285 , n10284 );
or ( n10286 , n10269 , n10285 );
buf ( n10287 , n2342 );
not ( n10288 , n10287 );
nand ( n10289 , n10288 , n10213 );
not ( n10290 , n10289 );
nand ( n10291 , n2282 , n2485 );
not ( n10292 , n10291 );
or ( n10293 , n10290 , n10292 );
nand ( n10294 , n10293 , n2424 );
and ( n10295 , n2302 , n2270 );
not ( n10296 , n10295 );
not ( n10297 , n10296 );
nand ( n10298 , n10297 , n2377 );
nand ( n10299 , n10190 , n2324 );
and ( n10300 , n10298 , n10299 , n2471 );
not ( n10301 , n133 );
nor ( n10302 , n10301 , n131 );
not ( n10303 , n10302 );
or ( n10304 , n2380 , n10303 );
and ( n10305 , n10294 , n10300 , n10304 );
nand ( n10306 , n10286 , n10305 );
nand ( n10307 , n10306 , n2316 );
nor ( n10308 , n2382 , n128 );
nand ( n10309 , n10308 , n132 );
not ( n10310 , n10309 );
nand ( n10311 , n10310 , n10258 );
nand ( n10312 , n10185 , n2461 );
not ( n10313 , n10261 );
nor ( n10314 , n130 , n132 );
nand ( n10315 , n10313 , n10314 );
nand ( n10316 , n10311 , n10312 , n10315 );
not ( n10317 , n10224 );
not ( n10318 , n130 );
nand ( n10319 , n10318 , n2342 );
not ( n10320 , n10319 );
or ( n10321 , n10317 , n10320 );
nand ( n10322 , n10321 , n2324 );
not ( n10323 , n2310 );
not ( n10324 , n10323 );
nand ( n10325 , n10324 , n2403 );
nand ( n10326 , n10322 , n10325 );
nand ( n10327 , n10326 , n2507 );
nand ( n10328 , n2308 , n2485 , n133 );
nand ( n10329 , n10327 , n10328 );
nor ( n10330 , n10316 , n10329 );
nand ( n10331 , n10268 , n10307 , n10330 );
not ( n10332 , n10331 );
not ( n10333 , n10332 );
not ( n10334 , n215 );
and ( n10335 , n10333 , n10334 );
not ( n10336 , n10331 );
and ( n10337 , n10336 , n215 );
nor ( n10338 , n10335 , n10337 );
not ( n10339 , n10338 );
not ( n10340 , n3435 );
and ( n10341 , n10339 , n10340 );
and ( n10342 , n3435 , n10338 );
nor ( n10343 , n10341 , n10342 );
and ( n10344 , n10172 , n10343 );
not ( n10345 , n10172 );
not ( n10346 , n10343 );
and ( n10347 , n10345 , n10346 );
nor ( n10348 , n10344 , n10347 );
or ( n10349 , n10348 , n1 );
xnor ( n10350 , n215 , n216 );
or ( n10351 , n2246 , n10350 );
nand ( n10352 , n10349 , n10351 );
nand ( n10353 , n1476 , n1378 );
not ( n10354 , n1283 );
nand ( n10355 , n10354 , n1493 );
nand ( n10356 , n10353 , n10355 );
or ( n10357 , n10356 , n176 );
nand ( n10358 , n10357 , n177 );
and ( n10359 , n1289 , n1298 );
not ( n10360 , n10359 );
nand ( n10361 , n1347 , n173 );
not ( n10362 , n175 );
nor ( n10363 , n10362 , n1377 );
nand ( n10364 , n10363 , n1285 );
and ( n10365 , n10360 , n10361 , n10364 , n1469 );
nand ( n10366 , n10358 , n10365 );
not ( n10367 , n10366 );
not ( n10368 , n1336 );
not ( n10369 , n1284 );
nand ( n10370 , n1525 , n172 );
nand ( n10371 , n10368 , n10369 , n10370 , n176 );
not ( n10372 , n10371 );
or ( n10373 , n10367 , n10372 );
not ( n10374 , n1382 );
not ( n10375 , n10374 );
not ( n10376 , n174 );
nand ( n10377 , n10376 , n175 );
buf ( n10378 , n10377 );
nor ( n10379 , n10378 , n172 );
not ( n10380 , n10379 );
or ( n10381 , n10375 , n10380 );
nand ( n10382 , n10381 , n1469 );
nand ( n10383 , n1467 , n172 );
nand ( n10384 , n1484 , n173 );
nor ( n10385 , n10383 , n10384 );
or ( n10386 , n10382 , n10385 );
nand ( n10387 , n10386 , n1370 );
not ( n10388 , n10387 );
or ( n10389 , n176 , n177 );
not ( n10390 , n10389 );
not ( n10391 , n10390 );
not ( n10392 , n1397 );
nand ( n10393 , n10392 , n172 );
not ( n10394 , n10393 );
not ( n10395 , n10394 );
or ( n10396 , n10391 , n10395 );
nand ( n10397 , n10396 , n178 );
not ( n10398 , n171 );
not ( n10399 , n10398 );
not ( n10400 , n10377 );
not ( n10401 , n173 );
nor ( n10402 , n10401 , n172 );
nand ( n10403 , n10400 , n10402 );
not ( n10404 , n10403 );
not ( n10405 , n10404 );
or ( n10406 , n10399 , n10405 );
nand ( n10407 , n1512 , n1493 );
nor ( n10408 , n173 , n176 );
or ( n10409 , n10407 , n10408 );
nand ( n10410 , n10406 , n10409 );
nor ( n10411 , n10388 , n10397 , n10410 );
nand ( n10412 , n10373 , n10411 );
not ( n10413 , n10412 );
nor ( n10414 , n1402 , n175 );
and ( n10415 , n10414 , n173 );
nand ( n10416 , n1441 , n1315 );
nand ( n10417 , n10416 , n10390 );
or ( n10418 , n10415 , n10417 );
not ( n10419 , n1375 );
nand ( n10420 , n1526 , n10419 );
or ( n10421 , n10420 , n10359 );
nand ( n10422 , n10418 , n10421 );
not ( n10423 , n1296 );
nand ( n10424 , n10423 , n1524 );
and ( n10425 , n10424 , n1486 );
nand ( n10426 , n10422 , n10425 );
not ( n10427 , n10426 );
nand ( n10428 , n172 , n1289 );
nand ( n10429 , n10428 , n1529 );
not ( n10430 , n10429 );
nand ( n10431 , n173 , n177 );
nor ( n10432 , n10431 , n176 );
not ( n10433 , n10432 );
not ( n10434 , n1487 );
or ( n10435 , n10433 , n10434 );
nand ( n10436 , n1409 , n10408 , n177 );
nand ( n10437 , n10435 , n10436 );
not ( n10438 , n174 );
nand ( n10439 , n10438 , n1510 );
nand ( n10440 , n10437 , n10439 );
nor ( n10441 , n1531 , n172 );
nand ( n10442 , n10441 , n174 );
not ( n10443 , n1531 );
nand ( n10444 , n10443 , n173 );
nand ( n10445 , n10442 , n10444 , n1435 );
nand ( n10446 , n10440 , n10445 );
nand ( n10447 , n1328 , n1444 );
nand ( n10448 , n10430 , n10446 , n10447 );
not ( n10449 , n10448 );
or ( n10450 , n10427 , n10449 );
not ( n10451 , n1329 );
nor ( n10452 , n171 , n173 );
not ( n10453 , n10452 );
not ( n10454 , n10453 );
or ( n10455 , n10451 , n10454 );
nand ( n10456 , n10455 , n1306 );
not ( n10457 , n1448 );
not ( n10458 , n10457 );
and ( n10459 , n10456 , n10458 , n1350 );
nand ( n10460 , n1460 , n173 );
not ( n10461 , n1486 );
not ( n10462 , n173 );
nor ( n10463 , n10439 , n10462 );
nand ( n10464 , n10463 , n175 );
not ( n10465 , n10464 );
or ( n10466 , n10461 , n10465 );
nand ( n10467 , n10466 , n1280 );
and ( n10468 , n10459 , n10460 , n10467 );
nand ( n10469 , n10450 , n10468 );
not ( n10470 , n10469 );
or ( n10471 , n10413 , n10470 );
or ( n10472 , n10447 , n1417 );
and ( n10473 , n1398 , n1459 );
nand ( n10474 , n10473 , n173 );
nand ( n10475 , n10472 , n10474 );
nor ( n10476 , n1321 , n174 );
not ( n10477 , n175 );
nor ( n10478 , n10477 , n171 );
not ( n10479 , n10478 );
not ( n10480 , n10479 );
nand ( n10481 , n10476 , n10480 );
not ( n10482 , n10481 );
not ( n10483 , n1505 );
or ( n10484 , n10482 , n10483 );
nand ( n10485 , n10484 , n1370 );
not ( n10486 , n10444 );
not ( n10487 , n10379 );
or ( n10488 , n10486 , n10487 );
nand ( n10489 , n10488 , n10447 );
not ( n10490 , n1409 );
nand ( n10491 , n10490 , n10452 );
not ( n10492 , n1288 );
nor ( n10493 , n171 , n173 );
nand ( n10494 , n10492 , n10493 );
buf ( n10495 , n10494 );
nand ( n10496 , n10491 , n10495 );
or ( n10497 , n10489 , n10496 );
nand ( n10498 , n10497 , n1446 );
nand ( n10499 , n10485 , n10498 );
not ( n10500 , n1476 );
not ( n10501 , n10500 );
not ( n10502 , n10355 );
or ( n10503 , n10501 , n10502 );
nand ( n10504 , n10503 , n172 );
not ( n10505 , n10504 );
not ( n10506 , n1336 );
not ( n10507 , n10506 );
nand ( n10508 , n10507 , n1512 );
not ( n10509 , n10508 );
or ( n10510 , n10505 , n10509 );
nand ( n10511 , n10510 , n1435 );
not ( n10512 , n1512 );
not ( n10513 , n10490 );
or ( n10514 , n10512 , n10513 );
nand ( n10515 , n10514 , n10458 );
nand ( n10516 , n173 , n175 );
nor ( n10517 , n1484 , n10516 );
nand ( n10518 , n10517 , n1298 );
not ( n10519 , n10518 );
or ( n10520 , n10515 , n10519 );
nand ( n10521 , n10520 , n10419 );
nand ( n10522 , n10511 , n10521 );
nand ( n10523 , n10363 , n10462 );
nand ( n10524 , n1524 , n1357 );
and ( n10525 , n1414 , n10523 , n10524 );
nor ( n10526 , n10525 , n10389 );
nor ( n10527 , n10475 , n10499 , n10522 , n10526 );
nand ( n10528 , n10471 , n10527 );
not ( n10529 , n10528 );
nand ( n10530 , n1180 , n1120 );
not ( n10531 , n10530 );
not ( n10532 , n1016 );
nor ( n10533 , n10532 , n737 );
nand ( n10534 , n746 , n737 );
not ( n10535 , n165 );
nand ( n10536 , n10535 , n815 );
nand ( n10537 , n10534 , n10536 );
or ( n10538 , n10533 , n10537 );
nand ( n10539 , n10538 , n805 );
not ( n10540 , n1139 );
nor ( n10541 , n10540 , n779 );
nand ( n10542 , n10531 , n10539 , n10541 );
not ( n10543 , n10542 );
nand ( n10544 , n1062 , n892 );
not ( n10545 , n10544 );
nand ( n10546 , n836 , n165 );
not ( n10547 , n10546 );
or ( n10548 , n10545 , n10547 );
nand ( n10549 , n10548 , n920 );
not ( n10550 , n1258 );
and ( n10551 , n10550 , n950 , n779 );
nand ( n10552 , n10549 , n10551 );
not ( n10553 , n10552 );
or ( n10554 , n10543 , n10553 );
not ( n10555 , n1217 );
not ( n10556 , n753 );
or ( n10557 , n10555 , n10556 );
nand ( n10558 , n10557 , n1019 );
and ( n10559 , n10558 , n785 , n1050 );
nand ( n10560 , n10554 , n10559 );
not ( n10561 , n767 );
or ( n10562 , n793 , n166 );
not ( n10563 , n10562 );
or ( n10564 , n10561 , n10563 );
nand ( n10565 , n10564 , n779 );
nand ( n10566 , n1010 , n788 );
nand ( n10567 , n10566 , n167 );
not ( n10568 , n10567 );
not ( n10569 , n900 );
or ( n10570 , n863 , n10569 );
nand ( n10571 , n10570 , n169 );
and ( n10572 , n10565 , n10568 , n10571 );
and ( n10573 , n1259 , n843 );
nor ( n10574 , n10572 , n10573 );
or ( n10575 , n10560 , n10574 );
nand ( n10576 , n1013 , n920 );
not ( n10577 , n804 );
and ( n10578 , n10576 , n10577 );
not ( n10579 , n1040 );
nor ( n10580 , n10578 , n10579 );
not ( n10581 , n10580 );
not ( n10582 , n1007 );
not ( n10583 , n10562 );
or ( n10584 , n10582 , n10583 , n1265 );
nand ( n10585 , n10584 , n805 );
not ( n10586 , n10585 );
or ( n10587 , n10581 , n10586 );
nand ( n10588 , n10587 , n952 );
not ( n10589 , n169 );
nand ( n10590 , n861 , n957 );
not ( n10591 , n10590 );
or ( n10592 , n10589 , n10591 );
not ( n10593 , n847 );
not ( n10594 , n1219 );
or ( n10595 , n10593 , n10594 );
not ( n10596 , n909 );
nand ( n10597 , n831 , n10596 );
nand ( n10598 , n10595 , n10597 );
not ( n10599 , n933 );
not ( n10600 , n948 );
or ( n10601 , n10599 , n10600 );
nand ( n10602 , n10601 , n895 );
or ( n10603 , n10598 , n10602 );
nand ( n10604 , n10603 , n779 );
nand ( n10605 , n10592 , n10604 );
nand ( n10606 , n765 , n760 );
nand ( n10607 , n1134 , n10606 );
or ( n10608 , n10607 , n1016 );
not ( n10609 , n749 );
nand ( n10610 , n10608 , n10609 );
nand ( n10611 , n10610 , n170 );
nor ( n10612 , n10605 , n10611 );
nand ( n10613 , n10588 , n10612 );
nand ( n10614 , n10575 , n10613 );
not ( n10615 , n990 );
not ( n10616 , n1037 );
nor ( n10617 , n10616 , n807 );
not ( n10618 , n10617 );
or ( n10619 , n10615 , n10618 );
nand ( n10620 , n10619 , n945 );
nor ( n10621 , n738 , n1042 );
nand ( n10622 , n894 , n777 );
nand ( n10623 , n1139 , n10622 );
nor ( n10624 , n903 , n168 );
or ( n10625 , n10621 , n10623 , n10624 );
nand ( n10626 , n10625 , n756 );
nand ( n10627 , n10624 , n953 );
nand ( n10628 , n10620 , n10626 , n10627 );
not ( n10629 , n167 );
not ( n10630 , n914 );
or ( n10631 , n10629 , n10630 );
nand ( n10632 , n913 , n894 );
not ( n10633 , n10632 );
not ( n10634 , n830 );
or ( n10635 , n10633 , n10634 );
nand ( n10636 , n10635 , n1019 );
nand ( n10637 , n10631 , n10636 );
nand ( n10638 , n10566 , n817 );
or ( n10639 , n10637 , n10638 );
nand ( n10640 , n10639 , n779 );
not ( n10641 , n917 );
not ( n10642 , n776 );
and ( n10643 , n10641 , n10642 );
not ( n10644 , n165 );
nand ( n10645 , n10644 , n797 );
not ( n10646 , n10645 );
and ( n10647 , n10646 , n803 );
nor ( n10648 , n10643 , n10647 );
and ( n10649 , n1013 , n10648 );
nor ( n10650 , n10649 , n749 );
nor ( n10651 , n970 , n10650 );
nand ( n10652 , n10640 , n10651 );
nor ( n10653 , n10628 , n10652 );
nand ( n10654 , n10614 , n10653 );
not ( n10655 , n10654 );
not ( n10656 , n10655 );
or ( n10657 , n10529 , n10656 );
not ( n10658 , n10528 );
nand ( n10659 , n10654 , n10658 );
nand ( n10660 , n10657 , n10659 );
not ( n10661 , n10660 );
not ( n10662 , n779 );
nor ( n10663 , n10534 , n1036 );
or ( n10664 , n10663 , n167 );
nand ( n10665 , n10664 , n1166 );
nand ( n10666 , n782 , n801 );
nand ( n10667 , n1015 , n1042 );
nand ( n10668 , n10666 , n10667 , n10645 );
nor ( n10669 , n1060 , n10668 );
or ( n10670 , n10665 , n10669 );
nand ( n10671 , n790 , n737 );
and ( n10672 , n1227 , n10671 );
nand ( n10673 , n10670 , n10672 );
not ( n10674 , n10673 );
or ( n10675 , n10662 , n10674 );
nor ( n10676 , n10546 , n779 );
nand ( n10677 , n10562 , n170 );
nor ( n10678 , n1228 , n10676 , n10677 );
nand ( n10679 , n10675 , n10678 );
and ( n10680 , n843 , n1209 , n1037 );
and ( n10681 , n10680 , n10568 );
nor ( n10682 , n777 , n167 );
not ( n10683 , n10682 );
not ( n10684 , n753 );
or ( n10685 , n10683 , n10684 );
nand ( n10686 , n10685 , n946 );
not ( n10687 , n1217 );
not ( n10688 , n891 );
or ( n10689 , n10687 , n10688 );
nand ( n10690 , n10689 , n166 );
and ( n10691 , n10690 , n1075 , n1043 );
nand ( n10692 , n10686 , n10691 );
not ( n10693 , n10692 );
nor ( n10694 , n10681 , n10693 );
or ( n10695 , n10679 , n10694 );
and ( n10696 , n741 , n771 );
not ( n10697 , n917 );
not ( n10698 , n782 );
or ( n10699 , n10697 , n10698 );
nand ( n10700 , n10699 , n169 );
nor ( n10701 , n10696 , n10700 );
not ( n10702 , n10701 );
not ( n10703 , n1042 );
not ( n10704 , n10703 );
not ( n10705 , n1194 );
or ( n10706 , n10704 , n10705 );
nand ( n10707 , n10706 , n765 );
not ( n10708 , n10707 );
or ( n10709 , n10702 , n10708 );
not ( n10710 , n737 );
not ( n10711 , n1115 );
or ( n10712 , n10710 , n10711 );
nand ( n10713 , n10712 , n1173 );
nand ( n10714 , n10709 , n10713 );
nand ( n10715 , n843 , n10606 );
nor ( n10716 , n10536 , n166 );
or ( n10717 , n10715 , n10716 );
nand ( n10718 , n10717 , n805 );
nand ( n10719 , n1073 , n1127 );
and ( n10720 , n10719 , n953 );
or ( n10721 , n762 , n994 );
nand ( n10722 , n10721 , n1050 );
nor ( n10723 , n10720 , n10722 );
nand ( n10724 , n10714 , n10718 , n10723 );
nand ( n10725 , n10695 , n10724 );
nor ( n10726 , n738 , n1217 );
not ( n10727 , n737 );
not ( n10728 , n836 );
or ( n10729 , n10727 , n10728 );
nand ( n10730 , n10729 , n945 );
nor ( n10731 , n10726 , n1239 , n10730 );
nand ( n10732 , n1062 , n815 );
nand ( n10733 , n780 , n10732 );
nor ( n10734 , n10733 , n10567 );
or ( n10735 , n10731 , n10734 );
nand ( n10736 , n933 , n872 );
or ( n10737 , n10736 , n974 );
nand ( n10738 , n10735 , n10737 );
not ( n10739 , n10738 );
not ( n10740 , n1189 );
nand ( n10741 , n836 , n1140 );
not ( n10742 , n10741 );
or ( n10743 , n10740 , n10742 );
nand ( n10744 , n912 , n805 );
nand ( n10745 , n10743 , n10744 );
and ( n10746 , n1177 , n1158 , n169 );
nand ( n10747 , n10745 , n10746 );
not ( n10748 , n10747 );
or ( n10749 , n10739 , n10748 );
not ( n10750 , n802 );
not ( n10751 , n1018 );
or ( n10752 , n10750 , n10751 );
nand ( n10753 , n872 , n1042 );
and ( n10754 , n10622 , n10753 );
not ( n10755 , n10754 );
nand ( n10756 , n10752 , n10755 );
nand ( n10757 , n10749 , n10756 );
not ( n10758 , n10757 );
nand ( n10759 , n10725 , n10758 );
not ( n10760 , n10759 );
not ( n10761 , n10760 );
not ( n10762 , n1053 );
not ( n10763 , n1111 );
or ( n10764 , n10762 , n10763 );
nand ( n10765 , n10764 , n1149 );
not ( n10766 , n10765 );
and ( n10767 , n10761 , n10766 );
and ( n10768 , n1150 , n10760 );
nor ( n10769 , n10767 , n10768 );
not ( n10770 , n10769 );
not ( n10771 , n10770 );
or ( n10772 , n10661 , n10771 );
or ( n10773 , n10770 , n10660 );
nand ( n10774 , n10772 , n10773 );
not ( n10775 , n1841 );
nand ( n10776 , n1952 , n1971 );
not ( n10777 , n10776 );
or ( n10778 , n10775 , n10777 );
not ( n10779 , n2154 );
nand ( n10780 , n10778 , n10779 );
not ( n10781 , n2125 );
nand ( n10782 , n10781 , n2001 );
or ( n10783 , n10780 , n10782 );
not ( n10784 , n2187 );
nor ( n10785 , n1971 , n158 );
not ( n10786 , n10785 );
nand ( n10787 , n10784 , n10786 , n2006 );
nand ( n10788 , n10783 , n10787 );
not ( n10789 , n10788 );
and ( n10790 , n1834 , n1810 );
not ( n10791 , n10790 );
not ( n10792 , n1850 );
not ( n10793 , n10792 );
nand ( n10794 , n1834 , n10793 );
and ( n10795 , n10791 , n10794 );
not ( n10796 , n10795 );
or ( n10797 , n10789 , n10796 );
nor ( n10798 , n1868 , n1930 );
nand ( n10799 , n1952 , n10798 );
nand ( n10800 , n159 , n160 );
nand ( n10801 , n10799 , n10800 );
nand ( n10802 , n2137 , n1810 );
nand ( n10803 , n10801 , n10802 );
nand ( n10804 , n10797 , n10803 );
nor ( n10805 , n1855 , n154 );
not ( n10806 , n10805 );
nand ( n10807 , n10806 , n159 );
buf ( n10808 , n1820 );
not ( n10809 , n10808 );
not ( n10810 , n1834 );
or ( n10811 , n10809 , n10810 );
nand ( n10812 , n2073 , n1940 );
nand ( n10813 , n10811 , n10812 );
or ( n10814 , n10807 , n1826 , n10813 );
nor ( n10815 , n2063 , n1841 );
nor ( n10816 , n10815 , n159 );
not ( n10817 , n2029 );
not ( n10818 , n157 );
nand ( n10819 , n10817 , n10818 );
nand ( n10820 , n10816 , n2098 , n1941 , n10819 );
nand ( n10821 , n10814 , n10820 );
not ( n10822 , n2210 );
nand ( n10823 , n10822 , n1825 );
not ( n10824 , n10823 );
not ( n10825 , n2124 );
nor ( n10826 , n10825 , n158 );
nor ( n10827 , n10824 , n10826 , n1905 );
nand ( n10828 , n10804 , n10821 , n10827 );
not ( n10829 , n10828 );
not ( n10830 , n1947 );
nand ( n10831 , n10830 , n1979 );
not ( n10832 , n10831 );
nand ( n10833 , n10832 , n1841 );
nand ( n10834 , n1865 , n2190 );
nand ( n10835 , n1905 , n10834 , n1812 );
not ( n10836 , n10835 );
not ( n10837 , n1906 );
or ( n10838 , n10836 , n10837 );
nand ( n10839 , n1883 , n1921 , n1890 );
nand ( n10840 , n10838 , n10839 );
and ( n10841 , n1877 , n2001 );
nor ( n10842 , n10840 , n2133 , n10841 );
nand ( n10843 , n2009 , n154 );
nand ( n10844 , n1959 , n1897 );
nand ( n10845 , n1816 , n2052 );
and ( n10846 , n10843 , n10844 , n10845 );
not ( n10847 , n10846 );
or ( n10848 , n2192 , n2004 );
nand ( n10849 , n10848 , n1845 );
not ( n10850 , n10849 );
or ( n10851 , n10847 , n10850 );
nand ( n10852 , n2178 , n1841 );
nand ( n10853 , n10852 , n2215 , n1868 );
nand ( n10854 , n10851 , n10853 );
nand ( n10855 , n10833 , n10842 , n10854 );
not ( n10856 , n10855 );
or ( n10857 , n10829 , n10856 );
nor ( n10858 , n2179 , n1920 );
nand ( n10859 , n10858 , n10818 );
nand ( n10860 , n10859 , n2004 );
not ( n10861 , n10860 );
not ( n10862 , n2218 );
buf ( n10863 , n1971 );
nand ( n10864 , n10862 , n10863 );
not ( n10865 , n1931 );
not ( n10866 , n10865 );
not ( n10867 , n1910 );
nand ( n10868 , n1856 , n10867 );
not ( n10869 , n10868 );
or ( n10870 , n10866 , n10869 );
nand ( n10871 , n10870 , n159 );
nand ( n10872 , n10861 , n10864 , n10871 );
and ( n10873 , n2191 , n1835 );
nor ( n10874 , n10873 , n159 );
or ( n10875 , n10872 , n10874 );
not ( n10876 , n1956 );
nor ( n10877 , n2136 , n10876 );
not ( n10878 , n1986 );
or ( n10879 , n10877 , n10878 );
nand ( n10880 , n10879 , n1810 );
and ( n10881 , n1856 , n1921 );
nand ( n10882 , n10808 , n154 );
not ( n10883 , n159 );
nand ( n10884 , n10883 , n1841 );
or ( n10885 , n10882 , n10884 );
nand ( n10886 , n10885 , n160 );
nor ( n10887 , n10881 , n10886 );
not ( n10888 , n10819 );
nand ( n10889 , n10888 , n2046 );
nand ( n10890 , n10880 , n10887 , n10889 );
nand ( n10891 , n10875 , n10890 );
not ( n10892 , n10843 );
nand ( n10893 , n1831 , n1956 );
not ( n10894 , n10893 );
or ( n10895 , n10892 , n10894 );
nand ( n10896 , n10895 , n1858 );
and ( n10897 , n10891 , n10896 );
nand ( n10898 , n10857 , n10897 );
not ( n10899 , n10898 );
not ( n10900 , n2228 );
or ( n10901 , n10899 , n10900 );
not ( n10902 , n10855 );
not ( n10903 , n10828 );
or ( n10904 , n10902 , n10903 );
nand ( n10905 , n10904 , n10897 );
not ( n10906 , n10905 );
nand ( n10907 , n10906 , n2232 );
nand ( n10908 , n10901 , n10907 );
not ( n10909 , n10908 );
not ( n10910 , n1764 );
not ( n10911 , n1779 );
nand ( n10912 , n10911 , n148 );
not ( n10913 , n1662 );
not ( n10914 , n10913 );
nand ( n10915 , n1778 , n1631 );
not ( n10916 , n10915 );
or ( n10917 , n10914 , n10916 );
nand ( n10918 , n10917 , n150 );
and ( n10919 , n10912 , n10918 , n1699 );
nand ( n10920 , n1786 , n1603 );
nand ( n10921 , n10920 , n149 );
or ( n10922 , n10921 , n1702 );
not ( n10923 , n1660 );
nand ( n10924 , n10922 , n10923 );
not ( n10925 , n147 );
nor ( n10926 , n10925 , n151 );
not ( n10927 , n146 );
nand ( n10928 , n10926 , n10927 , n1793 );
nand ( n10929 , n1768 , n1662 );
and ( n10930 , n10924 , n10928 , n10929 , n1752 );
or ( n10931 , n10919 , n10930 );
not ( n10932 , n1783 );
nor ( n10933 , n1707 , n10932 );
nand ( n10934 , n10933 , n10927 );
nand ( n10935 , n10931 , n10934 );
nand ( n10936 , n1570 , n1603 );
and ( n10937 , n10928 , n10936 );
nor ( n10938 , n149 , n152 );
and ( n10939 , n1608 , n1654 , n10938 );
nand ( n10940 , n10937 , n10939 );
nand ( n10941 , n10935 , n10940 );
not ( n10942 , n10941 );
or ( n10943 , n10910 , n10942 );
not ( n10944 , n1729 );
nand ( n10945 , n10944 , n1620 );
nand ( n10946 , n10945 , n152 );
nand ( n10947 , n1683 , n1726 );
nand ( n10948 , n10947 , n1711 );
nor ( n10949 , n10946 , n10948 );
nand ( n10950 , n1682 , n1631 );
or ( n10951 , n10950 , n150 );
not ( n10952 , n1614 );
nand ( n10953 , n10949 , n10951 , n1771 , n10952 );
nand ( n10954 , n10943 , n10953 );
nor ( n10955 , n10915 , n150 );
not ( n10956 , n10938 );
nor ( n10957 , n10955 , n10956 );
not ( n10958 , n10957 );
not ( n10959 , n151 );
nand ( n10960 , n10959 , n146 , n148 , n1599 );
not ( n10961 , n10960 );
or ( n10962 , n10958 , n10961 );
nand ( n10963 , n1695 , n1615 );
not ( n10964 , n1621 );
nor ( n10965 , n10964 , n1560 );
nand ( n10966 , n10963 , n10965 );
nand ( n10967 , n10962 , n10966 );
not ( n10968 , n10967 );
nor ( n10969 , n1615 , n10960 );
nor ( n10970 , n10969 , n1776 );
not ( n10971 , n10970 );
or ( n10972 , n10968 , n10971 );
not ( n10973 , n149 );
nor ( n10974 , n1767 , n1725 );
not ( n10975 , n10974 );
or ( n10976 , n10973 , n10975 );
nand ( n10977 , n10976 , n1626 );
nor ( n10978 , n10977 , n10946 );
not ( n10979 , n1793 );
not ( n10980 , n1778 );
or ( n10981 , n10979 , n10980 );
buf ( n10982 , n1583 );
nand ( n10983 , n10982 , n1615 );
nand ( n10984 , n10981 , n10983 );
buf ( n10985 , n1613 );
not ( n10986 , n10985 );
or ( n10987 , n10984 , n10986 );
nand ( n10988 , n10987 , n1711 );
nand ( n10989 , n1723 , n1573 );
nand ( n10990 , n10978 , n10988 , n1760 , n10989 );
nand ( n10991 , n10972 , n10990 );
not ( n10992 , n10991 );
not ( n10993 , n1683 );
not ( n10994 , n10993 );
not ( n10995 , n1687 );
or ( n10996 , n10994 , n10995 );
not ( n10997 , n149 );
nor ( n10998 , n10997 , n150 );
buf ( n10999 , n10998 );
nand ( n11000 , n10996 , n10999 );
and ( n11001 , n11000 , n1788 , n1735 );
not ( n11002 , n1705 );
nand ( n11003 , n11002 , n1646 );
not ( n11004 , n11003 );
or ( n11005 , n11004 , n1776 );
nand ( n11006 , n11005 , n1711 );
nand ( n11007 , n11001 , n11006 );
and ( n11008 , n1642 , n1682 , n1660 , n148 );
nor ( n11009 , n11007 , n11008 );
not ( n11010 , n11009 );
or ( n11011 , n10992 , n11010 );
nand ( n11012 , n1774 , n1793 );
and ( n11013 , n11012 , n10915 );
not ( n11014 , n150 );
nor ( n11015 , n11014 , n1565 );
or ( n11016 , n1754 , n11015 );
nand ( n11017 , n11016 , n149 );
and ( n11018 , n11017 , n152 );
nand ( n11019 , n1778 , n1723 );
nand ( n11020 , n11013 , n11018 , n11019 );
nand ( n11021 , n1778 , n1683 );
nand ( n11022 , n10926 , n1793 );
and ( n11023 , n11021 , n11022 , n1752 );
not ( n11024 , n1748 );
not ( n11025 , n149 );
nand ( n11026 , n11025 , n150 );
not ( n11027 , n11026 );
or ( n11028 , n11024 , n11027 );
not ( n11029 , n1584 );
nand ( n11030 , n11028 , n11029 );
nand ( n11031 , n10951 , n11023 , n11030 );
and ( n11032 , n11020 , n11031 );
and ( n11033 , n10911 , n1656 );
nor ( n11034 , n11032 , n11033 );
nand ( n11035 , n10963 , n153 );
nand ( n11036 , n1590 , n148 );
nand ( n11037 , n1570 , n10927 );
buf ( n11038 , n11037 );
nand ( n11039 , n11036 , n11021 , n11038 );
or ( n11040 , n11035 , n11039 );
not ( n11041 , n1579 );
not ( n11042 , n150 );
nand ( n11043 , n11042 , n10944 );
nand ( n11044 , n11041 , n11043 );
nand ( n11045 , n11040 , n11044 );
nand ( n11046 , n11034 , n11045 );
nand ( n11047 , n11011 , n11046 );
nand ( n11048 , n10954 , n11047 );
not ( n11049 , n11048 );
not ( n11050 , n258 );
not ( n11051 , n11050 );
and ( n11052 , n11049 , n11051 );
buf ( n11053 , n11048 );
and ( n11054 , n11053 , n11050 );
nor ( n11055 , n11052 , n11054 );
not ( n11056 , n11055 );
or ( n11057 , n10909 , n11056 );
or ( n11058 , n11055 , n10908 );
nand ( n11059 , n11057 , n11058 );
not ( n11060 , n11059 );
and ( n11061 , n10774 , n11060 );
not ( n11062 , n10774 );
and ( n11063 , n11062 , n11059 );
nor ( n11064 , n11061 , n11063 );
or ( n11065 , n11064 , n1 );
and ( n11066 , n259 , n11050 );
not ( n11067 , n259 );
and ( n11068 , n11067 , n258 );
nor ( n11069 , n11066 , n11068 );
or ( n11070 , n2246 , n11069 );
nand ( n11071 , n11065 , n11070 );
not ( n11072 , n9474 );
not ( n11073 , n9575 );
not ( n11074 , n11073 );
or ( n11075 , n11072 , n11074 );
buf ( n11076 , n9474 );
not ( n11077 , n9575 );
or ( n11078 , n11076 , n11077 );
nand ( n11079 , n11075 , n11078 );
and ( n11080 , n11079 , n8406 );
not ( n11081 , n11079 );
not ( n11082 , n8406 );
and ( n11083 , n11081 , n11082 );
nor ( n11084 , n11080 , n11083 );
not ( n11085 , n7486 );
not ( n11086 , n75 );
and ( n11087 , n11085 , n11086 );
not ( n11088 , n7485 );
and ( n11089 , n11088 , n75 );
nor ( n11090 , n11087 , n11089 );
and ( n11091 , n8630 , n8894 );
not ( n11092 , n8630 );
and ( n11093 , n11092 , n8897 );
or ( n11094 , n11091 , n11093 );
and ( n11095 , n11090 , n11094 );
not ( n11096 , n11090 );
not ( n11097 , n11094 );
and ( n11098 , n11096 , n11097 );
nor ( n11099 , n11095 , n11098 );
not ( n11100 , n11099 );
and ( n11101 , n11084 , n11100 );
not ( n11102 , n11084 );
and ( n11103 , n11102 , n11099 );
nor ( n11104 , n11101 , n11103 );
or ( n11105 , n11104 , n1 );
xnor ( n11106 , n75 , n76 );
or ( n11107 , n2246 , n11106 );
nand ( n11108 , n11105 , n11107 );
not ( n11109 , n3957 );
not ( n11110 , n4954 );
and ( n11111 , n11109 , n11110 );
not ( n11112 , n11109 );
and ( n11113 , n11112 , n4954 );
nor ( n11114 , n11111 , n11113 );
not ( n11115 , n11114 );
not ( n11116 , n11115 );
not ( n11117 , n6019 );
or ( n11118 , n11116 , n11117 );
nand ( n11119 , n6022 , n11114 );
nand ( n11120 , n11118 , n11119 );
not ( n11121 , n104 );
not ( n11122 , n4650 );
or ( n11123 , n11121 , n11122 );
not ( n11124 , n4648 );
not ( n11125 , n104 );
nand ( n11126 , n11124 , n11125 );
nand ( n11127 , n11123 , n11126 );
and ( n11128 , n11127 , n6274 );
not ( n11129 , n11127 );
not ( n11130 , n6274 );
and ( n11131 , n11129 , n11130 );
nor ( n11132 , n11128 , n11131 );
and ( n11133 , n11120 , n11132 );
not ( n11134 , n11120 );
not ( n11135 , n11132 );
and ( n11136 , n11134 , n11135 );
nor ( n11137 , n11133 , n11136 );
or ( n11138 , n11137 , n1 );
and ( n11139 , n267 , n11125 );
not ( n11140 , n267 );
and ( n11141 , n11140 , n104 );
nor ( n11142 , n11139 , n11141 );
or ( n11143 , n2246 , n11142 );
nand ( n11144 , n11138 , n11143 );
not ( n11145 , n322 );
not ( n11146 , n4648 );
or ( n11147 , n11145 , n11146 );
not ( n11148 , n322 );
nand ( n11149 , n4649 , n11148 );
nand ( n11150 , n11147 , n11149 );
not ( n11151 , n6017 );
not ( n11152 , n4830 );
not ( n11153 , n11152 );
or ( n11154 , n11151 , n11153 );
nand ( n11155 , n4830 , n6012 );
nand ( n11156 , n11154 , n11155 );
not ( n11157 , n11156 );
and ( n11158 , n11150 , n11157 );
not ( n11159 , n11150 );
and ( n11160 , n11159 , n11156 );
nor ( n11161 , n11158 , n11160 );
not ( n11162 , n4367 );
not ( n11163 , n3709 );
and ( n11164 , n11162 , n11163 );
buf ( n11165 , n5395 );
and ( n11166 , n11165 , n3709 );
nor ( n11167 , n11164 , n11166 );
not ( n11168 , n11167 );
not ( n11169 , n5895 );
or ( n11170 , n11168 , n11169 );
or ( n11171 , n5895 , n11167 );
nand ( n11172 , n11170 , n11171 );
and ( n11173 , n11161 , n11172 );
not ( n11174 , n11161 );
not ( n11175 , n11172 );
and ( n11176 , n11174 , n11175 );
nor ( n11177 , n11173 , n11176 );
or ( n11178 , n11177 , n1 );
and ( n11179 , n323 , n11148 );
not ( n11180 , n323 );
and ( n11181 , n11180 , n322 );
nor ( n11182 , n11179 , n11181 );
or ( n11183 , n2246 , n11182 );
nand ( n11184 , n11178 , n11183 );
not ( n11185 , n99 );
not ( n11186 , n11185 );
not ( n11187 , n6271 );
and ( n11188 , n5611 , n4413 );
nand ( n11189 , n6035 , n5520 );
nor ( n11190 , n11188 , n11189 );
not ( n11191 , n11190 );
not ( n11192 , n4548 );
nand ( n11193 , n11192 , n4393 );
not ( n11194 , n4467 );
nand ( n11195 , n11194 , n4437 , n190 );
and ( n11196 , n11193 , n11195 , n4576 );
not ( n11197 , n11196 );
or ( n11198 , n11191 , n11197 );
not ( n11199 , n4514 );
not ( n11200 , n4547 );
or ( n11201 , n11199 , n11200 );
nand ( n11202 , n5494 , n4631 );
nand ( n11203 , n11201 , n11202 );
nand ( n11204 , n11203 , n193 );
and ( n11205 , n4564 , n4590 , n194 );
not ( n11206 , n4569 );
nand ( n11207 , n11206 , n4529 );
nand ( n11208 , n11204 , n11205 , n11207 , n4504 );
nand ( n11209 , n11198 , n11208 );
not ( n11210 , n11209 );
nand ( n11211 , n4428 , n4615 );
and ( n11212 , n4390 , n11211 );
nor ( n11213 , n6197 , n190 );
or ( n11214 , n11213 , n4410 );
nand ( n11215 , n11214 , n193 );
and ( n11216 , n4534 , n4393 );
nor ( n11217 , n11216 , n195 );
nand ( n11218 , n11215 , n11217 );
nor ( n11219 , n11212 , n11218 );
not ( n11220 , n11219 );
or ( n11221 , n11210 , n11220 );
nor ( n11222 , n6082 , n4383 );
not ( n11223 , n11222 );
not ( n11224 , n6160 );
or ( n11225 , n11223 , n11224 );
not ( n11226 , n5502 );
and ( n11227 , n4569 , n6140 );
nand ( n11228 , n11226 , n11227 , n4598 , n4539 );
nand ( n11229 , n11225 , n11228 );
not ( n11230 , n5586 );
nor ( n11231 , n11230 , n5611 );
nand ( n11232 , n11229 , n11231 );
not ( n11233 , n11232 );
nand ( n11234 , n4433 , n6043 );
or ( n11235 , n5580 , n11234 );
or ( n11236 , n4641 , n193 );
nand ( n11237 , n11235 , n11236 );
not ( n11238 , n4628 );
nand ( n11239 , n6174 , n4604 );
nor ( n11240 , n11238 , n5531 , n11239 , n4617 );
nand ( n11241 , n11237 , n11240 );
not ( n11242 , n11241 );
or ( n11243 , n11233 , n11242 );
not ( n11244 , n6209 );
not ( n11245 , n11193 );
or ( n11246 , n11244 , n11245 );
nand ( n11247 , n11246 , n4390 );
not ( n11248 , n6257 );
nand ( n11249 , n6166 , n195 );
nor ( n11250 , n11248 , n11249 );
not ( n11251 , n6108 );
not ( n11252 , n11251 );
and ( n11253 , n190 , n193 );
not ( n11254 , n11253 );
or ( n11255 , n11252 , n11254 );
nand ( n11256 , n4423 , n4430 );
not ( n11257 , n11256 );
not ( n11258 , n4573 );
or ( n11259 , n11257 , n11258 );
nand ( n11260 , n11259 , n4494 );
nand ( n11261 , n11255 , n11260 );
not ( n11262 , n11261 );
and ( n11263 , n11247 , n11250 , n11262 );
nand ( n11264 , n11243 , n11263 );
nand ( n11265 , n11221 , n11264 );
not ( n11266 , n4452 );
nand ( n11267 , n11266 , n4633 );
and ( n11268 , n11267 , n4431 , n4592 );
not ( n11269 , n6167 );
not ( n11270 , n4545 );
or ( n11271 , n11269 , n11270 );
nand ( n11272 , n11271 , n6242 );
nand ( n11273 , n5612 , n11272 );
not ( n11274 , n6214 );
nand ( n11275 , n4462 , n4404 );
nand ( n11276 , n6108 , n11275 , n5594 );
nand ( n11277 , n11274 , n11276 );
not ( n11278 , n5497 );
nand ( n11279 , n11278 , n4413 );
nand ( n11280 , n11277 , n11279 );
or ( n11281 , n11273 , n11280 );
nand ( n11282 , n11281 , n194 );
nor ( n11283 , n4412 , n4541 , n194 );
or ( n11284 , n4456 , n11283 );
nand ( n11285 , n11284 , n4547 );
nand ( n11286 , n4621 , n4534 );
and ( n11287 , n11268 , n11282 , n11285 , n11286 );
nand ( n11288 , n11265 , n11287 );
not ( n11289 , n11288 );
not ( n11290 , n11289 );
or ( n11291 , n11187 , n11290 );
nand ( n11292 , n11288 , n6154 );
nand ( n11293 , n11291 , n11292 );
not ( n11294 , n11293 );
not ( n11295 , n11294 );
or ( n11296 , n11186 , n11295 );
nand ( n11297 , n11293 , n99 );
nand ( n11298 , n11296 , n11297 );
nand ( n11299 , n5636 , n2246 );
and ( n11300 , n269 , n99 );
not ( n11301 , n269 );
and ( n11302 , n11301 , n11185 );
nor ( n11303 , n11300 , n11302 );
nand ( n11304 , n11303 , n1 );
and ( n11305 , n11299 , n11304 );
and ( n11306 , n11298 , n11305 );
not ( n11307 , n11298 );
not ( n11308 , n11304 );
nor ( n11309 , n5636 , n1 );
nor ( n11310 , n11308 , n11309 );
and ( n11311 , n11307 , n11310 );
or ( n11312 , n11306 , n11311 );
not ( n11313 , n5245 );
nand ( n11314 , n4215 , n3525 );
not ( n11315 , n11314 );
and ( n11316 , n5262 , n4303 , n209 );
nand ( n11317 , n11315 , n11316 );
not ( n11318 , n3650 );
or ( n11319 , n11317 , n11318 , n9642 );
not ( n11320 , n205 );
not ( n11321 , n3678 );
or ( n11322 , n11320 , n11321 );
nand ( n11323 , n11322 , n5323 );
nor ( n11324 , n5928 , n11323 );
not ( n11325 , n5937 );
not ( n11326 , n4258 );
or ( n11327 , n11324 , n11325 , n11326 );
nand ( n11328 , n11319 , n11327 );
nand ( n11329 , n9642 , n3462 );
and ( n11330 , n11329 , n4217 );
nand ( n11331 , n11328 , n11330 );
not ( n11332 , n9623 );
not ( n11333 , n3511 );
nor ( n11334 , n11332 , n4309 , n4293 , n11333 );
not ( n11335 , n3693 );
nand ( n11336 , n3689 , n3678 );
and ( n11337 , n5329 , n11336 );
not ( n11338 , n11337 );
or ( n11339 , n11335 , n11338 );
nand ( n11340 , n11339 , n3485 );
nand ( n11341 , n11334 , n11340 );
nand ( n11342 , n11331 , n11341 );
and ( n11343 , n4336 , n3602 );
nor ( n11344 , n11343 , n212 );
and ( n11345 , n11329 , n11344 );
not ( n11346 , n11345 );
not ( n11347 , n9694 );
not ( n11348 , n3619 );
not ( n11349 , n5901 );
or ( n11350 , n11348 , n11349 );
not ( n11351 , n209 );
not ( n11352 , n3622 );
not ( n11353 , n3642 );
or ( n11354 , n11352 , n11353 );
nand ( n11355 , n11354 , n209 );
not ( n11356 , n11355 );
or ( n11357 , n11351 , n11356 );
nand ( n11358 , n11357 , n3629 );
not ( n11359 , n4333 );
nor ( n11360 , n4254 , n11359 );
nand ( n11361 , n11358 , n11360 );
nand ( n11362 , n11350 , n11361 );
not ( n11363 , n11362 );
or ( n11364 , n11347 , n11363 );
not ( n11365 , n3697 );
not ( n11366 , n4255 );
not ( n11367 , n11366 );
or ( n11368 , n11365 , n11367 );
nand ( n11369 , n11368 , n211 );
not ( n11370 , n3599 );
and ( n11371 , n3587 , n11370 );
nor ( n11372 , n11371 , n3597 );
nor ( n11373 , n11369 , n11372 );
not ( n11374 , n210 );
not ( n11375 , n3519 );
or ( n11376 , n11374 , n11375 );
not ( n11377 , n11355 );
nand ( n11378 , n11376 , n11377 );
and ( n11379 , n4241 , n3506 );
or ( n11380 , n11379 , n3470 );
nand ( n11381 , n11380 , n3485 );
nand ( n11382 , n11373 , n11378 , n11381 );
nand ( n11383 , n11364 , n11382 );
not ( n11384 , n11383 );
or ( n11385 , n11346 , n11384 );
and ( n11386 , n4263 , n207 );
nor ( n11387 , n4318 , n3593 );
nor ( n11388 , n11386 , n11387 , n3461 );
nand ( n11389 , n11388 , n3626 , n5348 );
not ( n11390 , n11389 );
not ( n11391 , n5912 );
nand ( n11392 , n11391 , n209 );
nor ( n11393 , n3699 , n3525 );
or ( n11394 , n5387 , n5356 );
nand ( n11395 , n11394 , n4304 );
nand ( n11396 , n5368 , n11392 , n11393 , n11395 );
not ( n11397 , n11396 );
or ( n11398 , n11390 , n11397 );
and ( n11399 , n5278 , n5947 );
and ( n11400 , n3693 , n11399 );
nor ( n11401 , n11400 , n209 );
not ( n11402 , n3506 );
not ( n11403 , n205 );
and ( n11404 , n11402 , n11403 );
and ( n11405 , n3564 , n5972 );
nor ( n11406 , n11404 , n11405 );
and ( n11407 , n3679 , n11406 , n3611 );
or ( n11408 , n11407 , n3485 );
nand ( n11409 , n11408 , n212 );
nor ( n11410 , n11401 , n11409 );
nand ( n11411 , n11398 , n11410 );
nand ( n11412 , n11385 , n11411 );
and ( n11413 , n5363 , n3503 );
and ( n11414 , n11359 , n3630 );
nor ( n11415 , n11413 , n11414 );
and ( n11416 , n11342 , n11412 , n11415 );
not ( n11417 , n11416 );
or ( n11418 , n11313 , n11417 );
not ( n11419 , n11416 );
nand ( n11420 , n11419 , n5244 );
nand ( n11421 , n11418 , n11420 );
not ( n11422 , n11421 );
buf ( n11423 , n11422 );
not ( n11424 , n5645 );
not ( n11425 , n5087 );
or ( n11426 , n11424 , n11425 );
not ( n11427 , n11110 );
nand ( n11428 , n5248 , n11427 );
nand ( n11429 , n11426 , n11428 );
not ( n11430 , n11429 );
not ( n11431 , n11304 );
or ( n11432 , n11423 , n11430 , n11431 );
nand ( n11433 , n11423 , n11430 , n11304 );
nand ( n11434 , n11432 , n11433 );
or ( n11435 , n11312 , n11434 );
not ( n11436 , n11309 );
not ( n11437 , n11298 );
or ( n11438 , n11436 , n11437 );
or ( n11439 , n11299 , n11298 );
nand ( n11440 , n11438 , n11439 );
not ( n11441 , n11423 );
and ( n11442 , n11430 , n11441 );
not ( n11443 , n11430 );
and ( n11444 , n11443 , n11423 );
nor ( n11445 , n11442 , n11444 );
nand ( n11446 , n11440 , n11445 );
nand ( n11447 , n11435 , n11446 );
not ( n11448 , n10936 );
not ( n11449 , n1728 );
or ( n11450 , n11448 , n11449 );
nand ( n11451 , n11450 , n1752 );
and ( n11452 , n1631 , n10938 );
nor ( n11453 , n11452 , n153 );
nand ( n11454 , n11451 , n11453 );
not ( n11455 , n11454 );
not ( n11456 , n1752 );
not ( n11457 , n1670 );
or ( n11458 , n11456 , n11457 );
nand ( n11459 , n1774 , n148 );
nand ( n11460 , n11458 , n11459 );
not ( n11461 , n11036 );
or ( n11462 , n11460 , n11461 , n1614 );
nand ( n11463 , n11462 , n1660 );
nor ( n11464 , n1687 , n1603 );
not ( n11465 , n10974 );
not ( n11466 , n147 );
nor ( n11467 , n11466 , n151 );
nand ( n11468 , n11467 , n1787 );
nand ( n11469 , n11465 , n11468 );
nor ( n11470 , n11464 , n11469 );
not ( n11471 , n11470 );
not ( n11472 , n1794 );
or ( n11473 , n11471 , n11472 );
nand ( n11474 , n11473 , n1617 );
not ( n11475 , n1556 );
not ( n11476 , n1654 );
or ( n11477 , n11475 , n11476 );
nand ( n11478 , n11477 , n1617 );
nand ( n11479 , n1768 , n148 );
not ( n11480 , n11479 );
nand ( n11481 , n10998 , n148 );
not ( n11482 , n11481 );
or ( n11483 , n11480 , n11482 );
nand ( n11484 , n11483 , n1778 );
nand ( n11485 , n11478 , n11038 , n11484 );
nand ( n11486 , n11485 , n152 );
nand ( n11487 , n11455 , n11463 , n11474 , n11486 );
not ( n11488 , n11043 );
not ( n11489 , n148 );
nand ( n11490 , n11489 , n146 );
nand ( n11491 , n11490 , n1597 );
nor ( n11492 , n11488 , n11491 );
or ( n11493 , n11492 , n1617 );
not ( n11494 , n1701 );
not ( n11495 , n1714 );
or ( n11496 , n11494 , n11495 );
nand ( n11497 , n11496 , n1721 );
nand ( n11498 , n11493 , n11497 );
or ( n11499 , n1676 , n1750 );
nand ( n11500 , n1625 , n1660 );
nand ( n11501 , n11499 , n11500 , n152 );
or ( n11502 , n11498 , n11501 );
and ( n11503 , n1754 , n1615 );
or ( n11504 , n11503 , n1560 );
not ( n11505 , n1630 );
nand ( n11506 , n1701 , n1725 );
not ( n11507 , n11506 );
or ( n11508 , n11505 , n11507 );
nand ( n11509 , n1783 , n148 );
and ( n11510 , n11509 , n10938 );
nand ( n11511 , n11508 , n11510 );
nand ( n11512 , n11504 , n11511 );
not ( n11513 , n1722 );
and ( n11514 , n11513 , n1743 , n1761 );
nand ( n11515 , n11512 , n11514 );
nand ( n11516 , n11502 , n11515 );
not ( n11517 , n1767 );
not ( n11518 , n11490 );
and ( n11519 , n11517 , n11518 );
nor ( n11520 , n11519 , n1735 );
nand ( n11521 , n1564 , n1778 );
nand ( n11522 , n1682 , n1646 );
and ( n11523 , n11520 , n11521 , n11522 );
not ( n11524 , n11523 );
nand ( n11525 , n1695 , n148 );
not ( n11526 , n11525 );
or ( n11527 , n11524 , n11526 );
nor ( n11528 , n1735 , n149 );
not ( n11529 , n11528 );
nand ( n11530 , n11527 , n11529 );
nand ( n11531 , n1646 , n10926 );
nand ( n11532 , n11516 , n11530 , n11531 );
and ( n11533 , n11487 , n11532 );
nand ( n11534 , n11021 , n1634 );
and ( n11535 , n1682 , n1630 );
nor ( n11536 , n11534 , n11535 );
or ( n11537 , n11536 , n11026 );
not ( n11538 , n151 );
not ( n11539 , n11491 );
or ( n11540 , n11538 , n11539 );
nand ( n11541 , n11540 , n1684 );
nand ( n11542 , n11541 , n10999 );
nand ( n11543 , n11537 , n11542 );
nand ( n11544 , n11543 , n152 );
not ( n11545 , n1615 );
not ( n11546 , n1662 );
or ( n11547 , n11545 , n11546 );
nand ( n11548 , n11547 , n10945 );
or ( n11549 , n1751 , n11548 );
not ( n11550 , n1560 );
nand ( n11551 , n11549 , n11550 );
nand ( n11552 , n1762 , n1783 );
not ( n11553 , n11552 );
nand ( n11554 , n1787 , n1633 );
not ( n11555 , n11554 );
nand ( n11556 , n11555 , n1642 );
not ( n11557 , n11556 );
or ( n11558 , n11553 , n11557 );
nand ( n11559 , n11558 , n1617 );
nand ( n11560 , n11469 , n10938 );
and ( n11561 , n11551 , n11559 , n11560 );
not ( n11562 , n10915 );
not ( n11563 , n11562 );
not ( n11564 , n11563 );
not ( n11565 , n1760 );
or ( n11566 , n11564 , n11565 );
nand ( n11567 , n11566 , n1699 );
not ( n11568 , n1754 );
or ( n11569 , n11568 , n11026 );
and ( n11570 , n1644 , n1572 );
buf ( n11571 , n11570 );
not ( n11572 , n11571 );
nand ( n11573 , n11569 , n11572 );
nand ( n11574 , n11573 , n1752 );
nand ( n11575 , n11544 , n11561 , n11567 , n11574 );
nor ( n11576 , n11533 , n11575 );
buf ( n11577 , n11576 );
not ( n11578 , n11577 );
nor ( n11579 , n147 , n150 );
nand ( n11580 , n1594 , n11579 );
nor ( n11581 , n1789 , n10956 );
and ( n11582 , n11580 , n11581 , n1743 );
and ( n11583 , n11506 , n1787 );
nor ( n11584 , n11583 , n1560 );
or ( n11585 , n11582 , n11584 );
not ( n11586 , n11026 );
nand ( n11587 , n11586 , n10926 );
nor ( n11588 , n11587 , n11490 );
not ( n11589 , n11588 );
nand ( n11590 , n11585 , n11589 );
or ( n11591 , n11590 , n11008 );
nand ( n11592 , n10982 , n1620 );
not ( n11593 , n11592 );
not ( n11594 , n1785 );
or ( n11595 , n11593 , n11594 );
nand ( n11596 , n11595 , n149 );
nand ( n11597 , n11571 , n1711 );
nand ( n11598 , n11596 , n1592 , n1616 , n11597 );
nand ( n11599 , n11591 , n11598 );
not ( n11600 , n151 );
nor ( n11601 , n11600 , n1748 );
and ( n11602 , n11601 , n1617 , n146 );
and ( n11603 , n1787 , n149 );
and ( n11604 , n1695 , n11603 );
nor ( n11605 , n11602 , n11604 );
nand ( n11606 , n11599 , n11605 );
not ( n11607 , n11606 );
not ( n11608 , n11531 );
not ( n11609 , n11459 );
or ( n11610 , n11608 , n11609 );
nand ( n11611 , n11610 , n1617 );
not ( n11612 , n10993 );
not ( n11613 , n1676 );
or ( n11614 , n11612 , n11613 );
nand ( n11615 , n11614 , n11586 );
nand ( n11616 , n11611 , n11615 , n1755 );
not ( n11617 , n1703 );
nor ( n11618 , n11617 , n11004 );
and ( n11619 , n10937 , n11618 );
nor ( n11620 , n11619 , n1711 );
nor ( n11621 , n11616 , n11035 , n11620 );
not ( n11622 , n11621 );
not ( n11623 , n11043 );
nand ( n11624 , n11623 , n1599 );
nand ( n11625 , n11525 , n11624 , n1671 );
not ( n11626 , n11625 );
not ( n11627 , n149 );
or ( n11628 , n11626 , n11627 );
nand ( n11629 , n1702 , n148 );
not ( n11630 , n11629 );
not ( n11631 , n1721 );
not ( n11632 , n11631 );
and ( n11633 , n11630 , n11632 );
nand ( n11634 , n11468 , n1752 );
not ( n11635 , n11634 );
not ( n11636 , n147 );
not ( n11637 , n1584 );
or ( n11638 , n11636 , n11637 );
nand ( n11639 , n11638 , n1564 );
nand ( n11640 , n11635 , n11639 );
nor ( n11641 , n11633 , n11640 );
nand ( n11642 , n11628 , n11641 );
nor ( n11643 , n1600 , n1752 , n1726 );
or ( n11644 , n11643 , n1699 );
nand ( n11645 , n11644 , n10960 );
nand ( n11646 , n11642 , n11645 );
not ( n11647 , n11646 );
or ( n11648 , n11622 , n11647 );
not ( n11649 , n1660 );
not ( n11650 , n1695 );
or ( n11651 , n11649 , n11650 );
or ( n11652 , n11601 , n1730 );
nand ( n11653 , n11652 , n1556 );
nand ( n11654 , n1763 , n1721 );
and ( n11655 , n11653 , n11654 , n152 );
nand ( n11656 , n11651 , n11655 );
not ( n11657 , n1615 );
not ( n11658 , n11534 );
or ( n11659 , n11657 , n11658 );
nand ( n11660 , n11659 , n1561 );
nand ( n11661 , n11656 , n11660 );
not ( n11662 , n1573 );
or ( n11663 , n11662 , n150 );
not ( n11664 , n1706 );
nand ( n11665 , n11663 , n11664 );
and ( n11666 , n11665 , n11550 );
not ( n11667 , n1590 );
and ( n11668 , n1676 , n11667 );
nand ( n11669 , n1564 , n149 );
nor ( n11670 , n11668 , n11669 );
nor ( n11671 , n11666 , n11670 , n153 );
and ( n11672 , n10985 , n1615 );
not ( n11673 , n1774 );
and ( n11674 , n11673 , n150 );
nor ( n11675 , n11672 , n11674 );
or ( n11676 , n11004 , n11675 );
nand ( n11677 , n11676 , n1711 );
nand ( n11678 , n11661 , n11671 , n11677 );
nand ( n11679 , n11648 , n11678 );
nand ( n11680 , n11607 , n11679 );
not ( n11681 , n11680 );
not ( n11682 , n11681 );
or ( n11683 , n11578 , n11682 );
or ( n11684 , n11681 , n11577 );
nand ( n11685 , n11683 , n11684 );
not ( n11686 , n11685 );
not ( n11687 , n10660 );
not ( n11688 , n11687 );
or ( n11689 , n11686 , n11688 );
not ( n11690 , n11685 );
nand ( n11691 , n11690 , n10660 );
nand ( n11692 , n11689 , n11691 );
not ( n11693 , n10908 );
not ( n11694 , n1989 );
nor ( n11695 , n1976 , n10813 , n2005 );
not ( n11696 , n11695 );
not ( n11697 , n1993 );
or ( n11698 , n11696 , n11697 );
not ( n11699 , n1984 );
not ( n11700 , n1855 );
or ( n11701 , n11699 , n11700 );
nand ( n11702 , n11701 , n1841 );
nand ( n11703 , n1902 , n11702 , n10812 , n159 );
nand ( n11704 , n11698 , n11703 );
not ( n11705 , n11704 );
or ( n11706 , n11694 , n11705 );
nand ( n11707 , n2103 , n160 );
not ( n11708 , n11707 );
not ( n11709 , n154 );
nand ( n11710 , n11709 , n2046 );
nand ( n11711 , n10844 , n11710 );
not ( n11712 , n11711 );
and ( n11713 , n2176 , n154 );
nor ( n11714 , n2032 , n11713 );
not ( n11715 , n11714 );
or ( n11716 , n11712 , n11715 );
and ( n11717 , n2124 , n1890 );
not ( n11718 , n11717 );
nand ( n11719 , n11716 , n11718 );
not ( n11720 , n11719 );
and ( n11721 , n11708 , n11720 );
not ( n11722 , n10800 );
nor ( n11723 , n11721 , n11722 );
nand ( n11724 , n11706 , n11723 );
not ( n11725 , n2108 );
not ( n11726 , n1862 );
and ( n11727 , n2066 , n2029 );
not ( n11728 , n11727 );
not ( n11729 , n11728 );
or ( n11730 , n11726 , n11729 );
nand ( n11731 , n11730 , n2118 );
not ( n11732 , n11731 );
not ( n11733 , n11722 );
or ( n11734 , n11732 , n11733 );
nand ( n11735 , n11734 , n2021 );
nor ( n11736 , n11725 , n11735 );
and ( n11737 , n11724 , n11736 );
and ( n11738 , n10882 , n159 );
not ( n11739 , n11738 );
not ( n11740 , n1874 );
or ( n11741 , n11739 , n11740 );
not ( n11742 , n155 );
not ( n11743 , n2067 );
or ( n11744 , n11742 , n11743 );
nand ( n11745 , n11744 , n2043 );
nand ( n11746 , n1810 , n2167 );
or ( n11747 , n11745 , n11746 );
not ( n11748 , n1841 );
not ( n11749 , n10793 );
or ( n11750 , n11748 , n11749 );
nand ( n11751 , n11750 , n1979 );
not ( n11752 , n11751 );
nand ( n11753 , n11747 , n11752 );
nand ( n11754 , n11741 , n11753 );
not ( n11755 , n10819 );
nand ( n11756 , n11755 , n155 );
nand ( n11757 , n11756 , n2193 );
nor ( n11758 , n11707 , n11757 );
and ( n11759 , n11754 , n11758 );
nor ( n11760 , n2013 , n160 );
nand ( n11761 , n1873 , n1834 );
and ( n11762 , n10893 , n11760 , n2018 , n11761 );
and ( n11763 , n1862 , n2190 );
not ( n11764 , n11763 );
not ( n11765 , n11764 );
not ( n11766 , n10802 );
or ( n11767 , n11765 , n11766 );
nand ( n11768 , n11767 , n2000 );
and ( n11769 , n11762 , n11768 );
nor ( n11770 , n11759 , n11769 );
not ( n11771 , n2107 );
not ( n11772 , n10818 );
or ( n11773 , n11771 , n11772 );
nand ( n11774 , n11773 , n10831 );
not ( n11775 , n11774 );
not ( n11776 , n1841 );
or ( n11777 , n11775 , n11776 );
and ( n11778 , n1915 , n1950 );
nor ( n11779 , n11778 , n161 );
nand ( n11780 , n1953 , n2190 );
nand ( n11781 , n1953 , n1956 );
and ( n11782 , n11780 , n11781 );
and ( n11783 , n10859 , n11779 , n11782 , n2191 );
nand ( n11784 , n11777 , n11783 );
or ( n11785 , n11770 , n11784 );
not ( n11786 , n2177 );
or ( n11787 , n2061 , n10826 , n11786 );
nand ( n11788 , n11787 , n1979 );
and ( n11789 , n1933 , n2194 );
nand ( n11790 , n11788 , n11789 );
not ( n11791 , n154 );
not ( n11792 , n2064 );
or ( n11793 , n11791 , n11792 );
nand ( n11794 , n11793 , n160 );
not ( n11795 , n11794 );
nand ( n11796 , n11795 , n2210 );
not ( n11797 , n11796 );
not ( n11798 , n1818 );
and ( n11799 , n11797 , n11798 );
nor ( n11800 , n11799 , n1846 );
or ( n11801 , n11790 , n11800 );
not ( n11802 , n2190 );
nor ( n11803 , n11802 , n1876 );
nor ( n11804 , n1851 , n2107 );
not ( n11805 , n1898 );
not ( n11806 , n1940 );
or ( n11807 , n11805 , n11806 );
nand ( n11808 , n11807 , n2177 );
nor ( n11809 , n11803 , n11804 , n11808 );
not ( n11810 , n2004 );
not ( n11811 , n10826 );
not ( n11812 , n11811 );
or ( n11813 , n11810 , n11812 );
nand ( n11814 , n11813 , n2000 );
nand ( n11815 , n11809 , n11814 );
nand ( n11816 , n11801 , n11815 );
not ( n11817 , n1978 );
and ( n11818 , n11817 , n2084 );
not ( n11819 , n1920 );
not ( n11820 , n2097 );
not ( n11821 , n11820 );
or ( n11822 , n11819 , n11821 );
nand ( n11823 , n11822 , n161 );
nor ( n11824 , n11818 , n11823 );
nand ( n11825 , n11816 , n11824 );
nand ( n11826 , n11785 , n11825 );
nand ( n11827 , n11737 , n11826 );
not ( n11828 , n11827 );
not ( n11829 , n11828 );
not ( n11830 , n288 );
and ( n11831 , n11829 , n11830 );
not ( n11832 , n11827 );
and ( n11833 , n11832 , n288 );
nor ( n11834 , n11831 , n11833 );
not ( n11835 , n11834 );
or ( n11836 , n11693 , n11835 );
or ( n11837 , n11834 , n10908 );
nand ( n11838 , n11836 , n11837 );
not ( n11839 , n11838 );
and ( n11840 , n11692 , n11839 );
not ( n11841 , n11692 );
and ( n11842 , n11841 , n11838 );
nor ( n11843 , n11840 , n11842 );
or ( n11844 , n11843 , n1 );
xnor ( n11845 , n288 , n289 );
or ( n11846 , n2246 , n11845 );
nand ( n11847 , n11844 , n11846 );
not ( n11848 , n1337 );
or ( n11849 , n10429 , n11848 );
nand ( n11850 , n11849 , n1280 );
not ( n11851 , n10518 );
and ( n11852 , n10414 , n1343 );
not ( n11853 , n11852 );
not ( n11854 , n11853 );
or ( n11855 , n11851 , n11854 );
nand ( n11856 , n11855 , n176 );
nand ( n11857 , n1466 , n173 );
nand ( n11858 , n1482 , n11857 );
or ( n11859 , n11858 , n1508 );
nand ( n11860 , n11859 , n1446 );
buf ( n11861 , n10480 );
nand ( n11862 , n11861 , n10408 );
nand ( n11863 , n11850 , n11856 , n11860 , n11862 );
not ( n11864 , n177 );
not ( n11865 , n10393 );
or ( n11866 , n11864 , n11865 );
nand ( n11867 , n11866 , n10431 );
and ( n11868 , n1414 , n10481 );
and ( n11869 , n10464 , n11867 , n11868 );
not ( n11870 , n176 );
nor ( n11871 , n11870 , n172 );
not ( n11872 , n11871 );
and ( n11873 , n1289 , n11872 );
nor ( n11874 , n11873 , n177 );
nand ( n11875 , n1326 , n11874 );
not ( n11876 , n1473 );
not ( n11877 , n1398 );
or ( n11878 , n11876 , n11877 );
nand ( n11879 , n11878 , n10518 );
nor ( n11880 , n11875 , n11879 );
or ( n11881 , n11869 , n11880 );
or ( n11882 , n10494 , n1298 );
and ( n11883 , n11882 , n178 );
nand ( n11884 , n11881 , n11883 );
or ( n11885 , n11863 , n11884 );
nand ( n11886 , n10403 , n10393 );
not ( n11887 , n1343 );
not ( n11888 , n1357 );
or ( n11889 , n11887 , n11888 );
nand ( n11890 , n11889 , n1280 );
or ( n11891 , n11886 , n11890 );
nand ( n11892 , n1289 , n173 );
not ( n11893 , n11892 );
not ( n11894 , n11893 );
nor ( n11895 , n10363 , n1280 );
nand ( n11896 , n11894 , n11895 );
nand ( n11897 , n11891 , n11896 );
not ( n11898 , n10378 );
nand ( n11899 , n11898 , n10374 );
or ( n11900 , n1531 , n1503 );
and ( n11901 , n10407 , n10447 , n11899 , n11900 );
and ( n11902 , n1361 , n1343 );
nand ( n11903 , n11902 , n10398 );
nand ( n11904 , n11903 , n177 );
not ( n11905 , n11904 );
nand ( n11906 , n11897 , n11901 , n11905 );
not ( n11907 , n11906 );
and ( n11908 , n10490 , n1537 );
nor ( n11909 , n11908 , n177 );
not ( n11910 , n11909 );
nand ( n11911 , n1365 , n1298 );
not ( n11912 , n11911 );
or ( n11913 , n11910 , n11912 );
nand ( n11914 , n11913 , n10389 );
buf ( n11915 , n1398 );
and ( n11916 , n11915 , n10402 );
not ( n11917 , n1442 );
nor ( n11918 , n11916 , n11917 );
nand ( n11919 , n11914 , n11918 );
not ( n11920 , n11919 );
or ( n11921 , n11907 , n11920 );
not ( n11922 , n1280 );
not ( n11923 , n1275 );
nand ( n11924 , n11923 , n173 );
not ( n11925 , n11924 );
or ( n11926 , n11922 , n11925 );
not ( n11927 , n10493 );
not ( n11928 , n174 );
and ( n11929 , n11927 , n11928 );
and ( n11930 , n1412 , n174 );
nor ( n11931 , n11929 , n11930 );
or ( n11932 , n11931 , n1537 );
nor ( n11933 , n10453 , n174 );
or ( n11934 , n11933 , n1468 );
nand ( n11935 , n11932 , n11934 );
nand ( n11936 , n11935 , n11900 , n176 );
nand ( n11937 , n11926 , n11936 );
not ( n11938 , n1493 );
not ( n11939 , n1383 );
or ( n11940 , n11938 , n11939 );
not ( n11941 , n11857 );
nand ( n11942 , n11941 , n1473 );
nand ( n11943 , n11940 , n11942 );
nand ( n11944 , n10491 , n1350 );
nor ( n11945 , n11943 , n11944 );
and ( n11946 , n11937 , n11945 );
nand ( n11947 , n11921 , n11946 );
nand ( n11948 , n11885 , n11947 );
not ( n11949 , n1280 );
not ( n11950 , n11924 );
not ( n11951 , n11950 );
or ( n11952 , n11949 , n11951 );
nand ( n11953 , n1524 , n11933 );
nand ( n11954 , n11952 , n11953 );
not ( n11955 , n11954 );
not ( n11956 , n177 );
or ( n11957 , n11955 , n11956 );
not ( n11958 , n1337 );
nand ( n11959 , n10462 , n10441 );
and ( n11960 , n1428 , n11959 );
not ( n11961 , n11960 );
or ( n11962 , n11958 , n11961 );
nand ( n11963 , n11962 , n1370 );
nand ( n11964 , n11957 , n11963 );
and ( n11965 , n11964 , n1375 );
nor ( n11966 , n11894 , n172 );
nand ( n11967 , n11966 , n1435 );
nor ( n11968 , n1339 , n175 );
and ( n11969 , n11968 , n1485 );
not ( n11970 , n10378 );
nand ( n11971 , n11970 , n10452 );
nor ( n11972 , n11971 , n1472 );
nor ( n11973 , n11969 , n11972 );
nand ( n11974 , n10460 , n11967 , n11973 );
nor ( n11975 , n11965 , n11974 );
not ( n11976 , n10517 );
not ( n11977 , n11976 );
not ( n11978 , n10414 );
nand ( n11979 , n10393 , n11978 );
or ( n11980 , n11979 , n11915 );
nand ( n11981 , n11980 , n1391 );
not ( n11982 , n11981 );
or ( n11983 , n11977 , n11982 );
nand ( n11984 , n11983 , n1306 );
not ( n11985 , n11984 );
not ( n11986 , n1285 );
not ( n11987 , n1524 );
or ( n11988 , n11986 , n11987 );
nand ( n11989 , n11988 , n176 );
not ( n11990 , n11989 );
not ( n11991 , n10476 );
not ( n11992 , n11991 );
and ( n11993 , n11990 , n11992 );
not ( n11994 , n10458 );
nor ( n11995 , n11993 , n11994 );
not ( n11996 , n11995 );
or ( n11997 , n11985 , n11996 );
nand ( n11998 , n11997 , n1370 );
nand ( n11999 , n11948 , n11975 , n11998 );
not ( n12000 , n11999 );
not ( n12001 , n12000 );
not ( n12002 , n11003 );
nand ( n12003 , n10982 , n1564 );
and ( n12004 , n10928 , n12003 , n1608 );
not ( n12005 , n12004 );
or ( n12006 , n12002 , n12005 );
nand ( n12007 , n12006 , n152 );
nor ( n12008 , n1696 , n1615 );
not ( n12009 , n1669 );
nand ( n12010 , n12009 , n146 );
nand ( n12011 , n11467 , n1603 );
nand ( n12012 , n12010 , n1626 , n12011 , n11528 );
or ( n12013 , n12008 , n12012 );
not ( n12014 , n11580 );
or ( n12015 , n12014 , n1579 );
nand ( n12016 , n12013 , n12015 );
not ( n12017 , n147 );
not ( n12018 , n1564 );
or ( n12019 , n12017 , n12018 );
not ( n12020 , n1613 );
not ( n12021 , n11509 );
nor ( n12022 , n12020 , n12021 );
nand ( n12023 , n12019 , n12022 );
nand ( n12024 , n12023 , n1712 );
not ( n12025 , n11481 );
nand ( n12026 , n12025 , n1774 );
nand ( n12027 , n1564 , n1695 );
and ( n12028 , n12024 , n12026 , n12027 );
not ( n12029 , n11586 );
not ( n12030 , n1702 );
or ( n12031 , n12029 , n12030 );
nand ( n12032 , n12031 , n1679 );
not ( n12033 , n10999 );
not ( n12034 , n12033 );
not ( n12035 , n1695 );
or ( n12036 , n12034 , n12035 );
nand ( n12037 , n12036 , n10929 );
or ( n12038 , n12032 , n12037 );
nand ( n12039 , n12038 , n1752 );
nand ( n12040 , n12007 , n12016 , n12028 , n12039 );
not ( n12041 , n10911 );
not ( n12042 , n11522 );
nand ( n12043 , n1583 , n150 );
not ( n12044 , n12043 );
or ( n12045 , n12042 , n12044 );
nand ( n12046 , n12045 , n1617 );
nand ( n12047 , n1594 , n1721 );
nand ( n12048 , n12041 , n12046 , n12047 , n10950 );
not ( n12049 , n10946 );
nand ( n12050 , n11601 , n147 );
nand ( n12051 , n12049 , n11556 , n12050 );
nor ( n12052 , n12048 , n12051 );
not ( n12053 , n1571 );
not ( n12054 , n11525 );
or ( n12055 , n12053 , n12054 );
nand ( n12056 , n12055 , n149 );
and ( n12057 , n12052 , n12056 );
nand ( n12058 , n10986 , n1660 );
nand ( n12059 , n1740 , n12058 , n1752 );
nand ( n12060 , n11629 , n1728 );
and ( n12061 , n12060 , n1615 );
nor ( n12062 , n12059 , n12061 );
nor ( n12063 , n12057 , n12062 );
nand ( n12064 , n12040 , n12063 );
nand ( n12065 , n12007 , n12039 );
nand ( n12066 , n12016 , n12028 );
or ( n12067 , n12065 , n12066 );
not ( n12068 , n1785 );
not ( n12069 , n1683 );
nand ( n12070 , n1653 , n1625 );
not ( n12071 , n12070 );
or ( n12072 , n12069 , n12071 );
nand ( n12073 , n12072 , n149 );
not ( n12074 , n12050 );
or ( n12075 , n12068 , n12073 , n12074 );
not ( n12076 , n1585 );
nand ( n12077 , n10982 , n12076 );
nand ( n12078 , n12077 , n1711 );
nand ( n12079 , n12075 , n12078 );
and ( n12080 , n11562 , n1711 );
and ( n12081 , n12021 , n11586 );
nor ( n12082 , n12080 , n12081 );
nor ( n12083 , n1614 , n153 );
nand ( n12084 , n12079 , n12082 , n12083 );
nand ( n12085 , n12067 , n12084 );
nand ( n12086 , n1660 , n1682 , n148 );
and ( n12087 , n1788 , n1752 );
and ( n12088 , n12026 , n12086 , n12087 );
not ( n12089 , n1575 );
nand ( n12090 , n1625 , n1599 );
nand ( n12091 , n12090 , n12043 );
or ( n12092 , n12091 , n1702 );
nand ( n12093 , n12092 , n1723 );
not ( n12094 , n12093 );
or ( n12095 , n12089 , n12094 );
nand ( n12096 , n12095 , n1615 );
not ( n12097 , n1671 );
not ( n12098 , n1794 );
or ( n12099 , n12097 , n12098 );
nand ( n12100 , n12099 , n1617 );
nand ( n12101 , n12088 , n12096 , n12100 );
not ( n12102 , n1699 );
not ( n12103 , n12102 );
nand ( n12104 , n12077 , n152 );
not ( n12105 , n12104 );
or ( n12106 , n12103 , n12105 );
nand ( n12107 , n12106 , n10934 );
and ( n12108 , n12101 , n12107 );
nand ( n12109 , n1695 , n1646 );
not ( n12110 , n12109 );
not ( n12111 , n149 );
or ( n12112 , n12110 , n12111 );
nand ( n12113 , n12112 , n1560 );
or ( n12114 , n1780 , n12113 );
nor ( n12115 , n1591 , n149 );
nor ( n12116 , n11008 , n12115 );
nand ( n12117 , n12114 , n12116 );
nor ( n12118 , n12108 , n12117 );
and ( n12119 , n12064 , n12085 , n12118 );
not ( n12120 , n12119 );
or ( n12121 , n12001 , n12120 );
not ( n12122 , n12119 );
nand ( n12123 , n12122 , n11999 );
nand ( n12124 , n12121 , n12123 );
xor ( n12125 , n12124 , n1547 );
not ( n12126 , n290 );
not ( n12127 , n12126 );
and ( n12128 , n10790 , n1959 );
nor ( n12129 , n12128 , n1868 );
not ( n12130 , n12129 );
not ( n12131 , n12130 );
not ( n12132 , n10808 );
not ( n12133 , n10867 );
or ( n12134 , n12132 , n12133 );
nand ( n12135 , n12134 , n10779 );
nand ( n12136 , n1831 , n1898 );
nand ( n12137 , n12136 , n2004 );
or ( n12138 , n12135 , n12137 );
nand ( n12139 , n12138 , n2000 );
not ( n12140 , n1902 );
not ( n12141 , n1860 );
or ( n12142 , n12140 , n12141 );
nand ( n12143 , n12142 , n1956 );
nor ( n12144 , n10878 , n10858 );
nand ( n12145 , n12139 , n12143 , n12144 );
not ( n12146 , n12145 );
or ( n12147 , n12131 , n12146 );
nand ( n12148 , n1865 , n158 );
or ( n12149 , n12148 , n2106 );
nand ( n12150 , n12149 , n2004 );
nor ( n12151 , n2187 , n12150 );
nand ( n12152 , n12151 , n1932 , n11781 );
not ( n12153 , n12152 );
not ( n12154 , n11707 );
buf ( n12155 , n2163 );
or ( n12156 , n12155 , n2084 );
or ( n12157 , n2179 , n159 );
nand ( n12158 , n12156 , n12157 );
or ( n12159 , n12158 , n11717 , n1862 );
nand ( n12160 , n12159 , n1841 );
not ( n12161 , n10808 );
nor ( n12162 , n1841 , n12161 );
or ( n12163 , n2125 , n12162 );
nand ( n12164 , n12163 , n159 );
and ( n12165 , n1988 , n156 );
not ( n12166 , n1851 );
and ( n12167 , n12166 , n1828 );
nor ( n12168 , n12165 , n12167 , n2050 );
nand ( n12169 , n12154 , n12160 , n12164 , n12168 );
not ( n12170 , n12169 );
or ( n12171 , n12153 , n12170 );
not ( n12172 , n1984 );
not ( n12173 , n1810 );
not ( n12174 , n11727 );
or ( n12175 , n12173 , n12174 );
nand ( n12176 , n1909 , n1987 );
nand ( n12177 , n12175 , n12176 );
not ( n12178 , n12177 );
or ( n12179 , n12172 , n12178 );
nand ( n12180 , n12179 , n159 );
not ( n12181 , n12180 );
not ( n12182 , n1950 );
not ( n12183 , n11713 );
or ( n12184 , n12182 , n12183 );
nand ( n12185 , n1862 , n1892 );
nand ( n12186 , n12184 , n12185 );
nor ( n12187 , n1984 , n156 );
nor ( n12188 , n12186 , n12187 , n161 );
nand ( n12189 , n10831 , n12188 );
nor ( n12190 , n12181 , n12189 );
nand ( n12191 , n12171 , n12190 );
not ( n12192 , n12191 );
nand ( n12193 , n12147 , n12192 );
not ( n12194 , n12193 );
nand ( n12195 , n10831 , n12129 );
not ( n12196 , n12195 );
not ( n12197 , n12145 );
or ( n12198 , n12196 , n12197 );
not ( n12199 , n1826 );
and ( n12200 , n12199 , n10794 , n10812 , n160 );
nand ( n12201 , n1993 , n12200 );
not ( n12202 , n2000 );
not ( n12203 , n1969 );
or ( n12204 , n12202 , n12203 );
not ( n12205 , n1960 );
nand ( n12206 , n2064 , n1890 );
not ( n12207 , n12206 );
or ( n12208 , n12205 , n12207 );
not ( n12209 , n1841 );
not ( n12210 , n1959 );
or ( n12211 , n12209 , n12210 );
nand ( n12212 , n12211 , n159 );
not ( n12213 , n12212 );
nand ( n12214 , n12208 , n12213 );
and ( n12215 , n1902 , n12214 , n2193 , n2004 );
nand ( n12216 , n12204 , n12215 );
and ( n12217 , n12201 , n12216 );
not ( n12218 , n1874 );
not ( n12219 , n1858 );
and ( n12220 , n12218 , n12219 );
and ( n12221 , n1995 , n159 );
nor ( n12222 , n12220 , n12221 );
nand ( n12223 , n10779 , n10863 );
or ( n12224 , n12223 , n11757 );
nand ( n12225 , n12224 , n1828 );
not ( n12226 , n11714 );
nor ( n12227 , n1957 , n154 );
or ( n12228 , n12226 , n12227 );
nand ( n12229 , n12228 , n1846 );
and ( n12230 , n12229 , n1836 );
nand ( n12231 , n12222 , n12225 , n12230 );
nor ( n12232 , n12217 , n12231 );
nand ( n12233 , n12198 , n12232 );
not ( n12234 , n12233 );
or ( n12235 , n12194 , n12234 );
not ( n12236 , n11817 );
nand ( n12237 , n12236 , n10889 );
and ( n12238 , n12237 , n2078 );
not ( n12239 , n11722 );
not ( n12240 , n1942 );
or ( n12241 , n12239 , n12240 );
nand ( n12242 , n12241 , n10859 );
nor ( n12243 , n12238 , n12242 );
nand ( n12244 , n12235 , n12243 );
not ( n12245 , n12244 );
or ( n12246 , n12127 , n12245 );
or ( n12247 , n12126 , n12244 );
nand ( n12248 , n12246 , n12247 );
not ( n12249 , n12248 );
and ( n12250 , n12125 , n12249 );
not ( n12251 , n12125 );
and ( n12252 , n12251 , n12248 );
nor ( n12253 , n12250 , n12252 );
or ( n12254 , n12253 , n1 );
and ( n12255 , n291 , n12126 );
not ( n12256 , n291 );
and ( n12257 , n12256 , n290 );
nor ( n12258 , n12255 , n12257 );
or ( n12259 , n2246 , n12258 );
nand ( n12260 , n12254 , n12259 );
nor ( n12261 , n8787 , n8881 );
nand ( n12262 , n7786 , n7240 );
not ( n12263 , n12262 );
not ( n12264 , n7683 );
or ( n12265 , n12263 , n12264 );
nand ( n12266 , n12265 , n7316 );
nand ( n12267 , n7288 , n2 );
nand ( n12268 , n7703 , n7733 );
and ( n12269 , n12261 , n12266 , n12267 , n12268 );
not ( n12270 , n12269 );
not ( n12271 , n7290 );
or ( n12272 , n12271 , n4 );
nand ( n12273 , n12272 , n7697 );
nand ( n12274 , n12273 , n7696 );
nor ( n12275 , n7817 , n7 );
nor ( n12276 , n7674 , n12271 );
nor ( n12277 , n12275 , n12276 );
nand ( n12278 , n7810 , n7765 , n8 );
or ( n12279 , n12278 , n9366 );
nand ( n12280 , n12279 , n8889 );
nand ( n12281 , n12274 , n12277 , n12280 );
nor ( n12282 , n12270 , n12281 );
not ( n12283 , n12282 );
or ( n12284 , n7410 , n3 );
nand ( n12285 , n12284 , n7 );
not ( n12286 , n7375 );
nor ( n12287 , n12285 , n12286 );
not ( n12288 , n7696 );
and ( n12289 , n7322 , n12287 , n12288 );
nand ( n12290 , n9397 , n4 );
not ( n12291 , n7671 );
not ( n12292 , n7818 );
and ( n12293 , n12290 , n12291 , n12292 );
or ( n12294 , n12289 , n12293 );
nand ( n12295 , n12294 , n7765 );
not ( n12296 , n7233 );
or ( n12297 , n12296 , n9409 );
nand ( n12298 , n12297 , n7265 );
nand ( n12299 , n7678 , n3 );
nand ( n12300 , n7715 , n12299 );
or ( n12301 , n12300 , n7779 );
nand ( n12302 , n12301 , n7698 );
nand ( n12303 , n12298 , n12302 , n9365 , n9 );
or ( n12304 , n12295 , n12303 );
nor ( n12305 , n9090 , n7 );
nor ( n12306 , n7821 , n9457 );
nor ( n12307 , n12306 , n7768 );
or ( n12308 , n12305 , n12307 );
not ( n12309 , n12262 );
nor ( n12310 , n12309 , n9 );
nand ( n12311 , n12308 , n12310 );
not ( n12312 , n12311 );
not ( n12313 , n7806 );
not ( n12314 , n9045 );
or ( n12315 , n12313 , n12314 );
nand ( n12316 , n12315 , n7 );
nand ( n12317 , n7690 , n7411 );
and ( n12318 , n7826 , n8839 , n12317 , n8880 );
nand ( n12319 , n12312 , n12316 , n12318 );
nand ( n12320 , n12304 , n12319 );
not ( n12321 , n12320 );
or ( n12322 , n12283 , n12321 );
nand ( n12323 , n7733 , n8822 , n7801 );
not ( n12324 , n12323 );
nand ( n12325 , n7354 , n8880 , n7325 , n7316 );
not ( n12326 , n12325 );
or ( n12327 , n12324 , n12326 );
and ( n12328 , n7798 , n8794 , n9027 );
nand ( n12329 , n12327 , n12328 );
nor ( n12330 , n12303 , n12329 );
not ( n12331 , n7265 );
not ( n12332 , n7364 );
or ( n12333 , n12331 , n12332 );
nand ( n12334 , n7336 , n4 );
nand ( n12335 , n8822 , n12334 , n9396 );
nand ( n12336 , n12333 , n12335 );
nor ( n12337 , n12296 , n8 );
nand ( n12338 , n9116 , n12336 , n12337 );
nor ( n12339 , n12338 , n12311 );
or ( n12340 , n12330 , n12339 );
nand ( n12341 , n12340 , n12269 );
nand ( n12342 , n12322 , n12341 );
not ( n12343 , n12342 );
nand ( n12344 , n6379 , n6356 );
not ( n12345 , n12344 );
not ( n12346 , n9483 );
nor ( n12347 , n12346 , n9506 );
nand ( n12348 , n12345 , n12347 );
not ( n12349 , n6308 );
and ( n12350 , n6467 , n6430 );
nor ( n12351 , n12350 , n8471 );
nand ( n12352 , n12349 , n12351 );
and ( n12353 , n12348 , n12352 );
nor ( n12354 , n12353 , n6397 );
not ( n12355 , n12354 );
and ( n12356 , n6327 , n6348 , n25 );
not ( n12357 , n12356 );
not ( n12358 , n8039 );
nand ( n12359 , n12358 , n9512 , n6339 );
nand ( n12360 , n12357 , n12359 , n8109 , n6355 );
or ( n12361 , n12360 , n6320 );
not ( n12362 , n6604 );
nor ( n12363 , n12362 , n6473 , n26 );
nand ( n12364 , n6291 , n25 );
nand ( n12365 , n12363 , n8487 , n8023 , n12364 );
nand ( n12366 , n12361 , n12365 );
not ( n12367 , n12366 );
or ( n12368 , n12355 , n12367 );
not ( n12369 , n6299 );
not ( n12370 , n6563 );
or ( n12371 , n12369 , n12370 );
not ( n12372 , n6634 );
nor ( n12373 , n12372 , n6356 );
not ( n12374 , n12373 );
not ( n12375 , n8107 );
or ( n12376 , n12374 , n12375 );
nand ( n12377 , n12376 , n6470 );
not ( n12378 , n6620 );
nor ( n12379 , n12378 , n23 );
nor ( n12380 , n6642 , n12379 );
nand ( n12381 , n12377 , n12380 );
nand ( n12382 , n12371 , n12381 );
not ( n12383 , n6299 );
not ( n12384 , n8470 );
not ( n12385 , n8065 );
not ( n12386 , n12385 );
or ( n12387 , n12384 , n12386 );
nand ( n12388 , n12387 , n8476 );
not ( n12389 , n12388 );
or ( n12390 , n12383 , n12389 );
nand ( n12391 , n12390 , n6432 );
nor ( n12392 , n8073 , n6493 );
or ( n12393 , n12391 , n12392 );
nand ( n12394 , n12393 , n26 );
and ( n12395 , n8425 , n6539 );
and ( n12396 , n6313 , n6320 , n23 );
not ( n12397 , n6320 );
not ( n12398 , n6521 );
or ( n12399 , n12397 , n12398 );
nand ( n12400 , n12399 , n6339 );
and ( n12401 , n6519 , n12400 );
nor ( n12402 , n12396 , n12401 );
nand ( n12403 , n12382 , n12394 , n12395 , n12402 );
nand ( n12404 , n12368 , n12403 );
nand ( n12405 , n6404 , n6299 );
not ( n12406 , n12405 );
not ( n12407 , n8410 );
nand ( n12408 , n12406 , n12407 , n9492 );
not ( n12409 , n12408 );
not ( n12410 , n8093 );
nor ( n12411 , n12410 , n8432 );
not ( n12412 , n6667 );
nor ( n12413 , n12412 , n6356 );
nand ( n12414 , n9482 , n12411 , n12413 , n6441 );
not ( n12415 , n12414 );
or ( n12416 , n12409 , n12415 );
and ( n12417 , n8425 , n6498 , n6447 );
nand ( n12418 , n12416 , n12417 );
or ( n12419 , n8019 , n12344 , n6527 );
not ( n12420 , n6470 );
nand ( n12421 , n12420 , n6660 );
nand ( n12422 , n12419 , n12421 );
and ( n12423 , n8472 , n6631 , n6501 );
nand ( n12424 , n12422 , n12423 );
nand ( n12425 , n12418 , n12424 );
not ( n12426 , n6356 );
not ( n12427 , n6674 );
or ( n12428 , n12426 , n12427 );
or ( n12429 , n9545 , n6679 );
nand ( n12430 , n12428 , n12429 );
nand ( n12431 , n12404 , n12425 , n12430 );
not ( n12432 , n12431 );
not ( n12433 , n12432 );
and ( n12434 , n12343 , n12433 );
not ( n12435 , n12432 );
not ( n12436 , n12435 );
and ( n12437 , n12436 , n12342 );
nor ( n12438 , n12434 , n12437 );
not ( n12439 , n8274 );
and ( n12440 , n12438 , n12439 );
not ( n12441 , n12438 );
and ( n12442 , n12441 , n8274 );
nor ( n12443 , n12440 , n12442 );
not ( n12444 , n7486 );
not ( n12445 , n7664 );
or ( n12446 , n12444 , n12445 );
or ( n12447 , n7490 , n7668 );
nand ( n12448 , n12446 , n12447 );
xor ( n12449 , n7834 , n84 );
not ( n12450 , n12449 );
and ( n12451 , n12448 , n12450 );
not ( n12452 , n12448 );
and ( n12453 , n12452 , n12449 );
nor ( n12454 , n12451 , n12453 );
not ( n12455 , n12454 );
and ( n12456 , n12443 , n12455 );
not ( n12457 , n12443 );
and ( n12458 , n12457 , n12454 );
nor ( n12459 , n12456 , n12458 );
or ( n12460 , n12459 , n1 );
xnor ( n12461 , n84 , n85 );
or ( n12462 , n2246 , n12461 );
nand ( n12463 , n12460 , n12462 );
not ( n12464 , n4305 );
nor ( n12465 , n12464 , n5350 );
not ( n12466 , n5336 );
nor ( n12467 , n11314 , n12466 );
nand ( n12468 , n12465 , n12467 , n11355 );
not ( n12469 , n12468 );
not ( n12470 , n5912 );
not ( n12471 , n3605 );
and ( n12472 , n12470 , n12471 );
nor ( n12473 , n12472 , n3525 );
nand ( n12474 , n12473 , n5368 , n3481 , n3458 );
not ( n12475 , n12474 );
or ( n12476 , n12469 , n12475 );
nand ( n12477 , n12466 , n209 );
and ( n12478 , n5299 , n12477 , n5364 );
nand ( n12479 , n12476 , n12478 );
not ( n12480 , n4215 );
not ( n12481 , n5919 );
or ( n12482 , n12480 , n12481 );
nand ( n12483 , n12482 , n11314 );
and ( n12484 , n4232 , n9636 , n5947 );
and ( n12485 , n12483 , n12484 );
nor ( n12486 , n12485 , n5288 );
or ( n12487 , n12479 , n12486 );
nand ( n12488 , n5367 , n206 );
not ( n12489 , n5951 );
nand ( n12490 , n12489 , n3630 );
and ( n12491 , n5329 , n12488 , n12490 );
nand ( n12492 , n12491 , n3526 );
not ( n12493 , n12492 );
not ( n12494 , n3665 );
not ( n12495 , n4356 );
or ( n12496 , n12494 , n12495 );
nand ( n12497 , n12496 , n5291 );
or ( n12498 , n9676 , n12497 );
not ( n12499 , n3535 );
not ( n12500 , n3461 );
nand ( n12501 , n12500 , n209 );
or ( n12502 , n12499 , n12501 );
nand ( n12503 , n12498 , n12502 );
nand ( n12504 , n3457 , n3638 );
nand ( n12505 , n9663 , n12504 );
nor ( n12506 , n4357 , n5946 , n12505 , n5253 );
nand ( n12507 , n12503 , n12506 );
not ( n12508 , n12507 );
or ( n12509 , n12493 , n12508 );
not ( n12510 , n3506 );
not ( n12511 , n3487 );
nand ( n12512 , n12511 , n205 );
not ( n12513 , n12512 );
or ( n12514 , n12510 , n12513 );
nand ( n12515 , n12514 , n5322 );
and ( n12516 , n12515 , n5990 , n12504 );
nor ( n12517 , n12516 , n3471 );
nand ( n12518 , n5302 , n3485 );
nor ( n12519 , n4225 , n212 );
nand ( n12520 , n12518 , n12519 );
nor ( n12521 , n12517 , n12520 , n9657 );
nand ( n12522 , n12509 , n12521 );
nand ( n12523 , n12487 , n12522 );
not ( n12524 , n5296 );
nand ( n12525 , n12524 , n3605 );
not ( n12526 , n12477 );
or ( n12527 , n3670 , n11370 );
nand ( n12528 , n12527 , n3691 , n3619 );
nor ( n12529 , n12526 , n12528 );
and ( n12530 , n12525 , n12529 );
not ( n12531 , n3462 );
not ( n12532 , n5946 );
or ( n12533 , n12531 , n12532 );
nand ( n12534 , n12533 , n12518 );
nand ( n12535 , n5312 , n209 );
and ( n12536 , n12535 , n211 );
nor ( n12537 , n12536 , n3462 );
nor ( n12538 , n12534 , n12537 );
nor ( n12539 , n12530 , n12538 );
not ( n12540 , n5252 );
not ( n12541 , n3700 );
or ( n12542 , n12540 , n12541 );
nand ( n12543 , n12542 , n3471 );
not ( n12544 , n4217 );
not ( n12545 , n3582 );
not ( n12546 , n3637 );
and ( n12547 , n12545 , n12546 );
nor ( n12548 , n12547 , n4336 );
not ( n12549 , n12548 );
or ( n12550 , n12544 , n12549 );
nand ( n12551 , n12550 , n4258 );
nand ( n12552 , n12543 , n12551 , n3672 );
nor ( n12553 , n12539 , n12552 );
nand ( n12554 , n12523 , n12553 );
not ( n12555 , n12554 );
not ( n12556 , n12555 );
not ( n12557 , n9755 );
nand ( n12558 , n4812 , n12557 , n4704 , n3741 );
not ( n12559 , n12558 );
nand ( n12560 , n4916 , n3862 , n3749 );
nor ( n12561 , n9772 , n12560 );
nand ( n12562 , n4995 , n3858 );
nor ( n12563 , n5013 , n12562 );
or ( n12564 , n12561 , n12563 );
not ( n12565 , n3879 );
or ( n12566 , n3949 , n12565 );
nand ( n12567 , n12564 , n12566 );
not ( n12568 , n12567 );
or ( n12569 , n12559 , n12568 );
nand ( n12570 , n12569 , n5025 );
not ( n12571 , n3786 );
nand ( n12572 , n4916 , n186 );
or ( n12573 , n12572 , n183 );
not ( n12574 , n5043 );
nand ( n12575 , n12573 , n12574 );
not ( n12576 , n12575 );
or ( n12577 , n12571 , n12576 );
and ( n12578 , n3719 , n3811 );
nand ( n12579 , n12577 , n12578 );
not ( n12580 , n12579 );
not ( n12581 , n4675 );
not ( n12582 , n12581 );
not ( n12583 , n12572 );
or ( n12584 , n12583 , n5043 );
or ( n12585 , n5067 , n4789 );
nand ( n12586 , n12584 , n12585 );
nand ( n12587 , n12582 , n4678 , n12586 );
not ( n12588 , n12587 );
and ( n12589 , n12580 , n12588 );
and ( n12590 , n9773 , n3905 );
nor ( n12591 , n12589 , n12590 );
or ( n12592 , n12570 , n12591 );
and ( n12593 , n5048 , n186 );
nand ( n12594 , n4881 , n5073 );
nor ( n12595 , n12594 , n4756 );
not ( n12596 , n4669 );
not ( n12597 , n3755 );
or ( n12598 , n12596 , n12597 );
nand ( n12599 , n12598 , n184 );
nand ( n12600 , n12593 , n12595 , n12599 );
not ( n12601 , n3732 );
not ( n12602 , n3868 );
or ( n12603 , n12601 , n12602 );
not ( n12604 , n4760 );
not ( n12605 , n12604 );
not ( n12606 , n3723 );
or ( n12607 , n12605 , n12606 );
nand ( n12608 , n12607 , n185 );
nand ( n12609 , n12603 , n12608 );
and ( n12610 , n12609 , n4840 );
nor ( n12611 , n3772 , n185 );
nor ( n12612 , n12600 , n12610 , n12611 );
nor ( n12613 , n5014 , n186 );
not ( n12614 , n3731 );
nand ( n12615 , n12614 , n3715 );
nand ( n12616 , n3849 , n3829 );
and ( n12617 , n12613 , n12615 , n4697 , n12616 );
or ( n12618 , n12612 , n12617 );
nand ( n12619 , n9781 , n9746 );
not ( n12620 , n184 );
not ( n12621 , n9738 );
or ( n12622 , n12620 , n12621 );
nand ( n12623 , n4805 , n185 );
nor ( n12624 , n3928 , n12623 );
nand ( n12625 , n12622 , n12624 );
and ( n12626 , n12619 , n12625 );
nand ( n12627 , n4946 , n5007 );
nor ( n12628 , n12626 , n12627 );
nand ( n12629 , n12618 , n12628 );
nand ( n12630 , n12592 , n12629 );
not ( n12631 , n4805 );
not ( n12632 , n5029 );
or ( n12633 , n12631 , n12632 );
nand ( n12634 , n12633 , n3854 );
not ( n12635 , n3916 );
not ( n12636 , n4723 );
or ( n12637 , n12635 , n12636 );
nand ( n12638 , n12637 , n181 );
or ( n12639 , n12638 , n4708 );
nand ( n12640 , n12639 , n4873 );
nand ( n12641 , n12640 , n3811 );
not ( n12642 , n4995 );
and ( n12643 , n12642 , n185 );
or ( n12644 , n3778 , n4835 );
nand ( n12645 , n12644 , n3749 );
nor ( n12646 , n12643 , n12645 );
nand ( n12647 , n12634 , n12641 , n12646 );
not ( n12648 , n3824 );
or ( n12649 , n12648 , n4820 );
not ( n12650 , n4792 );
nand ( n12651 , n12649 , n12650 , n186 );
and ( n12652 , n12647 , n12651 );
not ( n12653 , n3923 );
not ( n12654 , n186 );
not ( n12655 , n4978 );
or ( n12656 , n12654 , n12655 );
nand ( n12657 , n12656 , n5048 );
nand ( n12658 , n12657 , n3811 );
nand ( n12659 , n12653 , n12658 , n9795 );
nor ( n12660 , n12652 , n12659 );
nand ( n12661 , n12630 , n12660 );
not ( n12662 , n12661 );
not ( n12663 , n12662 );
or ( n12664 , n12556 , n12663 );
nand ( n12665 , n12554 , n12661 );
nand ( n12666 , n12664 , n12665 );
not ( n12667 , n4413 );
nand ( n12668 , n4514 , n192 );
not ( n12669 , n12668 );
not ( n12670 , n12669 );
or ( n12671 , n12667 , n12670 );
nand ( n12672 , n4454 , n4529 );
nand ( n12673 , n12671 , n12672 );
not ( n12674 , n12673 );
and ( n12675 , n5583 , n188 );
not ( n12676 , n6212 );
nor ( n12677 , n12675 , n12676 , n4390 );
nand ( n12678 , n4600 , n4415 );
nor ( n12679 , n12677 , n12678 );
nand ( n12680 , n4597 , n5554 );
nand ( n12681 , n12674 , n12679 , n4391 , n12680 );
not ( n12682 , n12681 );
not ( n12683 , n192 );
nand ( n12684 , n12683 , n4521 );
nand ( n12685 , n6209 , n4643 , n12684 );
nor ( n12686 , n5600 , n12685 );
nand ( n12687 , n4590 , n4604 );
or ( n12688 , n12687 , n6147 );
nand ( n12689 , n12688 , n4452 );
not ( n12690 , n4615 );
nor ( n12691 , n12690 , n5562 );
nand ( n12692 , n12689 , n12691 );
nor ( n12693 , n12692 , n5524 );
or ( n12694 , n12686 , n12693 );
not ( n12695 , n11249 );
not ( n12696 , n4468 );
and ( n12697 , n5566 , n12668 );
not ( n12698 , n12697 );
or ( n12699 , n12696 , n12698 );
nand ( n12700 , n12699 , n4605 );
nand ( n12701 , n12695 , n12700 );
not ( n12702 , n6188 );
not ( n12703 , n6043 );
nor ( n12704 , n4481 , n12703 );
not ( n12705 , n12704 );
or ( n12706 , n12702 , n12705 );
nand ( n12707 , n12706 , n6038 );
not ( n12708 , n4515 );
not ( n12709 , n6029 );
or ( n12710 , n12708 , n12709 );
nand ( n12711 , n12710 , n4437 );
nand ( n12712 , n12707 , n12711 );
nor ( n12713 , n12701 , n12712 );
nand ( n12714 , n12694 , n12713 );
not ( n12715 , n12714 );
or ( n12716 , n12682 , n12715 );
not ( n12717 , n4496 );
not ( n12718 , n4503 );
or ( n12719 , n12717 , n12718 );
nand ( n12720 , n12719 , n6188 );
or ( n12721 , n12720 , n5626 );
nand ( n12722 , n12721 , n4452 );
not ( n12723 , n6029 );
or ( n12724 , n11261 , n12723 );
nand ( n12725 , n12724 , n4437 );
nor ( n12726 , n4418 , n4617 );
nand ( n12727 , n12722 , n12725 , n12726 );
or ( n12728 , n6198 , n4604 );
nand ( n12729 , n12728 , n6248 );
nand ( n12730 , n4391 , n12729 );
and ( n12731 , n12727 , n12730 );
nor ( n12732 , n5591 , n193 );
not ( n12733 , n12732 );
not ( n12734 , n11202 );
not ( n12735 , n4538 );
and ( n12736 , n12734 , n12735 );
nor ( n12737 , n12736 , n5531 );
nand ( n12738 , n12733 , n12737 , n4419 );
nor ( n12739 , n12731 , n12738 );
nand ( n12740 , n12716 , n12739 );
not ( n12741 , n12740 );
or ( n12742 , n4607 , n4576 );
not ( n12743 , n12742 );
not ( n12744 , n6096 );
or ( n12745 , n4390 , n4496 );
nand ( n12746 , n12745 , n4436 );
not ( n12747 , n12746 );
or ( n12748 , n12744 , n12747 );
and ( n12749 , n6113 , n4503 );
and ( n12750 , n4496 , n4427 );
nor ( n12751 , n12749 , n12750 );
nor ( n12752 , n6208 , n193 );
nand ( n12753 , n12751 , n12752 , n4573 );
nand ( n12754 , n12748 , n12753 );
and ( n12755 , n4434 , n4503 );
not ( n12756 , n11275 );
nor ( n12757 , n12755 , n4493 , n12756 );
nand ( n12758 , n12743 , n12754 , n12757 );
nand ( n12759 , n4383 , n4437 );
not ( n12760 , n4629 );
not ( n12761 , n188 );
nand ( n12762 , n12761 , n190 );
nor ( n12763 , n12760 , n12762 );
or ( n12764 , n5543 , n12763 );
nor ( n12765 , n4529 , n189 );
nand ( n12766 , n12764 , n12765 );
nand ( n12767 , n12759 , n12766 , n4504 , n4576 );
nand ( n12768 , n12714 , n12758 , n12767 );
nand ( n12769 , n12741 , n12768 );
not ( n12770 , n12769 );
not ( n12771 , n12770 );
not ( n12772 , n270 );
and ( n12773 , n12771 , n12772 );
and ( n12774 , n12770 , n270 );
nor ( n12775 , n12773 , n12774 );
and ( n12776 , n11421 , n12775 );
not ( n12777 , n11421 );
not ( n12778 , n12775 );
and ( n12779 , n12777 , n12778 );
nor ( n12780 , n12776 , n12779 );
and ( n12781 , n12666 , n12780 );
not ( n12782 , n12666 );
not ( n12783 , n12780 );
and ( n12784 , n12782 , n12783 );
nor ( n12785 , n12781 , n12784 );
or ( n12786 , n12785 , n1 );
xnor ( n12787 , n270 , n271 );
or ( n12788 , n2246 , n12787 );
nand ( n12789 , n12786 , n12788 );
nand ( n12790 , n1940 , n1950 );
not ( n12791 , n12790 );
not ( n12792 , n2198 );
or ( n12793 , n12791 , n12792 );
nand ( n12794 , n12793 , n1868 );
and ( n12795 , n1947 , n12794 );
nand ( n12796 , n2147 , n1864 );
not ( n12797 , n10779 );
nand ( n12798 , n12797 , n1921 );
nand ( n12799 , n12795 , n12796 , n12798 );
not ( n12800 , n12213 );
not ( n12801 , n11756 );
or ( n12802 , n12800 , n12801 );
nor ( n12803 , n1919 , n2009 );
nand ( n12804 , n10816 , n12803 );
nand ( n12805 , n12802 , n12804 );
not ( n12806 , n2061 );
and ( n12807 , n12805 , n12806 );
nor ( n12808 , n12807 , n1868 );
or ( n12809 , n12799 , n12808 );
nand ( n12810 , n12809 , n1905 );
not ( n12811 , n2026 );
and ( n12812 , n1882 , n1815 );
nor ( n12813 , n12812 , n2106 , n158 );
nor ( n12814 , n12811 , n12813 );
and ( n12815 , n12810 , n12814 );
and ( n12816 , n11717 , n1950 );
not ( n12817 , n11745 );
and ( n12818 , n12817 , n1846 );
and ( n12819 , n1984 , n11722 );
nor ( n12820 , n12818 , n12819 );
nor ( n12821 , n12816 , n12820 );
not ( n12822 , n1986 );
not ( n12823 , n10779 );
or ( n12824 , n12822 , n12823 );
nand ( n12825 , n12824 , n1828 );
not ( n12826 , n12825 );
or ( n12827 , n10792 , n154 );
not ( n12828 , n12827 );
or ( n12829 , n1843 , n1967 , n12828 );
nand ( n12830 , n12829 , n159 );
buf ( n12831 , n1884 );
not ( n12832 , n2008 );
or ( n12833 , n1833 , n12832 );
nand ( n12834 , n12833 , n2004 );
nor ( n12835 , n10785 , n12834 );
nand ( n12836 , n12830 , n12831 , n12835 );
nor ( n12837 , n12826 , n12836 );
or ( n12838 , n12821 , n12837 );
not ( n12839 , n10802 );
or ( n12840 , n12839 , n11820 , n1873 );
nand ( n12841 , n12840 , n1921 );
not ( n12842 , n10893 );
not ( n12843 , n10868 );
not ( n12844 , n2191 );
nor ( n12845 , n12842 , n12843 , n12844 );
and ( n12846 , n12841 , n12845 );
nand ( n12847 , n12838 , n12846 );
nand ( n12848 , n12847 , n161 );
not ( n12849 , n1868 );
or ( n12850 , n12828 , n2073 );
nand ( n12851 , n12850 , n1810 );
not ( n12852 , n12851 );
or ( n12853 , n12849 , n12852 );
not ( n12854 , n12155 );
not ( n12855 , n12854 );
not ( n12856 , n10790 );
or ( n12857 , n12855 , n12856 );
and ( n12858 , n1817 , n11722 );
nand ( n12859 , n12857 , n12858 );
or ( n12860 , n12135 , n12859 );
not ( n12861 , n2084 );
not ( n12862 , n11751 );
or ( n12863 , n12861 , n12862 );
nand ( n12864 , n12863 , n160 );
not ( n12865 , n12864 );
nand ( n12866 , n12865 , n11789 );
nand ( n12867 , n12860 , n12866 );
nand ( n12868 , n12867 , n12236 );
nand ( n12869 , n12853 , n12868 );
not ( n12870 , n10844 );
and ( n12871 , n12870 , n156 );
nand ( n12872 , n10793 , n1898 );
not ( n12873 , n159 );
nand ( n12874 , n12872 , n12873 );
nor ( n12875 , n12871 , n12874 );
and ( n12876 , n12875 , n12136 );
not ( n12877 , n12148 );
nor ( n12878 , n2199 , n12877 , n1979 );
and ( n12879 , n12878 , n11761 );
nor ( n12880 , n12876 , n12879 );
nand ( n12881 , n12868 , n12880 );
nand ( n12882 , n12815 , n12848 , n12869 , n12881 );
xor ( n12883 , n334 , n12882 );
not ( n12884 , n12883 );
not ( n12885 , n2235 );
or ( n12886 , n12884 , n12885 );
not ( n12887 , n12883 );
nand ( n12888 , n12887 , n2234 );
nand ( n12889 , n12886 , n12888 );
not ( n12890 , n999 );
not ( n12891 , n11577 );
or ( n12892 , n12890 , n12891 );
not ( n12893 , n11577 );
nand ( n12894 , n12893 , n998 );
nand ( n12895 , n12892 , n12894 );
not ( n12896 , n152 );
and ( n12897 , n1781 , n1597 , n1711 );
not ( n12898 , n12897 );
or ( n12899 , n12896 , n12898 );
nand ( n12900 , n10920 , n1699 );
nand ( n12901 , n12899 , n12900 );
nand ( n12902 , n12901 , n1790 );
or ( n12903 , n12902 , n11588 );
and ( n12904 , n149 , n12070 );
not ( n12905 , n149 );
and ( n12906 , n12905 , n12010 );
or ( n12907 , n12904 , n12906 );
not ( n12908 , n1567 );
nor ( n12909 , n12908 , n11634 , n1604 );
not ( n12910 , n1656 );
not ( n12911 , n1599 );
or ( n12912 , n12910 , n12911 );
nand ( n12913 , n12912 , n11623 );
nand ( n12914 , n12907 , n12909 , n12913 );
nand ( n12915 , n12903 , n12914 );
not ( n12916 , n1774 );
nand ( n12917 , n12916 , n10960 );
or ( n12918 , n12917 , n11461 );
nand ( n12919 , n12918 , n1660 );
and ( n12920 , n1695 , n10999 );
not ( n12921 , n1769 );
nor ( n12922 , n12920 , n12921 );
and ( n12923 , n12919 , n12922 );
nand ( n12924 , n12915 , n12923 );
nand ( n12925 , n12924 , n153 );
not ( n12926 , n10983 );
nand ( n12927 , n12926 , n148 );
not ( n12928 , n12927 );
not ( n12929 , n11013 );
or ( n12930 , n12928 , n12929 );
nand ( n12931 , n12930 , n1617 );
nand ( n12932 , n1594 , n1620 );
not ( n12933 , n12932 );
not ( n12934 , n1671 );
or ( n12935 , n12933 , n12934 );
nand ( n12936 , n12935 , n149 );
nand ( n12937 , n1631 , n10998 );
and ( n12938 , n1779 , n12937 , n152 );
nand ( n12939 , n12931 , n12936 , n12938 );
not ( n12940 , n1617 );
nand ( n12941 , n10982 , n1793 );
nand ( n12942 , n1794 , n1684 , n12941 );
not ( n12943 , n12942 );
or ( n12944 , n12940 , n12943 );
not ( n12945 , n1752 );
not ( n12946 , n1771 );
or ( n12947 , n12945 , n12946 );
nand ( n12948 , n12947 , n1560 );
and ( n12949 , n1703 , n11552 );
not ( n12950 , n1775 );
nor ( n12951 , n1639 , n147 );
nor ( n12952 , n11570 , n12951 );
not ( n12953 , n12952 );
or ( n12954 , n12950 , n12953 );
nand ( n12955 , n12954 , n149 );
and ( n12956 , n12948 , n12949 , n12955 );
nand ( n12957 , n12944 , n12956 );
and ( n12958 , n12939 , n12957 );
not ( n12959 , n1703 );
nand ( n12960 , n12959 , n11586 );
or ( n12961 , n1590 , n1763 );
nand ( n12962 , n12961 , n11603 );
nand ( n12963 , n12960 , n12962 );
nor ( n12964 , n12958 , n12963 );
nand ( n12965 , n11043 , n11037 );
not ( n12966 , n12965 );
and ( n12967 , n12966 , n1626 );
not ( n12968 , n11037 );
nor ( n12969 , n12968 , n149 );
nor ( n12970 , n12967 , n12969 );
not ( n12971 , n11015 );
nand ( n12972 , n12971 , n10932 );
not ( n12973 , n12972 );
not ( n12974 , n12897 );
or ( n12975 , n12973 , n12974 );
nand ( n12976 , n12975 , n152 );
or ( n12977 , n12970 , n12976 );
nand ( n12978 , n11572 , n11587 , n1752 );
nand ( n12979 , n12977 , n12978 );
not ( n12980 , n12979 );
nor ( n12981 , n12010 , n1659 );
nor ( n12982 , n12981 , n12115 , n1586 );
not ( n12983 , n12982 );
or ( n12984 , n12980 , n12983 );
nand ( n12985 , n12984 , n1735 );
and ( n12986 , n12925 , n12964 , n12985 );
not ( n12987 , n12986 );
not ( n12988 , n11902 );
nand ( n12989 , n1505 , n10458 , n12988 );
nor ( n12990 , n12989 , n10473 );
and ( n12991 , n11861 , n10462 );
nand ( n12992 , n1290 , n1370 , n176 );
or ( n12993 , n12991 , n12992 );
nand ( n12994 , n10524 , n10407 , n10390 );
nand ( n12995 , n12993 , n12994 );
and ( n12996 , n12990 , n12995 );
not ( n12997 , n1275 );
not ( n12998 , n10379 );
and ( n12999 , n1303 , n12998 , n1435 );
not ( n13000 , n12999 );
or ( n13001 , n12997 , n13000 );
nand ( n13002 , n1329 , n1446 );
nand ( n13003 , n13001 , n13002 );
nand ( n13004 , n10402 , n1532 );
not ( n13005 , n13004 );
not ( n13006 , n13005 );
nand ( n13007 , n13006 , n1526 , n1358 );
nor ( n13008 , n13007 , n11950 );
and ( n13009 , n13003 , n13008 );
nor ( n13010 , n12996 , n13009 );
and ( n13011 , n11981 , n11882 );
nand ( n13012 , n1302 , n1343 );
nand ( n13013 , n13012 , n178 );
not ( n13014 , n174 );
not ( n13015 , n10363 );
or ( n13016 , n13014 , n13015 );
nand ( n13017 , n13016 , n10464 );
or ( n13018 , n13013 , n13017 );
nand ( n13019 , n176 , n178 );
nand ( n13020 , n13018 , n13019 );
nand ( n13021 , n13011 , n13020 );
or ( n13022 , n13010 , n13021 );
not ( n13023 , n1489 );
not ( n13024 , n11966 );
not ( n13025 , n13024 );
or ( n13026 , n13023 , n13025 );
nand ( n13027 , n13026 , n1435 );
nand ( n13028 , n1383 , n11970 );
nand ( n13029 , n13028 , n1536 );
not ( n13030 , n10353 );
or ( n13031 , n13029 , n11917 , n13030 );
nand ( n13032 , n13031 , n177 );
nand ( n13033 , n13027 , n13032 );
not ( n13034 , n1370 );
nand ( n13035 , n11950 , n1473 );
nand ( n13036 , n1365 , n173 );
not ( n13037 , n1391 );
not ( n13038 , n1363 );
or ( n13039 , n13037 , n13038 );
nand ( n13040 , n11871 , n171 );
or ( n13041 , n13040 , n10490 );
nand ( n13042 , n13039 , n13041 );
not ( n13043 , n13012 );
nor ( n13044 , n13042 , n13043 );
nand ( n13045 , n13035 , n13036 , n13044 );
not ( n13046 , n13045 );
or ( n13047 , n13034 , n13046 );
not ( n13048 , n10518 );
nor ( n13049 , n1296 , n1298 );
nor ( n13050 , n13048 , n13049 );
nand ( n13051 , n13050 , n1280 );
not ( n13052 , n10453 );
nand ( n13053 , n13052 , n1524 );
nand ( n13054 , n13053 , n1533 , n176 );
and ( n13055 , n13051 , n13054 );
nand ( n13056 , n11853 , n1350 );
nor ( n13057 , n13055 , n13056 );
nand ( n13058 , n13047 , n13057 );
or ( n13059 , n13033 , n13058 );
nand ( n13060 , n13022 , n13059 );
nand ( n13061 , n11853 , n1414 );
and ( n13062 , n13061 , n10419 );
or ( n13063 , n1482 , n1434 , n1285 );
nor ( n13064 , n1435 , n1418 );
or ( n13065 , n1526 , n13064 );
nand ( n13066 , n13063 , n13065 );
nor ( n13067 , n13062 , n13066 );
not ( n13068 , n10474 );
or ( n13069 , n1387 , n10389 );
nand ( n13070 , n13069 , n10424 );
nor ( n13071 , n13068 , n13070 );
nand ( n13072 , n1286 , n1473 );
nand ( n13073 , n13072 , n1392 );
buf ( n13074 , n11899 );
nand ( n13075 , n1408 , n173 );
and ( n13076 , n13074 , n1404 , n13075 );
nor ( n13077 , n13076 , n1339 );
or ( n13078 , n13073 , n13077 );
nand ( n13079 , n13078 , n177 );
and ( n13080 , n13067 , n13071 , n13079 );
nand ( n13081 , n13060 , n13080 );
not ( n13082 , n13081 );
and ( n13083 , n12987 , n13082 );
not ( n13084 , n12987 );
and ( n13085 , n13084 , n13081 );
nor ( n13086 , n13083 , n13085 );
xor ( n13087 , n12895 , n13086 );
and ( n13088 , n12889 , n13087 );
not ( n13089 , n12889 );
not ( n13090 , n13087 );
and ( n13091 , n13089 , n13090 );
nor ( n13092 , n13088 , n13091 );
or ( n13093 , n13092 , n1 );
xnor ( n13094 , n334 , n335 );
or ( n13095 , n2246 , n13094 );
nand ( n13096 , n13093 , n13095 );
not ( n13097 , n200 );
nor ( n13098 , n13097 , n5703 , n201 );
or ( n13099 , n4132 , n13098 );
nand ( n13100 , n13099 , n202 );
not ( n13101 , n5217 );
nand ( n13102 , n13101 , n4107 );
not ( n13103 , n4026 );
nor ( n13104 , n13103 , n203 );
nand ( n13105 , n5687 , n13100 , n13102 , n13104 );
not ( n13106 , n13105 );
nor ( n13107 , n5739 , n4027 );
not ( n13108 , n4097 );
nor ( n13109 , n13108 , n199 );
or ( n13110 , n13107 , n13109 );
nand ( n13111 , n13110 , n202 );
and ( n13112 , n5211 , n5731 );
nand ( n13113 , n5875 , n203 );
nor ( n13114 , n13112 , n13113 );
nor ( n13115 , n5180 , n5783 );
nand ( n13116 , n13111 , n13114 , n13115 );
not ( n13117 , n13116 );
or ( n13118 , n13106 , n13117 );
not ( n13119 , n5867 );
nand ( n13120 , n13118 , n13119 );
not ( n13121 , n4058 );
nor ( n13122 , n5089 , n202 );
not ( n13123 , n13122 );
not ( n13124 , n4182 );
or ( n13125 , n13123 , n13124 );
nand ( n13126 , n13125 , n4085 );
not ( n13127 , n13126 );
or ( n13128 , n13121 , n13127 );
and ( n13129 , n199 , n4072 );
not ( n13130 , n199 );
and ( n13131 , n13130 , n13108 );
nor ( n13132 , n13129 , n13131 );
nand ( n13133 , n13132 , n5671 );
not ( n13134 , n5189 );
nor ( n13135 , n13134 , n5691 );
nand ( n13136 , n13133 , n13135 );
nand ( n13137 , n13128 , n13136 );
not ( n13138 , n13137 );
nor ( n13139 , n13120 , n13138 );
nand ( n13140 , n3982 , n4126 , n4026 );
and ( n13141 , n13140 , n4160 );
nand ( n13142 , n5092 , n5875 , n5135 );
nand ( n13143 , n4159 , n4141 , n5185 );
and ( n13144 , n13142 , n13143 );
nand ( n13145 , n5178 , n4067 );
nor ( n13146 , n13145 , n4054 );
nand ( n13147 , n4186 , n13146 );
nor ( n13148 , n13144 , n13147 );
nand ( n13149 , n5768 , n4062 , n5724 , n5217 );
not ( n13150 , n4049 );
not ( n13151 , n4120 );
and ( n13152 , n13150 , n13151 );
not ( n13153 , n4009 );
not ( n13154 , n5731 );
or ( n13155 , n13153 , n13154 );
nand ( n13156 , n13155 , n5669 );
nor ( n13157 , n13156 , n4077 );
nor ( n13158 , n13152 , n13157 );
nor ( n13159 , n13149 , n13158 );
or ( n13160 , n13148 , n13159 );
nand ( n13161 , n4158 , n4036 );
nand ( n13162 , n3966 , n201 );
nand ( n13163 , n13161 , n13162 );
or ( n13164 , n13163 , n4207 );
nand ( n13165 , n13164 , n4086 );
not ( n13166 , n4193 );
and ( n13167 , n13166 , n201 );
nor ( n13168 , n13167 , n4058 );
and ( n13169 , n13165 , n13168 );
nand ( n13170 , n13160 , n13169 );
nor ( n13171 , n13141 , n13170 );
or ( n13172 , n13139 , n13171 );
not ( n13173 , n4121 );
not ( n13174 , n5173 );
or ( n13175 , n13173 , n13174 );
nand ( n13176 , n5217 , n4078 );
nand ( n13177 , n13175 , n13176 );
not ( n13178 , n5704 );
not ( n13179 , n13178 );
not ( n13180 , n4033 );
not ( n13181 , n5103 );
or ( n13182 , n13180 , n13181 );
nand ( n13183 , n13182 , n3996 );
nand ( n13184 , n13179 , n13183 );
nand ( n13185 , n13184 , n5125 );
and ( n13186 , n13177 , n13185 );
nand ( n13187 , n13119 , n4068 );
or ( n13188 , n13187 , n5233 );
nand ( n13189 , n5158 , n5213 );
nand ( n13190 , n13188 , n13189 );
nor ( n13191 , n13186 , n13190 );
not ( n13192 , n197 );
not ( n13193 , n5151 );
or ( n13194 , n13192 , n13193 );
nand ( n13195 , n13194 , n4062 );
nand ( n13196 , n13195 , n203 );
not ( n13197 , n13196 );
not ( n13198 , n4199 );
or ( n13199 , n13197 , n13198 );
nand ( n13200 , n13199 , n202 );
not ( n13201 , n4030 );
nand ( n13202 , n13200 , n4208 , n13201 );
nor ( n13203 , n13191 , n13202 );
nand ( n13204 , n13172 , n13203 );
not ( n13205 , n13204 );
not ( n13206 , n13205 );
not ( n13207 , n9599 );
not ( n13208 , n13207 );
or ( n13209 , n13206 , n13208 );
buf ( n13210 , n13204 );
nand ( n13211 , n9599 , n13210 );
nand ( n13212 , n13209 , n13211 );
not ( n13213 , n13212 );
not ( n13214 , n5400 );
or ( n13215 , n13213 , n13214 );
or ( n13216 , n5400 , n13212 );
nand ( n13217 , n13215 , n13216 );
not ( n13218 , n5491 );
not ( n13219 , n11416 );
or ( n13220 , n13218 , n13219 );
nand ( n13221 , n11419 , n5490 );
nand ( n13222 , n13220 , n13221 );
nand ( n13223 , n5617 , n5577 );
nand ( n13224 , n13223 , n5635 );
not ( n13225 , n13224 );
not ( n13226 , n342 );
not ( n13227 , n13226 );
and ( n13228 , n13225 , n13227 );
and ( n13229 , n5636 , n13226 );
nor ( n13230 , n13228 , n13229 );
xor ( n13231 , n13222 , n13230 );
and ( n13232 , n13217 , n13231 );
not ( n13233 , n13217 );
not ( n13234 , n13231 );
and ( n13235 , n13233 , n13234 );
nor ( n13236 , n13232 , n13235 );
or ( n13237 , n13236 , n1 );
and ( n13238 , n343 , n13226 );
not ( n13239 , n343 );
and ( n13240 , n13239 , n342 );
nor ( n13241 , n13238 , n13240 );
or ( n13242 , n2246 , n13241 );
nand ( n13243 , n13237 , n13242 );
not ( n13244 , n9578 );
not ( n13245 , n8510 );
or ( n13246 , n13244 , n13245 );
or ( n13247 , n9578 , n8510 );
nand ( n13248 , n13246 , n13247 );
not ( n13249 , n71 );
xnor ( n13250 , n8894 , n13249 );
and ( n13251 , n9357 , n13250 );
not ( n13252 , n9357 );
not ( n13253 , n13250 );
and ( n13254 , n13252 , n13253 );
nor ( n13255 , n13251 , n13254 );
and ( n13256 , n13248 , n13255 );
not ( n13257 , n13248 );
not ( n13258 , n13255 );
and ( n13259 , n13257 , n13258 );
nor ( n13260 , n13256 , n13259 );
or ( n13261 , n13260 , n1 );
and ( n13262 , n72 , n13249 );
not ( n13263 , n72 );
and ( n13264 , n13263 , n71 );
nor ( n13265 , n13262 , n13264 );
or ( n13266 , n2246 , n13265 );
nand ( n13267 , n13261 , n13266 );
not ( n13268 , n10815 );
nand ( n13269 , n13268 , n1936 );
nand ( n13270 , n1932 , n11780 );
or ( n13271 , n13269 , n13270 );
nand ( n13272 , n13271 , n1979 );
not ( n13273 , n13272 );
not ( n13274 , n10877 );
or ( n13275 , n1882 , n1920 );
nand ( n13276 , n13274 , n10823 , n13275 );
nor ( n13277 , n13276 , n2156 );
not ( n13278 , n13277 );
or ( n13279 , n13273 , n13278 );
nand ( n13280 , n11761 , n2068 );
or ( n13281 , n13280 , n11817 );
nand ( n13282 , n13281 , n1979 );
not ( n13283 , n156 );
not ( n13284 , n2165 );
or ( n13285 , n13283 , n13284 );
or ( n13286 , n11728 , n1855 );
nand ( n13287 , n13285 , n13286 );
or ( n13288 , n13287 , n2147 );
nand ( n13289 , n13288 , n159 );
nor ( n13290 , n12844 , n12137 );
nand ( n13291 , n13282 , n13289 , n13290 );
nand ( n13292 , n13279 , n13291 );
not ( n13293 , n161 );
not ( n13294 , n1959 );
not ( n13295 , n13294 );
not ( n13296 , n2044 );
or ( n13297 , n13295 , n13296 );
nand ( n13298 , n13297 , n1846 );
not ( n13299 , n13298 );
nand ( n13300 , n12827 , n11722 );
not ( n13301 , n13300 );
or ( n13302 , n13299 , n13301 );
nand ( n13303 , n13302 , n10889 );
not ( n13304 , n13303 );
not ( n13305 , n13304 );
not ( n13306 , n1993 );
or ( n13307 , n13305 , n13306 );
and ( n13308 , n1841 , n2084 );
nor ( n13309 , n13308 , n12161 );
nor ( n13310 , n12834 , n13309 );
nand ( n13311 , n2038 , n13310 , n2215 );
nand ( n13312 , n13307 , n13311 );
not ( n13313 , n13312 );
or ( n13314 , n13293 , n13313 );
not ( n13315 , n1899 );
not ( n13316 , n13315 );
or ( n13317 , n1876 , n1834 );
nand ( n13318 , n13317 , n1846 );
or ( n13319 , n13318 , n10805 );
nand ( n13320 , n2186 , n11722 );
or ( n13321 , n13320 , n1967 );
nand ( n13322 , n13319 , n13321 );
not ( n13323 , n13322 );
or ( n13324 , n13316 , n13323 );
nand ( n13325 , n11755 , n1825 );
nand ( n13326 , n2092 , n13325 );
not ( n13327 , n13326 );
nand ( n13328 , n13327 , n2221 );
nand ( n13329 , n13324 , n13328 );
not ( n13330 , n2186 );
nand ( n13331 , n13330 , n155 );
nand ( n13332 , n1905 , n13331 );
and ( n13333 , n13332 , n1906 );
nor ( n13334 , n1953 , n1841 );
or ( n13335 , n12214 , n13334 );
nand ( n13336 , n13335 , n2191 );
nor ( n13337 , n13333 , n13336 );
nand ( n13338 , n13329 , n13337 );
nand ( n13339 , n13314 , n13338 );
and ( n13340 , n1863 , n11780 , n11756 , n12873 );
not ( n13341 , n1825 );
not ( n13342 , n1834 );
or ( n13343 , n13341 , n13342 );
not ( n13344 , n1915 );
nand ( n13345 , n13343 , n13344 );
not ( n13346 , n10818 );
not ( n13347 , n2067 );
or ( n13348 , n13346 , n13347 );
nand ( n13349 , n13348 , n159 );
nor ( n13350 , n13345 , n13349 );
and ( n13351 , n13350 , n1936 );
nor ( n13352 , n13340 , n13351 );
nand ( n13353 , n13338 , n13352 );
not ( n13354 , n1977 );
and ( n13355 , n13354 , n1892 );
and ( n13356 , n1921 , n2117 );
nor ( n13357 , n13355 , n13356 );
nand ( n13358 , n13292 , n13339 , n13353 , n13357 );
not ( n13359 , n13358 );
not ( n13360 , n13359 );
not ( n13361 , n386 );
or ( n13362 , n13360 , n13361 );
or ( n13363 , n13359 , n386 );
nand ( n13364 , n13362 , n13363 );
not ( n13365 , n1543 );
not ( n13366 , n1800 );
or ( n13367 , n13365 , n13366 );
nand ( n13368 , n1799 , n1542 );
nand ( n13369 , n13367 , n13368 );
not ( n13370 , n13369 );
and ( n13371 , n13364 , n13370 );
not ( n13372 , n13364 );
and ( n13373 , n13372 , n13369 );
nor ( n13374 , n13371 , n13373 );
nand ( n13375 , n13374 , n2246 );
not ( n13376 , n10447 );
not ( n13377 , n1417 );
and ( n13378 , n13376 , n13377 );
not ( n13379 , n178 );
not ( n13380 , n11976 );
not ( n13381 , n10361 );
or ( n13382 , n13380 , n13381 );
nand ( n13383 , n13382 , n1459 );
nand ( n13384 , n1343 , n10478 );
not ( n13385 , n13384 );
not ( n13386 , n10442 );
or ( n13387 , n13385 , n13386 );
nand ( n13388 , n13387 , n1280 );
nand ( n13389 , n13379 , n13383 , n13388 );
nor ( n13390 , n13378 , n13389 );
not ( n13391 , n1428 );
not ( n13392 , n13036 );
or ( n13393 , n13391 , n13392 );
nand ( n13394 , n13393 , n1280 );
nand ( n13395 , n13390 , n13394 );
nand ( n13396 , n1304 , n1459 );
nand ( n13397 , n13396 , n1366 , n10523 , n1384 );
or ( n13398 , n13395 , n13397 );
not ( n13399 , n1456 );
nand ( n13400 , n1453 , n1338 );
not ( n13401 , n13400 );
or ( n13402 , n13399 , n13401 );
nand ( n13403 , n13402 , n177 );
not ( n13404 , n11892 );
not ( n13405 , n1440 );
nand ( n13406 , n13405 , n1438 );
not ( n13407 , n13019 );
and ( n13408 , n10403 , n13406 , n13407 );
not ( n13409 , n13408 );
or ( n13410 , n13404 , n13409 );
nor ( n13411 , n1350 , n176 );
nand ( n13412 , n1432 , n13411 );
nand ( n13413 , n13410 , n13412 );
nand ( n13414 , n13403 , n13413 );
nand ( n13415 , n13075 , n1313 );
not ( n13416 , n13415 );
not ( n13417 , n13416 );
not ( n13418 , n1500 );
or ( n13419 , n13417 , n13418 );
nand ( n13420 , n13419 , n1435 );
nor ( n13421 , n1487 , n1417 );
nor ( n13422 , n10479 , n1412 );
nor ( n13423 , n13421 , n13422 );
nand ( n13424 , n13420 , n13423 );
nor ( n13425 , n13414 , n13424 );
nor ( n13426 , n13012 , n1280 );
nor ( n13427 , n1515 , n13426 );
not ( n13428 , n1357 );
not ( n13429 , n1523 );
or ( n13430 , n13428 , n13429 );
nand ( n13431 , n13430 , n10500 );
nor ( n13432 , n10384 , n11970 );
or ( n13433 , n13431 , n13432 );
nand ( n13434 , n13433 , n1280 );
and ( n13435 , n13427 , n13434 , n1432 );
nand ( n13436 , n13425 , n13435 );
nand ( n13437 , n13398 , n13436 );
not ( n13438 , n13437 );
nand ( n13439 , n1476 , n1298 );
nand ( n13440 , n13439 , n10447 , n1456 );
not ( n13441 , n13440 );
not ( n13442 , n10419 );
or ( n13443 , n13441 , n13442 );
not ( n13444 , n1315 );
not ( n13445 , n1323 );
not ( n13446 , n13445 );
or ( n13447 , n13444 , n13446 );
nand ( n13448 , n13447 , n11903 );
nand ( n13449 , n13448 , n1280 );
nand ( n13450 , n13443 , n13449 );
and ( n13451 , n13004 , n1370 );
nand ( n13452 , n1284 , n1473 );
nand ( n13453 , n13388 , n13451 , n13452 );
nor ( n13454 , n13450 , n13453 );
not ( n13455 , n13454 );
or ( n13456 , n13438 , n13455 );
not ( n13457 , n10364 );
not ( n13458 , n13457 );
not ( n13459 , n11991 );
not ( n13460 , n10524 );
or ( n13461 , n13459 , n13460 );
nand ( n13462 , n13461 , n1280 );
nand ( n13463 , n1336 , n1306 );
nand ( n13464 , n13458 , n13462 , n13463 , n10508 );
or ( n13465 , n13395 , n13464 );
not ( n13466 , n13425 );
nand ( n13467 , n13465 , n13466 );
not ( n13468 , n171 );
not ( n13469 , n13415 );
or ( n13470 , n13468 , n13469 );
nand ( n13471 , n13470 , n11971 );
nand ( n13472 , n13471 , n1306 );
not ( n13473 , n11970 );
not ( n13474 , n1382 );
or ( n13475 , n13473 , n13474 );
nand ( n13476 , n13475 , n1533 );
or ( n13477 , n13476 , n1470 );
nand ( n13478 , n13477 , n1473 );
not ( n13479 , n10355 );
not ( n13480 , n10428 );
or ( n13481 , n13479 , n13480 );
nand ( n13482 , n13481 , n176 );
nand ( n13483 , n13472 , n13478 , n13482 , n177 );
nor ( n13484 , n13483 , n13450 );
nand ( n13485 , n13467 , n13484 );
nand ( n13486 , n13456 , n13485 );
buf ( n13487 , n13486 );
not ( n13488 , n13487 );
not ( n13489 , n13488 );
not ( n13490 , n13082 );
not ( n13491 , n1156 );
or ( n13492 , n13490 , n13491 );
nand ( n13493 , n1155 , n13081 );
nand ( n13494 , n13492 , n13493 );
not ( n13495 , n13494 );
or ( n13496 , n13489 , n13495 );
or ( n13497 , n13488 , n13494 );
nand ( n13498 , n13496 , n13497 );
or ( n13499 , n13375 , n13498 );
xnor ( n13500 , n386 , n387 );
or ( n13501 , n13500 , n2246 );
nor ( n13502 , n13374 , n1 );
nand ( n13503 , n13498 , n13502 );
nand ( n13504 , n13499 , n13501 , n13503 );
not ( n13505 , n11577 );
not ( n13506 , n1723 );
nand ( n13507 , n13506 , n1784 );
nand ( n13508 , n12109 , n13507 );
and ( n13509 , n13508 , n149 );
nand ( n13510 , n1740 , n11592 , n11012 );
nor ( n13511 , n13509 , n13510 );
not ( n13512 , n13511 );
nand ( n13513 , n1716 , n10929 );
or ( n13514 , n13513 , n149 );
or ( n13515 , n10933 , n1635 );
nand ( n13516 , n13514 , n13515 );
nor ( n13517 , n12014 , n153 );
nand ( n13518 , n13516 , n13517 );
nor ( n13519 , n10950 , n149 );
nor ( n13520 , n13518 , n13519 );
not ( n13521 , n13520 );
or ( n13522 , n13512 , n13521 );
and ( n13523 , n12027 , n12093 );
nand ( n13524 , n11664 , n1669 );
or ( n13525 , n13524 , n1772 );
not ( n13526 , n1601 );
nand ( n13527 , n13525 , n13526 );
nand ( n13528 , n11003 , n153 );
nand ( n13529 , n1754 , n1615 );
nand ( n13530 , n1774 , n150 );
nand ( n13531 , n13529 , n13530 );
or ( n13532 , n13528 , n13531 );
nand ( n13533 , n13532 , n1579 );
nor ( n13534 , n1722 , n11571 , n1586 , n10964 );
nand ( n13535 , n13523 , n13527 , n13533 , n13534 );
nand ( n13536 , n13522 , n13535 );
not ( n13537 , n13536 );
not ( n13538 , n10950 );
or ( n13539 , n1598 , n13538 );
nand ( n13540 , n13539 , n1721 );
or ( n13541 , n1707 , n1725 );
nand ( n13542 , n13541 , n1621 );
or ( n13543 , n13542 , n12104 );
not ( n13544 , n1712 );
nand ( n13545 , n13543 , n13544 );
and ( n13546 , n13540 , n13545 , n12960 );
not ( n13547 , n13546 );
or ( n13548 , n13537 , n13547 );
not ( n13549 , n13529 );
nor ( n13550 , n1767 , n1711 , n1596 );
nor ( n13551 , n13549 , n13550 );
not ( n13552 , n11026 );
nand ( n13553 , n13552 , n1586 );
not ( n13554 , n11464 );
nand ( n13555 , n1723 , n1730 );
nand ( n13556 , n13551 , n13553 , n13554 , n13555 );
nor ( n13557 , n13518 , n13556 );
nand ( n13558 , n13523 , n13533 );
not ( n13559 , n1654 );
not ( n13560 , n1780 );
or ( n13561 , n13559 , n13560 );
not ( n13562 , n1711 );
nand ( n13563 , n13562 , n1696 , n12011 , n11592 );
nand ( n13564 , n13561 , n13563 );
not ( n13565 , n1764 );
nand ( n13566 , n11554 , n1788 );
nor ( n13567 , n13565 , n13566 );
nand ( n13568 , n13564 , n13567 );
nor ( n13569 , n13558 , n13568 );
or ( n13570 , n13557 , n13569 );
nand ( n13571 , n13570 , n1752 );
nand ( n13572 , n13548 , n13571 );
or ( n13573 , n11000 , n13566 );
or ( n13574 , n12971 , n1656 );
nand ( n13575 , n13573 , n13574 );
and ( n13576 , n13575 , n1752 );
not ( n13577 , n10969 );
not ( n13578 , n11563 );
not ( n13579 , n11629 );
or ( n13580 , n13578 , n13579 );
nand ( n13581 , n13580 , n1660 );
nand ( n13582 , n13577 , n13581 );
nor ( n13583 , n13576 , n13582 );
nand ( n13584 , n13572 , n13583 );
not ( n13585 , n13584 );
not ( n13586 , n13585 );
or ( n13587 , n13505 , n13586 );
nand ( n13588 , n13584 , n12893 );
nand ( n13589 , n13587 , n13588 );
xor ( n13590 , n1547 , n13589 );
xor ( n13591 , n390 , n13359 );
and ( n13592 , n13591 , n2234 );
not ( n13593 , n13591 );
and ( n13594 , n13593 , n2235 );
nor ( n13595 , n13592 , n13594 );
xnor ( n13596 , n13590 , n13595 );
or ( n13597 , n13596 , n1 );
xnor ( n13598 , n390 , n391 );
or ( n13599 , n2246 , n13598 );
nand ( n13600 , n13597 , n13599 );
not ( n13601 , n13486 );
and ( n13602 , n1271 , n13601 );
not ( n13603 , n1271 );
and ( n13604 , n13603 , n13487 );
nor ( n13605 , n13602 , n13604 );
not ( n13606 , n13081 );
not ( n13607 , n13584 );
not ( n13608 , n13607 );
or ( n13609 , n13606 , n13608 );
not ( n13610 , n13081 );
nand ( n13611 , n13610 , n13584 );
nand ( n13612 , n13609 , n13611 );
xor ( n13613 , n13605 , n13612 );
xor ( n13614 , n13359 , n1800 );
not ( n13615 , n286 );
and ( n13616 , n13615 , n12893 );
not ( n13617 , n13615 );
and ( n13618 , n13617 , n11577 );
nor ( n13619 , n13616 , n13618 );
not ( n13620 , n13619 );
and ( n13621 , n13614 , n13620 );
not ( n13622 , n13614 );
and ( n13623 , n13622 , n13619 );
nor ( n13624 , n13621 , n13623 );
xor ( n13625 , n13613 , n13624 );
or ( n13626 , n13625 , n1 );
and ( n13627 , n287 , n13615 );
not ( n13628 , n287 );
and ( n13629 , n13628 , n286 );
nor ( n13630 , n13627 , n13629 );
or ( n13631 , n2246 , n13630 );
nand ( n13632 , n13626 , n13631 );
and ( n13633 , n7926 , n8221 , n6807 );
not ( n13634 , n13633 );
nor ( n13635 , n7997 , n6943 );
not ( n13636 , n13635 );
not ( n13637 , n32 );
nand ( n13638 , n6724 , n7885 , n6787 );
nand ( n13639 , n13637 , n13638 );
not ( n13640 , n13639 );
or ( n13641 , n13636 , n13640 );
not ( n13642 , n7859 );
nand ( n13643 , n13641 , n13642 );
not ( n13644 , n13643 );
or ( n13645 , n13634 , n13644 );
not ( n13646 , n8321 );
not ( n13647 , n7870 );
not ( n13648 , n8694 );
or ( n13649 , n13647 , n13648 );
nand ( n13650 , n13649 , n33 );
nor ( n13651 , n13646 , n8323 , n13650 );
nand ( n13652 , n13639 , n13651 , n8748 );
nand ( n13653 , n13645 , n13652 );
nand ( n13654 , n6908 , n8649 , n8929 );
and ( n13655 , n13654 , n8141 );
nor ( n13656 , n13655 , n8178 );
or ( n13657 , n6825 , n8698 );
nand ( n13658 , n13657 , n6912 );
nand ( n13659 , n7933 , n6782 );
and ( n13660 , n13656 , n13658 , n13659 );
nand ( n13661 , n13653 , n13660 );
not ( n13662 , n13661 );
and ( n13663 , n31 , n8292 );
not ( n13664 , n31 );
and ( n13665 , n13664 , n7953 );
nor ( n13666 , n13663 , n13665 );
or ( n13667 , n8949 , n13666 , n32 );
nand ( n13668 , n6944 , n6873 , n32 );
nand ( n13669 , n13667 , n13668 );
not ( n13670 , n13669 );
and ( n13671 , n31 , n8655 );
not ( n13672 , n31 );
and ( n13673 , n13672 , n6776 );
nor ( n13674 , n13671 , n13673 );
nor ( n13675 , n8658 , n13674 , n8154 , n8253 );
not ( n13676 , n13675 );
or ( n13677 , n13670 , n13676 );
not ( n13678 , n8289 );
not ( n13679 , n13678 );
not ( n13680 , n6887 );
or ( n13681 , n13679 , n13680 );
nand ( n13682 , n13681 , n6719 );
not ( n13683 , n8649 );
nand ( n13684 , n13683 , n6828 );
and ( n13685 , n8208 , n13684 , n6807 );
nand ( n13686 , n13682 , n13685 );
nand ( n13687 , n13677 , n13686 );
not ( n13688 , n8655 );
and ( n13689 , n13688 , n31 );
not ( n13690 , n6819 );
nor ( n13691 , n13689 , n13690 );
not ( n13692 , n13691 );
or ( n13693 , n8377 , n8196 );
nand ( n13694 , n13693 , n8158 );
not ( n13695 , n13694 );
or ( n13696 , n13692 , n13695 );
nand ( n13697 , n13696 , n32 );
not ( n13698 , n6882 );
not ( n13699 , n8146 );
or ( n13700 , n13698 , n13699 );
nor ( n13701 , n6820 , n34 );
nand ( n13702 , n13700 , n13701 );
nor ( n13703 , n8932 , n13702 );
nand ( n13704 , n13697 , n13703 );
not ( n13705 , n13704 );
nand ( n13706 , n13687 , n13705 );
not ( n13707 , n13706 );
or ( n13708 , n13662 , n13707 );
not ( n13709 , n8221 );
not ( n13710 , n8173 );
or ( n13711 , n13709 , n13710 );
nand ( n13712 , n13711 , n6912 );
and ( n13713 , n8369 , n6779 );
nor ( n13714 , n13713 , n8161 );
and ( n13715 , n13712 , n13714 );
nor ( n13716 , n13715 , n33 );
nand ( n13717 , n7932 , n8690 );
or ( n13718 , n13717 , n7875 );
nand ( n13719 , n13718 , n8140 );
nand ( n13720 , n13719 , n7961 , n7872 );
not ( n13721 , n13720 );
and ( n13722 , n8387 , n6899 );
not ( n13723 , n13722 );
or ( n13724 , n13721 , n13723 );
nand ( n13725 , n8731 , n33 );
nand ( n13726 , n8933 , n8141 );
and ( n13727 , n13725 , n8370 , n13726 );
nand ( n13728 , n13724 , n13727 );
nor ( n13729 , n13716 , n13728 );
nand ( n13730 , n13708 , n13729 );
not ( n13731 , n13730 );
not ( n13732 , n13731 );
not ( n13733 , n6688 );
nor ( n13734 , n6542 , n6314 );
nor ( n13735 , n13733 , n6385 , n13734 , n26 );
and ( n13736 , n6637 , n6399 );
and ( n13737 , n6640 , n13736 , n6404 );
nor ( n13738 , n6473 , n6299 );
not ( n13739 , n13738 );
not ( n13740 , n6520 );
or ( n13741 , n13739 , n13740 );
not ( n13742 , n6608 );
nand ( n13743 , n13742 , n6468 , n8045 , n6299 );
nand ( n13744 , n13741 , n13743 );
nand ( n13745 , n13737 , n13744 );
nor ( n13746 , n13745 , n9528 );
or ( n13747 , n13735 , n13746 );
not ( n13748 , n23 );
not ( n13749 , n6492 );
or ( n13750 , n13748 , n13749 );
not ( n13751 , n6313 );
nand ( n13752 , n13750 , n13751 );
or ( n13753 , n13752 , n8410 );
nand ( n13754 , n13753 , n25 );
nand ( n13755 , n6291 , n6299 );
and ( n13756 , n6421 , n6539 );
and ( n13757 , n13754 , n13755 , n13756 , n6464 );
nand ( n13758 , n13747 , n13757 );
not ( n13759 , n13758 );
not ( n13760 , n6579 );
nor ( n13761 , n13760 , n6562 );
not ( n13762 , n13761 );
nor ( n13763 , n9484 , n13762 );
or ( n13764 , n13763 , n25 );
not ( n13765 , n8052 );
not ( n13766 , n9560 );
or ( n13767 , n13765 , n13766 );
nand ( n13768 , n13767 , n6417 );
nand ( n13769 , n13764 , n13768 );
not ( n13770 , n9484 );
not ( n13771 , n6451 );
nor ( n13772 , n13771 , n25 );
and ( n13773 , n13761 , n6353 , n13772 );
nand ( n13774 , n13770 , n13773 , n6542 );
nand ( n13775 , n13769 , n13774 );
nor ( n13776 , n9538 , n24 );
nor ( n13777 , n6494 , n6518 );
or ( n13778 , n13776 , n13777 , n9559 );
nand ( n13779 , n13778 , n6447 );
not ( n13780 , n8109 );
not ( n13781 , n6483 );
not ( n13782 , n8471 );
nor ( n13783 , n13782 , n6430 );
nor ( n13784 , n13781 , n8478 , n13783 );
not ( n13785 , n13784 );
or ( n13786 , n13780 , n13785 );
nand ( n13787 , n13786 , n26 );
nand ( n13788 , n6342 , n6330 );
and ( n13789 , n13788 , n12378 );
nor ( n13790 , n13789 , n6448 );
nor ( n13791 , n8099 , n13790 );
nand ( n13792 , n13775 , n13779 , n13787 , n13791 );
not ( n13793 , n13792 );
or ( n13794 , n13759 , n13793 );
nand ( n13795 , n8102 , n6343 );
and ( n13796 , n6606 , n6428 );
nor ( n13797 , n13796 , n6546 );
not ( n13798 , n13797 );
nand ( n13799 , n6498 , n6356 );
not ( n13800 , n13799 );
not ( n13801 , n13800 );
or ( n13802 , n13798 , n13801 );
nand ( n13803 , n13802 , n9561 );
nor ( n13804 , n6477 , n6287 );
nand ( n13805 , n13799 , n13804 );
nand ( n13806 , n13795 , n13803 , n13805 , n8092 );
and ( n13807 , n6447 , n13806 );
not ( n13808 , n6637 );
nand ( n13809 , n13808 , n6348 );
nand ( n13810 , n13755 , n13809 );
nor ( n13811 , n8469 , n6375 );
or ( n13812 , n13810 , n13811 );
nand ( n13813 , n13812 , n26 );
or ( n13814 , n8437 , n12405 );
nand ( n13815 , n13814 , n8430 );
nand ( n13816 , n13813 , n13815 );
nor ( n13817 , n13807 , n13816 );
nand ( n13818 , n13794 , n13817 );
not ( n13819 , n13818 );
not ( n13820 , n13819 );
or ( n13821 , n13732 , n13820 );
nand ( n13822 , n13818 , n13730 );
nand ( n13823 , n13821 , n13822 );
not ( n13824 , n9123 );
not ( n13825 , n7224 );
not ( n13826 , n39 );
and ( n13827 , n13825 , n13826 );
and ( n13828 , n7224 , n39 );
nor ( n13829 , n13827 , n13828 );
not ( n13830 , n13829 );
and ( n13831 , n13824 , n13830 );
and ( n13832 , n9123 , n13829 );
nor ( n13833 , n13831 , n13832 );
and ( n13834 , n13823 , n13833 );
not ( n13835 , n13823 );
not ( n13836 , n13833 );
and ( n13837 , n13835 , n13836 );
nor ( n13838 , n13834 , n13837 );
or ( n13839 , n13838 , n1 );
not ( n13840 , n38 );
not ( n13841 , n39 );
and ( n13842 , n13840 , n13841 );
and ( n13843 , n38 , n39 );
nor ( n13844 , n13842 , n13843 );
or ( n13845 , n2246 , n13844 );
nand ( n13846 , n13839 , n13845 );
nand ( n13847 , n7143 , n6985 );
nand ( n13848 , n7197 , n7036 );
or ( n13849 , n13847 , n13848 );
nand ( n13850 , n13849 , n7170 );
not ( n13851 , n7530 );
not ( n13852 , n9151 );
or ( n13853 , n13851 , n13852 );
nand ( n13854 , n13853 , n16 );
not ( n13855 , n7605 );
not ( n13856 , n7644 );
and ( n13857 , n13855 , n13856 );
not ( n13858 , n9320 );
nor ( n13859 , n13857 , n13858 );
and ( n13860 , n13854 , n13859 );
nand ( n13861 , n7009 , n7018 );
nand ( n13862 , n13850 , n13860 , n13861 );
and ( n13863 , n13862 , n6978 );
not ( n13864 , n7545 );
and ( n13865 , n8543 , n13864 );
nand ( n13866 , n7517 , n7206 );
and ( n13867 , n13866 , n7552 );
nor ( n13868 , n13865 , n13867 );
not ( n13869 , n8604 );
nand ( n13870 , n13869 , n7026 , n7048 );
not ( n13871 , n13870 );
or ( n13872 , n7615 , n7080 );
nand ( n13873 , n13872 , n7108 );
not ( n13874 , n7193 );
and ( n13875 , n13874 , n7009 , n14 );
nor ( n13876 , n13873 , n13875 );
not ( n13877 , n13876 );
or ( n13878 , n13871 , n13877 );
nand ( n13879 , n13878 , n17 );
nand ( n13880 , n13868 , n13879 );
nor ( n13881 , n13863 , n13880 );
not ( n13882 , n9182 );
nand ( n13883 , n13882 , n8532 );
not ( n13884 , n13883 );
not ( n13885 , n9341 );
not ( n13886 , n13885 );
or ( n13887 , n13884 , n13886 );
not ( n13888 , n16 );
nand ( n13889 , n13887 , n13888 );
not ( n13890 , n13889 );
and ( n13891 , n7015 , n16 );
nor ( n13892 , n13891 , n7131 );
not ( n13893 , n13892 );
or ( n13894 , n13890 , n13893 );
nor ( n13895 , n9302 , n7587 );
not ( n13896 , n9184 );
not ( n13897 , n7205 );
or ( n13898 , n13896 , n13897 );
nand ( n13899 , n13898 , n16 );
nand ( n13900 , n7162 , n6976 );
nand ( n13901 , n13900 , n7206 );
nand ( n13902 , n13901 , n7170 );
nand ( n13903 , n13895 , n13899 , n7143 , n13902 );
nand ( n13904 , n13894 , n13903 );
not ( n13905 , n8559 );
not ( n13906 , n7003 );
nor ( n13907 , n8520 , n7155 );
not ( n13908 , n13907 );
or ( n13909 , n13906 , n13908 );
nand ( n13910 , n13909 , n7009 );
not ( n13911 , n7518 );
and ( n13912 , n13910 , n13911 , n10 );
nand ( n13913 , n13904 , n13905 , n7537 , n13912 );
not ( n13914 , n7650 );
not ( n13915 , n7023 );
or ( n13916 , n13914 , n13915 );
nand ( n13917 , n13916 , n16 );
not ( n13918 , n13917 );
not ( n13919 , n8546 );
nor ( n13920 , n8588 , n13919 , n16 );
not ( n13921 , n9165 );
nor ( n13922 , n13920 , n13921 );
not ( n13923 , n13922 );
or ( n13924 , n13918 , n13923 );
or ( n13925 , n7038 , n8546 );
nand ( n13926 , n13925 , n9151 , n6978 );
nand ( n13927 , n13924 , n13926 );
not ( n13928 , n7039 );
not ( n13929 , n7206 );
and ( n13930 , n13929 , n7009 );
nor ( n13931 , n13930 , n6992 , n10 );
nand ( n13932 , n13927 , n13928 , n13931 );
nand ( n13933 , n13913 , n13932 );
or ( n13934 , n7106 , n12 );
nand ( n13935 , n13934 , n7036 );
nand ( n13936 , n13935 , n7052 );
nand ( n13937 , n13881 , n13933 , n13936 );
not ( n13938 , n13937 );
not ( n13939 , n13938 );
not ( n13940 , n9221 );
and ( n13941 , n13939 , n13940 );
and ( n13942 , n13938 , n9221 );
nor ( n13943 , n13941 , n13942 );
not ( n13944 , n13943 );
not ( n13945 , n65 );
buf ( n13946 , n12342 );
not ( n13947 , n13946 );
or ( n13948 , n13945 , n13947 );
or ( n13949 , n65 , n13946 );
nand ( n13950 , n13948 , n13949 );
not ( n13951 , n13950 );
or ( n13952 , n13944 , n13951 );
or ( n13953 , n13943 , n13950 );
nand ( n13954 , n13952 , n13953 );
nand ( n13955 , n13954 , n2246 );
not ( n13956 , n8917 );
not ( n13957 , n13956 );
nand ( n13958 , n6288 , n6588 , n8491 );
and ( n13959 , n13958 , n6315 );
nand ( n13960 , n6519 , n6384 );
nand ( n13961 , n8433 , n13960 , n8425 );
nor ( n13962 , n13959 , n13961 );
nand ( n13963 , n6604 , n6447 );
not ( n13964 , n8461 );
nor ( n13965 , n13963 , n13964 );
or ( n13966 , n6378 , n6546 );
nand ( n13967 , n13966 , n6356 );
and ( n13968 , n6284 , n6526 , n25 );
nor ( n13969 , n12356 , n13968 );
nand ( n13970 , n13965 , n13967 , n13969 , n6441 );
not ( n13971 , n8038 );
and ( n13972 , n6426 , n13971 , n26 );
nand ( n13973 , n8098 , n13972 , n6299 );
nand ( n13974 , n13751 , n6340 );
nand ( n13975 , n13970 , n13973 , n13974 );
nand ( n13976 , n13962 , n13975 );
and ( n13977 , n19 , n13976 );
not ( n13978 , n19 );
not ( n13979 , n6632 );
not ( n13980 , n6357 );
or ( n13981 , n13979 , n13980 );
nand ( n13982 , n13981 , n6292 );
not ( n13983 , n13982 );
not ( n13984 , n6340 );
not ( n13985 , n8454 );
or ( n13986 , n13984 , n13985 );
nand ( n13987 , n6491 , n8061 , n26 );
or ( n13988 , n8084 , n13987 );
nand ( n13989 , n13986 , n13988 );
not ( n13990 , n13989 );
not ( n13991 , n6298 );
or ( n13992 , n13990 , n13991 );
not ( n13993 , n6482 );
or ( n13994 , n13993 , n6454 );
nand ( n13995 , n13994 , n6650 , n6447 );
nand ( n13996 , n13992 , n13995 );
nand ( n13997 , n13983 , n13996 );
and ( n13998 , n13978 , n13997 );
nor ( n13999 , n13977 , n13998 );
and ( n14000 , n9563 , n22 );
not ( n14001 , n6693 );
nor ( n14002 , n14000 , n14001 );
not ( n14003 , n14002 );
not ( n14004 , n9527 );
or ( n14005 , n14003 , n14004 );
nand ( n14006 , n14005 , n6356 );
not ( n14007 , n6621 );
nand ( n14008 , n14007 , n6543 );
and ( n14009 , n6606 , n21 );
nor ( n14010 , n14009 , n6546 );
nand ( n14011 , n14008 , n14010 );
nand ( n14012 , n14011 , n12405 );
nand ( n14013 , n14006 , n14012 , n26 );
not ( n14014 , n6330 );
and ( n14015 , n6440 , n14014 );
nor ( n14016 , n14015 , n6332 );
nand ( n14017 , n13800 , n14016 );
not ( n14018 , n14017 );
nor ( n14019 , n6308 , n6535 );
or ( n14020 , n14019 , n6384 );
nand ( n14021 , n14020 , n6650 );
not ( n14022 , n14021 );
or ( n14023 , n14018 , n14022 );
not ( n14024 , n13971 );
nand ( n14025 , n14024 , n23 );
and ( n14026 , n14025 , n8476 , n6447 );
nand ( n14027 , n14023 , n14026 );
and ( n14028 , n14013 , n14027 );
not ( n14029 , n6656 );
not ( n14030 , n8425 );
or ( n14031 , n14029 , n14030 );
nand ( n14032 , n14031 , n25 );
nand ( n14033 , n8047 , n14032 );
nor ( n14034 , n14028 , n14033 );
nand ( n14035 , n13999 , n14034 );
not ( n14036 , n14035 );
and ( n14037 , n13957 , n14036 );
not ( n14038 , n14035 );
not ( n14039 , n14038 );
and ( n14040 , n8918 , n14039 );
nor ( n14041 , n14037 , n14040 );
not ( n14042 , n14041 );
xor ( n14043 , n8264 , n8127 );
buf ( n14044 , n14043 );
not ( n14045 , n14044 );
or ( n14046 , n14042 , n14045 );
or ( n14047 , n14044 , n14041 );
nand ( n14048 , n14046 , n14047 );
or ( n14049 , n13955 , n14048 );
xnor ( n14050 , n65 , n66 );
or ( n14051 , n14050 , n2246 );
not ( n14052 , n13954 );
nand ( n14053 , n14048 , n14052 , n2246 );
nand ( n14054 , n14049 , n14051 , n14053 );
nand ( n14055 , n7887 , n8188 );
nor ( n14056 , n14055 , n13717 );
or ( n14057 , n14056 , n6882 );
and ( n14058 , n7872 , n33 );
nand ( n14059 , n14057 , n14058 );
not ( n14060 , n8674 );
nor ( n14061 , n8646 , n6706 );
not ( n14062 , n14061 );
and ( n14063 , n14060 , n14062 );
nor ( n14064 , n14063 , n32 );
or ( n14065 , n14059 , n14064 );
not ( n14066 , n6779 );
nand ( n14067 , n14066 , n7849 );
not ( n14068 , n14067 );
not ( n14069 , n6704 );
or ( n14070 , n14068 , n14069 );
nand ( n14071 , n14070 , n6807 );
not ( n14072 , n14071 );
not ( n14073 , n7960 );
nand ( n14074 , n6838 , n8993 , n14073 );
or ( n14075 , n8923 , n14074 );
nand ( n14076 , n7871 , n8369 , n8148 );
nand ( n14077 , n14075 , n14076 );
nand ( n14078 , n14072 , n14077 );
nand ( n14079 , n14065 , n14078 );
not ( n14080 , n8252 );
and ( n14081 , n14073 , n8682 );
not ( n14082 , n6912 );
nor ( n14083 , n14081 , n14082 );
nor ( n14084 , n14080 , n14083 );
nand ( n14085 , n14079 , n14084 );
not ( n14086 , n14085 );
and ( n14087 , n8169 , n6817 , n6791 );
nor ( n14088 , n14087 , n6827 );
not ( n14089 , n32 );
not ( n14090 , n8315 );
not ( n14091 , n14090 );
or ( n14092 , n14089 , n14091 );
nor ( n14093 , n7862 , n7879 , n6812 );
nand ( n14094 , n14092 , n14093 );
nor ( n14095 , n14088 , n14094 );
not ( n14096 , n14095 );
nand ( n14097 , n7838 , n7899 );
nand ( n14098 , n6903 , n6912 );
and ( n14099 , n8922 , n14098 );
nand ( n14100 , n8298 , n7974 );
nor ( n14101 , n7963 , n14100 );
nand ( n14102 , n14097 , n14099 , n14101 , n13659 );
nand ( n14103 , n8706 , n6924 );
or ( n14104 , n14103 , n8140 );
or ( n14105 , n13690 , n6868 );
nand ( n14106 , n14104 , n14105 );
nand ( n14107 , n14106 , n8373 );
nand ( n14108 , n14102 , n14107 );
not ( n14109 , n14108 );
or ( n14110 , n14096 , n14109 );
not ( n14111 , n8653 );
nand ( n14112 , n6902 , n8195 , n8683 );
not ( n14113 , n14112 );
or ( n14114 , n14111 , n14113 );
not ( n14115 , n8302 );
not ( n14116 , n6858 );
or ( n14117 , n14115 , n14116 );
and ( n14118 , n6848 , n33 );
nand ( n14119 , n14117 , n14118 );
not ( n14120 , n14119 );
nand ( n14121 , n14114 , n14120 );
not ( n14122 , n8199 );
or ( n14123 , n6750 , n14122 );
nand ( n14124 , n14123 , n8148 , n6807 );
nand ( n14125 , n14121 , n14124 );
not ( n14126 , n8667 );
not ( n14127 , n7961 );
or ( n14128 , n14126 , n14127 );
nand ( n14129 , n14128 , n8692 );
nor ( n14130 , n8933 , n34 );
nand ( n14131 , n14125 , n14129 , n14130 );
nand ( n14132 , n14110 , n14131 );
nand ( n14133 , n14086 , n14132 );
not ( n14134 , n14133 );
not ( n14135 , n14134 );
nand ( n14136 , n13999 , n14034 );
not ( n14137 , n14136 );
not ( n14138 , n14137 );
and ( n14139 , n14135 , n14138 );
and ( n14140 , n14134 , n14137 );
nor ( n14141 , n14139 , n14140 );
not ( n14142 , n14141 );
not ( n14143 , n6963 );
or ( n14144 , n14142 , n14143 );
or ( n14145 , n14141 , n6963 );
nand ( n14146 , n14144 , n14145 );
xor ( n14147 , n67 , n8263 );
not ( n14148 , n7222 );
nand ( n14149 , n7161 , n7170 );
nand ( n14150 , n13874 , n7009 );
nand ( n14151 , n9246 , n14149 , n6973 , n14150 );
not ( n14152 , n14151 );
or ( n14153 , n14148 , n14152 );
not ( n14154 , n7565 );
not ( n14155 , n9246 );
or ( n14156 , n14154 , n14155 );
nand ( n14157 , n14156 , n7132 );
and ( n14158 , n7552 , n6992 );
not ( n14159 , n9157 );
and ( n14160 , n7649 , n7626 );
not ( n14161 , n14160 );
or ( n14162 , n14159 , n14161 );
nand ( n14163 , n14162 , n8557 );
nor ( n14164 , n14158 , n14163 );
not ( n14165 , n7568 );
not ( n14166 , n14165 );
not ( n14167 , n7124 );
or ( n14168 , n14166 , n14167 );
nand ( n14169 , n14168 , n7009 );
and ( n14170 , n14157 , n14164 , n14169 );
nand ( n14171 , n14153 , n14170 );
not ( n14172 , n6979 );
not ( n14173 , n13900 );
nor ( n14174 , n14172 , n7506 , n14173 );
not ( n14175 , n7620 );
nand ( n14176 , n14175 , n7033 );
or ( n14177 , n7153 , n14176 );
nand ( n14178 , n7060 , n7108 , n7170 );
nand ( n14179 , n14177 , n14178 );
nand ( n14180 , n14174 , n14179 );
and ( n14181 , n7185 , n7651 , n17 );
not ( n14182 , n9151 );
not ( n14183 , n11 );
nor ( n14184 , n14183 , n7163 );
and ( n14185 , n14184 , n7636 );
nor ( n14186 , n14185 , n7175 );
not ( n14187 , n14186 );
or ( n14188 , n14182 , n14187 );
nand ( n14189 , n14188 , n9274 );
not ( n14190 , n8591 );
nand ( n14191 , n7657 , n7097 );
nand ( n14192 , n14181 , n14189 , n14190 , n14191 );
nand ( n14193 , n14180 , n14192 , n10 );
nand ( n14194 , n7107 , n7046 );
and ( n14195 , n14194 , n9289 );
nor ( n14196 , n14195 , n16 );
nand ( n14197 , n7134 , n8604 );
or ( n14198 , n14197 , n6996 );
nand ( n14199 , n14198 , n7063 );
nand ( n14200 , n14199 , n13885 );
or ( n14201 , n14196 , n14200 );
nand ( n14202 , n14201 , n10 );
nand ( n14203 , n14193 , n14202 );
nor ( n14204 , n14171 , n14203 );
and ( n14205 , n14194 , n6978 );
or ( n14206 , n8536 , n7063 );
nand ( n14207 , n14206 , n7013 );
and ( n14208 , n7049 , n14205 , n14207 );
not ( n14209 , n7623 );
nand ( n14210 , n14209 , n7073 );
and ( n14211 , n14208 , n14210 );
not ( n14212 , n9208 );
not ( n14213 , n7643 );
or ( n14214 , n14212 , n14213 );
nand ( n14215 , n14214 , n17 );
not ( n14216 , n14215 );
and ( n14217 , n9157 , n8551 );
nor ( n14218 , n14217 , n8541 );
nand ( n14219 , n14216 , n14218 );
not ( n14220 , n7193 );
not ( n14221 , n7116 );
and ( n14222 , n14220 , n14221 );
nor ( n14223 , n6988 , n7058 );
nor ( n14224 , n14222 , n14223 );
nand ( n14225 , n7543 , n14224 );
or ( n14226 , n14219 , n14225 );
nand ( n14227 , n14226 , n7222 );
nor ( n14228 , n14211 , n14227 );
not ( n14229 , n7169 );
not ( n14230 , n8564 );
not ( n14231 , n14230 );
or ( n14232 , n14229 , n14231 );
nand ( n14233 , n14232 , n7009 );
nand ( n14234 , n7026 , n7657 , n7097 );
and ( n14235 , n14233 , n13870 , n14234 );
not ( n14236 , n9201 );
not ( n14237 , n7114 );
or ( n14238 , n14236 , n14237 );
nand ( n14239 , n14238 , n7097 );
and ( n14240 , n14235 , n14239 );
nor ( n14241 , n14240 , n7131 );
nor ( n14242 , n14228 , n14241 );
nand ( n14243 , n14204 , n14242 );
not ( n14244 , n14243 );
xnor ( n14245 , n14147 , n14244 );
buf ( n14246 , n13946 );
and ( n14247 , n14245 , n14246 );
not ( n14248 , n14245 );
not ( n14249 , n13946 );
and ( n14250 , n14248 , n14249 );
nor ( n14251 , n14247 , n14250 );
not ( n14252 , n14251 );
and ( n14253 , n14146 , n14252 );
not ( n14254 , n14146 );
and ( n14255 , n14254 , n14251 );
nor ( n14256 , n14253 , n14255 );
or ( n14257 , n14256 , n1 );
not ( n14258 , n67 );
and ( n14259 , n68 , n14258 );
not ( n14260 , n68 );
and ( n14261 , n14260 , n67 );
nor ( n14262 , n14259 , n14261 );
or ( n14263 , n2246 , n14262 );
nand ( n14264 , n14257 , n14263 );
not ( n14265 , n8132 );
not ( n14266 , n14265 );
not ( n14267 , n8002 );
not ( n14268 , n12432 );
and ( n14269 , n14267 , n14268 );
and ( n14270 , n8002 , n12432 );
nor ( n14271 , n14269 , n14270 );
not ( n14272 , n14271 );
not ( n14273 , n14272 );
or ( n14274 , n14266 , n14273 );
nand ( n14275 , n14271 , n8132 );
nand ( n14276 , n14274 , n14275 );
xor ( n14277 , n86 , n7834 );
xor ( n14278 , n14243 , n9215 );
xnor ( n14279 , n14277 , n14278 );
and ( n14280 , n14276 , n14279 );
not ( n14281 , n14276 );
not ( n14282 , n14279 );
and ( n14283 , n14281 , n14282 );
nor ( n14284 , n14280 , n14283 );
or ( n14285 , n14284 , n1 );
xnor ( n14286 , n86 , n87 );
or ( n14287 , n2246 , n14286 );
nand ( n14288 , n14285 , n14287 );
and ( n14289 , n14244 , n79 );
not ( n14290 , n14244 );
not ( n14291 , n79 );
and ( n14292 , n14290 , n14291 );
nor ( n14293 , n14289 , n14292 );
not ( n14294 , n12342 );
not ( n14295 , n9218 );
or ( n14296 , n14294 , n14295 );
or ( n14297 , n12342 , n9218 );
nand ( n14298 , n14296 , n14297 );
xor ( n14299 , n14293 , n14298 );
not ( n14300 , n8404 );
not ( n14301 , n14300 );
not ( n14302 , n8127 );
not ( n14303 , n14302 );
or ( n14304 , n14301 , n14303 );
not ( n14305 , n8127 );
buf ( n14306 , n8267 );
or ( n14307 , n14305 , n14306 );
nand ( n14308 , n14304 , n14307 );
not ( n14309 , n14134 );
not ( n14310 , n7399 );
nor ( n14311 , n7759 , n7 );
not ( n14312 , n14311 );
or ( n14313 , n14310 , n14312 );
nand ( n14314 , n7 , n7679 , n7256 );
nand ( n14315 , n14313 , n14314 );
nor ( n14316 , n7704 , n7743 );
nand ( n14317 , n14315 , n7793 , n14316 );
not ( n14318 , n7338 );
not ( n14319 , n7828 );
and ( n14320 , n14318 , n14319 );
not ( n14321 , n8889 );
not ( n14322 , n3 );
nand ( n14323 , n14322 , n4 , n5 );
nand ( n14324 , n14321 , n14323 , n7672 );
not ( n14325 , n14324 );
and ( n14326 , n9365 , n14325 );
nor ( n14327 , n14320 , n14326 );
nand ( n14328 , n14317 , n14327 );
nand ( n14329 , n7355 , n7438 );
and ( n14330 , n7795 , n14329 , n7744 , n9 );
not ( n14331 , n8807 );
or ( n14332 , n7448 , n14331 );
nand ( n14333 , n14332 , n7457 );
nand ( n14334 , n14328 , n14330 , n14333 );
not ( n14335 , n7687 );
not ( n14336 , n7 );
and ( n14337 , n14335 , n14336 );
nor ( n14338 , n14337 , n9023 );
not ( n14339 , n7315 );
not ( n14340 , n7322 );
not ( n14341 , n14340 );
or ( n14342 , n14339 , n14341 );
not ( n14343 , n7396 );
and ( n14344 , n14343 , n8 );
nor ( n14345 , n14344 , n9 );
nand ( n14346 , n14342 , n14345 );
nor ( n14347 , n7807 , n8889 );
nor ( n14348 , n14346 , n14347 );
not ( n14349 , n7240 );
not ( n14350 , n7336 );
or ( n14351 , n14349 , n14350 );
nand ( n14352 , n14351 , n7763 );
and ( n14353 , n14352 , n8863 );
and ( n14354 , n7313 , n7 );
nor ( n14355 , n14353 , n14354 );
nand ( n14356 , n7350 , n7279 );
nand ( n14357 , n14338 , n14348 , n14355 , n14356 );
nand ( n14358 , n14334 , n14357 );
and ( n14359 , n7275 , n9457 , n7682 );
nor ( n14360 , n14359 , n8 );
not ( n14361 , n14360 );
nand ( n14362 , n7793 , n7436 , n7265 );
or ( n14363 , n8832 , n14362 );
not ( n14364 , n7251 );
not ( n14365 , n7310 );
or ( n14366 , n14364 , n14365 );
nand ( n14367 , n14366 , n7 );
not ( n14368 , n14367 );
nand ( n14369 , n14368 , n7322 );
or ( n14370 , n8779 , n14369 );
nand ( n14371 , n14363 , n14370 );
not ( n14372 , n14371 );
or ( n14373 , n14361 , n14372 );
nor ( n14374 , n8777 , n7337 );
or ( n14375 , n14374 , n8840 );
nand ( n14376 , n14375 , n7265 );
and ( n14377 , n8822 , n8 );
nand ( n14378 , n14376 , n14377 );
nand ( n14379 , n14373 , n14378 );
not ( n14380 , n12275 );
or ( n14381 , n9367 , n7347 );
nand ( n14382 , n14381 , n7438 );
not ( n14383 , n7473 );
or ( n14384 , n12306 , n12286 );
nand ( n14385 , n14384 , n5 );
not ( n14386 , n14385 );
or ( n14387 , n14383 , n14386 );
nand ( n14388 , n14387 , n8863 );
and ( n14389 , n14380 , n14382 , n14388 );
nand ( n14390 , n14358 , n14379 , n14389 );
not ( n14391 , n14390 );
not ( n14392 , n14391 );
or ( n14393 , n14309 , n14392 );
nand ( n14394 , n14390 , n14133 );
nand ( n14395 , n14393 , n14394 );
not ( n14396 , n14395 );
and ( n14397 , n14308 , n14396 );
not ( n14398 , n14308 );
and ( n14399 , n14398 , n14395 );
nor ( n14400 , n14397 , n14399 );
xnor ( n14401 , n14299 , n14400 );
or ( n14402 , n14401 , n1 );
and ( n14403 , n89 , n14291 );
not ( n14404 , n89 );
and ( n14405 , n14404 , n79 );
nor ( n14406 , n14403 , n14405 );
or ( n14407 , n2246 , n14406 );
nand ( n14408 , n14402 , n14407 );
not ( n14409 , n9218 );
nand ( n14410 , n14358 , n14379 , n14389 );
not ( n14411 , n14410 );
not ( n14412 , n14411 );
and ( n14413 , n14409 , n14412 );
not ( n14414 , n14410 );
and ( n14415 , n7490 , n14414 );
nor ( n14416 , n14413 , n14415 );
xor ( n14417 , n14043 , n14416 );
not ( n14418 , n95 );
and ( n14419 , n14418 , n14244 );
not ( n14420 , n14418 );
not ( n14421 , n14244 );
and ( n14422 , n14420 , n14421 );
or ( n14423 , n14419 , n14422 );
xnor ( n14424 , n14423 , n13943 );
and ( n14425 , n14417 , n14424 );
not ( n14426 , n14417 );
xor ( n14427 , n14423 , n13943 );
and ( n14428 , n14426 , n14427 );
nor ( n14429 , n14425 , n14428 );
or ( n14430 , n14429 , n1 );
and ( n14431 , n96 , n14418 );
not ( n14432 , n96 );
and ( n14433 , n14432 , n95 );
nor ( n14434 , n14431 , n14433 );
or ( n14435 , n2246 , n14434 );
nand ( n14436 , n14430 , n14435 );
buf ( n14437 , n9810 );
not ( n14438 , n14437 );
not ( n14439 , n6183 );
nand ( n14440 , n14439 , n11256 , n193 );
not ( n14441 , n14440 );
nand ( n14442 , n5563 , n4390 );
not ( n14443 , n14442 );
or ( n14444 , n14441 , n14443 );
not ( n14445 , n5611 );
nand ( n14446 , n14444 , n14445 );
nor ( n14447 , n14446 , n12673 );
not ( n14448 , n4442 );
not ( n14449 , n4522 );
or ( n14450 , n14448 , n14449 );
not ( n14451 , n193 );
nand ( n14452 , n14450 , n14451 );
nor ( n14453 , n12762 , n4426 );
nor ( n14454 , n11239 , n14453 );
not ( n14455 , n4409 );
not ( n14456 , n5511 );
or ( n14457 , n14455 , n14456 );
nand ( n14458 , n14457 , n193 );
nand ( n14459 , n14452 , n4391 , n14454 , n14458 );
not ( n14460 , n14459 );
nand ( n14461 , n14447 , n14460 );
not ( n14462 , n4605 );
not ( n14463 , n14462 );
not ( n14464 , n4447 );
nand ( n14465 , n14464 , n5556 , n11275 , n194 );
not ( n14466 , n14465 );
or ( n14467 , n14463 , n14466 );
and ( n14468 , n4430 , n6046 , n6088 );
nor ( n14469 , n4638 , n14468 );
nand ( n14470 , n14467 , n14469 );
nand ( n14471 , n14461 , n14470 );
nand ( n14472 , n5579 , n4600 );
or ( n14473 , n14472 , n11211 );
nand ( n14474 , n4556 , n4601 , n4390 );
nand ( n14475 , n14473 , n14474 );
nand ( n14476 , n14475 , n195 );
not ( n14477 , n14476 );
nand ( n14478 , n14471 , n14477 );
not ( n14479 , n4445 );
not ( n14480 , n4462 );
or ( n14481 , n14479 , n14480 );
nand ( n14482 , n4546 , n4584 );
nand ( n14483 , n14481 , n14482 );
not ( n14484 , n4601 );
nor ( n14485 , n14483 , n14484 );
nand ( n14486 , n6183 , n4390 );
nand ( n14487 , n4608 , n5555 , n14485 , n14486 );
nor ( n14488 , n14459 , n14487 );
not ( n14489 , n4468 );
nand ( n14490 , n14489 , n5604 );
nand ( n14491 , n4597 , n4437 );
and ( n14492 , n14490 , n14491 , n5625 , n194 );
or ( n14493 , n14488 , n14492 );
nand ( n14494 , n4503 , n4467 );
not ( n14495 , n14494 );
not ( n14496 , n4608 );
or ( n14497 , n14495 , n14496 );
nand ( n14498 , n14497 , n193 );
not ( n14499 , n14498 );
not ( n14500 , n195 );
not ( n14501 , n5546 );
nand ( n14502 , n4541 , n192 );
nand ( n14503 , n14501 , n14502 );
not ( n14504 , n6108 );
not ( n14505 , n4433 );
or ( n14506 , n14504 , n14505 );
nor ( n14507 , n4630 , n193 );
nand ( n14508 , n14506 , n14507 );
nand ( n14509 , n14500 , n14503 , n14508 );
nor ( n14510 , n14499 , n14509 );
nand ( n14511 , n14493 , n14510 );
nand ( n14512 , n14478 , n14511 );
not ( n14513 , n4386 );
nor ( n14514 , n14513 , n11188 );
nand ( n14515 , n6108 , n11275 );
not ( n14516 , n14515 );
not ( n14517 , n12697 );
not ( n14518 , n14517 );
or ( n14519 , n14516 , n14518 );
nand ( n14520 , n14519 , n4618 );
nand ( n14521 , n14520 , n4539 );
and ( n14522 , n5592 , n4605 );
and ( n14523 , n6242 , n12669 );
nor ( n14524 , n14522 , n14523 );
and ( n14525 , n14514 , n14521 , n14524 );
nand ( n14526 , n14512 , n14525 );
not ( n14527 , n221 );
xor ( n14528 , n14526 , n14527 );
not ( n14529 , n12554 );
not ( n14530 , n13165 );
nand ( n14531 , n14530 , n3986 );
nand ( n14532 , n4071 , n4086 );
and ( n14533 , n14532 , n4055 );
nand ( n14534 , n4087 , n5731 );
nand ( n14535 , n14531 , n14533 , n14534 );
not ( n14536 , n5185 );
not ( n14537 , n4092 );
not ( n14538 , n4073 );
or ( n14539 , n14537 , n14538 );
nand ( n14540 , n14539 , n5815 );
not ( n14541 , n14540 );
or ( n14542 , n14536 , n14541 );
and ( n14543 , n5689 , n4160 );
nor ( n14544 , n14543 , n203 );
nand ( n14545 , n14542 , n14544 );
nor ( n14546 , n14535 , n14545 );
and ( n14547 , n4086 , n4139 );
not ( n14548 , n4018 );
not ( n14549 , n5800 );
or ( n14550 , n14548 , n14549 );
nand ( n14551 , n13101 , n5185 );
nand ( n14552 , n14550 , n14551 );
nor ( n14553 , n14547 , n14552 );
or ( n14554 , n14546 , n14553 );
nand ( n14555 , n4096 , n4016 , n4107 , n198 );
not ( n14556 , n5709 );
nand ( n14557 , n14556 , n197 );
and ( n14558 , n14555 , n4088 , n14557 );
nand ( n14559 , n14554 , n14558 );
not ( n14560 , n14559 );
buf ( n14561 , n4011 );
nand ( n14562 , n5815 , n5135 );
or ( n14563 , n14561 , n14562 );
nand ( n14564 , n14563 , n5185 );
not ( n14565 , n202 );
not ( n14566 , n5867 );
or ( n14567 , n14565 , n14566 );
nand ( n14568 , n14567 , n14532 );
not ( n14569 , n199 );
not ( n14570 , n4097 );
or ( n14571 , n14569 , n14570 );
nand ( n14572 , n14571 , n5150 );
or ( n14573 , n14572 , n3997 );
nand ( n14574 , n14573 , n4121 );
nand ( n14575 , n13168 , n14574 );
nor ( n14576 , n14568 , n14575 );
not ( n14577 , n4182 );
nand ( n14578 , n5094 , n5741 );
or ( n14579 , n5149 , n14578 );
nand ( n14580 , n5875 , n4003 );
or ( n14581 , n14580 , n5159 );
nand ( n14582 , n14579 , n14581 );
not ( n14583 , n14582 );
or ( n14584 , n14577 , n14583 );
nand ( n14585 , n5827 , n203 );
not ( n14586 , n14585 );
nand ( n14587 , n14586 , n4167 , n5234 , n3973 );
nand ( n14588 , n14584 , n14587 );
nand ( n14589 , n14564 , n14576 , n14588 );
and ( n14590 , n5181 , n4067 );
nand ( n14591 , n3997 , n5671 );
nand ( n14592 , n14590 , n5747 , n4052 , n14591 );
not ( n14593 , n14592 );
nor ( n14594 , n5730 , n4170 );
nand ( n14595 , n5732 , n4160 );
nand ( n14596 , n13162 , n5096 );
nor ( n14597 , n14595 , n14596 );
or ( n14598 , n14594 , n14597 );
nand ( n14599 , n5731 , n4127 );
nand ( n14600 , n3992 , n4073 );
and ( n14601 , n14599 , n14600 , n4141 );
not ( n14602 , n4018 );
and ( n14603 , n14601 , n14602 , n5775 );
nand ( n14604 , n14598 , n14603 );
not ( n14605 , n14604 );
or ( n14606 , n14593 , n14605 );
nand ( n14607 , n5676 , n13133 );
and ( n14608 , n3996 , n4015 , n202 );
nor ( n14609 , n14608 , n204 );
not ( n14610 , n4128 );
nand ( n14611 , n3992 , n4097 );
not ( n14612 , n14611 );
or ( n14613 , n14610 , n14612 );
nand ( n14614 , n14613 , n5185 );
nand ( n14615 , n14609 , n14614 , n4191 , n14551 );
nor ( n14616 , n14607 , n14615 );
nand ( n14617 , n14606 , n14616 );
nand ( n14618 , n14589 , n14617 );
nand ( n14619 , n14560 , n14618 );
not ( n14620 , n14619 );
not ( n14621 , n14620 );
or ( n14622 , n14529 , n14621 );
nand ( n14623 , n14619 , n12555 );
nand ( n14624 , n14622 , n14623 );
xor ( n14625 , n14528 , n14624 );
not ( n14626 , n14625 );
or ( n14627 , n14438 , n14626 );
or ( n14628 , n14625 , n14437 );
nand ( n14629 , n14627 , n14628 );
or ( n14630 , n14629 , n1 );
and ( n14631 , n220 , n14527 );
not ( n14632 , n220 );
and ( n14633 , n14632 , n221 );
nor ( n14634 , n14631 , n14633 );
or ( n14635 , n2246 , n14634 );
nand ( n14636 , n14630 , n14635 );
not ( n14637 , n2512 );
not ( n14638 , n14637 );
nand ( n14639 , n2464 , n2324 );
not ( n14640 , n14639 );
not ( n14641 , n2272 );
nor ( n14642 , n2380 , n2301 );
nor ( n14643 , n14641 , n14642 );
not ( n14644 , n14643 );
or ( n14645 , n14640 , n14644 );
nand ( n14646 , n14645 , n2424 );
nand ( n14647 , n10175 , n132 );
not ( n14648 , n14647 );
and ( n14649 , n2325 , n2486 );
not ( n14650 , n14649 );
or ( n14651 , n14648 , n14650 );
nand ( n14652 , n131 , n133 );
not ( n14653 , n14652 );
nand ( n14654 , n14651 , n14653 );
not ( n14655 , n129 );
nand ( n14656 , n2287 , n2293 );
not ( n14657 , n14656 );
not ( n14658 , n14657 );
or ( n14659 , n14655 , n14658 );
nand ( n14660 , n14659 , n135 );
not ( n14661 , n14660 );
and ( n14662 , n14646 , n14654 , n14661 );
not ( n14663 , n14662 );
not ( n14664 , n2289 );
nor ( n14665 , n14664 , n10185 );
nand ( n14666 , n2441 , n131 );
nand ( n14667 , n2339 , n14666 );
or ( n14668 , n14667 , n10213 );
nand ( n14669 , n14668 , n133 );
not ( n14670 , n2464 );
not ( n14671 , n2345 );
nand ( n14672 , n14671 , n2415 );
and ( n14673 , n14670 , n14672 , n134 );
buf ( n14674 , n2366 );
not ( n14675 , n14674 );
nand ( n14676 , n14675 , n2424 );
nand ( n14677 , n14665 , n14669 , n14673 , n14676 );
nand ( n14678 , n10176 , n2332 );
nand ( n14679 , n2382 , n133 );
or ( n14680 , n14678 , n14679 );
not ( n14681 , n2416 );
or ( n14682 , n14681 , n133 );
nand ( n14683 , n14680 , n14682 );
nand ( n14684 , n2469 , n10250 );
and ( n14685 , n2471 , n14684 , n2316 );
nand ( n14686 , n10190 , n10254 );
nand ( n14687 , n2499 , n2327 );
and ( n14688 , n14685 , n14686 , n14687 );
nand ( n14689 , n14683 , n14688 );
nand ( n14690 , n14677 , n14689 );
not ( n14691 , n14690 );
or ( n14692 , n14663 , n14691 );
nand ( n14693 , n14653 , n10250 );
and ( n14694 , n10325 , n14693 , n2316 );
not ( n14695 , n14641 );
not ( n14696 , n10254 );
nand ( n14697 , n14696 , n2285 , n130 );
nand ( n14698 , n10312 , n14694 , n14695 , n14697 );
not ( n14699 , n10239 );
not ( n14700 , n10247 );
or ( n14701 , n14699 , n14700 );
nand ( n14702 , n14701 , n133 );
not ( n14703 , n2471 );
nand ( n14704 , n14703 , n130 );
nand ( n14705 , n2372 , n2408 );
and ( n14706 , n14704 , n14705 );
not ( n14707 , n2435 );
nand ( n14708 , n14707 , n10213 );
and ( n14709 , n14708 , n10176 , n134 );
nand ( n14710 , n14702 , n14706 , n14709 );
nand ( n14711 , n14698 , n14710 );
nor ( n14712 , n10239 , n2376 );
nor ( n14713 , n14712 , n135 );
not ( n14714 , n10319 );
nand ( n14715 , n14714 , n2336 );
nand ( n14716 , n10180 , n2424 );
and ( n14717 , n14713 , n14715 , n14716 , n10304 );
nand ( n14718 , n14711 , n14717 );
nand ( n14719 , n14692 , n14718 );
nand ( n14720 , n2326 , n2270 );
not ( n14721 , n14720 );
nand ( n14722 , n14721 , n2461 );
nand ( n14723 , n10213 , n14653 );
nand ( n14724 , n10302 , n132 );
not ( n14725 , n14724 );
nand ( n14726 , n14725 , n2470 );
nand ( n14727 , n14722 , n14723 , n14726 );
buf ( n14728 , n10214 );
and ( n14729 , n131 , n10323 );
not ( n14730 , n131 );
and ( n14731 , n14730 , n2279 );
nor ( n14732 , n14729 , n14731 );
not ( n14733 , n14732 );
and ( n14734 , n14728 , n14733 );
not ( n14735 , n2327 );
nor ( n14736 , n14734 , n14735 );
or ( n14737 , n14727 , n14736 );
nand ( n14738 , n14737 , n134 );
not ( n14739 , n14686 );
not ( n14740 , n2424 );
and ( n14741 , n14739 , n14740 );
nand ( n14742 , n2346 , n132 );
buf ( n14743 , n14742 );
or ( n14744 , n14743 , n2435 , n134 );
not ( n14745 , n2307 );
nand ( n14746 , n14745 , n2485 );
nand ( n14747 , n14744 , n14746 );
nor ( n14748 , n14741 , n14747 );
not ( n14749 , n14715 );
nand ( n14750 , n2367 , n2357 );
not ( n14751 , n14750 );
or ( n14752 , n14749 , n14751 );
nand ( n14753 , n14752 , n2275 );
not ( n14754 , n14724 );
nand ( n14755 , n14754 , n2499 );
and ( n14756 , n14748 , n14753 , n14755 );
not ( n14757 , n14672 );
nand ( n14758 , n14757 , n2507 );
nand ( n14759 , n14719 , n14738 , n14756 , n14758 );
not ( n14760 , n14759 );
not ( n14761 , n14760 );
or ( n14762 , n14638 , n14761 );
nand ( n14763 , n2512 , n14759 );
nand ( n14764 , n14762 , n14763 );
xor ( n14765 , n14764 , n228 );
not ( n14766 , n3018 );
nand ( n14767 , n9947 , n2942 );
nand ( n14768 , n2939 , n2942 );
and ( n14769 , n14767 , n14768 );
and ( n14770 , n9904 , n2843 );
and ( n14771 , n9905 , n120 );
nor ( n14772 , n14769 , n14770 , n14771 );
not ( n14773 , n14772 );
nor ( n14774 , n2911 , n2972 );
not ( n14775 , n14774 );
not ( n14776 , n2949 );
or ( n14777 , n14775 , n14776 );
not ( n14778 , n2866 );
nor ( n14779 , n14778 , n123 );
not ( n14780 , n121 );
nand ( n14781 , n14780 , n9960 );
nand ( n14782 , n2924 , n2843 );
nand ( n14783 , n14779 , n9893 , n14781 , n14782 );
not ( n14784 , n126 );
nor ( n14785 , n14784 , n120 );
nand ( n14786 , n14783 , n14785 );
nand ( n14787 , n14777 , n14786 );
not ( n14788 , n14787 );
nand ( n14789 , n9961 , n2987 );
and ( n14790 , n3002 , n14789 , n2827 );
not ( n14791 , n14790 );
or ( n14792 , n14788 , n14791 );
not ( n14793 , n9928 );
not ( n14794 , n9962 );
or ( n14795 , n14793 , n14794 );
nor ( n14796 , n3011 , n125 );
nand ( n14797 , n9947 , n2861 );
or ( n14798 , n14796 , n14797 );
nand ( n14799 , n14795 , n14798 );
not ( n14800 , n14783 );
and ( n14801 , n14800 , n2905 );
nand ( n14802 , n9846 , n3007 );
nand ( n14803 , n9857 , n14802 );
nor ( n14804 , n14801 , n14803 );
nand ( n14805 , n14799 , n14804 );
nand ( n14806 , n14792 , n14805 );
not ( n14807 , n14806 );
or ( n14808 , n14773 , n14807 );
not ( n14809 , n2922 );
nand ( n14810 , n2778 , n14809 );
nand ( n14811 , n9982 , n14810 , n2970 );
buf ( n14812 , n3010 );
not ( n14813 , n14812 );
and ( n14814 , n2934 , n14802 , n120 );
and ( n14815 , n14813 , n14814 );
not ( n14816 , n2902 );
nor ( n14817 , n14816 , n2911 , n120 );
nor ( n14818 , n14815 , n14817 );
or ( n14819 , n14811 , n14818 );
not ( n14820 , n2861 );
not ( n14821 , n2990 );
not ( n14822 , n2947 );
or ( n14823 , n14821 , n14822 );
nand ( n14824 , n14823 , n2897 );
not ( n14825 , n14824 );
or ( n14826 , n14820 , n14825 );
nand ( n14827 , n2925 , n9928 );
nand ( n14828 , n14826 , n14827 );
not ( n14829 , n9962 );
nand ( n14830 , n2791 , n9865 );
nor ( n14831 , n14829 , n2979 , n14830 );
nand ( n14832 , n14828 , n14831 );
nand ( n14833 , n14819 , n14832 );
not ( n14834 , n2942 );
buf ( n14835 , n2790 );
nand ( n14836 , n14835 , n124 );
not ( n14837 , n14836 );
nand ( n14838 , n2824 , n9846 );
not ( n14839 , n14838 );
or ( n14840 , n14837 , n14839 );
nand ( n14841 , n14840 , n122 );
nand ( n14842 , n14834 , n14841 , n2827 );
nand ( n14843 , n120 , n127 );
and ( n14844 , n14842 , n14843 );
nand ( n14845 , n2815 , n2924 );
nand ( n14846 , n14845 , n9847 );
or ( n14847 , n14846 , n2779 );
nand ( n14848 , n14847 , n9951 );
nand ( n14849 , n14848 , n9879 );
nor ( n14850 , n14844 , n14849 );
nand ( n14851 , n14833 , n14850 );
nand ( n14852 , n14808 , n14851 );
not ( n14853 , n2972 );
not ( n14854 , n123 );
not ( n14855 , n14854 );
not ( n14856 , n9836 );
not ( n14857 , n14856 );
or ( n14858 , n14855 , n14857 );
nand ( n14859 , n14858 , n126 );
not ( n14860 , n14859 );
or ( n14861 , n14853 , n14860 );
nand ( n14862 , n2965 , n2850 , n9907 );
nand ( n14863 , n14861 , n14862 );
and ( n14864 , n9844 , n9950 );
nand ( n14865 , n14864 , n122 );
nand ( n14866 , n14865 , n2785 );
not ( n14867 , n14866 );
not ( n14868 , n14810 );
nand ( n14869 , n14868 , n2905 );
not ( n14870 , n9962 );
nand ( n14871 , n2832 , n2976 );
not ( n14872 , n14871 );
or ( n14873 , n14870 , n14872 );
nand ( n14874 , n14873 , n9987 );
nand ( n14875 , n14867 , n14869 , n14874 );
nand ( n14876 , n14863 , n14875 );
not ( n14877 , n2959 );
not ( n14878 , n2951 );
or ( n14879 , n14877 , n14878 );
nand ( n14880 , n14879 , n2940 );
not ( n14881 , n2968 );
not ( n14882 , n2791 );
or ( n14883 , n14881 , n14882 );
nand ( n14884 , n14883 , n2861 );
not ( n14885 , n14884 );
buf ( n14886 , n2791 );
nand ( n14887 , n14886 , n2922 );
nand ( n14888 , n14885 , n14887 );
not ( n14889 , n2902 );
nand ( n14890 , n14889 , n125 );
and ( n14891 , n14880 , n14888 , n14890 );
and ( n14892 , n14876 , n14891 );
nand ( n14893 , n14852 , n14892 );
not ( n14894 , n14893 );
not ( n14895 , n14894 );
or ( n14896 , n14766 , n14895 );
or ( n14897 , n3018 , n14894 );
nand ( n14898 , n14896 , n14897 );
not ( n14899 , n14898 );
not ( n14900 , n2715 );
not ( n14901 , n139 );
nand ( n14902 , n14900 , n14901 );
and ( n14903 , n2745 , n138 );
nand ( n14904 , n14903 , n2672 );
and ( n14905 , n14902 , n14904 );
nor ( n14906 , n14905 , n141 );
not ( n14907 , n2626 );
not ( n14908 , n3380 );
and ( n14909 , n14907 , n14908 );
nor ( n14910 , n14909 , n2564 );
nand ( n14911 , n2540 , n141 );
nand ( n14912 , n14910 , n14911 , n3323 );
or ( n14913 , n14906 , n14912 );
nand ( n14914 , n140 , n141 );
not ( n14915 , n14914 );
not ( n14916 , n2755 );
or ( n14917 , n14915 , n14916 );
nand ( n14918 , n14917 , n2558 );
nand ( n14919 , n14918 , n2670 , n3336 );
nand ( n14920 , n14913 , n14919 );
not ( n14921 , n14920 );
not ( n14922 , n2753 );
not ( n14923 , n2579 );
nand ( n14924 , n14923 , n14901 );
not ( n14925 , n14924 );
or ( n14926 , n14922 , n14925 );
nand ( n14927 , n14926 , n2517 );
not ( n14928 , n14927 );
not ( n14929 , n2639 );
not ( n14930 , n2679 );
or ( n14931 , n14929 , n14930 );
nand ( n14932 , n14931 , n2642 );
nand ( n14933 , n3274 , n140 );
nor ( n14934 , n14933 , n2584 );
nor ( n14935 , n14928 , n14932 , n14934 );
not ( n14936 , n14935 );
or ( n14937 , n14921 , n14936 );
nand ( n14938 , n2673 , n3322 );
nand ( n14939 , n2648 , n2575 );
and ( n14940 , n14938 , n14939 , n2686 );
not ( n14941 , n14940 );
not ( n14942 , n3387 );
or ( n14943 , n14941 , n14942 );
not ( n14944 , n14901 );
not ( n14945 , n2673 );
or ( n14946 , n14944 , n14945 );
not ( n14947 , n143 );
nand ( n14948 , n14947 , n2761 );
nand ( n14949 , n14946 , n14948 );
not ( n14950 , n2559 );
nor ( n14951 , n14949 , n14950 );
nand ( n14952 , n14951 , n3321 );
nand ( n14953 , n14943 , n14952 );
and ( n14954 , n14953 , n137 );
nand ( n14955 , n3347 , n141 );
not ( n14956 , n14955 );
not ( n14957 , n2618 );
not ( n14958 , n2611 );
or ( n14959 , n14957 , n14958 );
nand ( n14960 , n14959 , n2564 );
not ( n14961 , n14960 );
not ( n14962 , n3367 );
not ( n14963 , n2693 );
nand ( n14964 , n14962 , n14963 );
nand ( n14965 , n2568 , n138 );
nand ( n14966 , n14961 , n14964 , n2659 , n14965 );
or ( n14967 , n14956 , n14966 );
nor ( n14968 , n2746 , n2519 );
nand ( n14969 , n3322 , n2578 );
nand ( n14970 , n14969 , n144 );
or ( n14971 , n14968 , n14970 );
nand ( n14972 , n14971 , n2654 );
not ( n14973 , n143 );
nand ( n14974 , n14973 , n2588 , n3384 );
nand ( n14975 , n2745 , n2752 );
nand ( n14976 , n14974 , n14975 );
nor ( n14977 , n14976 , n3357 );
nand ( n14978 , n14972 , n14977 );
nand ( n14979 , n14967 , n14978 );
nand ( n14980 , n14954 , n14979 );
nand ( n14981 , n14937 , n14980 );
not ( n14982 , n2529 );
not ( n14983 , n14982 );
nand ( n14984 , n14983 , n2611 );
and ( n14985 , n14984 , n2609 );
nand ( n14986 , n14963 , n138 );
not ( n14987 , n14986 );
not ( n14988 , n2717 );
or ( n14989 , n14987 , n14988 );
nand ( n14990 , n14989 , n14901 );
nand ( n14991 , n14985 , n14990 );
nand ( n14992 , n3298 , n2541 );
nor ( n14993 , n14991 , n14992 );
nand ( n14994 , n3274 , n2517 );
nand ( n14995 , n14994 , n2686 );
buf ( n14996 , n14995 );
not ( n14997 , n2576 );
nand ( n14998 , n2673 , n14997 );
not ( n14999 , n2656 );
and ( n15000 , n14999 , n2564 );
nand ( n15001 , n14998 , n15000 );
nor ( n15002 , n14996 , n15001 );
or ( n15003 , n14993 , n15002 );
buf ( n15004 , n2527 );
not ( n15005 , n15004 );
and ( n15006 , n2683 , n15005 );
nand ( n15007 , n15003 , n15006 );
and ( n15008 , n2525 , n143 );
and ( n15009 , n15008 , n2558 );
or ( n15010 , n3388 , n15009 );
nand ( n15011 , n15010 , n2686 );
not ( n15012 , n3395 );
nor ( n15013 , n15012 , n2743 );
nand ( n15014 , n3279 , n3381 );
nor ( n15015 , n3339 , n138 );
nand ( n15016 , n2673 , n15015 );
not ( n15017 , n3366 );
and ( n15018 , n15014 , n15016 , n15017 );
nand ( n15019 , n15011 , n15013 , n15018 );
nand ( n15020 , n15007 , n15019 );
and ( n15021 , n14963 , n3410 );
not ( n15022 , n141 );
nand ( n15023 , n15022 , n139 );
not ( n15024 , n15023 );
and ( n15025 , n15021 , n15024 );
not ( n15026 , n140 );
nor ( n15027 , n15026 , n2604 );
and ( n15028 , n2639 , n15027 );
nor ( n15029 , n15025 , n15028 );
and ( n15030 , n14981 , n15020 , n15029 );
not ( n15031 , n15030 );
not ( n15032 , n15031 );
and ( n15033 , n14899 , n15032 );
and ( n15034 , n15031 , n14898 );
nor ( n15035 , n15033 , n15034 );
not ( n15036 , n9903 );
not ( n15037 , n14835 );
or ( n15038 , n15036 , n15037 );
not ( n15039 , n2829 );
nand ( n15040 , n15038 , n15039 );
nand ( n15041 , n14812 , n120 );
not ( n15042 , n15041 );
nor ( n15043 , n15040 , n15042 );
not ( n15044 , n15043 );
nand ( n15045 , n2938 , n2828 );
not ( n15046 , n15045 );
nand ( n15047 , n2948 , n2780 );
not ( n15048 , n15047 );
or ( n15049 , n15046 , n15048 );
nand ( n15050 , n15049 , n123 );
not ( n15051 , n15050 );
or ( n15052 , n15044 , n15051 );
nand ( n15053 , n15052 , n2785 );
not ( n15054 , n9938 );
nand ( n15055 , n15054 , n9853 );
not ( n15056 , n120 );
nor ( n15057 , n15056 , n122 );
and ( n15058 , n15055 , n15057 );
nand ( n15059 , n3006 , n14809 );
not ( n15060 , n15059 );
not ( n15061 , n9867 );
or ( n15062 , n15060 , n15061 );
nand ( n15063 , n15062 , n126 );
nand ( n15064 , n2969 , n125 );
not ( n15065 , n15064 );
not ( n15066 , n2925 );
or ( n15067 , n15065 , n15066 );
nand ( n15068 , n15067 , n2973 );
nand ( n15069 , n15063 , n15068 );
nor ( n15070 , n15058 , n15069 );
not ( n15071 , n9981 );
nand ( n15072 , n15071 , n122 );
not ( n15073 , n15072 );
nor ( n15074 , n2912 , n120 );
nor ( n15075 , n15073 , n15074 , n127 );
nand ( n15076 , n15053 , n15070 , n15075 );
not ( n15077 , n15045 );
nand ( n15078 , n2807 , n124 );
and ( n15079 , n15077 , n15078 );
nor ( n15080 , n15079 , n14864 );
nand ( n15081 , n9992 , n9843 , n15080 );
not ( n15082 , n2857 );
not ( n15083 , n9837 );
or ( n15084 , n15082 , n15083 );
nand ( n15085 , n9988 , n9924 );
not ( n15086 , n14865 );
nor ( n15087 , n14859 , n15085 , n15086 );
nand ( n15088 , n15084 , n15087 );
nand ( n15089 , n15076 , n15081 , n15088 );
not ( n15090 , n14771 );
not ( n15091 , n14802 );
and ( n15092 , n2967 , n2854 );
not ( n15093 , n2897 );
nor ( n15094 , n15092 , n15093 , n2905 );
not ( n15095 , n15094 );
or ( n15096 , n15091 , n15095 );
and ( n15097 , n9895 , n14886 , n2905 );
nand ( n15098 , n15097 , n9841 );
nand ( n15099 , n15096 , n15098 );
nand ( n15100 , n15090 , n15099 , n127 );
nand ( n15101 , n15076 , n15100 );
nand ( n15102 , n3000 , n126 );
nor ( n15103 , n15073 , n15102 );
nand ( n15104 , n2948 , n2843 );
not ( n15105 , n15104 );
nand ( n15106 , n2957 , n2968 );
not ( n15107 , n15106 );
nand ( n15108 , n15107 , n3006 , n2850 );
not ( n15109 , n15108 );
or ( n15110 , n15105 , n15109 );
nand ( n15111 , n15110 , n120 );
nor ( n15112 , n2835 , n2854 );
and ( n15113 , n2805 , n9840 );
or ( n15114 , n15112 , n15113 );
nand ( n15115 , n15114 , n2857 );
nand ( n15116 , n15103 , n15111 , n15115 );
not ( n15117 , n2798 );
not ( n15118 , n2940 );
not ( n15119 , n2948 );
or ( n15120 , n15118 , n15119 );
nand ( n15121 , n15120 , n14810 );
nor ( n15122 , n15117 , n15121 );
not ( n15123 , n9987 );
not ( n15124 , n15123 );
not ( n15125 , n14886 );
or ( n15126 , n15124 , n15125 );
not ( n15127 , n9858 );
nand ( n15128 , n15126 , n15127 );
not ( n15129 , n9841 );
or ( n15130 , n15128 , n15129 );
nand ( n15131 , n15130 , n2819 );
nand ( n15132 , n15122 , n15131 );
and ( n15133 , n15116 , n15132 );
or ( n15134 , n2922 , n2968 );
nand ( n15135 , n15134 , n2986 );
not ( n15136 , n15135 );
nor ( n15137 , n9904 , n120 );
nor ( n15138 , n15136 , n15137 );
nor ( n15139 , n15133 , n15138 );
nand ( n15140 , n15089 , n15101 , n15139 );
not ( n15141 , n15140 );
not ( n15142 , n15141 );
not ( n15143 , n116 );
nand ( n15144 , n15143 , n10003 );
not ( n15145 , n15144 );
nand ( n15146 , n15145 , n3113 );
nand ( n15147 , n15146 , n10035 );
nor ( n15148 , n15147 , n3175 );
not ( n15149 , n15148 );
nand ( n15150 , n10104 , n3164 );
nor ( n15151 , n15150 , n3183 );
not ( n15152 , n15151 );
not ( n15153 , n113 );
nand ( n15154 , n15153 , n114 );
nor ( n15155 , n15154 , n3084 );
and ( n15156 , n15155 , n3037 );
nand ( n15157 , n15156 , n112 );
not ( n15158 , n15157 );
or ( n15159 , n15152 , n15158 );
nand ( n15160 , n3052 , n3025 );
nand ( n15161 , n15160 , n117 );
not ( n15162 , n15161 );
not ( n15163 , n116 );
not ( n15164 , n10091 );
or ( n15165 , n15163 , n15164 );
nand ( n15166 , n15165 , n3226 );
nand ( n15167 , n15166 , n112 );
and ( n15168 , n3193 , n115 );
and ( n15169 , n15168 , n3113 );
nand ( n15170 , n15169 , n116 );
and ( n15171 , n3152 , n3026 );
nand ( n15172 , n15171 , n3071 );
nand ( n15173 , n15162 , n15167 , n15170 , n15172 );
nand ( n15174 , n15159 , n15173 );
not ( n15175 , n15174 );
or ( n15176 , n15149 , n15175 );
nand ( n15177 , n3090 , n3174 , n3251 );
nand ( n15178 , n15177 , n118 );
nor ( n15179 , n10051 , n3051 );
nor ( n15180 , n15178 , n15179 );
nor ( n15181 , n3258 , n115 );
not ( n15182 , n3126 );
not ( n15183 , n10124 );
or ( n15184 , n15182 , n15183 );
nand ( n15185 , n15184 , n10121 );
or ( n15186 , n15181 , n15185 );
nand ( n15187 , n15186 , n3164 );
nand ( n15188 , n15180 , n15187 );
nand ( n15189 , n15176 , n15188 );
nand ( n15190 , n3118 , n3111 );
not ( n15191 , n15190 );
not ( n15192 , n3200 );
or ( n15193 , n15191 , n15192 );
nand ( n15194 , n15193 , n3235 );
not ( n15195 , n113 );
nor ( n15196 , n15195 , n115 );
nand ( n15197 , n3090 , n15196 );
not ( n15198 , n15197 );
and ( n15199 , n15198 , n3266 );
and ( n15200 , n3248 , n115 );
and ( n15201 , n15200 , n3199 );
nor ( n15202 , n15199 , n15201 );
and ( n15203 , n15194 , n15202 );
nand ( n15204 , n15189 , n15203 );
not ( n15205 , n15204 );
not ( n15206 , n15171 );
not ( n15207 , n15206 );
and ( n15208 , n3229 , n3051 );
nor ( n15209 , n15208 , n117 );
not ( n15210 , n15209 );
or ( n15211 , n15207 , n15210 );
not ( n15212 , n116 );
nand ( n15213 , n15212 , n15168 );
and ( n15214 , n10039 , n117 );
nand ( n15215 , n15213 , n15214 );
nand ( n15216 , n15211 , n15215 );
not ( n15217 , n15216 );
not ( n15218 , n3119 );
or ( n15219 , n15217 , n15218 );
nand ( n15220 , n15219 , n118 );
nand ( n15221 , n15200 , n10037 );
and ( n15222 , n15146 , n15221 );
nor ( n15223 , n117 , n119 );
not ( n15224 , n15223 );
nand ( n15225 , n3183 , n3251 );
not ( n15226 , n15225 );
or ( n15227 , n15224 , n15226 );
and ( n15228 , n3144 , n3061 , n10030 );
not ( n15229 , n15228 );
and ( n15230 , n3059 , n3257 );
nand ( n15231 , n3137 , n117 );
nor ( n15232 , n15230 , n15231 );
nand ( n15233 , n15229 , n15232 );
nand ( n15234 , n15227 , n15233 );
nand ( n15235 , n10076 , n117 );
nand ( n15236 , n15235 , n3219 );
nor ( n15237 , n10039 , n3064 );
or ( n15238 , n15236 , n15237 );
nand ( n15239 , n15238 , n3106 );
nand ( n15240 , n15220 , n15222 , n15234 , n15239 );
and ( n15241 , n3134 , n113 );
nor ( n15242 , n15241 , n3128 );
nand ( n15243 , n3241 , n15242 );
not ( n15244 , n15181 );
and ( n15245 , n3149 , n10009 , n10145 );
nand ( n15246 , n15244 , n15245 );
and ( n15247 , n15243 , n15246 );
nand ( n15248 , n15240 , n15247 );
not ( n15249 , n10142 );
not ( n15250 , n15169 );
not ( n15251 , n10014 );
and ( n15252 , n15250 , n15251 , n118 );
nor ( n15253 , n15252 , n3235 );
nor ( n15254 , n15249 , n15253 );
not ( n15255 , n10077 );
not ( n15256 , n3026 );
not ( n15257 , n15256 );
not ( n15258 , n117 );
nor ( n15259 , n15258 , n114 );
and ( n15260 , n15257 , n15259 );
nor ( n15261 , n15255 , n15260 );
and ( n15262 , n15254 , n15261 );
not ( n15263 , n15156 );
nand ( n15264 , n3095 , n112 );
nand ( n15265 , n3055 , n116 );
nand ( n15266 , n15263 , n15264 , n15265 );
not ( n15267 , n3099 );
not ( n15268 , n3144 );
or ( n15269 , n15267 , n15268 );
nand ( n15270 , n15269 , n3106 );
not ( n15271 , n15270 );
nand ( n15272 , n10133 , n117 );
nand ( n15273 , n15271 , n15272 );
nor ( n15274 , n15266 , n15273 );
nor ( n15275 , n15262 , n15274 );
nand ( n15276 , n15240 , n15275 );
nand ( n15277 , n15240 , n3137 );
nand ( n15278 , n15205 , n15248 , n15276 , n15277 );
not ( n15279 , n15278 );
not ( n15280 , n15279 );
and ( n15281 , n15142 , n15280 );
and ( n15282 , n15279 , n15141 );
nor ( n15283 , n15281 , n15282 );
not ( n15284 , n15283 );
and ( n15285 , n15035 , n15284 );
not ( n15286 , n15035 );
and ( n15287 , n15286 , n15283 );
nor ( n15288 , n15285 , n15287 );
and ( n15289 , n14765 , n15288 );
not ( n15290 , n14765 );
not ( n15291 , n15288 );
and ( n15292 , n15290 , n15291 );
nor ( n15293 , n15289 , n15292 );
or ( n15294 , n15293 , n1 );
xnor ( n15295 , n228 , n229 );
or ( n15296 , n2246 , n15295 );
nand ( n15297 , n15294 , n15296 );
not ( n15298 , n100 );
not ( n15299 , n15298 );
not ( n15300 , n13224 );
or ( n15301 , n15299 , n15300 );
not ( n15302 , n13224 );
nand ( n15303 , n15302 , n100 );
nand ( n15304 , n15301 , n15303 );
buf ( n15305 , n12770 );
not ( n15306 , n15305 );
and ( n15307 , n15304 , n15306 );
not ( n15308 , n15304 );
not ( n15309 , n12770 );
not ( n15310 , n15309 );
and ( n15311 , n15308 , n15310 );
nor ( n15312 , n15307 , n15311 );
not ( n15313 , n14624 );
not ( n15314 , n5492 );
and ( n15315 , n15313 , n15314 );
and ( n15316 , n14624 , n5492 );
nor ( n15317 , n15315 , n15316 );
not ( n15318 , n15317 );
and ( n15319 , n15312 , n15318 );
not ( n15320 , n15312 );
and ( n15321 , n15320 , n15317 );
nor ( n15322 , n15319 , n15321 );
or ( n15323 , n15322 , n1 );
and ( n15324 , n268 , n15298 );
not ( n15325 , n268 );
and ( n15326 , n15325 , n100 );
nor ( n15327 , n15324 , n15326 );
or ( n15328 , n2246 , n15327 );
nand ( n15329 , n15323 , n15328 );
nand ( n15330 , n2779 , n2940 );
and ( n15331 , n15330 , n9988 );
not ( n15332 , n15331 );
not ( n15333 , n9838 );
nor ( n15334 , n15333 , n9842 );
not ( n15335 , n15334 );
or ( n15336 , n15332 , n15335 );
nor ( n15337 , n2865 , n121 );
nor ( n15338 , n2956 , n9874 );
nand ( n15339 , n15337 , n15338 );
not ( n15340 , n15339 );
not ( n15341 , n9879 );
or ( n15342 , n15340 , n15341 );
nand ( n15343 , n15342 , n2905 );
not ( n15344 , n9860 );
nand ( n15345 , n15344 , n9938 );
not ( n15346 , n15345 );
not ( n15347 , n9838 );
or ( n15348 , n15346 , n15347 );
nand ( n15349 , n15348 , n120 );
nand ( n15350 , n15343 , n126 , n15349 );
nand ( n15351 , n15336 , n15350 );
not ( n15352 , n14836 );
and ( n15353 , n15077 , n15352 );
nor ( n15354 , n15353 , n9978 );
nand ( n15355 , n15351 , n15354 );
not ( n15356 , n15355 );
not ( n15357 , n9943 );
not ( n15358 , n9875 );
not ( n15359 , n2857 );
and ( n15360 , n15358 , n15359 );
not ( n15361 , n2843 );
not ( n15362 , n9898 );
or ( n15363 , n15361 , n15362 );
not ( n15364 , n2900 );
not ( n15365 , n125 );
and ( n15366 , n15364 , n15365 );
nor ( n15367 , n15366 , n2785 );
nand ( n15368 , n15363 , n15367 );
nor ( n15369 , n15360 , n15368 );
nand ( n15370 , n15357 , n15369 , n9849 );
or ( n15371 , n15106 , n9846 , n126 );
nand ( n15372 , n15371 , n2860 );
nand ( n15373 , n2832 , n9884 );
nand ( n15374 , n15372 , n15373 );
and ( n15375 , n15370 , n15374 );
not ( n15376 , n3011 );
nor ( n15377 , n2808 , n9903 );
nor ( n15378 , n15377 , n2986 );
nor ( n15379 , n15376 , n15378 );
or ( n15380 , n2880 , n9905 );
nand ( n15381 , n15380 , n14843 );
nand ( n15382 , n15379 , n15381 );
nor ( n15383 , n15375 , n15382 );
not ( n15384 , n15383 );
not ( n15385 , n2951 );
or ( n15386 , n9839 , n15385 );
nand ( n15387 , n15386 , n120 );
not ( n15388 , n15387 );
or ( n15389 , n15384 , n15388 );
not ( n15390 , n14770 );
not ( n15391 , n15390 );
not ( n15392 , n9859 );
or ( n15393 , n15391 , n15392 );
not ( n15394 , n2797 );
not ( n15395 , n15337 );
nand ( n15396 , n15394 , n15041 , n15395 , n15123 );
nand ( n15397 , n15393 , n15396 );
nand ( n15398 , n15397 , n120 );
not ( n15399 , n15398 );
nor ( n15400 , n14770 , n9837 );
not ( n15401 , n15400 );
not ( n15402 , n9859 );
or ( n15403 , n15401 , n15402 );
nand ( n15404 , n15403 , n15396 );
not ( n15405 , n14841 );
and ( n15406 , n2832 , n2909 );
nor ( n15407 , n15405 , n15406 );
nand ( n15408 , n15404 , n15407 );
not ( n15409 , n15408 );
or ( n15410 , n15399 , n15409 );
and ( n15411 , n2845 , n2942 );
not ( n15412 , n15411 );
and ( n15413 , n2948 , n125 );
not ( n15414 , n15413 );
not ( n15415 , n15414 );
or ( n15416 , n15412 , n15415 );
nand ( n15417 , n15416 , n14768 );
not ( n15418 , n14835 );
nand ( n15419 , n2973 , n2977 , n15418 );
and ( n15420 , n15417 , n15419 );
nand ( n15421 , n15410 , n15420 );
nand ( n15422 , n15389 , n15421 );
nand ( n15423 , n15356 , n15422 );
not ( n15424 , n15423 );
and ( n15425 , n15249 , n117 );
nand ( n15426 , n10033 , n3199 );
nand ( n15427 , n15426 , n3137 );
nor ( n15428 , n15425 , n15427 );
not ( n15429 , n15428 );
not ( n15430 , n3205 );
not ( n15431 , n117 );
and ( n15432 , n15430 , n15431 );
nand ( n15433 , n3239 , n15197 );
nor ( n15434 , n15432 , n15433 );
or ( n15435 , n15434 , n116 );
not ( n15436 , n3229 );
and ( n15437 , n10161 , n15436 );
nor ( n15438 , n15437 , n3164 );
nor ( n15439 , n15270 , n15438 );
nand ( n15440 , n15435 , n15439 );
nand ( n15441 , n3160 , n3199 );
nand ( n15442 , n3148 , n10030 );
and ( n15443 , n15442 , n118 );
nand ( n15444 , n3144 , n10116 );
nand ( n15445 , n3063 , n3194 );
nand ( n15446 , n15441 , n15443 , n15444 , n15445 );
and ( n15447 , n15440 , n15446 );
not ( n15448 , n3164 );
not ( n15449 , n10073 );
or ( n15450 , n15448 , n15449 );
nand ( n15451 , n3266 , n3055 , n114 );
nand ( n15452 , n15450 , n15451 );
nor ( n15453 , n15447 , n15452 );
not ( n15454 , n15453 );
or ( n15455 , n15429 , n15454 );
nor ( n15456 , n3259 , n10002 );
and ( n15457 , n15456 , n10084 );
nor ( n15458 , n15457 , n3164 );
and ( n15459 , n15144 , n10035 );
nand ( n15460 , n15169 , n3063 );
nor ( n15461 , n10078 , n10156 );
nand ( n15462 , n15459 , n15460 , n15461 );
or ( n15463 , n15458 , n15462 );
not ( n15464 , n3248 );
nand ( n15465 , n15464 , n10075 , n118 );
and ( n15466 , n15465 , n3234 );
buf ( n15467 , n3243 );
or ( n15468 , n15466 , n15467 );
nand ( n15469 , n15463 , n15468 );
nand ( n15470 , n15206 , n3130 );
or ( n15471 , n3057 , n10073 , n15470 );
nand ( n15472 , n3134 , n3048 );
nand ( n15473 , n15472 , n10046 , n3138 );
nand ( n15474 , n15471 , n15473 );
nand ( n15475 , n3160 , n3111 );
not ( n15476 , n15475 );
not ( n15477 , n15179 );
not ( n15478 , n15196 );
not ( n15479 , n15478 );
not ( n15480 , n10032 );
or ( n15481 , n15479 , n15480 );
nand ( n15482 , n15481 , n3266 );
nand ( n15483 , n15477 , n15482 );
nor ( n15484 , n15476 , n15483 );
nand ( n15485 , n15469 , n15474 , n15484 );
nand ( n15486 , n15455 , n15485 );
not ( n15487 , n10000 );
nand ( n15488 , n10091 , n3257 );
nand ( n15489 , n15488 , n15190 );
nor ( n15490 , n15489 , n15147 );
not ( n15491 , n15490 );
or ( n15492 , n15487 , n15491 );
nand ( n15493 , n15492 , n10036 );
not ( n15494 , n15493 );
not ( n15495 , n10148 );
or ( n15496 , n15494 , n15495 );
not ( n15497 , n3171 );
and ( n15498 , n15497 , n3063 );
nor ( n15499 , n15498 , n15181 );
not ( n15500 , n15488 );
not ( n15501 , n10054 );
and ( n15502 , n15500 , n15501 );
nor ( n15503 , n15502 , n3106 );
nand ( n15504 , n10052 , n3199 );
nand ( n15505 , n15499 , n10142 , n15503 , n15504 );
nand ( n15506 , n15496 , n15505 );
not ( n15507 , n15442 );
nand ( n15508 , n3160 , n3212 );
not ( n15509 , n15508 );
or ( n15510 , n15507 , n15509 );
nand ( n15511 , n15510 , n10054 );
not ( n15512 , n3249 );
not ( n15513 , n15512 );
not ( n15514 , n15172 );
or ( n15515 , n15513 , n15514 );
nand ( n15516 , n15515 , n10037 );
nand ( n15517 , n15486 , n15506 , n15511 , n15516 );
not ( n15518 , n15517 );
and ( n15519 , n15424 , n15518 );
not ( n15520 , n15424 );
and ( n15521 , n15520 , n15517 );
or ( n15522 , n15519 , n15521 );
not ( n15523 , n15522 );
not ( n15524 , n2771 );
or ( n15525 , n15523 , n15524 );
not ( n15526 , n15522 );
not ( n15527 , n2771 );
nand ( n15528 , n15526 , n15527 );
nand ( n15529 , n15525 , n15528 );
not ( n15530 , n2417 );
not ( n15531 , n2474 );
or ( n15532 , n15530 , n15531 );
or ( n15533 , n2488 , n132 );
nand ( n15534 , n15532 , n15533 );
not ( n15535 , n15534 );
not ( n15536 , n2316 );
or ( n15537 , n15535 , n15536 );
not ( n15538 , n2394 );
not ( n15539 , n15538 );
nand ( n15540 , n2333 , n133 );
not ( n15541 , n15540 );
or ( n15542 , n15539 , n15541 );
nand ( n15543 , n15542 , n2284 );
not ( n15544 , n15543 );
not ( n15545 , n10250 );
not ( n15546 , n15545 );
not ( n15547 , n10191 );
or ( n15548 , n15546 , n15547 );
nand ( n15549 , n15548 , n2418 );
not ( n15550 , n15549 );
or ( n15551 , n15544 , n15550 );
nand ( n15552 , n15551 , n134 );
nand ( n15553 , n15537 , n15552 );
not ( n15554 , n2301 );
and ( n15555 , n10184 , n2424 );
not ( n15556 , n15555 );
or ( n15557 , n15554 , n15556 );
nand ( n15558 , n15557 , n2359 );
not ( n15559 , n15558 );
or ( n15560 , n10261 , n132 );
not ( n15561 , n14642 );
nand ( n15562 , n15560 , n15561 );
and ( n15563 , n15562 , n2424 );
nand ( n15564 , n128 , n132 );
not ( n15565 , n15564 );
or ( n15566 , n2274 , n15565 , n2463 );
nor ( n15567 , n2489 , n2336 );
or ( n15568 , n15567 , n14724 );
nand ( n15569 , n15566 , n15568 );
nor ( n15570 , n15563 , n15569 );
nand ( n15571 , n15559 , n15570 );
or ( n15572 , n15553 , n15571 );
nand ( n15573 , n10226 , n14639 );
not ( n15574 , n15573 );
not ( n15575 , n10224 );
nor ( n15576 , n15575 , n14721 );
nand ( n15577 , n15574 , n15576 );
and ( n15578 , n15577 , n133 );
not ( n15579 , n2336 );
not ( n15580 , n15579 );
not ( n15581 , n2460 );
and ( n15582 , n15580 , n15581 );
not ( n15583 , n2353 );
not ( n15584 , n10253 );
or ( n15585 , n15583 , n15584 );
nand ( n15586 , n15585 , n135 );
nor ( n15587 , n15582 , n15586 );
not ( n15588 , n130 );
nand ( n15589 , n15588 , n2461 );
not ( n15590 , n15589 );
not ( n15591 , n2325 );
or ( n15592 , n15590 , n15591 );
not ( n15593 , n2293 );
not ( n15594 , n15593 );
nand ( n15595 , n15592 , n15594 );
not ( n15596 , n2373 );
nand ( n15597 , n15596 , n2424 );
nand ( n15598 , n2333 , n2301 );
nand ( n15599 , n15587 , n15595 , n15597 , n15598 );
nor ( n15600 , n15578 , n15599 );
not ( n15601 , n2382 );
nand ( n15602 , n15601 , n2301 );
nor ( n15603 , n14647 , n131 );
nor ( n15604 , n15603 , n134 );
not ( n15605 , n2415 );
not ( n15606 , n15605 );
not ( n15607 , n2328 );
or ( n15608 , n15606 , n15607 );
buf ( n15609 , n10276 );
nand ( n15610 , n15608 , n15609 );
nand ( n15611 , n15602 , n15604 , n15610 );
and ( n15612 , n2367 , n2301 );
not ( n15613 , n15612 );
and ( n15614 , n2334 , n15613 , n10263 );
nor ( n15615 , n15614 , n2424 );
or ( n15616 , n15611 , n15615 );
not ( n15617 , n2506 );
not ( n15618 , n2470 );
nand ( n15619 , n15618 , n14674 , n134 );
not ( n15620 , n15619 );
or ( n15621 , n15617 , n15620 );
nand ( n15622 , n15621 , n10291 );
nand ( n15623 , n15616 , n15622 );
nand ( n15624 , n15600 , n15623 );
nand ( n15625 , n15572 , n15624 );
not ( n15626 , n134 );
not ( n15627 , n10177 );
or ( n15628 , n15626 , n15627 );
nand ( n15629 , n14670 , n10258 );
nand ( n15630 , n15628 , n15629 );
not ( n15631 , n14684 );
buf ( n15632 , n2286 );
not ( n15633 , n15632 );
or ( n15634 , n15631 , n15633 );
nand ( n15635 , n15634 , n2485 );
and ( n15636 , n15630 , n10309 , n15635 );
not ( n15637 , n2471 );
nand ( n15638 , n14641 , n2324 );
not ( n15639 , n15638 );
or ( n15640 , n15637 , n15639 );
nand ( n15641 , n15640 , n2435 );
nand ( n15642 , n2491 , n2389 , n2377 );
not ( n15643 , n10210 );
nand ( n15644 , n15643 , n2461 );
and ( n15645 , n15642 , n15644 , n2316 );
nor ( n15646 , n10187 , n2282 );
not ( n15647 , n15646 );
not ( n15648 , n10308 );
not ( n15649 , n15648 );
or ( n15650 , n15647 , n15649 );
nand ( n15651 , n15650 , n2327 );
and ( n15652 , n15641 , n15645 , n15651 );
nor ( n15653 , n15636 , n15652 );
not ( n15654 , n10235 );
not ( n15655 , n15643 );
or ( n15656 , n15654 , n15655 );
or ( n15657 , n10283 , n2324 );
nand ( n15658 , n15656 , n15657 );
nor ( n15659 , n15653 , n15658 );
nand ( n15660 , n15625 , n15659 );
buf ( n15661 , n15660 );
not ( n15662 , n15661 );
not ( n15663 , n274 );
and ( n15664 , n15662 , n15663 );
and ( n15665 , n15661 , n274 );
nor ( n15666 , n15664 , n15665 );
not ( n15667 , n15666 );
and ( n15668 , n15529 , n15667 );
not ( n15669 , n15529 );
and ( n15670 , n15669 , n15666 );
nor ( n15671 , n15668 , n15670 );
or ( n15672 , n15671 , n1 );
xnor ( n15673 , n274 , n275 );
or ( n15674 , n2246 , n15673 );
nand ( n15675 , n15672 , n15674 );
not ( n15676 , n10216 );
not ( n15677 , n15676 );
not ( n15678 , n10291 );
or ( n15679 , n15677 , n15678 );
nand ( n15680 , n15679 , n2424 );
nor ( n15681 , n14742 , n131 );
nand ( n15682 , n15681 , n129 );
not ( n15683 , n15682 );
nand ( n15684 , n14757 , n133 );
nand ( n15685 , n14746 , n15684 , n2316 );
nor ( n15686 , n15683 , n15685 );
nand ( n15687 , n2333 , n2285 );
nand ( n15688 , n15680 , n15686 , n15687 );
or ( n15689 , n2398 , n2301 );
nand ( n15690 , n15689 , n10278 , n134 );
not ( n15691 , n10261 );
or ( n15692 , n15690 , n15691 );
nand ( n15693 , n15692 , n2506 );
and ( n15694 , n2451 , n14656 );
nand ( n15695 , n2380 , n10241 );
nand ( n15696 , n10224 , n15695 , n133 );
nand ( n15697 , n15693 , n15694 , n15696 , n2497 );
nand ( n15698 , n15688 , n15697 );
not ( n15699 , n15698 );
and ( n15700 , n15683 , n2424 );
not ( n15701 , n14684 );
nor ( n15702 , n15700 , n15701 );
nand ( n15703 , n10226 , n10319 );
or ( n15704 , n15703 , n15612 );
nand ( n15705 , n15704 , n133 );
nand ( n15706 , n15702 , n15705 );
nor ( n15707 , n15558 , n15706 );
not ( n15708 , n15707 );
or ( n15709 , n15699 , n15708 );
not ( n15710 , n2370 );
and ( n15711 , n15710 , n2376 );
nor ( n15712 , n15711 , n2359 );
not ( n15713 , n10237 );
nand ( n15714 , n15713 , n2315 );
not ( n15715 , n15714 );
not ( n15716 , n2391 );
or ( n15717 , n15715 , n15716 );
nand ( n15718 , n15717 , n2424 );
not ( n15719 , n2424 );
not ( n15720 , n2333 );
or ( n15721 , n15719 , n15720 );
nand ( n15722 , n2499 , n2435 );
nand ( n15723 , n15721 , n15722 );
nand ( n15724 , n15723 , n2301 );
and ( n15725 , n15712 , n15718 , n15724 );
not ( n15726 , n2256 );
not ( n15727 , n2407 );
and ( n15728 , n15726 , n15727 );
not ( n15729 , n15714 );
nor ( n15730 , n15728 , n15729 );
nand ( n15731 , n10213 , n10287 );
not ( n15732 , n14647 );
nand ( n15733 , n15732 , n10303 );
nand ( n15734 , n15730 , n15731 , n15733 );
and ( n15735 , n15734 , n2316 );
not ( n15736 , n134 );
nand ( n15737 , n2500 , n14705 );
not ( n15738 , n15737 );
or ( n15739 , n15736 , n15738 );
buf ( n15740 , n2457 );
nand ( n15741 , n15740 , n14743 );
or ( n15742 , n15741 , n2399 );
nand ( n15743 , n15742 , n2507 );
nand ( n15744 , n15739 , n15743 );
nor ( n15745 , n15735 , n15744 );
nand ( n15746 , n15725 , n15745 );
nand ( n15747 , n15709 , n15746 );
or ( n15748 , n10242 , n2339 );
nand ( n15749 , n15748 , n10210 );
not ( n15750 , n2451 );
or ( n15751 , n15749 , n2368 , n15750 );
nand ( n15752 , n10298 , n2321 );
nand ( n15753 , n15751 , n15752 );
not ( n15754 , n14686 );
nand ( n15755 , n2408 , n2470 );
not ( n15756 , n15755 );
not ( n15757 , n10277 );
or ( n15758 , n15756 , n15757 );
nand ( n15759 , n15758 , n134 );
not ( n15760 , n15759 );
or ( n15761 , n15754 , n15760 );
nand ( n15762 , n15761 , n2321 );
and ( n15763 , n10224 , n2416 );
not ( n15764 , n15763 );
not ( n15765 , n14750 );
or ( n15766 , n15764 , n15765 );
nand ( n15767 , n15766 , n2265 );
not ( n15768 , n15767 );
not ( n15769 , n2316 );
not ( n15770 , n10226 );
not ( n15771 , n15770 );
or ( n15772 , n15769 , n15771 );
nand ( n15773 , n10296 , n2325 );
or ( n15774 , n15773 , n15596 );
nand ( n15775 , n15774 , n2476 );
nand ( n15776 , n15772 , n15775 );
nor ( n15777 , n15768 , n15776 );
and ( n15778 , n15753 , n15762 , n15777 );
nand ( n15779 , n15747 , n15778 );
not ( n15780 , n15779 );
not ( n15781 , n15780 );
not ( n15782 , n278 );
and ( n15783 , n15781 , n15782 );
buf ( n15784 , n15779 );
not ( n15785 , n15784 );
and ( n15786 , n15785 , n278 );
nor ( n15787 , n15783 , n15786 );
not ( n15788 , n15660 );
and ( n15789 , n15788 , n2512 );
not ( n15790 , n15788 );
and ( n15791 , n15790 , n2513 );
nor ( n15792 , n15789 , n15791 );
xnor ( n15793 , n15787 , n15792 );
not ( n15794 , n14933 );
nand ( n15795 , n3333 , n2517 );
not ( n15796 , n15795 );
not ( n15797 , n138 );
and ( n15798 , n15796 , n15797 );
buf ( n15799 , n2721 );
not ( n15800 , n15799 );
nor ( n15801 , n15798 , n15800 );
not ( n15802 , n15801 );
or ( n15803 , n15794 , n15802 );
nand ( n15804 , n15803 , n141 );
and ( n15805 , n2747 , n140 );
nand ( n15806 , n3339 , n138 );
not ( n15807 , n15806 );
not ( n15808 , n2673 );
or ( n15809 , n15807 , n15808 );
and ( n15810 , n2526 , n2564 );
nand ( n15811 , n15809 , n15810 );
nor ( n15812 , n15805 , n15811 );
nand ( n15813 , n15804 , n15812 );
not ( n15814 , n2654 );
nand ( n15815 , n2665 , n2604 , n144 );
not ( n15816 , n15815 );
or ( n15817 , n15814 , n15816 );
nand ( n15818 , n15817 , n3345 );
nand ( n15819 , n15813 , n15818 );
nand ( n15820 , n3325 , n143 );
nand ( n15821 , n15820 , n3293 );
nand ( n15822 , n14902 , n2674 );
or ( n15823 , n15821 , n15822 );
nand ( n15824 , n15823 , n141 );
nand ( n15825 , n2540 , n2517 );
not ( n15826 , n2763 );
not ( n15827 , n3316 );
or ( n15828 , n15826 , n15827 );
nand ( n15829 , n15828 , n2686 );
or ( n15830 , n2555 , n2554 );
and ( n15831 , n15830 , n2562 );
nor ( n15832 , n15831 , n2642 );
and ( n15833 , n15825 , n15829 , n15016 , n15832 );
nand ( n15834 , n15819 , n15824 , n15833 );
not ( n15835 , n15834 );
not ( n15836 , n142 );
not ( n15837 , n14997 );
or ( n15838 , n15836 , n15837 );
nand ( n15839 , n15838 , n15820 );
not ( n15840 , n3385 );
or ( n15841 , n15839 , n15840 );
nand ( n15842 , n15841 , n2686 );
not ( n15843 , n2517 );
nand ( n15844 , n2556 , n2559 );
not ( n15845 , n15844 );
or ( n15846 , n15843 , n15845 );
not ( n15847 , n142 );
nor ( n15848 , n15847 , n3367 );
not ( n15849 , n15848 );
nand ( n15850 , n15849 , n2590 , n141 );
nand ( n15851 , n15846 , n15850 );
or ( n15852 , n15851 , n14960 );
nand ( n15853 , n2540 , n2639 );
not ( n15854 , n3310 );
not ( n15855 , n3334 );
or ( n15856 , n15854 , n15855 );
not ( n15857 , n2652 );
nand ( n15858 , n15856 , n15857 );
nand ( n15859 , n3288 , n143 );
nand ( n15860 , n15853 , n15858 , n15859 , n144 );
nand ( n15861 , n15852 , n15860 );
not ( n15862 , n2753 );
not ( n15863 , n3395 );
or ( n15864 , n15862 , n15863 );
nand ( n15865 , n15864 , n2673 );
nand ( n15866 , n15842 , n15861 , n15865 , n2642 );
not ( n15867 , n15866 );
or ( n15868 , n15835 , n15867 );
nor ( n15869 , n14999 , n143 );
or ( n15870 , n15869 , n3320 );
not ( n15871 , n2591 );
or ( n15872 , n15871 , n141 );
nand ( n15873 , n15870 , n15872 );
not ( n15874 , n3357 );
nand ( n15875 , n15873 , n3387 , n15874 , n144 );
not ( n15876 , n2707 );
nand ( n15877 , n15876 , n2668 );
nor ( n15878 , n15004 , n15877 );
not ( n15879 , n15878 );
not ( n15880 , n3311 );
nand ( n15881 , n15880 , n2758 );
not ( n15882 , n15881 );
nor ( n15883 , n14986 , n2706 );
nor ( n15884 , n15882 , n15883 );
not ( n15885 , n15884 );
or ( n15886 , n15879 , n15885 );
not ( n15887 , n2604 );
not ( n15888 , n2746 );
or ( n15889 , n15887 , n15888 );
nand ( n15890 , n15889 , n2758 );
nand ( n15891 , n15890 , n2609 );
nand ( n15892 , n15886 , n15891 );
nor ( n15893 , n3301 , n2640 );
nand ( n15894 , n15893 , n2595 );
nand ( n15895 , n15892 , n15894 );
and ( n15896 , n15875 , n15895 );
not ( n15897 , n2752 );
or ( n15898 , n15825 , n15897 );
or ( n15899 , n3310 , n15023 );
nand ( n15900 , n15898 , n15899 );
nor ( n15901 , n15896 , n15900 );
nand ( n15902 , n15868 , n15901 );
not ( n15903 , n15902 );
not ( n15904 , n15903 );
not ( n15905 , n2767 );
or ( n15906 , n15904 , n15905 );
or ( n15907 , n15903 , n2767 );
nand ( n15908 , n15906 , n15907 );
nor ( n15909 , n15112 , n126 );
not ( n15910 , n15909 );
not ( n15911 , n2959 );
nor ( n15912 , n15910 , n15911 );
nand ( n15913 , n9861 , n14809 );
not ( n15914 , n9904 );
and ( n15915 , n15913 , n15914 , n126 );
or ( n15916 , n15912 , n15915 );
and ( n15917 , n15072 , n127 );
not ( n15918 , n2888 );
nand ( n15919 , n14836 , n15918 , n2990 );
and ( n15920 , n15919 , n2861 );
nor ( n15921 , n2988 , n2893 );
nor ( n15922 , n15920 , n15921 );
nand ( n15923 , n15916 , n15917 , n15922 );
not ( n15924 , n9921 );
not ( n15925 , n15914 );
or ( n15926 , n15924 , n15925 );
nand ( n15927 , n15137 , n2816 );
nand ( n15928 , n15926 , n15927 );
not ( n15929 , n2894 );
nand ( n15930 , n3011 , n15929 );
nor ( n15931 , n15413 , n15930 );
and ( n15932 , n15928 , n15931 );
and ( n15933 , n9921 , n120 );
nor ( n15934 , n15932 , n15933 );
or ( n15935 , n15923 , n15934 );
or ( n15936 , n2900 , n2802 );
or ( n15937 , n2893 , n121 );
nand ( n15938 , n15936 , n15937 );
nor ( n15939 , n9889 , n15938 );
not ( n15940 , n15939 );
not ( n15941 , n15909 );
or ( n15942 , n15940 , n15941 );
nand ( n15943 , n15942 , n2860 );
and ( n15944 , n2966 , n9896 );
nand ( n15945 , n15943 , n15944 );
not ( n15946 , n15945 );
not ( n15947 , n15112 );
nand ( n15948 , n14812 , n2886 );
and ( n15949 , n15947 , n14890 , n15948 );
nor ( n15950 , n2910 , n125 );
nand ( n15951 , n15373 , n14785 );
or ( n15952 , n15950 , n15951 );
not ( n15953 , n14886 );
or ( n15954 , n15953 , n2972 );
nand ( n15955 , n15952 , n15954 );
nand ( n15956 , n15949 , n15955 );
not ( n15957 , n15956 );
or ( n15958 , n15946 , n15957 );
or ( n15959 , n2861 , n14768 );
nand ( n15960 , n2949 , n2942 );
and ( n15961 , n15959 , n15960 );
nand ( n15962 , n2965 , n9907 );
nand ( n15963 , n2886 , n9903 );
and ( n15964 , n9981 , n15963 );
nand ( n15965 , n15962 , n15964 );
nor ( n15966 , n15961 , n15965 );
nand ( n15967 , n15958 , n15966 );
nand ( n15968 , n15935 , n15967 );
nand ( n15969 , n2966 , n9965 , n15104 , n2855 );
and ( n15970 , n15969 , n9928 );
not ( n15971 , n9951 );
or ( n15972 , n2966 , n15971 );
not ( n15973 , n2909 );
not ( n15974 , n9846 );
or ( n15975 , n15973 , n15974 );
nand ( n15976 , n15975 , n9981 );
and ( n15977 , n15976 , n2973 );
nor ( n15978 , n15977 , n2913 );
nand ( n15979 , n15972 , n15978 , n14888 );
nor ( n15980 , n15970 , n15979 );
nand ( n15981 , n2920 , n2902 );
nor ( n15982 , n15129 , n15981 );
not ( n15983 , n15982 );
not ( n15984 , n14785 );
not ( n15985 , n15984 );
and ( n15986 , n15983 , n15985 );
nand ( n15987 , n9992 , n14810 );
and ( n15988 , n15987 , n126 );
nor ( n15989 , n15986 , n15988 );
and ( n15990 , n15968 , n15980 , n15989 );
not ( n15991 , n15990 );
not ( n15992 , n15157 );
nor ( n15993 , n15992 , n3256 );
not ( n15994 , n15993 );
nand ( n15995 , n3244 , n10035 );
not ( n15996 , n3038 );
or ( n15997 , n15995 , n15996 );
nand ( n15998 , n3149 , n10037 );
or ( n15999 , n15476 , n15998 );
nand ( n16000 , n15997 , n15999 );
not ( n16001 , n16000 );
or ( n16002 , n15994 , n16001 );
nand ( n16003 , n10160 , n114 );
not ( n16004 , n16003 );
or ( n16005 , n16004 , n15497 );
nand ( n16006 , n16005 , n117 );
not ( n16007 , n115 );
nand ( n16008 , n116 , n114 );
nor ( n16009 , n16007 , n16008 , n112 );
nand ( n16010 , n3205 , n3190 );
or ( n16011 , n16009 , n16010 );
nand ( n16012 , n16011 , n10145 );
nand ( n16013 , n16006 , n16012 , n10101 , n10010 );
nand ( n16014 , n16002 , n16013 );
nand ( n16015 , n15157 , n10074 );
and ( n16016 , n16015 , n3094 );
not ( n16017 , n15478 );
not ( n16018 , n10075 );
or ( n16019 , n16017 , n16018 );
nand ( n16020 , n16019 , n3212 );
nand ( n16021 , n10148 , n10061 , n16020 , n3137 );
nor ( n16022 , n16016 , n16021 );
nand ( n16023 , n16014 , n16022 );
not ( n16024 , n16023 );
not ( n16025 , n3082 );
nand ( n16026 , n16025 , n115 );
nand ( n16027 , n16026 , n15197 );
not ( n16028 , n10048 );
not ( n16029 , n3027 );
or ( n16030 , n16028 , n16029 );
nand ( n16031 , n16030 , n3198 );
not ( n16032 , n16031 );
nand ( n16033 , n3176 , n3252 );
or ( n16034 , n16027 , n16032 , n16033 );
nand ( n16035 , n16034 , n3106 );
nand ( n16036 , n10045 , n116 );
nand ( n16037 , n15257 , n3092 );
nand ( n16038 , n16036 , n16037 );
nand ( n16039 , n16038 , n118 );
not ( n16040 , n3095 );
not ( n16041 , n16040 );
not ( n16042 , n16041 );
not ( n16043 , n10104 );
and ( n16044 , n16042 , n16043 );
not ( n16045 , n113 );
not ( n16046 , n3135 );
not ( n16047 , n16046 );
or ( n16048 , n16045 , n16047 );
nand ( n16049 , n16048 , n119 );
nor ( n16050 , n16044 , n16049 );
nand ( n16051 , n15257 , n3061 );
not ( n16052 , n16051 );
and ( n16053 , n3090 , n115 );
nor ( n16054 , n16053 , n15155 );
not ( n16055 , n16054 );
or ( n16056 , n16052 , n16055 );
nand ( n16057 , n16056 , n3235 );
and ( n16058 , n16039 , n16050 , n16057 );
nand ( n16059 , n15475 , n3230 );
or ( n16060 , n16027 , n16059 );
nand ( n16061 , n16060 , n3164 );
nand ( n16062 , n16035 , n16058 , n16061 );
not ( n16063 , n16062 );
or ( n16064 , n16024 , n16063 );
nand ( n16065 , n10046 , n10051 );
or ( n16066 , n10125 , n16065 );
nand ( n16067 , n16066 , n3212 );
not ( n16068 , n16067 );
not ( n16069 , n3106 );
or ( n16070 , n16068 , n16069 );
nor ( n16071 , n10101 , n3235 );
nand ( n16072 , n16070 , n16071 );
nor ( n16073 , n10064 , n116 );
and ( n16074 , n16073 , n10020 );
not ( n16075 , n3136 );
nor ( n16076 , n16074 , n16075 );
and ( n16077 , n16076 , n3124 );
nor ( n16078 , n16077 , n3042 );
nand ( n16079 , n15169 , n3199 );
and ( n16080 , n3052 , n3100 );
nand ( n16081 , n16080 , n15259 );
nand ( n16082 , n16079 , n16081 );
nor ( n16083 , n16078 , n16082 );
nor ( n16084 , n10099 , n3028 );
not ( n16085 , n16084 );
nand ( n16086 , n16085 , n10077 , n3056 );
and ( n16087 , n16086 , n10040 );
nand ( n16088 , n15170 , n3049 );
and ( n16089 , n16088 , n3106 );
nor ( n16090 , n16087 , n16089 );
not ( n16091 , n15225 );
not ( n16092 , n15200 );
not ( n16093 , n16092 );
not ( n16094 , n16037 );
or ( n16095 , n16093 , n16094 );
nand ( n16096 , n16095 , n116 );
not ( n16097 , n16096 );
or ( n16098 , n16091 , n16097 );
nand ( n16099 , n16098 , n3235 );
and ( n16100 , n16072 , n16083 , n16090 , n16099 );
nand ( n16101 , n16064 , n16100 );
not ( n16102 , n16101 );
and ( n16103 , n15991 , n16102 );
not ( n16104 , n15991 );
and ( n16105 , n16104 , n16101 );
nor ( n16106 , n16103 , n16105 );
and ( n16107 , n15908 , n16106 );
not ( n16108 , n15908 );
not ( n16109 , n16106 );
and ( n16110 , n16108 , n16109 );
nor ( n16111 , n16107 , n16110 );
and ( n16112 , n15793 , n16111 );
not ( n16113 , n15793 );
not ( n16114 , n16111 );
and ( n16115 , n16113 , n16114 );
nor ( n16116 , n16112 , n16115 );
or ( n16117 , n16116 , n1 );
xnor ( n16118 , n278 , n279 );
or ( n16119 , n2246 , n16118 );
nand ( n16120 , n16117 , n16119 );
and ( n16121 , n2541 , n14938 );
nand ( n16122 , n14933 , n2580 , n16121 );
not ( n16123 , n16122 );
not ( n16124 , n2686 );
or ( n16125 , n16123 , n16124 );
nor ( n16126 , n15883 , n2642 );
not ( n16127 , n16126 );
and ( n16128 , n14986 , n2635 , n2678 );
or ( n16129 , n16128 , n3284 );
or ( n16130 , n3416 , n14901 );
nand ( n16131 , n16129 , n16130 );
nor ( n16132 , n16127 , n16131 );
nand ( n16133 , n16125 , n16132 );
not ( n16134 , n14914 );
nand ( n16135 , n3333 , n16134 );
nand ( n16136 , n2539 , n16135 );
nor ( n16137 , n2746 , n141 );
or ( n16138 , n16136 , n16137 );
nand ( n16139 , n16138 , n142 );
not ( n16140 , n2753 );
nor ( n16141 , n16140 , n3317 );
and ( n16142 , n16139 , n16141 , n2712 );
not ( n16143 , n15821 );
nand ( n16144 , n2516 , n142 );
not ( n16145 , n16144 );
not ( n16146 , n140 );
and ( n16147 , n16145 , n16146 );
nand ( n16148 , n14974 , n144 );
nor ( n16149 , n16147 , n16148 );
and ( n16150 , n16143 , n16149 );
nor ( n16151 , n16142 , n16150 );
or ( n16152 , n16133 , n16151 );
nand ( n16153 , n14994 , n144 );
not ( n16154 , n2595 );
not ( n16155 , n2616 );
or ( n16156 , n16154 , n16155 );
or ( n16157 , n2589 , n2596 );
nand ( n16158 , n3277 , n16157 );
nor ( n16159 , n16158 , n2601 );
nand ( n16160 , n16156 , n16159 );
nor ( n16161 , n16153 , n16160 );
not ( n16162 , n16161 );
not ( n16163 , n16144 );
nor ( n16164 , n16163 , n141 );
not ( n16165 , n16164 );
not ( n16166 , n3301 );
not ( n16167 , n14969 );
or ( n16168 , n16166 , n16167 );
nand ( n16169 , n16168 , n2517 );
not ( n16170 , n16169 );
or ( n16171 , n16165 , n16170 );
nand ( n16172 , n15799 , n2659 , n141 );
nand ( n16173 , n16171 , n16172 );
not ( n16174 , n16173 );
or ( n16175 , n16162 , n16174 );
not ( n16176 , n15009 );
and ( n16177 , n2636 , n2639 );
nor ( n16178 , n16177 , n144 );
nand ( n16179 , n2522 , n3382 , n16176 , n16178 );
nand ( n16180 , n16175 , n16179 );
nor ( n16181 , n137 , n141 );
not ( n16182 , n16181 );
not ( n16183 , n3307 );
not ( n16184 , n16183 );
or ( n16185 , n16182 , n16184 );
not ( n16186 , n15869 );
nand ( n16187 , n3364 , n2578 );
nor ( n16188 , n15021 , n3425 );
nand ( n16189 , n16186 , n16187 , n16188 , n16157 );
nand ( n16190 , n16185 , n16189 );
nand ( n16191 , n16180 , n16190 , n2637 );
nand ( n16192 , n16152 , n16191 );
not ( n16193 , n2654 );
nand ( n16194 , n3362 , n16193 );
not ( n16195 , n3367 );
nand ( n16196 , n16195 , n3288 );
nand ( n16197 , n3358 , n16194 , n15894 , n16196 );
nand ( n16198 , n15008 , n138 );
and ( n16199 , n3404 , n2683 , n16198 );
nor ( n16200 , n16199 , n2669 );
nor ( n16201 , n16197 , n16200 );
not ( n16202 , n3316 );
nand ( n16203 , n142 , n143 );
or ( n16204 , n16203 , n139 );
nand ( n16205 , n16204 , n3311 );
or ( n16206 , n16205 , n15015 );
nand ( n16207 , n16206 , n16134 );
not ( n16208 , n16207 );
or ( n16209 , n16202 , n16208 );
nand ( n16210 , n16209 , n3381 );
not ( n16211 , n3352 );
nor ( n16212 , n16211 , n15893 , n144 );
nand ( n16213 , n16210 , n16212 );
not ( n16214 , n14901 );
not ( n16215 , n15021 );
or ( n16216 , n16214 , n16215 );
or ( n16217 , n3347 , n2564 );
nand ( n16218 , n16217 , n2654 );
nand ( n16219 , n16216 , n16218 );
nand ( n16220 , n16213 , n16219 );
and ( n16221 , n16192 , n16201 , n16220 );
not ( n16222 , n16221 );
not ( n16223 , n10168 );
or ( n16224 , n16222 , n16223 );
not ( n16225 , n16221 );
nand ( n16226 , n10167 , n16225 );
nand ( n16227 , n16224 , n16226 );
not ( n16228 , n16227 );
not ( n16229 , n132 );
not ( n16230 , n10242 );
or ( n16231 , n16229 , n16230 );
not ( n16232 , n2486 );
nand ( n16233 , n16232 , n2357 );
not ( n16234 , n16233 );
nor ( n16235 , n16234 , n10297 );
nand ( n16236 , n16231 , n16235 );
not ( n16237 , n16236 );
not ( n16238 , n133 );
or ( n16239 , n16237 , n16238 );
not ( n16240 , n10204 );
nand ( n16241 , n16239 , n16240 );
not ( n16242 , n15555 );
nand ( n16243 , n16242 , n10182 , n2359 );
nor ( n16244 , n16241 , n16243 );
not ( n16245 , n16244 );
and ( n16246 , n2395 , n134 );
nand ( n16247 , n16246 , n14728 , n2451 );
not ( n16248 , n10223 );
not ( n16249 , n16248 );
not ( n16250 , n2334 );
or ( n16251 , n16249 , n16250 );
nand ( n16252 , n16251 , n133 );
not ( n16253 , n16252 );
nand ( n16254 , n2287 , n2342 );
not ( n16255 , n16254 );
not ( n16256 , n14647 );
or ( n16257 , n16255 , n16256 );
nand ( n16258 , n16257 , n2424 );
not ( n16259 , n16248 );
not ( n16260 , n10210 );
or ( n16261 , n16259 , n16260 );
nand ( n16262 , n16261 , n2292 );
nand ( n16263 , n10253 , n2294 );
nand ( n16264 , n16258 , n16262 , n16263 );
or ( n16265 , n16247 , n16253 , n16264 );
not ( n16266 , n10302 );
not ( n16267 , n2449 );
or ( n16268 , n16266 , n16267 );
nand ( n16269 , n16268 , n2496 );
not ( n16270 , n16269 );
or ( n16271 , n15612 , n134 );
nand ( n16272 , n16271 , n2431 );
nand ( n16273 , n16270 , n14704 , n16272 );
nand ( n16274 , n16265 , n16273 );
not ( n16275 , n16274 );
or ( n16276 , n16245 , n16275 );
not ( n16277 , n15573 );
not ( n16278 , n14750 );
nor ( n16279 , n16278 , n15603 , n2316 );
nand ( n16280 , n16277 , n16279 );
not ( n16281 , n16280 );
or ( n16282 , n14678 , n134 );
nand ( n16283 , n16282 , n2274 );
nand ( n16284 , n10250 , n2408 );
not ( n16285 , n16284 );
not ( n16286 , n2337 );
or ( n16287 , n16285 , n16286 );
nand ( n16288 , n16287 , n133 );
and ( n16289 , n16288 , n10179 );
nand ( n16290 , n16283 , n16289 , n2497 );
not ( n16291 , n16290 );
or ( n16292 , n16281 , n16291 );
not ( n16293 , n2298 );
nor ( n16294 , n16293 , n133 );
and ( n16295 , n10261 , n2437 , n10201 );
or ( n16296 , n16295 , n2321 );
not ( n16297 , n2353 );
not ( n16298 , n16297 );
not ( n16299 , n14656 );
or ( n16300 , n16298 , n16299 );
nand ( n16301 , n15564 , n131 );
and ( n16302 , n16301 , n2424 );
nand ( n16303 , n16300 , n16302 );
nand ( n16304 , n16296 , n16303 );
nand ( n16305 , n2373 , n15714 );
and ( n16306 , n16305 , n2285 );
nor ( n16307 , n16294 , n16304 , n16306 , n14660 );
nand ( n16308 , n16292 , n16307 );
nand ( n16309 , n16276 , n16308 );
and ( n16310 , n2410 , n2265 );
not ( n16311 , n16310 );
not ( n16312 , n10240 );
not ( n16313 , n10287 );
or ( n16314 , n16312 , n16313 );
nand ( n16315 , n16314 , n10263 );
not ( n16316 , n16315 );
not ( n16317 , n16316 );
or ( n16318 , n16311 , n16317 );
not ( n16319 , n2487 );
not ( n16320 , n2357 );
or ( n16321 , n16319 , n16320 );
nand ( n16322 , n16321 , n2275 );
nand ( n16323 , n16318 , n16322 );
and ( n16324 , n2491 , n2377 );
nor ( n16325 , n16324 , n15701 );
nand ( n16326 , n16323 , n16325 );
not ( n16327 , n15642 );
not ( n16328 , n2293 );
not ( n16329 , n14675 );
or ( n16330 , n16328 , n16329 );
nand ( n16331 , n16330 , n134 );
nor ( n16332 , n16327 , n16331 );
nand ( n16333 , n16242 , n16332 );
and ( n16334 , n16326 , n16333 );
not ( n16335 , n15540 );
nand ( n16336 , n16335 , n2357 , n134 );
nand ( n16337 , n2295 , n2474 );
nand ( n16338 , n16336 , n16337 , n14687 );
nor ( n16339 , n16334 , n16338 );
nand ( n16340 , n16309 , n16339 );
not ( n16341 , n16340 );
not ( n16342 , n16341 );
not ( n16343 , n280 );
and ( n16344 , n16342 , n16343 );
and ( n16345 , n16341 , n280 );
nor ( n16346 , n16344 , n16345 );
not ( n16347 , n16346 );
or ( n16348 , n16228 , n16347 );
or ( n16349 , n16346 , n16227 );
nand ( n16350 , n16348 , n16349 );
buf ( n16351 , n15283 );
and ( n16352 , n16350 , n16351 );
not ( n16353 , n16350 );
not ( n16354 , n16351 );
and ( n16355 , n16353 , n16354 );
nor ( n16356 , n16352 , n16355 );
or ( n16357 , n16356 , n1 );
xnor ( n16358 , n280 , n281 );
or ( n16359 , n2246 , n16358 );
nand ( n16360 , n16357 , n16359 );
not ( n16361 , n8606 );
not ( n16362 , n14199 );
or ( n16363 , n16361 , n16362 );
nand ( n16364 , n16363 , n7052 );
not ( n16365 , n8533 );
not ( n16366 , n13866 );
or ( n16367 , n16365 , n16366 );
nand ( n16368 , n16367 , n7197 );
and ( n16369 , n16368 , n7170 );
not ( n16370 , n7513 );
or ( n16371 , n9161 , n16370 );
nand ( n16372 , n16371 , n13900 , n6978 );
nor ( n16373 , n16369 , n16372 );
nand ( n16374 , n16364 , n16373 );
not ( n16375 , n16374 );
nor ( n16376 , n14215 , n8591 );
nand ( n16377 , n8619 , n16376 );
not ( n16378 , n16377 );
or ( n16379 , n16375 , n16378 );
nand ( n16380 , n7610 , n14 );
and ( n16381 , n13928 , n16380 , n9337 );
nand ( n16382 , n16379 , n16381 );
not ( n16383 , n16382 );
nor ( n16384 , n7205 , n7142 );
nor ( n16385 , n16384 , n7089 , n9288 );
not ( n16386 , n16385 );
not ( n16387 , n7566 );
not ( n16388 , n16387 );
or ( n16389 , n16386 , n16388 );
not ( n16390 , n9300 );
not ( n16391 , n7076 );
or ( n16392 , n16390 , n16391 );
nand ( n16393 , n16392 , n8569 );
and ( n16394 , n7156 , n7511 );
nand ( n16395 , n13869 , n7048 );
nand ( n16396 , n16393 , n16394 , n16395 , n7603 );
nand ( n16397 , n16389 , n16396 );
not ( n16398 , n7215 );
not ( n16399 , n7096 );
or ( n16400 , n16398 , n16399 );
nand ( n16401 , n16400 , n7616 );
nand ( n16402 , n16401 , n13864 );
and ( n16403 , n16402 , n13885 , n10 );
not ( n16404 , n7156 );
not ( n16405 , n9246 );
or ( n16406 , n16404 , n16405 );
nand ( n16407 , n16406 , n16 );
not ( n16408 , n8579 );
not ( n16409 , n7033 );
or ( n16410 , n16408 , n16409 , n13929 );
nand ( n16411 , n16410 , n7170 );
nand ( n16412 , n16397 , n16403 , n16407 , n16411 );
nor ( n16413 , n7165 , n10 );
and ( n16414 , n16413 , n14190 , n7128 );
nand ( n16415 , n7194 , n13 );
not ( n16416 , n16415 );
nor ( n16417 , n7525 , n7015 );
not ( n16418 , n16417 );
or ( n16419 , n16416 , n16418 );
nand ( n16420 , n16419 , n16 );
nand ( n16421 , n16414 , n16420 );
not ( n16422 , n16421 );
and ( n16423 , n9327 , n7108 , n7062 );
nand ( n16424 , n9134 , n7114 , n16423 );
or ( n16425 , n8585 , n16424 );
nand ( n16426 , n7543 , n7053 );
not ( n16427 , n9140 );
and ( n16428 , n9206 , n7018 );
nor ( n16429 , n16428 , n17 );
nand ( n16430 , n16427 , n16429 );
or ( n16431 , n16426 , n16430 );
nand ( n16432 , n16425 , n16431 );
nand ( n16433 , n16422 , n16432 );
nand ( n16434 , n16412 , n16433 );
nand ( n16435 , n16383 , n16434 );
not ( n16436 , n53 );
xor ( n16437 , n16435 , n16436 );
not ( n16438 , n13731 );
not ( n16439 , n7 );
not ( n16440 , n7447 );
or ( n16441 , n16439 , n16440 );
nand ( n16442 , n16441 , n7403 );
not ( n16443 , n16442 );
not ( n16444 , n7472 );
or ( n16445 , n16443 , n16444 );
nand ( n16446 , n7818 , n7337 );
and ( n16447 , n12299 , n7265 );
nand ( n16448 , n16446 , n16447 , n9096 );
nand ( n16449 , n16445 , n16448 );
not ( n16450 , n7295 );
not ( n16451 , n7679 );
or ( n16452 , n16450 , n16451 );
nand ( n16453 , n16452 , n6 );
not ( n16454 , n16453 );
nor ( n16455 , n16454 , n7343 );
nand ( n16456 , n16449 , n16455 , n14377 );
nand ( n16457 , n14374 , n7714 );
and ( n16458 , n7826 , n7271 );
nand ( n16459 , n7461 , n7457 );
nand ( n16460 , n16457 , n16458 , n9108 , n16459 );
nand ( n16461 , n16456 , n16460 );
nand ( n16462 , n9023 , n7265 );
nor ( n16463 , n9092 , n9 );
and ( n16464 , n9076 , n16463 );
not ( n16465 , n7416 );
not ( n16466 , n8770 );
or ( n16467 , n16465 , n16466 );
not ( n16468 , n7338 );
nand ( n16469 , n16467 , n16468 );
nand ( n16470 , n16469 , n7 );
not ( n16471 , n9051 );
nand ( n16472 , n16471 , n7457 );
and ( n16473 , n16462 , n16464 , n16470 , n16472 );
or ( n16474 , n12302 , n3 );
nor ( n16475 , n8875 , n7265 );
or ( n16476 , n14367 , n7385 );
nand ( n16477 , n16476 , n8794 , n7271 );
nor ( n16478 , n16475 , n16477 );
nand ( n16479 , n16474 , n16478 );
nand ( n16480 , n16479 , n7271 );
and ( n16481 , n16461 , n16473 , n16480 );
and ( n16482 , n9092 , n3 );
nor ( n16483 , n16482 , n7315 );
nand ( n16484 , n16483 , n16462 );
not ( n16485 , n16484 );
not ( n16486 , n16479 );
or ( n16487 , n16485 , n16486 );
nand ( n16488 , n7355 , n7403 );
nand ( n16489 , n7750 , n16488 , n8875 );
and ( n16490 , n7271 , n16489 );
not ( n16491 , n7271 );
nand ( n16492 , n7773 , n2 );
nand ( n16493 , n9463 , n7683 , n16492 );
and ( n16494 , n16491 , n16493 );
nor ( n16495 , n16490 , n16494 );
nand ( n16496 , n16487 , n16495 );
not ( n16497 , n7248 );
and ( n16498 , n7416 , n4 );
nor ( n16499 , n16498 , n7461 );
not ( n16500 , n16499 );
or ( n16501 , n16497 , n16500 );
nand ( n16502 , n16501 , n8 );
and ( n16503 , n7399 , n7325 , n9097 );
nand ( n16504 , n16502 , n16503 );
nor ( n16505 , n8760 , n16504 );
not ( n16506 , n8819 );
nor ( n16507 , n16506 , n12309 );
or ( n16508 , n16505 , n16507 );
not ( n16509 , n16475 );
nand ( n16510 , n7779 , n7350 );
and ( n16511 , n16509 , n9365 , n16510 );
nand ( n16512 , n16508 , n16511 );
nor ( n16513 , n16496 , n16512 );
or ( n16514 , n16481 , n16513 );
not ( n16515 , n8863 );
not ( n16516 , n9045 );
not ( n16517 , n16516 );
or ( n16518 , n16515 , n16517 );
not ( n16519 , n7814 );
nand ( n16520 , n7321 , n7232 );
and ( n16521 , n7399 , n16520 );
not ( n16522 , n16521 );
or ( n16523 , n16519 , n16522 );
nand ( n16524 , n16523 , n7811 );
nand ( n16525 , n16518 , n16524 );
not ( n16526 , n8822 );
not ( n16527 , n7687 );
or ( n16528 , n16526 , n16527 );
nand ( n16529 , n16528 , n7265 );
nand ( n16530 , n16529 , n8792 );
nor ( n16531 , n16525 , n16530 );
nand ( n16532 , n16514 , n16531 );
not ( n16533 , n16532 );
not ( n16534 , n16533 );
or ( n16535 , n16438 , n16534 );
nand ( n16536 , n16532 , n13730 );
nand ( n16537 , n16535 , n16536 );
xnor ( n16538 , n16437 , n16537 );
and ( n16539 , n14271 , n16538 );
not ( n16540 , n14271 );
not ( n16541 , n16538 );
and ( n16542 , n16540 , n16541 );
nor ( n16543 , n16539 , n16542 );
or ( n16544 , n16543 , n1 );
and ( n16545 , n54 , n16436 );
not ( n16546 , n54 );
and ( n16547 , n16546 , n53 );
nor ( n16548 , n16545 , n16547 );
or ( n16549 , n2246 , n16548 );
nand ( n16550 , n16544 , n16549 );
not ( n16551 , n3962 );
not ( n16552 , n5895 );
or ( n16553 , n16551 , n16552 );
or ( n16554 , n5895 , n3962 );
nand ( n16555 , n16553 , n16554 );
xor ( n16556 , n388 , n6271 );
not ( n16557 , n16556 );
and ( n16558 , n16555 , n16557 );
not ( n16559 , n16555 );
and ( n16560 , n16559 , n16556 );
nor ( n16561 , n16558 , n16560 );
or ( n16562 , n16561 , n1 );
xnor ( n16563 , n388 , n389 );
or ( n16564 , n2246 , n16563 );
nand ( n16565 , n16562 , n16564 );
nor ( n16566 , n4725 , n5003 );
and ( n16567 , n3812 , n16566 );
nor ( n16568 , n3714 , n12581 );
nor ( n16569 , n16567 , n16568 );
or ( n16570 , n16569 , n4930 );
not ( n16571 , n4841 );
not ( n16572 , n3806 );
or ( n16573 , n16571 , n16572 );
nand ( n16574 , n16573 , n4838 );
nand ( n16575 , n16570 , n16574 );
not ( n16576 , n16575 );
nand ( n16577 , n4797 , n4948 );
and ( n16578 , n9795 , n4977 , n16577 );
not ( n16579 , n16578 );
or ( n16580 , n16576 , n16579 );
nand ( n16581 , n16580 , n5007 );
not ( n16582 , n4889 );
nand ( n16583 , n16582 , n3949 );
nand ( n16584 , n3913 , n16583 );
not ( n16585 , n4994 );
and ( n16586 , n16585 , n3921 , n3765 );
nor ( n16587 , n16586 , n3922 );
or ( n16588 , n16584 , n16587 );
nand ( n16589 , n16588 , n187 );
not ( n16590 , n4722 );
nand ( n16591 , n16590 , n4855 );
and ( n16592 , n16591 , n3949 );
nor ( n16593 , n16592 , n5071 );
and ( n16594 , n16589 , n16593 );
not ( n16595 , n5052 );
not ( n16596 , n12578 );
or ( n16597 , n16595 , n16596 );
nand ( n16598 , n5436 , n12565 );
nand ( n16599 , n16597 , n16598 );
nor ( n16600 , n3750 , n4688 );
nand ( n16601 , n3949 , n3908 );
and ( n16602 , n4773 , n16600 , n16601 );
nand ( n16603 , n16599 , n16602 );
nor ( n16604 , n4660 , n3749 );
nand ( n16605 , n3903 , n16604 );
and ( n16606 , n4805 , n4727 );
nor ( n16607 , n16606 , n5007 );
nand ( n16608 , n16603 , n16605 , n16607 );
not ( n16609 , n4835 );
not ( n16610 , n185 );
not ( n16611 , n12581 );
or ( n16612 , n16610 , n16611 );
nand ( n16613 , n3731 , n4739 );
or ( n16614 , n16613 , n4741 );
nand ( n16615 , n16614 , n3811 );
nand ( n16616 , n16612 , n16615 );
not ( n16617 , n16616 );
or ( n16618 , n16609 , n16617 );
not ( n16619 , n12593 );
nor ( n16620 , n3733 , n12638 );
nor ( n16621 , n16619 , n16620 );
nand ( n16622 , n16618 , n16621 );
not ( n16623 , n3858 );
not ( n16624 , n4659 );
or ( n16625 , n16623 , n16624 );
nand ( n16626 , n3888 , n3749 );
nand ( n16627 , n16625 , n16626 );
nand ( n16628 , n3712 , n3860 , n180 );
nand ( n16629 , n4873 , n16627 , n9791 , n16628 );
or ( n16630 , n3811 , n4658 );
nand ( n16631 , n16630 , n3948 );
nand ( n16632 , n4838 , n4689 , n16631 );
nand ( n16633 , n16629 , n16632 );
not ( n16634 , n5461 );
nand ( n16635 , n16633 , n16634 );
nand ( n16636 , n16622 , n16635 );
nand ( n16637 , n16581 , n16594 , n16608 , n16636 );
xor ( n16638 , n16637 , n11427 );
not ( n16639 , n5392 );
not ( n16640 , n13210 );
or ( n16641 , n16639 , n16640 );
nand ( n16642 , n13205 , n5393 );
nand ( n16643 , n16641 , n16642 );
xnor ( n16644 , n16638 , n16643 );
not ( n16645 , n98 );
not ( n16646 , n195 );
nor ( n16647 , n6195 , n5609 );
not ( n16648 , n12765 );
nand ( n16649 , n16648 , n4402 );
nand ( n16650 , n6113 , n4437 );
nand ( n16651 , n5495 , n16647 , n16649 , n16650 );
not ( n16652 , n4390 );
not ( n16653 , n6187 );
or ( n16654 , n16652 , n16653 );
nand ( n16655 , n16654 , n5598 );
or ( n16656 , n16651 , n16655 );
and ( n16657 , n14484 , n4413 );
and ( n16658 , n5527 , n4379 );
nor ( n16659 , n16657 , n16658 );
or ( n16660 , n4396 , n4604 );
nand ( n16661 , n16660 , n6248 );
nand ( n16662 , n16659 , n16661 );
nand ( n16663 , n16656 , n16662 );
not ( n16664 , n4510 );
not ( n16665 , n4442 );
or ( n16666 , n16664 , n16665 , n4502 );
nand ( n16667 , n16666 , n5554 );
not ( n16668 , n4438 );
nor ( n16669 , n5621 , n16668 , n5569 );
nand ( n16670 , n16663 , n16667 , n16669 );
not ( n16671 , n16670 );
or ( n16672 , n16646 , n16671 );
not ( n16673 , n4415 );
not ( n16674 , n4475 );
not ( n16675 , n4401 );
or ( n16676 , n16674 , n16675 );
nand ( n16677 , n16676 , n193 );
nor ( n16678 , n4479 , n193 );
nand ( n16679 , n6093 , n16678 );
nand ( n16680 , n16677 , n16679 );
or ( n16681 , n16680 , n6052 );
nand ( n16682 , n4576 , n6140 );
nor ( n16683 , n4412 , n4478 );
or ( n16684 , n16682 , n16683 );
nand ( n16685 , n16681 , n16684 );
not ( n16686 , n5554 );
not ( n16687 , n6187 );
or ( n16688 , n16686 , n16687 );
nand ( n16689 , n16688 , n14445 );
nor ( n16690 , n12732 , n16689 );
nand ( n16691 , n16685 , n16690 );
not ( n16692 , n16691 );
or ( n16693 , n16673 , n16692 );
and ( n16694 , n5564 , n4396 );
and ( n16695 , n4397 , n4546 );
nor ( n16696 , n16694 , n16695 );
nand ( n16697 , n16693 , n16696 );
not ( n16698 , n5594 );
and ( n16699 , n16698 , n4639 );
nor ( n16700 , n16699 , n4390 );
nand ( n16701 , n11193 , n16700 );
or ( n16702 , n16701 , n12720 );
or ( n16703 , n4565 , n12763 , n193 );
nand ( n16704 , n16702 , n16703 );
not ( n16705 , n11279 );
nor ( n16706 , n16705 , n12742 );
and ( n16707 , n16704 , n16706 );
not ( n16708 , n4492 );
nand ( n16709 , n16708 , n192 );
not ( n16710 , n14453 );
nand ( n16711 , n16709 , n6124 , n5625 , n16710 );
or ( n16712 , n14442 , n16711 );
nand ( n16713 , n4439 , n4492 , n6140 , n193 );
nand ( n16714 , n16712 , n16713 );
nor ( n16715 , n5498 , n194 );
and ( n16716 , n16714 , n16715 );
nor ( n16717 , n16707 , n16716 );
nor ( n16718 , n16697 , n16717 );
nand ( n16719 , n16672 , n16718 );
not ( n16720 , n16719 );
not ( n16721 , n16720 );
or ( n16722 , n16645 , n16721 );
not ( n16723 , n98 );
nand ( n16724 , n16719 , n16723 );
nand ( n16725 , n16722 , n16724 );
and ( n16726 , n16725 , n11293 );
not ( n16727 , n16725 );
and ( n16728 , n16727 , n11294 );
nor ( n16729 , n16726 , n16728 );
and ( n16730 , n16644 , n16729 );
not ( n16731 , n16644 );
not ( n16732 , n16729 );
and ( n16733 , n16731 , n16732 );
nor ( n16734 , n16730 , n16733 );
or ( n16735 , n16734 , n1 );
and ( n16736 , n315 , n16723 );
not ( n16737 , n315 );
and ( n16738 , n16737 , n98 );
nor ( n16739 , n16736 , n16738 );
or ( n16740 , n2246 , n16739 );
nand ( n16741 , n16735 , n16740 );
not ( n16742 , n316 );
and ( n16743 , n11288 , n16742 );
not ( n16744 , n11288 );
and ( n16745 , n16744 , n316 );
nor ( n16746 , n16743 , n16745 );
xor ( n16747 , n16746 , n11429 );
not ( n16748 , n13205 );
not ( n16749 , n16748 );
not ( n16750 , n4363 );
or ( n16751 , n16749 , n16750 );
not ( n16752 , n5395 );
or ( n16753 , n16752 , n16748 );
nand ( n16754 , n16751 , n16753 );
not ( n16755 , n16754 );
and ( n16756 , n3691 , n9636 , n4258 );
nand ( n16757 , n3598 , n3677 );
and ( n16758 , n5912 , n16757 , n3636 );
nor ( n16759 , n16756 , n16758 );
not ( n16760 , n9642 );
not ( n16761 , n3547 );
nor ( n16762 , n16761 , n11387 );
nand ( n16763 , n16760 , n16762 );
or ( n16764 , n16759 , n16763 );
not ( n16765 , n5298 );
and ( n16766 , n12512 , n4273 , n5980 );
not ( n16767 , n16766 );
or ( n16768 , n16765 , n16767 );
nand ( n16769 , n5990 , n5376 );
nand ( n16770 , n16768 , n16769 );
not ( n16771 , n16770 );
nand ( n16772 , n16764 , n16771 );
not ( n16773 , n16772 );
nand ( n16774 , n3567 , n4229 , n4221 );
nand ( n16775 , n16774 , n3630 );
nor ( n16776 , n3704 , n4236 );
and ( n16777 , n3650 , n11329 , n16775 , n16776 );
not ( n16778 , n16777 );
or ( n16779 , n16773 , n16778 );
not ( n16780 , n3700 );
not ( n16781 , n209 );
and ( n16782 , n16780 , n16781 );
nand ( n16783 , n4337 , n9645 , n4236 );
nor ( n16784 , n16782 , n16783 );
not ( n16785 , n11323 );
and ( n16786 , n9699 , n3609 );
nor ( n16787 , n16786 , n3552 );
not ( n16788 , n16787 );
and ( n16789 , n16785 , n16788 );
not ( n16790 , n209 );
not ( n16791 , n3689 );
or ( n16792 , n16790 , n16791 );
nand ( n16793 , n16792 , n3629 );
and ( n16794 , n16793 , n5947 );
nor ( n16795 , n16789 , n16794 );
or ( n16796 , n16795 , n4243 );
and ( n16797 , n3489 , n3619 );
nor ( n16798 , n16797 , n3663 );
not ( n16799 , n4340 );
or ( n16800 , n16798 , n16799 );
nand ( n16801 , n16796 , n16800 );
nand ( n16802 , n16784 , n16801 );
nand ( n16803 , n16779 , n16802 );
not ( n16804 , n3657 );
nand ( n16805 , n16804 , n4217 , n9702 );
or ( n16806 , n16805 , n9642 );
nand ( n16807 , n5937 , n4340 , n5258 , n209 );
nand ( n16808 , n16806 , n16807 );
not ( n16809 , n3670 );
not ( n16810 , n5912 );
or ( n16811 , n16809 , n16810 );
nand ( n16812 , n16811 , n3468 );
and ( n16813 , n16808 , n16812 );
nor ( n16814 , n16813 , n211 );
not ( n16815 , n5351 );
and ( n16816 , n5939 , n3632 );
nor ( n16817 , n16816 , n3696 );
nor ( n16818 , n16815 , n16817 );
not ( n16819 , n210 );
not ( n16820 , n5363 );
or ( n16821 , n16819 , n16820 );
not ( n16822 , n3582 );
not ( n16823 , n5953 );
or ( n16824 , n16822 , n16823 );
nand ( n16825 , n16824 , n206 );
nand ( n16826 , n16821 , n16825 );
and ( n16827 , n16826 , n5376 );
nor ( n16828 , n5252 , n3619 );
nor ( n16829 , n16827 , n16828 );
not ( n16830 , n5932 );
nand ( n16831 , n5972 , n3467 );
and ( n16832 , n5318 , n16831 );
not ( n16833 , n16832 );
or ( n16834 , n16830 , n16833 );
nand ( n16835 , n16834 , n5980 );
nand ( n16836 , n16818 , n16829 , n16835 );
nor ( n16837 , n16814 , n16836 );
nand ( n16838 , n16803 , n16837 );
not ( n16839 , n16838 );
not ( n16840 , n16637 );
and ( n16841 , n16839 , n16840 );
and ( n16842 , n16838 , n16637 );
nor ( n16843 , n16841 , n16842 );
not ( n16844 , n16843 );
or ( n16845 , n16755 , n16844 );
not ( n16846 , n16754 );
not ( n16847 , n16843 );
nand ( n16848 , n16846 , n16847 );
nand ( n16849 , n16845 , n16848 );
xnor ( n16850 , n16747 , n16849 );
or ( n16851 , n16850 , n1 );
and ( n16852 , n317 , n16742 );
not ( n16853 , n317 );
and ( n16854 , n16853 , n316 );
nor ( n16855 , n16852 , n16854 );
or ( n16856 , n2246 , n16855 );
nand ( n16857 , n16851 , n16856 );
not ( n16858 , n11827 );
not ( n16859 , n11577 );
and ( n16860 , n16858 , n16859 );
and ( n16861 , n11827 , n11577 );
nor ( n16862 , n16860 , n16861 );
and ( n16863 , n11048 , n318 );
not ( n16864 , n11048 );
not ( n16865 , n318 );
and ( n16866 , n16864 , n16865 );
nor ( n16867 , n16863 , n16866 );
xor ( n16868 , n16862 , n16867 );
and ( n16869 , n10654 , n13487 );
not ( n16870 , n10654 );
and ( n16871 , n16870 , n13601 );
or ( n16872 , n16869 , n16871 );
not ( n16873 , n1344 );
nand ( n16874 , n16873 , n1408 );
nand ( n16875 , n1525 , n1504 );
nand ( n16876 , n16874 , n16875 );
not ( n16877 , n16876 );
not ( n16878 , n13017 );
and ( n16879 , n16877 , n16878 );
nor ( n16880 , n16879 , n176 );
nand ( n16881 , n1376 , n1442 );
or ( n16882 , n16881 , n11852 );
not ( n16883 , n1338 );
not ( n16884 , n1302 );
or ( n16885 , n16883 , n16884 );
nand ( n16886 , n16885 , n177 );
not ( n16887 , n16886 );
nand ( n16888 , n1363 , n1503 );
nand ( n16889 , n1459 , n1289 );
nand ( n16890 , n16887 , n16888 , n16889 , n16875 );
nand ( n16891 , n16882 , n16890 );
and ( n16892 , n1460 , n10462 );
not ( n16893 , n13421 );
not ( n16894 , n10441 );
not ( n16895 , n16894 );
not ( n16896 , n1275 );
or ( n16897 , n16895 , n16896 );
nand ( n16898 , n16897 , n10419 );
nand ( n16899 , n16893 , n16898 );
nor ( n16900 , n16892 , n16899 );
nand ( n16901 , n16891 , n16900 );
or ( n16902 , n16880 , n16901 );
and ( n16903 , n16875 , n178 );
nor ( n16904 , n16903 , n13407 );
nand ( n16905 , n16902 , n16904 );
nor ( n16906 , n10444 , n1339 );
nor ( n16907 , n10473 , n1422 , n16906 );
not ( n16908 , n16907 );
not ( n16909 , n1306 );
not ( n16910 , n10415 );
or ( n16911 , n16909 , n16910 );
nand ( n16912 , n16911 , n1521 );
not ( n16913 , n16912 );
not ( n16914 , n16913 );
or ( n16915 , n16908 , n16914 );
nand ( n16916 , n11882 , n1370 );
nand ( n16917 , n1349 , n1432 );
or ( n16918 , n16916 , n16917 , n11852 );
nand ( n16919 , n16918 , n1375 );
nand ( n16920 , n16919 , n10460 );
nand ( n16921 , n16915 , n16920 );
nand ( n16922 , n16905 , n16921 );
not ( n16923 , n16922 );
not ( n16924 , n12988 );
not ( n16925 , n1513 );
or ( n16926 , n16924 , n16925 );
nand ( n16927 , n16926 , n11904 );
not ( n16928 , n16927 );
not ( n16929 , n10464 );
nand ( n16930 , n10523 , n10481 );
nor ( n16931 , n16929 , n16930 , n1286 );
not ( n16932 , n16931 );
or ( n16933 , n16928 , n16932 );
nand ( n16934 , n16933 , n176 );
or ( n16935 , n13422 , n10517 );
nand ( n16936 , n16935 , n1280 );
or ( n16937 , n1493 , n10452 );
nand ( n16938 , n16937 , n1473 );
and ( n16939 , n1454 , n10360 , n16936 , n16938 );
nand ( n16940 , n16934 , n16939 );
nand ( n16941 , n11911 , n1337 , n11894 );
nand ( n16942 , n16941 , n176 );
not ( n16943 , n13400 );
and ( n16944 , n16943 , n173 );
not ( n16945 , n175 );
not ( n16946 , n1397 );
or ( n16947 , n16945 , n16946 );
nand ( n16948 , n16947 , n1278 );
nand ( n16949 , n16948 , n13384 , n1370 );
nor ( n16950 , n16944 , n16949 );
and ( n16951 , n16942 , n16950 );
nand ( n16952 , n1329 , n177 );
or ( n16953 , n16952 , n1361 );
nand ( n16954 , n16953 , n1434 );
not ( n16955 , n10415 );
and ( n16956 , n16954 , n16955 );
nor ( n16957 , n16951 , n16956 );
or ( n16958 , n16940 , n16957 );
or ( n16959 , n16927 , n1280 );
nand ( n16960 , n16959 , n1350 );
nand ( n16961 , n16958 , n16960 );
nand ( n16962 , n16923 , n16961 );
not ( n16963 , n16962 );
not ( n16964 , n16963 );
not ( n16965 , n11680 );
not ( n16966 , n16965 );
or ( n16967 , n16964 , n16966 );
nand ( n16968 , n11680 , n16962 );
nand ( n16969 , n16967 , n16968 );
not ( n16970 , n16969 );
and ( n16971 , n16872 , n16970 );
not ( n16972 , n16872 );
and ( n16973 , n16972 , n16969 );
nor ( n16974 , n16971 , n16973 );
and ( n16975 , n16868 , n16974 );
not ( n16976 , n16868 );
not ( n16977 , n16974 );
and ( n16978 , n16976 , n16977 );
nor ( n16979 , n16975 , n16978 );
or ( n16980 , n16979 , n1 );
and ( n16981 , n319 , n16865 );
not ( n16982 , n319 );
and ( n16983 , n16982 , n318 );
nor ( n16984 , n16981 , n16983 );
or ( n16985 , n2246 , n16984 );
nand ( n16986 , n16980 , n16985 );
not ( n16987 , n5889 );
not ( n16988 , n4366 );
or ( n16989 , n16987 , n16988 );
not ( n16990 , n5889 );
not ( n16991 , n16990 );
or ( n16992 , n16991 , n16752 );
nand ( n16993 , n16989 , n16992 );
not ( n16994 , n16993 );
not ( n16995 , n11115 );
or ( n16996 , n16994 , n16995 );
not ( n16997 , n16993 );
nand ( n16998 , n16997 , n11114 );
nand ( n16999 , n16996 , n16998 );
not ( n17000 , n6268 );
not ( n17001 , n328 );
and ( n17002 , n17000 , n17001 );
and ( n17003 , n6268 , n328 );
nor ( n17004 , n17002 , n17003 );
not ( n17005 , n17004 );
and ( n17006 , n16999 , n17005 );
not ( n17007 , n16999 );
and ( n17008 , n17007 , n17004 );
nor ( n17009 , n17006 , n17008 );
or ( n17010 , n17009 , n1 );
xnor ( n17011 , n328 , n329 );
or ( n17012 , n2246 , n17011 );
nand ( n17013 , n17010 , n17012 );
not ( n17014 , n12882 );
not ( n17015 , n17014 );
and ( n17016 , n1209 , n1145 );
not ( n17017 , n17016 );
and ( n17018 , n1127 , n805 );
nand ( n17019 , n916 , n746 );
and ( n17020 , n17019 , n779 );
nand ( n17021 , n17018 , n17020 );
nand ( n17022 , n1246 , n1001 );
or ( n17023 , n17021 , n17022 );
not ( n17024 , n167 );
not ( n17025 , n814 );
or ( n17026 , n17024 , n17025 );
nand ( n17027 , n17026 , n1018 );
nand ( n17028 , n1132 , n10550 , n17027 );
nand ( n17029 , n17023 , n17028 );
not ( n17030 , n17029 );
or ( n17031 , n17017 , n17030 );
or ( n17032 , n10590 , n10663 );
nand ( n17033 , n17032 , n805 );
nor ( n17034 , n10577 , n779 );
nand ( n17035 , n17033 , n17034 );
nand ( n17036 , n17031 , n17035 );
not ( n17037 , n1220 );
nor ( n17038 , n1180 , n164 );
not ( n17039 , n1062 );
nand ( n17040 , n10667 , n17039 );
or ( n17041 , n17038 , n17040 );
nand ( n17042 , n17041 , n881 );
not ( n17043 , n17042 );
or ( n17044 , n17037 , n17043 );
nand ( n17045 , n17044 , n167 );
and ( n17046 , n17045 , n981 );
and ( n17047 , n17036 , n17046 );
not ( n17048 , n1194 );
not ( n17049 , n1127 );
nor ( n17050 , n17049 , n980 );
not ( n17051 , n17050 );
or ( n17052 , n17048 , n17051 );
nand ( n17053 , n17052 , n737 );
not ( n17054 , n10546 );
nand ( n17055 , n1040 , n898 );
or ( n17056 , n17054 , n17055 );
nand ( n17057 , n17056 , n953 );
and ( n17058 , n17053 , n17057 , n170 );
nand ( n17059 , n1019 , n770 );
and ( n17060 , n944 , n17059 , n1159 , n779 );
not ( n17061 , n17060 );
nand ( n17062 , n1246 , n10671 );
not ( n17063 , n784 );
not ( n17064 , n10667 );
or ( n17065 , n17063 , n17064 );
nand ( n17066 , n17065 , n920 );
nand ( n17067 , n1194 , n17066 );
nor ( n17068 , n17062 , n17067 );
not ( n17069 , n17068 );
or ( n17070 , n17061 , n17069 );
not ( n17071 , n167 );
not ( n17072 , n10632 );
or ( n17073 , n17071 , n17072 );
nand ( n17074 , n931 , n972 , n920 );
nand ( n17075 , n17073 , n17074 );
nand ( n17076 , n17075 , n10737 , n169 );
nand ( n17077 , n17070 , n17076 );
nand ( n17078 , n17058 , n17077 );
not ( n17079 , n1132 );
not ( n17080 , n10736 );
not ( n17081 , n17018 );
or ( n17082 , n17080 , n17081 );
nand ( n17083 , n1105 , n873 );
nand ( n17084 , n17082 , n17083 );
not ( n17085 , n17084 );
or ( n17086 , n17079 , n17085 );
not ( n17087 , n17018 );
nand ( n17088 , n17087 , n17083 );
not ( n17089 , n737 );
not ( n17090 , n782 );
or ( n17091 , n17089 , n17090 );
nand ( n17092 , n17091 , n1180 );
or ( n17093 , n17092 , n749 );
not ( n17094 , n1254 );
not ( n17095 , n934 );
or ( n17096 , n17094 , n17095 );
nand ( n17097 , n17096 , n756 );
nand ( n17098 , n17093 , n17097 );
nand ( n17099 , n17088 , n17098 , n1007 );
nand ( n17100 , n17086 , n17099 );
not ( n17101 , n982 );
and ( n17102 , n17101 , n1050 );
nand ( n17103 , n17100 , n17102 );
nand ( n17104 , n17078 , n17103 );
nand ( n17105 , n17047 , n17104 );
buf ( n17106 , n17105 );
not ( n17107 , n17106 );
not ( n17108 , n17107 );
and ( n17109 , n17015 , n17108 );
buf ( n17110 , n17014 );
and ( n17111 , n17110 , n17107 );
nor ( n17112 , n17109 , n17111 );
not ( n17113 , n17112 );
not ( n17114 , n338 );
and ( n17115 , n17114 , n2228 );
not ( n17116 , n17114 );
and ( n17117 , n17116 , n2232 );
nor ( n17118 , n17115 , n17117 );
buf ( n17119 , n13584 );
xor ( n17120 , n17118 , n17119 );
not ( n17121 , n17120 );
or ( n17122 , n17113 , n17121 );
or ( n17123 , n17112 , n17120 );
nand ( n17124 , n17122 , n17123 );
not ( n17125 , n13494 );
nand ( n17126 , n17125 , n2246 );
or ( n17127 , n17124 , n17126 );
and ( n17128 , n339 , n17114 );
not ( n17129 , n339 );
and ( n17130 , n17129 , n338 );
nor ( n17131 , n17128 , n17130 );
or ( n17132 , n17131 , n2246 );
nor ( n17133 , n17125 , n1 );
nand ( n17134 , n17124 , n17133 );
nand ( n17135 , n17127 , n17132 , n17134 );
not ( n17136 , n16102 );
not ( n17137 , n2686 );
nor ( n17138 , n16157 , n14901 );
nor ( n17139 , n17138 , n3305 );
not ( n17140 , n17139 );
or ( n17141 , n17137 , n17140 );
nand ( n17142 , n17141 , n144 );
not ( n17143 , n17142 );
not ( n17144 , n2660 );
and ( n17145 , n2632 , n15825 , n17144 , n2556 );
not ( n17146 , n17145 );
or ( n17147 , n17143 , n17146 );
and ( n17148 , n2554 , n140 );
nor ( n17149 , n17148 , n15848 );
and ( n17150 , n17149 , n2715 , n141 );
nor ( n17151 , n17150 , n2609 );
nand ( n17152 , n17147 , n17151 );
nand ( n17153 , n3274 , n2569 );
not ( n17154 , n17153 );
not ( n17155 , n2632 );
or ( n17156 , n17154 , n17155 );
nand ( n17157 , n17156 , n2517 );
buf ( n17158 , n3277 );
nor ( n17159 , n17158 , n142 );
nor ( n17160 , n16144 , n2752 );
not ( n17161 , n2682 );
not ( n17162 , n2762 );
or ( n17163 , n17161 , n17162 );
nand ( n17164 , n17163 , n2556 );
or ( n17165 , n17159 , n17160 , n17164 );
nand ( n17166 , n17165 , n2564 );
and ( n17167 , n17157 , n17166 , n137 );
nand ( n17168 , n17152 , n17167 );
not ( n17169 , n17168 );
or ( n17170 , n3311 , n2651 );
and ( n17171 , n14998 , n17170 , n2564 );
not ( n17172 , n17171 );
nand ( n17173 , n3345 , n3275 );
nand ( n17174 , n15820 , n2686 );
or ( n17175 , n17173 , n17174 );
not ( n17176 , n15825 );
not ( n17177 , n14939 );
not ( n17178 , n17177 );
nand ( n17179 , n17178 , n141 );
or ( n17180 , n17176 , n17179 );
nand ( n17181 , n17175 , n17180 );
not ( n17182 , n17181 );
or ( n17183 , n17172 , n17182 );
not ( n17184 , n2601 );
nand ( n17185 , n17184 , n144 );
not ( n17186 , n17185 );
nand ( n17187 , n2554 , n2682 );
and ( n17188 , n2518 , n17187 , n2635 );
nand ( n17189 , n17188 , n14998 );
or ( n17190 , n17174 , n17189 );
nand ( n17191 , n3413 , n141 );
or ( n17192 , n15009 , n17191 );
nand ( n17193 , n17190 , n17192 );
nand ( n17194 , n17186 , n16121 , n17193 );
nand ( n17195 , n17183 , n17194 );
and ( n17196 , n3381 , n2555 );
nor ( n17197 , n17196 , n137 );
and ( n17198 , n15894 , n3382 , n17197 , n3352 );
nand ( n17199 , n17195 , n17198 );
not ( n17200 , n17199 );
or ( n17201 , n17169 , n17200 );
not ( n17202 , n3317 );
not ( n17203 , n2746 );
not ( n17204 , n16187 );
or ( n17205 , n17203 , n17204 );
nand ( n17206 , n17205 , n2517 );
nand ( n17207 , n17202 , n17206 );
not ( n17208 , n17207 );
not ( n17209 , n2609 );
or ( n17210 , n17208 , n17209 );
not ( n17211 , n14968 );
not ( n17212 , n17211 );
not ( n17213 , n2637 );
or ( n17214 , n17212 , n17213 );
nand ( n17215 , n17214 , n2639 );
nand ( n17216 , n17210 , n17215 );
not ( n17217 , n3293 );
not ( n17218 , n14984 );
or ( n17219 , n17217 , n17218 );
nand ( n17220 , n17219 , n2564 );
buf ( n17221 , n2649 );
nand ( n17222 , n14974 , n17221 , n2674 );
nand ( n17223 , n17222 , n2668 );
nand ( n17224 , n17220 , n17223 );
nor ( n17225 , n17216 , n17224 );
or ( n17226 , n3305 , n15027 );
nand ( n17227 , n17226 , n142 );
not ( n17228 , n17227 );
not ( n17229 , n3406 );
or ( n17230 , n17228 , n17229 );
nand ( n17231 , n17230 , n16193 );
not ( n17232 , n3284 );
nand ( n17233 , n17184 , n3327 );
nor ( n17234 , n17159 , n17233 );
nand ( n17235 , n17234 , n2637 , n3298 );
nand ( n17236 , n17232 , n17235 );
and ( n17237 , n17225 , n17231 , n17236 );
nand ( n17238 , n17201 , n17237 );
not ( n17239 , n17238 );
not ( n17240 , n17239 );
or ( n17241 , n17136 , n17240 );
nand ( n17242 , n17238 , n16101 );
nand ( n17243 , n17241 , n17242 );
buf ( n17244 , n14838 );
and ( n17245 , n15912 , n17244 );
or ( n17246 , n17245 , n2861 );
nand ( n17247 , n17246 , n9921 );
nand ( n17248 , n2948 , n2922 );
not ( n17249 , n17248 );
nand ( n17250 , n9932 , n14785 );
nor ( n17251 , n9848 , n17250 );
not ( n17252 , n17251 );
or ( n17253 , n17249 , n17252 );
and ( n17254 , n2958 , n121 );
nor ( n17255 , n17254 , n2972 );
nand ( n17256 , n15947 , n2980 , n17255 );
nand ( n17257 , n17253 , n17256 );
nand ( n17258 , n17257 , n2951 );
and ( n17259 , n17247 , n17258 );
not ( n17260 , n9875 );
not ( n17261 , n9887 );
not ( n17262 , n15418 );
and ( n17263 , n17261 , n17262 );
and ( n17264 , n2843 , n2956 );
nor ( n17265 , n17263 , n17264 );
not ( n17266 , n17265 );
or ( n17267 , n17260 , n17266 );
nand ( n17268 , n17267 , n2861 );
nand ( n17269 , n14869 , n17268 , n15039 );
nor ( n17270 , n17259 , n17269 );
and ( n17271 , n9912 , n2886 );
nor ( n17272 , n17271 , n14864 );
and ( n17273 , n9877 , n15104 , n17272 );
nor ( n17274 , n15042 , n14859 );
or ( n17275 , n15077 , n9898 );
nand ( n17276 , n17275 , n2843 );
nand ( n17277 , n17273 , n17274 , n17276 );
not ( n17278 , n17277 );
nor ( n17279 , n9889 , n126 );
nand ( n17280 , n9879 , n17279 , n9937 );
not ( n17281 , n17280 );
not ( n17282 , n2860 );
or ( n17283 , n17281 , n17282 );
nand ( n17284 , n17283 , n9952 );
not ( n17285 , n17284 );
or ( n17286 , n17278 , n17285 );
not ( n17287 , n2931 );
not ( n17288 , n15373 );
or ( n17289 , n17287 , n17288 );
nand ( n17290 , n17289 , n2940 );
and ( n17291 , n15917 , n17290 , n15948 );
nand ( n17292 , n17286 , n17291 );
not ( n17293 , n15929 );
not ( n17294 , n15395 );
not ( n17295 , n9895 );
or ( n17296 , n17294 , n17295 );
nand ( n17297 , n17296 , n120 );
not ( n17298 , n17297 );
or ( n17299 , n17293 , n17298 );
nand ( n17300 , n17299 , n2785 );
not ( n17301 , n2942 );
not ( n17302 , n9875 );
or ( n17303 , n17301 , n17302 );
nand ( n17304 , n17303 , n14768 );
not ( n17305 , n2988 );
nand ( n17306 , n17305 , n2876 );
nand ( n17307 , n17304 , n17306 , n9973 );
not ( n17308 , n126 );
not ( n17309 , n2979 );
or ( n17310 , n17308 , n17309 );
not ( n17311 , n9947 );
nor ( n17312 , n9862 , n9912 );
or ( n17313 , n17311 , n17312 );
nand ( n17314 , n17313 , n9928 );
nand ( n17315 , n17310 , n17314 );
nor ( n17316 , n17307 , n17315 );
or ( n17317 , n2949 , n2986 );
nand ( n17318 , n17300 , n17316 , n17317 );
nand ( n17319 , n17292 , n17318 );
nand ( n17320 , n17270 , n17319 );
not ( n17321 , n17320 );
not ( n17322 , n17321 );
xnor ( n17323 , n17243 , n17322 );
not ( n17324 , n353 );
not ( n17325 , n2392 );
not ( n17326 , n15565 );
not ( n17327 , n2256 );
or ( n17328 , n17326 , n17327 );
nand ( n17329 , n17328 , n10239 );
not ( n17330 , n17329 );
not ( n17331 , n2424 );
or ( n17332 , n17330 , n17331 );
not ( n17333 , n2303 );
not ( n17334 , n14656 );
or ( n17335 , n17333 , n17334 );
nand ( n17336 , n17335 , n133 );
nand ( n17337 , n17332 , n17336 );
or ( n17338 , n17325 , n17337 );
nand ( n17339 , n14670 , n2316 );
nor ( n17340 , n16297 , n2460 );
or ( n17341 , n17339 , n17340 );
nand ( n17342 , n17338 , n17341 );
and ( n17343 , n16337 , n10186 , n2359 );
nand ( n17344 , n2298 , n2377 );
nand ( n17345 , n17342 , n17343 , n17344 );
not ( n17346 , n17345 );
nor ( n17347 , n15681 , n134 );
and ( n17348 , n15602 , n17347 , n15540 );
not ( n17349 , n2288 );
not ( n17350 , n10295 );
or ( n17351 , n17349 , n17350 );
nand ( n17352 , n10175 , n10302 );
nand ( n17353 , n17351 , n17352 );
not ( n17354 , n17353 );
nand ( n17355 , n2287 , n2285 );
and ( n17356 , n10195 , n17354 , n17355 );
nand ( n17357 , n17348 , n17356 );
or ( n17358 , n17357 , n16294 );
or ( n17359 , n2294 , n16301 );
nand ( n17360 , n17359 , n134 );
and ( n17361 , n17360 , n2506 );
and ( n17362 , n10302 , n10250 );
nor ( n17363 , n17361 , n17362 );
nand ( n17364 , n17363 , n15644 );
nand ( n17365 , n17358 , n17364 );
not ( n17366 , n2359 );
nand ( n17367 , n17366 , n15638 , n2503 , n15687 );
and ( n17368 , n10291 , n2370 , n2380 );
nor ( n17369 , n17368 , n2376 );
nor ( n17370 , n17367 , n17369 );
nand ( n17371 , n17365 , n17370 );
not ( n17372 , n17371 );
or ( n17373 , n17346 , n17372 );
not ( n17374 , n15729 );
not ( n17375 , n132 );
or ( n17376 , n17374 , n17375 );
nand ( n17377 , n17376 , n133 );
nor ( n17378 , n17377 , n16315 );
not ( n17379 , n131 );
not ( n17380 , n10278 );
not ( n17381 , n17380 );
or ( n17382 , n17379 , n17381 );
nand ( n17383 , n17382 , n2424 );
nor ( n17384 , n15737 , n17383 );
or ( n17385 , n17378 , n17384 );
nand ( n17386 , n17385 , n16246 );
and ( n17387 , n10195 , n15648 , n10299 , n16310 );
not ( n17388 , n2449 );
nand ( n17389 , n17388 , n14670 , n2275 );
nor ( n17390 , n15683 , n17389 );
or ( n17391 , n17387 , n17390 );
and ( n17392 , n14720 , n2472 );
nand ( n17393 , n17391 , n17392 );
and ( n17394 , n17386 , n17393 );
not ( n17395 , n14695 );
not ( n17396 , n2503 );
or ( n17397 , n17395 , n17396 );
nand ( n17398 , n17397 , n133 );
nand ( n17399 , n17398 , n14722 );
nor ( n17400 , n17394 , n17399 );
nand ( n17401 , n17373 , n17400 );
not ( n17402 , n17401 );
not ( n17403 , n16153 );
not ( n17404 , n17403 );
not ( n17405 , n2520 );
not ( n17406 , n17405 );
not ( n17407 , n17139 );
or ( n17408 , n17406 , n17407 );
nand ( n17409 , n17408 , n2686 );
not ( n17410 , n17409 );
or ( n17411 , n17404 , n17410 );
nand ( n17412 , n2683 , n14924 , n3341 );
nor ( n17413 , n3299 , n17412 );
nand ( n17414 , n14901 , n2571 );
and ( n17415 , n14998 , n2591 , n17414 , n2609 );
or ( n17416 , n17413 , n17415 );
not ( n17417 , n14902 );
nor ( n17418 , n17417 , n2613 );
nand ( n17419 , n17416 , n17418 );
nand ( n17420 , n17411 , n17419 );
and ( n17421 , n15021 , n139 );
nor ( n17422 , n17421 , n15008 );
not ( n17423 , n17422 );
not ( n17424 , n3404 );
or ( n17425 , n17423 , n17424 );
nand ( n17426 , n17425 , n16193 );
not ( n17427 , n2631 );
not ( n17428 , n17427 );
not ( n17429 , n14982 );
or ( n17430 , n17428 , n17429 );
and ( n17431 , n2758 , n141 );
nand ( n17432 , n17430 , n17431 );
nand ( n17433 , n2573 , n14901 );
and ( n17434 , n17432 , n17433 );
and ( n17435 , n17426 , n17434 );
nand ( n17436 , n17420 , n17435 );
not ( n17437 , n17436 );
not ( n17438 , n14964 );
not ( n17439 , n3381 );
not ( n17440 , n3322 );
or ( n17441 , n17439 , n17440 );
nand ( n17442 , n17441 , n14975 );
nor ( n17443 , n17438 , n17442 );
nand ( n17444 , n14911 , n3298 , n17443 , n15810 );
and ( n17445 , n3404 , n3352 );
nor ( n17446 , n17445 , n141 );
or ( n17447 , n17444 , n17446 );
not ( n17448 , n139 );
not ( n17449 , n2761 );
or ( n17450 , n17448 , n17449 );
nand ( n17451 , n17450 , n2731 );
not ( n17452 , n17451 );
nand ( n17453 , n17452 , n144 );
or ( n17454 , n15883 , n17453 );
nand ( n17455 , n17454 , n2654 );
nand ( n17456 , n3335 , n2752 );
nand ( n17457 , n17455 , n17456 );
nand ( n17458 , n17447 , n17457 );
not ( n17459 , n17458 );
nand ( n17460 , n3345 , n2576 );
not ( n17461 , n2632 );
or ( n17462 , n17460 , n17461 );
nand ( n17463 , n17462 , n2639 );
nand ( n17464 , n14902 , n14924 , n14911 );
nand ( n17465 , n17464 , n2517 );
and ( n17466 , n17463 , n17465 , n137 );
not ( n17467 , n17466 );
or ( n17468 , n17459 , n17467 );
and ( n17469 , n3405 , n2639 );
nand ( n17470 , n3302 , n2642 );
nor ( n17471 , n17469 , n17470 );
not ( n17472 , n15848 );
not ( n17473 , n3410 );
and ( n17474 , n17472 , n17473 );
nor ( n17475 , n17474 , n17451 );
or ( n17476 , n17475 , n3284 );
nand ( n17477 , n15795 , n16193 );
not ( n17478 , n14938 );
or ( n17479 , n17477 , n17478 );
nand ( n17480 , n17476 , n17479 );
not ( n17481 , n17480 );
not ( n17482 , n17144 );
or ( n17483 , n17481 , n17482 );
not ( n17484 , n2562 );
not ( n17485 , n2762 );
or ( n17486 , n17484 , n17485 );
nand ( n17487 , n17486 , n2592 );
nand ( n17488 , n17483 , n17487 );
nand ( n17489 , n17471 , n17488 , n3358 );
nand ( n17490 , n17468 , n17489 );
nand ( n17491 , n17437 , n17490 );
not ( n17492 , n17491 );
not ( n17493 , n17492 );
or ( n17494 , n17402 , n17493 );
not ( n17495 , n17401 );
nand ( n17496 , n17495 , n17491 );
nand ( n17497 , n17494 , n17496 );
xnor ( n17498 , n17324 , n17497 );
not ( n17499 , n17498 );
and ( n17500 , n17323 , n17499 );
not ( n17501 , n17323 );
and ( n17502 , n17501 , n17498 );
nor ( n17503 , n17500 , n17502 );
or ( n17504 , n17503 , n1 );
and ( n17505 , n354 , n17324 );
not ( n17506 , n354 );
and ( n17507 , n17506 , n353 );
nor ( n17508 , n17505 , n17507 );
or ( n17509 , n2246 , n17508 );
nand ( n17510 , n17504 , n17509 );
not ( n17511 , n17014 );
not ( n17512 , n357 );
and ( n17513 , n17511 , n17512 );
and ( n17514 , n17110 , n357 );
nor ( n17515 , n17513 , n17514 );
not ( n17516 , n17515 );
not ( n17517 , n10660 );
and ( n17518 , n10490 , n10453 , n1412 );
nor ( n17519 , n17518 , n177 );
not ( n17520 , n17519 );
nand ( n17521 , n1378 , n173 );
or ( n17522 , n17521 , n174 );
nand ( n17523 , n17522 , n11971 );
nand ( n17524 , n1348 , n1298 );
nand ( n17525 , n17524 , n1280 );
not ( n17526 , n1428 );
or ( n17527 , n17523 , n17525 , n17526 );
nor ( n17528 , n11989 , n13005 );
nand ( n17529 , n1486 , n17528 );
nand ( n17530 , n17527 , n17529 );
not ( n17531 , n17530 );
or ( n17532 , n17520 , n17531 );
or ( n17533 , n10356 , n10463 , n1370 );
nand ( n17534 , n17533 , n1434 );
nand ( n17535 , n17534 , n10407 );
nand ( n17536 , n17532 , n17535 );
not ( n17537 , n1418 );
not ( n17538 , n1363 );
or ( n17539 , n17537 , n17538 );
not ( n17540 , n11882 );
nand ( n17541 , n10402 , n174 );
and ( n17542 , n17541 , n13075 , n177 );
not ( n17543 , n17542 );
or ( n17544 , n17540 , n17543 );
nand ( n17545 , n17544 , n1434 );
nand ( n17546 , n17539 , n17545 );
not ( n17547 , n17546 );
and ( n17548 , n17524 , n1419 , n1387 , n13384 );
nor ( n17549 , n10457 , n10389 );
not ( n17550 , n17549 );
not ( n17551 , n1337 );
or ( n17552 , n17550 , n17551 );
nand ( n17553 , n17552 , n12992 );
nand ( n17554 , n1357 , n11871 );
and ( n17555 , n17548 , n17553 , n17554 );
nor ( n17556 , n17547 , n17555 );
nand ( n17557 , n16955 , n10361 );
not ( n17558 , n1485 );
and ( n17559 , n10458 , n17554 , n17558 );
nor ( n17560 , n17559 , n1315 );
or ( n17561 , n17557 , n17560 );
not ( n17562 , n17554 );
not ( n17563 , n10458 );
or ( n17564 , n17562 , n17563 );
nand ( n17565 , n17564 , n175 );
nand ( n17566 , n17565 , n1458 );
nand ( n17567 , n17561 , n17566 );
not ( n17568 , n1513 );
nor ( n17569 , n17568 , n1350 );
nand ( n17570 , n17567 , n17569 );
or ( n17571 , n17556 , n17570 );
nor ( n17572 , n11972 , n178 );
not ( n17573 , n1526 );
nand ( n17574 , n17573 , n1391 );
and ( n17575 , n17572 , n11924 , n17574 );
and ( n17576 , n1363 , n1298 );
nor ( n17577 , n17576 , n1528 , n1434 );
nand ( n17578 , n10370 , n1446 );
nor ( n17579 , n17578 , n1490 );
nor ( n17580 , n17577 , n17579 );
or ( n17581 , n17580 , n13457 );
not ( n17582 , n11861 );
not ( n17583 , n1473 );
or ( n17584 , n17582 , n17583 );
nand ( n17585 , n17584 , n13451 );
nand ( n17586 , n17581 , n17585 );
nand ( n17587 , n17575 , n17586 );
nand ( n17588 , n17571 , n17587 );
not ( n17589 , n1403 );
not ( n17590 , n1524 );
or ( n17591 , n17589 , n17590 );
not ( n17592 , n1344 );
not ( n17593 , n10506 );
or ( n17594 , n17592 , n17593 );
nand ( n17595 , n17594 , n171 );
nand ( n17596 , n17591 , n17595 );
nand ( n17597 , n17596 , n1435 );
not ( n17598 , n1349 );
or ( n17599 , n17598 , n13043 );
nand ( n17600 , n17599 , n176 );
and ( n17601 , n17597 , n17600 , n13072 );
nand ( n17602 , n17536 , n17588 , n17601 );
not ( n17603 , n17602 );
nor ( n17604 , n12986 , n17603 );
not ( n17605 , n17604 );
not ( n17606 , n17602 );
nand ( n17607 , n17606 , n12986 );
nand ( n17608 , n17605 , n17607 );
not ( n17609 , n17608 );
not ( n17610 , n17609 );
or ( n17611 , n17517 , n17610 );
not ( n17612 , n11687 );
or ( n17613 , n17612 , n17609 );
nand ( n17614 , n17611 , n17613 );
not ( n17615 , n17614 );
or ( n17616 , n17516 , n17615 );
or ( n17617 , n17614 , n17515 );
nand ( n17618 , n17616 , n17617 );
or ( n17619 , n17618 , n1 );
xnor ( n17620 , n357 , n358 );
or ( n17621 , n2246 , n17620 );
nand ( n17622 , n17619 , n17621 );
not ( n17623 , n13487 );
not ( n17624 , n16963 );
and ( n17625 , n17623 , n17624 );
not ( n17626 , n16962 );
and ( n17627 , n13487 , n17626 );
nor ( n17628 , n17625 , n17627 );
and ( n17629 , n17628 , n10770 );
not ( n17630 , n17628 );
and ( n17631 , n17630 , n10769 );
or ( n17632 , n17629 , n17631 );
and ( n17633 , n346 , n11827 );
not ( n17634 , n346 );
and ( n17635 , n17634 , n11832 );
nor ( n17636 , n17633 , n17635 );
not ( n17637 , n11048 );
not ( n17638 , n10528 );
and ( n17639 , n17637 , n17638 );
and ( n17640 , n10528 , n11048 );
nor ( n17641 , n17639 , n17640 );
and ( n17642 , n17636 , n17641 );
not ( n17643 , n17636 );
not ( n17644 , n17641 );
and ( n17645 , n17643 , n17644 );
nor ( n17646 , n17642 , n17645 );
and ( n17647 , n17632 , n17646 );
not ( n17648 , n17632 );
not ( n17649 , n17646 );
and ( n17650 , n17648 , n17649 );
nor ( n17651 , n17647 , n17650 );
or ( n17652 , n17651 , n1 );
xnor ( n17653 , n346 , n347 );
or ( n17654 , n2246 , n17653 );
nand ( n17655 , n17652 , n17654 );
not ( n17656 , n16643 );
not ( n17657 , n3985 );
nor ( n17658 , n4096 , n17657 );
not ( n17659 , n17658 );
nand ( n17660 , n4096 , n4016 , n198 );
nand ( n17661 , n17659 , n17660 );
and ( n17662 , n17661 , n4160 );
not ( n17663 , n5156 );
not ( n17664 , n5757 );
or ( n17665 , n17663 , n17664 );
nand ( n17666 , n17665 , n4179 );
and ( n17667 , n17666 , n5703 );
nor ( n17668 , n17662 , n17667 );
not ( n17669 , n5768 );
not ( n17670 , n3980 );
or ( n17671 , n17669 , n17670 );
nand ( n17672 , n17671 , n202 );
nand ( n17673 , n14544 , n17668 , n17672 );
not ( n17674 , n3973 );
nor ( n17675 , n17674 , n4150 );
not ( n17676 , n17675 );
not ( n17677 , n4129 );
or ( n17678 , n17676 , n17677 );
nand ( n17679 , n17678 , n4142 );
nand ( n17680 , n17679 , n203 );
and ( n17681 , n17673 , n17680 );
not ( n17682 , n5185 );
not ( n17683 , n5173 );
not ( n17684 , n17683 );
or ( n17685 , n17682 , n17684 );
nand ( n17686 , n4103 , n5671 , n203 );
nand ( n17687 , n17685 , n17686 );
not ( n17688 , n17687 );
not ( n17689 , n4026 );
not ( n17690 , n5137 );
or ( n17691 , n17689 , n17690 );
nand ( n17692 , n17691 , n202 );
nand ( n17693 , n14540 , n4078 );
nand ( n17694 , n17688 , n17692 , n17693 );
nor ( n17695 , n17681 , n17694 );
nand ( n17696 , n4195 , n5826 , n4067 );
not ( n17697 , n4051 );
not ( n17698 , n4158 );
or ( n17699 , n17697 , n17698 );
nand ( n17700 , n17699 , n5213 );
nor ( n17701 , n17696 , n17700 );
not ( n17702 , n17701 );
not ( n17703 , n5224 );
not ( n17704 , n5092 );
or ( n17705 , n17703 , n17704 );
nand ( n17706 , n5815 , n4055 , n5185 );
nand ( n17707 , n17705 , n17706 );
not ( n17708 , n17707 );
or ( n17709 , n17702 , n17708 );
not ( n17710 , n197 );
not ( n17711 , n3971 );
not ( n17712 , n17711 );
or ( n17713 , n17710 , n17712 );
nand ( n17714 , n17713 , n5704 );
or ( n17715 , n17714 , n4067 );
nand ( n17716 , n17715 , n4077 );
nor ( n17717 , n5862 , n14608 );
nand ( n17718 , n17716 , n17717 );
nand ( n17719 , n17709 , n17718 );
not ( n17720 , n17719 );
or ( n17721 , n5675 , n5693 );
nand ( n17722 , n17721 , n5671 );
not ( n17723 , n4137 );
nand ( n17724 , n17723 , n5842 );
not ( n17725 , n5137 );
nor ( n17726 , n17725 , n5146 );
and ( n17727 , n17722 , n17724 , n17726 );
not ( n17728 , n17727 );
or ( n17729 , n17720 , n17728 );
not ( n17730 , n4136 );
not ( n17731 , n4078 );
buf ( n17732 , n5706 );
nor ( n17733 , n5199 , n17732 );
not ( n17734 , n17733 );
or ( n17735 , n17731 , n17734 );
nor ( n17736 , n4095 , n4097 );
or ( n17737 , n17714 , n17736 );
nand ( n17738 , n17737 , n4121 );
nand ( n17739 , n17735 , n17738 );
not ( n17740 , n17739 );
or ( n17741 , n17730 , n17740 );
not ( n17742 , n4166 );
not ( n17743 , n4107 );
or ( n17744 , n17742 , n17743 );
not ( n17745 , n5769 );
nand ( n17746 , n17744 , n17745 );
nand ( n17747 , n17741 , n17746 );
not ( n17748 , n14555 );
not ( n17749 , n5671 );
not ( n17750 , n5140 );
or ( n17751 , n17749 , n17750 );
nand ( n17752 , n17751 , n5217 );
nor ( n17753 , n17748 , n17752 , n204 );
nand ( n17754 , n17747 , n17753 );
nand ( n17755 , n17729 , n17754 );
nand ( n17756 , n17695 , n17755 );
not ( n17757 , n17756 );
xnor ( n17758 , n9599 , n17757 );
not ( n17759 , n17758 );
or ( n17760 , n17656 , n17759 );
or ( n17761 , n17758 , n16643 );
nand ( n17762 , n17760 , n17761 );
not ( n17763 , n16720 );
not ( n17764 , n5087 );
or ( n17765 , n17763 , n17764 );
nand ( n17766 , n5248 , n16719 );
nand ( n17767 , n17765 , n17766 );
not ( n17768 , n380 );
not ( n17769 , n17768 );
not ( n17770 , n6156 );
or ( n17771 , n17769 , n17770 );
or ( n17772 , n6272 , n17768 );
nand ( n17773 , n17771 , n17772 );
xor ( n17774 , n17767 , n17773 );
and ( n17775 , n17762 , n17774 );
not ( n17776 , n17762 );
not ( n17777 , n17774 );
and ( n17778 , n17776 , n17777 );
nor ( n17779 , n17775 , n17778 );
or ( n17780 , n17779 , n1 );
and ( n17781 , n381 , n17768 );
not ( n17782 , n381 );
and ( n17783 , n17782 , n380 );
nor ( n17784 , n17781 , n17783 );
or ( n17785 , n2246 , n17784 );
nand ( n17786 , n17780 , n17785 );
not ( n17787 , n382 );
xnor ( n17788 , n17787 , n2059 );
xor ( n17789 , n17788 , n13612 );
not ( n17790 , n13454 );
not ( n17791 , n13437 );
or ( n17792 , n17790 , n17791 );
nand ( n17793 , n17792 , n13485 );
not ( n17794 , n17793 );
not ( n17795 , n10765 );
not ( n17796 , n17795 );
or ( n17797 , n17794 , n17796 );
not ( n17798 , n17793 );
nand ( n17799 , n17798 , n10765 );
nand ( n17800 , n17797 , n17799 );
not ( n17801 , n17603 );
not ( n17802 , n17105 );
not ( n17803 , n17802 );
or ( n17804 , n17801 , n17803 );
nand ( n17805 , n17105 , n17602 );
nand ( n17806 , n17804 , n17805 );
xor ( n17807 , n17800 , n17806 );
xnor ( n17808 , n17789 , n17807 );
or ( n17809 , n17808 , n1 );
and ( n17810 , n383 , n17787 );
not ( n17811 , n383 );
and ( n17812 , n17811 , n382 );
nor ( n17813 , n17810 , n17812 );
or ( n17814 , n2246 , n17813 );
nand ( n17815 , n17809 , n17814 );
nand ( n17816 , n10039 , n3154 , n16092 );
nor ( n17817 , n15995 , n17816 );
nand ( n17818 , n15257 , n3257 );
and ( n17819 , n17818 , n10037 );
or ( n17820 , n17817 , n17819 );
nand ( n17821 , n10091 , n3063 );
and ( n17822 , n15190 , n15160 , n17821 );
nand ( n17823 , n17820 , n17822 );
nand ( n17824 , n3154 , n3060 );
not ( n17825 , n17824 );
not ( n17826 , n15166 );
nand ( n17827 , n17825 , n17826 , n15177 , n118 );
not ( n17828 , n17827 );
nand ( n17829 , n15177 , n10025 );
not ( n17830 , n17829 );
or ( n17831 , n17828 , n17830 );
or ( n17832 , n3118 , n10052 );
nand ( n17833 , n17832 , n3063 );
nand ( n17834 , n17831 , n17833 );
nand ( n17835 , n17823 , n17834 , n119 );
and ( n17836 , n112 , n3114 );
nor ( n17837 , n17836 , n10100 );
not ( n17838 , n17837 );
not ( n17839 , n15177 );
or ( n17840 , n17838 , n17839 );
nand ( n17841 , n17840 , n10037 );
not ( n17842 , n15472 );
not ( n17843 , n15426 );
or ( n17844 , n17842 , n17843 );
nand ( n17845 , n17844 , n119 );
or ( n17846 , n15228 , n10102 );
nand ( n17847 , n17846 , n3164 );
nand ( n17848 , n17841 , n17845 , n17847 );
not ( n17849 , n3130 );
nand ( n17850 , n3148 , n3247 );
nand ( n17851 , n10084 , n3135 , n17850 );
not ( n17852 , n17851 );
or ( n17853 , n17849 , n17852 );
nand ( n17854 , n16003 , n15144 );
or ( n17855 , n17854 , n3224 , n3175 );
nand ( n17856 , n17855 , n15223 );
nand ( n17857 , n17853 , n17856 );
nor ( n17858 , n17848 , n17857 );
not ( n17859 , n3230 );
nand ( n17860 , n3070 , n10145 );
not ( n17861 , n17860 );
not ( n17862 , n3183 );
or ( n17863 , n17861 , n17862 );
nor ( n17864 , n16084 , n3046 );
nand ( n17865 , n17863 , n17864 );
nand ( n17866 , n3184 , n117 );
nand ( n17867 , n17865 , n17866 );
not ( n17868 , n17867 );
or ( n17869 , n17859 , n17868 );
nand ( n17870 , n17869 , n118 );
not ( n17871 , n17870 );
not ( n17872 , n10063 );
nand ( n17873 , n3055 , n114 );
nand ( n17874 , n16026 , n17873 );
not ( n17875 , n17874 );
or ( n17876 , n17872 , n17875 );
nand ( n17877 , n17876 , n16081 );
or ( n17878 , n17871 , n17877 );
nand ( n17879 , n17878 , n3137 );
and ( n17880 , n17858 , n17879 );
not ( n17881 , n3251 );
not ( n17882 , n17824 );
or ( n17883 , n17881 , n17882 );
not ( n17884 , n15478 );
nand ( n17885 , n17884 , n3133 );
nand ( n17886 , n17883 , n17885 );
nand ( n17887 , n17886 , n3212 );
not ( n17888 , n16037 );
not ( n17889 , n9998 );
or ( n17890 , n17888 , n17889 );
nand ( n17891 , n17890 , n117 );
nand ( n17892 , n10110 , n10065 );
not ( n17893 , n17892 );
not ( n17894 , n15433 );
not ( n17895 , n17894 );
or ( n17896 , n17893 , n17895 );
nand ( n17897 , n17896 , n3266 );
nand ( n17898 , n17887 , n17891 , n17897 , n118 );
and ( n17899 , n3056 , n16040 );
nand ( n17900 , n10063 , n3194 );
and ( n17901 , n17899 , n15235 , n17900 );
nor ( n17902 , n17901 , n119 );
nand ( n17903 , n17898 , n17902 );
nand ( n17904 , n3134 , n3055 );
and ( n17905 , n17904 , n10035 );
not ( n17906 , n17905 );
not ( n17907 , n3195 );
or ( n17908 , n17854 , n17907 );
nand ( n17909 , n17908 , n3164 );
not ( n17910 , n17909 );
or ( n17911 , n17906 , n17910 );
nand ( n17912 , n17911 , n17898 );
nand ( n17913 , n17835 , n17880 , n17903 , n17912 );
and ( n17914 , n17913 , n3018 );
not ( n17915 , n17913 );
and ( n17916 , n17915 , n3019 );
nor ( n17917 , n17914 , n17916 );
not ( n17918 , n17917 );
not ( n17919 , n15903 );
not ( n17920 , n15518 );
or ( n17921 , n17919 , n17920 );
nand ( n17922 , n15517 , n15902 );
nand ( n17923 , n17921 , n17922 );
not ( n17924 , n17923 );
or ( n17925 , n17918 , n17924 );
not ( n17926 , n17923 );
not ( n17927 , n17917 );
nand ( n17928 , n17926 , n17927 );
nand ( n17929 , n17925 , n17928 );
not ( n17930 , n378 );
not ( n17931 , n15661 );
or ( n17932 , n17930 , n17931 );
or ( n17933 , n15661 , n378 );
nand ( n17934 , n17932 , n17933 );
not ( n17935 , n17934 );
and ( n17936 , n17929 , n17935 );
not ( n17937 , n17929 );
and ( n17938 , n17937 , n17934 );
nor ( n17939 , n17936 , n17938 );
or ( n17940 , n17939 , n1 );
xnor ( n17941 , n378 , n379 );
or ( n17942 , n2246 , n17941 );
nand ( n17943 , n17940 , n17942 );
not ( n17944 , n2059 );
not ( n17945 , n384 );
not ( n17946 , n17945 );
and ( n17947 , n17944 , n17946 );
and ( n17948 , n2059 , n17945 );
nor ( n17949 , n17947 , n17948 );
xor ( n17950 , n17949 , n13589 );
not ( n17951 , n17608 );
not ( n17952 , n999 );
not ( n17953 , n17793 );
and ( n17954 , n17952 , n17953 );
not ( n17955 , n13601 );
and ( n17956 , n17955 , n999 );
nor ( n17957 , n17954 , n17956 );
not ( n17958 , n17957 );
or ( n17959 , n17951 , n17958 );
or ( n17960 , n17608 , n17957 );
nand ( n17961 , n17959 , n17960 );
xnor ( n17962 , n17950 , n17961 );
or ( n17963 , n17962 , n1 );
and ( n17964 , n385 , n17945 );
not ( n17965 , n385 );
and ( n17966 , n17965 , n384 );
nor ( n17967 , n17964 , n17966 );
or ( n17968 , n2246 , n17967 );
nand ( n17969 , n17963 , n17968 );
not ( n17970 , n3164 );
not ( n17971 , n17818 );
not ( n17972 , n17971 );
or ( n17973 , n17970 , n17972 );
nand ( n17974 , n17973 , n10056 );
nor ( n17975 , n15452 , n17974 );
nand ( n17976 , n10001 , n17975 );
or ( n17977 , n15150 , n16084 );
not ( n17978 , n15214 );
or ( n17979 , n17978 , n10004 );
nand ( n17980 , n17977 , n17979 );
and ( n17981 , n10061 , n3250 , n15504 );
and ( n17982 , n17980 , n17981 , n15170 );
not ( n17983 , n16073 );
not ( n17984 , n15168 );
nand ( n17985 , n17983 , n17984 , n15436 , n3235 );
nand ( n17986 , n10075 , n10025 );
and ( n17987 , n17985 , n17986 );
nand ( n17988 , n3105 , n3149 , n17904 , n17821 );
nor ( n17989 , n17987 , n17988 );
nor ( n17990 , n17982 , n17989 );
or ( n17991 , n17976 , n17990 );
nor ( n17992 , n3169 , n3204 , n113 );
nor ( n17993 , n3224 , n17992 );
not ( n17994 , n17993 );
nand ( n17995 , n3144 , n10055 );
nand ( n17996 , n17995 , n17818 , n3106 );
nor ( n17997 , n17996 , n3268 );
not ( n17998 , n17997 );
or ( n17999 , n17994 , n17998 );
nand ( n18000 , n3095 , n10065 );
nand ( n18001 , n10121 , n18000 );
nor ( n18002 , n3128 , n3106 );
nand ( n18003 , n16036 , n18002 );
nor ( n18004 , n18001 , n18003 );
not ( n18005 , n3122 );
not ( n18006 , n3161 );
or ( n18007 , n18005 , n18006 );
nand ( n18008 , n18007 , n117 );
nand ( n18009 , n18004 , n18008 );
nand ( n18010 , n17999 , n18009 );
not ( n18011 , n15223 );
or ( n18012 , n18011 , n3120 );
not ( n18013 , n16080 );
not ( n18014 , n15231 );
nand ( n18015 , n18013 , n3240 , n18014 );
nand ( n18016 , n18012 , n18015 );
nand ( n18017 , n18010 , n18016 , n10015 );
nand ( n18018 , n17991 , n18017 );
not ( n18019 , n10015 );
not ( n18020 , n10077 );
or ( n18021 , n18019 , n18020 );
nand ( n18022 , n18021 , n10037 );
not ( n18023 , n18022 );
not ( n18024 , n10040 );
not ( n18025 , n15156 );
or ( n18026 , n18024 , n18025 );
nand ( n18027 , n18026 , n16079 );
nor ( n18028 , n15426 , n113 );
nor ( n18029 , n18023 , n18027 , n18028 , n3256 );
and ( n18030 , n3149 , n10023 );
or ( n18031 , n18030 , n15161 );
not ( n18032 , n10113 );
nand ( n18033 , n18032 , n3095 );
nand ( n18034 , n18031 , n18033 );
and ( n18035 , n3154 , n3027 , n15251 );
nor ( n18036 , n18035 , n3064 );
not ( n18037 , n15272 );
or ( n18038 , n18034 , n18036 , n18037 );
nand ( n18039 , n18038 , n118 );
and ( n18040 , n18029 , n18039 );
nand ( n18041 , n18018 , n18040 );
not ( n18042 , n18041 );
not ( n18043 , n18042 );
not ( n18044 , n14894 );
or ( n18045 , n18043 , n18044 );
nand ( n18046 , n18041 , n14893 );
nand ( n18047 , n18045 , n18046 );
not ( n18048 , n18047 );
not ( n18049 , n14764 );
or ( n18050 , n18048 , n18049 );
or ( n18051 , n14764 , n18047 );
nand ( n18052 , n18050 , n18051 );
not ( n18053 , n17491 );
nand ( n18054 , n2621 , n2766 );
not ( n18055 , n18054 );
or ( n18056 , n18053 , n18055 );
not ( n18057 , n18054 );
not ( n18058 , n18057 );
or ( n18059 , n18058 , n17491 );
nand ( n18060 , n18056 , n18059 );
xnor ( n18061 , n301 , n17401 );
not ( n18062 , n18061 );
and ( n18063 , n18060 , n18062 );
not ( n18064 , n18060 );
and ( n18065 , n18064 , n18061 );
nor ( n18066 , n18063 , n18065 );
not ( n18067 , n18066 );
and ( n18068 , n18052 , n18067 );
not ( n18069 , n18052 );
and ( n18070 , n18069 , n18066 );
nor ( n18071 , n18068 , n18070 );
or ( n18072 , n18071 , n1 );
xnor ( n18073 , n301 , n302 );
or ( n18074 , n2246 , n18073 );
nand ( n18075 , n18072 , n18074 );
or ( n18076 , n16481 , n16513 );
nand ( n18077 , n18076 , n16531 );
and ( n18078 , n12435 , n18077 );
not ( n18079 , n12435 );
and ( n18080 , n18079 , n16533 );
or ( n18081 , n18078 , n18080 );
not ( n18082 , n18081 );
not ( n18083 , n13823 );
or ( n18084 , n18082 , n18083 );
or ( n18085 , n13823 , n18081 );
nand ( n18086 , n18084 , n18085 );
not ( n18087 , n7668 );
not ( n18088 , n49 );
and ( n18089 , n18087 , n18088 );
and ( n18090 , n7668 , n49 );
nor ( n18091 , n18089 , n18090 );
not ( n18092 , n18091 );
and ( n18093 , n18086 , n18092 );
not ( n18094 , n18086 );
and ( n18095 , n18094 , n18091 );
nor ( n18096 , n18093 , n18095 );
or ( n18097 , n18096 , n1 );
xnor ( n18098 , n49 , n50 );
or ( n18099 , n2246 , n18098 );
nand ( n18100 , n18097 , n18099 );
not ( n18101 , n6553 );
not ( n18102 , n18101 );
not ( n18103 , n9017 );
or ( n18104 , n18102 , n18103 );
nand ( n18105 , n6553 , n9016 );
nand ( n18106 , n18104 , n18105 );
not ( n18107 , n18106 );
not ( n18108 , n8272 );
not ( n18109 , n55 );
and ( n18110 , n18108 , n18109 );
and ( n18111 , n14300 , n55 );
nor ( n18112 , n18110 , n18111 );
not ( n18113 , n18112 );
or ( n18114 , n18107 , n18113 );
or ( n18115 , n18112 , n18106 );
nand ( n18116 , n18114 , n18115 );
and ( n18117 , n18116 , n9224 );
not ( n18118 , n18116 );
and ( n18119 , n18118 , n9223 );
nor ( n18120 , n18117 , n18119 );
or ( n18121 , n18120 , n1 );
xnor ( n18122 , n55 , n56 );
or ( n18123 , n2246 , n18122 );
nand ( n18124 , n18121 , n18123 );
not ( n18125 , n14298 );
not ( n18126 , n14271 );
or ( n18127 , n18125 , n18126 );
or ( n18128 , n14298 , n14271 );
nand ( n18129 , n18127 , n18128 );
xnor ( n18130 , n81 , n7664 );
xnor ( n18131 , n14278 , n18130 );
and ( n18132 , n18129 , n18131 );
not ( n18133 , n18129 );
not ( n18134 , n18131 );
and ( n18135 , n18133 , n18134 );
nor ( n18136 , n18132 , n18135 );
or ( n18137 , n18136 , n1 );
xnor ( n18138 , n81 , n82 );
or ( n18139 , n2246 , n18138 );
nand ( n18140 , n18137 , n18139 );
not ( n18141 , n90 );
and ( n18142 , n9351 , n18141 );
not ( n18143 , n9351 );
and ( n18144 , n18143 , n90 );
nor ( n18145 , n18142 , n18144 );
not ( n18146 , n8505 );
and ( n18147 , n18146 , n14306 );
not ( n18148 , n18146 );
and ( n18149 , n18148 , n8268 );
nor ( n18150 , n18147 , n18149 );
xor ( n18151 , n18145 , n18150 );
xnor ( n18152 , n18151 , n9478 );
or ( n18153 , n18152 , n1 );
and ( n18154 , n91 , n18141 );
not ( n18155 , n91 );
and ( n18156 , n18155 , n90 );
nor ( n18157 , n18154 , n18156 );
or ( n18158 , n2246 , n18157 );
nand ( n18159 , n18153 , n18158 );
and ( n18160 , n136 , n2512 );
not ( n18161 , n136 );
and ( n18162 , n18161 , n2513 );
or ( n18163 , n18160 , n18162 );
not ( n18164 , n15330 );
nand ( n18165 , n15333 , n2785 );
not ( n18166 , n2855 );
not ( n18167 , n2844 );
or ( n18168 , n18166 , n18167 );
nand ( n18169 , n18168 , n2857 );
and ( n18170 , n2802 , n9928 , n9840 );
nor ( n18171 , n18170 , n2973 );
and ( n18172 , n18169 , n18171 );
and ( n18173 , n18165 , n18172 );
and ( n18174 , n9836 , n14845 , n2973 );
nor ( n18175 , n18173 , n18174 );
not ( n18176 , n14800 );
and ( n18177 , n9965 , n18176 , n126 );
nor ( n18178 , n18177 , n2857 );
not ( n18179 , n18178 );
nand ( n18180 , n9964 , n15047 );
not ( n18181 , n18180 );
and ( n18182 , n18179 , n18181 );
and ( n18183 , n2817 , n9962 , n2785 );
nand ( n18184 , n2911 , n2816 );
nand ( n18185 , n9965 , n18183 , n18184 , n18176 );
nand ( n18186 , n18185 , n9929 );
nor ( n18187 , n18182 , n18186 );
nor ( n18188 , n18164 , n18175 , n18187 );
not ( n18189 , n18188 );
not ( n18190 , n2942 );
and ( n18191 , n18189 , n18190 );
not ( n18192 , n2990 );
not ( n18193 , n2918 );
or ( n18194 , n18192 , n18193 );
nand ( n18195 , n18194 , n121 );
nand ( n18196 , n9925 , n18195 , n17244 );
or ( n18197 , n18196 , n2913 );
nand ( n18198 , n18197 , n126 );
not ( n18199 , n9907 );
not ( n18200 , n9948 );
or ( n18201 , n18199 , n18200 );
nand ( n18202 , n18201 , n3000 );
nor ( n18203 , n15045 , n122 );
or ( n18204 , n18202 , n18203 );
nand ( n18205 , n18204 , n2785 );
nand ( n18206 , n14886 , n14871 , n2922 );
and ( n18207 , n18206 , n2857 );
nor ( n18208 , n18207 , n15406 );
and ( n18209 , n18198 , n18205 , n18208 );
or ( n18210 , n18209 , n127 );
not ( n18211 , n9929 );
not ( n18212 , n15071 );
nand ( n18213 , n18212 , n3002 , n9962 , n2785 );
not ( n18214 , n18213 );
or ( n18215 , n18211 , n18214 );
nand ( n18216 , n18215 , n17317 );
or ( n18217 , n15951 , n2894 );
or ( n18218 , n9905 , n2972 );
nand ( n18219 , n18217 , n18218 );
not ( n18220 , n2941 );
nor ( n18221 , n18220 , n9833 );
nand ( n18222 , n18219 , n18221 , n9849 );
and ( n18223 , n18216 , n18222 );
not ( n18224 , n9981 );
not ( n18225 , n17297 );
or ( n18226 , n18224 , n18225 );
nand ( n18227 , n18226 , n2924 );
nand ( n18228 , n18227 , n14789 );
nor ( n18229 , n18223 , n18228 );
nand ( n18230 , n18210 , n18229 );
nor ( n18231 , n18191 , n18230 );
not ( n18232 , n18231 );
not ( n18233 , n18232 );
not ( n18234 , n3272 );
or ( n18235 , n18233 , n18234 );
nand ( n18236 , n3271 , n18231 );
nand ( n18237 , n18235 , n18236 );
xor ( n18238 , n18163 , n18237 );
buf ( n18239 , n2767 );
not ( n18240 , n17913 );
not ( n18241 , n18240 );
not ( n18242 , n18241 );
and ( n18243 , n18239 , n18242 );
not ( n18244 , n18239 );
and ( n18245 , n18244 , n18241 );
nor ( n18246 , n18243 , n18245 );
not ( n18247 , n18246 );
and ( n18248 , n18238 , n18247 );
not ( n18249 , n18238 );
and ( n18250 , n18249 , n18246 );
nor ( n18251 , n18248 , n18250 );
or ( n18252 , n18251 , n1 );
xnor ( n18253 , n136 , n145 );
or ( n18254 , n2246 , n18253 );
nand ( n18255 , n18252 , n18254 );
buf ( n18256 , n1150 );
not ( n18257 , n18256 );
nor ( n18258 , n13457 , n176 );
nand ( n18259 , n16955 , n18258 );
or ( n18260 , n18259 , n11950 );
not ( n18261 , n1364 );
or ( n18262 , n1534 , n18261 );
nand ( n18263 , n18260 , n18262 );
and ( n18264 , n17522 , n12988 );
nand ( n18265 , n18263 , n18264 );
and ( n18266 , n18265 , n1370 );
not ( n18267 , n10389 );
not ( n18268 , n1280 );
not ( n18269 , n1421 );
not ( n18270 , n18269 );
or ( n18271 , n18268 , n18270 );
not ( n18272 , n10424 );
not ( n18273 , n11911 );
or ( n18274 , n18272 , n18273 );
nand ( n18275 , n18274 , n176 );
nand ( n18276 , n18271 , n18275 );
not ( n18277 , n18276 );
or ( n18278 , n18267 , n18277 );
not ( n18279 , n11899 );
not ( n18280 , n13075 );
or ( n18281 , n18279 , n18280 );
nand ( n18282 , n18281 , n11858 );
not ( n18283 , n18282 );
not ( n18284 , n10458 );
or ( n18285 , n18283 , n18284 );
nand ( n18286 , n18285 , n1435 );
and ( n18287 , n18286 , n13035 , n1521 );
nand ( n18288 , n18278 , n18287 );
nor ( n18289 , n18266 , n18288 );
not ( n18290 , n1313 );
not ( n18291 , n11968 );
or ( n18292 , n18290 , n18291 );
not ( n18293 , n16930 );
nand ( n18294 , n18292 , n18293 );
and ( n18295 , n18294 , n177 );
and ( n18296 , n13074 , n10416 , n1296 );
nor ( n18297 , n18296 , n1434 );
nor ( n18298 , n18295 , n18297 );
nand ( n18299 , n11978 , n17521 , n176 );
not ( n18300 , n18299 );
not ( n18301 , n17525 );
or ( n18302 , n18300 , n18301 );
nor ( n18303 , n11950 , n11943 );
nand ( n18304 , n18302 , n18303 );
nand ( n18305 , n18304 , n1370 );
nand ( n18306 , n18298 , n18305 );
nand ( n18307 , n13050 , n1536 , n13407 , n10491 );
not ( n18308 , n10404 );
nand ( n18309 , n18308 , n10495 , n13411 );
and ( n18310 , n18307 , n18309 );
or ( n18311 , n18306 , n18310 );
not ( n18312 , n10508 );
nor ( n18313 , n18312 , n1460 );
not ( n18314 , n1524 );
nand ( n18315 , n18314 , n10439 );
and ( n18316 , n18315 , n10374 );
not ( n18317 , n10495 );
nor ( n18318 , n18316 , n18317 );
not ( n18319 , n1370 );
not ( n18320 , n17521 );
or ( n18321 , n18319 , n18320 );
nand ( n18322 , n18321 , n1375 );
nand ( n18323 , n18313 , n18318 , n18322 );
and ( n18324 , n1434 , n10431 );
not ( n18325 , n18324 );
not ( n18326 , n16952 );
or ( n18327 , n18325 , n18326 );
not ( n18328 , n1489 );
not ( n18329 , n10444 );
or ( n18330 , n18328 , n18329 );
nand ( n18331 , n18330 , n1306 );
and ( n18332 , n18331 , n1428 );
nand ( n18333 , n18327 , n18332 );
nand ( n18334 , n18323 , n18333 );
not ( n18335 , n16874 );
not ( n18336 , n10508 );
or ( n18337 , n18335 , n18336 );
nand ( n18338 , n18337 , n176 );
and ( n18339 , n18338 , n1350 );
nand ( n18340 , n18334 , n18339 );
not ( n18341 , n11966 );
not ( n18342 , n10384 );
or ( n18343 , n1445 , n18342 );
or ( n18344 , n1409 , n1412 );
nand ( n18345 , n18343 , n18344 );
not ( n18346 , n18345 );
and ( n18347 , n18341 , n18346 );
nor ( n18348 , n18347 , n176 );
or ( n18349 , n18340 , n18348 );
nand ( n18350 , n18311 , n18349 );
nand ( n18351 , n18289 , n18350 );
not ( n18352 , n11522 );
not ( n18353 , n10947 );
or ( n18354 , n18352 , n18353 , n11529 );
not ( n18355 , n1579 );
nand ( n18356 , n18355 , n10952 , n11592 );
or ( n18357 , n13513 , n18356 );
nand ( n18358 , n18354 , n18357 );
not ( n18359 , n18358 );
nand ( n18360 , n10960 , n11038 );
or ( n18361 , n12078 , n18360 );
nand ( n18362 , n1636 , n1731 );
nand ( n18363 , n18361 , n18362 );
and ( n18364 , n12941 , n11554 );
nand ( n18365 , n18363 , n18364 );
not ( n18366 , n12077 );
not ( n18367 , n12090 );
nor ( n18368 , n18367 , n11601 );
not ( n18369 , n18368 );
or ( n18370 , n18366 , n18369 );
nand ( n18371 , n18370 , n12078 );
nand ( n18372 , n12948 , n12082 , n18371 );
or ( n18373 , n18365 , n18372 );
or ( n18374 , n1715 , n13538 , n10955 );
nand ( n18375 , n18374 , n149 );
nand ( n18376 , n1599 , n11490 , n1721 );
nand ( n18377 , n18375 , n10937 , n18376 , n152 );
nand ( n18378 , n18373 , n18377 );
not ( n18379 , n18378 );
or ( n18380 , n18359 , n18379 );
not ( n18381 , n1653 );
not ( n18382 , n10983 );
or ( n18383 , n18381 , n18382 );
nand ( n18384 , n18383 , n1631 );
not ( n18385 , n1750 );
not ( n18386 , n149 );
and ( n18387 , n18385 , n18386 );
nand ( n18388 , n10947 , n1752 );
nor ( n18389 , n18387 , n18388 );
nand ( n18390 , n10912 , n18384 , n18389 , n1753 );
or ( n18391 , n18365 , n18390 );
nand ( n18392 , n1614 , n1711 );
or ( n18393 , n11481 , n11662 );
and ( n18394 , n1603 , n10999 , n1784 );
nor ( n18395 , n18394 , n1752 );
nand ( n18396 , n1794 , n18392 , n18393 , n18395 );
nand ( n18397 , n18391 , n18396 );
not ( n18398 , n148 );
not ( n18399 , n1565 );
or ( n18400 , n18398 , n18399 );
nand ( n18401 , n18400 , n1737 );
not ( n18402 , n18401 );
not ( n18403 , n12109 );
or ( n18404 , n18402 , n18403 );
nand ( n18405 , n18404 , n1617 );
not ( n18406 , n18405 );
not ( n18407 , n149 );
not ( n18408 , n10912 );
not ( n18409 , n18408 );
or ( n18410 , n18407 , n18409 );
not ( n18411 , n1597 );
nand ( n18412 , n18411 , n1721 );
nand ( n18413 , n18410 , n18412 );
not ( n18414 , n10999 );
not ( n18415 , n10986 );
or ( n18416 , n18414 , n18415 );
nand ( n18417 , n18416 , n1735 );
nor ( n18418 , n18406 , n18413 , n18417 );
nand ( n18419 , n18397 , n18418 );
nand ( n18420 , n18380 , n18419 );
not ( n18421 , n13553 );
and ( n18422 , n13577 , n11624 );
not ( n18423 , n1618 );
nor ( n18424 , n18422 , n18423 );
not ( n18425 , n152 );
not ( n18426 , n12115 );
or ( n18427 , n18425 , n18426 );
not ( n18428 , n1603 );
not ( n18429 , n12965 );
or ( n18430 , n18428 , n18429 );
nand ( n18431 , n18430 , n13554 );
nand ( n18432 , n18431 , n1699 );
nand ( n18433 , n18427 , n18432 );
nor ( n18434 , n18421 , n18424 , n18433 );
nand ( n18435 , n18420 , n18434 );
and ( n18436 , n18351 , n18435 );
not ( n18437 , n18351 );
not ( n18438 , n18435 );
and ( n18439 , n18437 , n18438 );
or ( n18440 , n18436 , n18439 );
not ( n18441 , n18440 );
or ( n18442 , n18257 , n18441 );
or ( n18443 , n18256 , n18440 );
nand ( n18444 , n18442 , n18443 );
not ( n18445 , n162 );
xor ( n18446 , n2232 , n11577 );
not ( n18447 , n18446 );
or ( n18448 , n18445 , n18447 );
or ( n18449 , n162 , n18446 );
nand ( n18450 , n18448 , n18449 );
and ( n18451 , n18444 , n18450 );
not ( n18452 , n18444 );
not ( n18453 , n18450 );
and ( n18454 , n18452 , n18453 );
nor ( n18455 , n18451 , n18454 );
or ( n18456 , n18455 , n1 );
xnor ( n18457 , n162 , n179 );
or ( n18458 , n2246 , n18457 );
nand ( n18459 , n18456 , n18458 );
xor ( n18460 , n18232 , n16227 );
xor ( n18461 , n109 , n3430 );
xnor ( n18462 , n18461 , n10331 );
xnor ( n18463 , n18460 , n18462 );
or ( n18464 , n18463 , n1 );
xnor ( n18465 , n109 , n214 );
or ( n18466 , n2246 , n18465 );
nand ( n18467 , n18464 , n18466 );
nor ( n18468 , n12187 , n1899 );
and ( n18469 , n1902 , n159 );
nand ( n18470 , n18468 , n1936 , n18469 );
not ( n18471 , n18470 );
nand ( n18472 , n11718 , n2129 , n2078 );
not ( n18473 , n18472 );
or ( n18474 , n18471 , n18473 );
not ( n18475 , n2001 );
not ( n18476 , n12176 );
or ( n18477 , n18475 , n18476 );
nand ( n18478 , n18477 , n161 );
not ( n18479 , n18478 );
not ( n18480 , n12831 );
nand ( n18481 , n18480 , n2006 );
not ( n18482 , n2050 );
nand ( n18483 , n18482 , n2136 );
or ( n18484 , n11763 , n18483 );
nand ( n18485 , n18484 , n11722 );
and ( n18486 , n18479 , n18481 , n18485 );
nand ( n18487 , n18474 , n18486 );
not ( n18488 , n160 );
nor ( n18489 , n11746 , n10884 );
or ( n18490 , n10813 , n18489 );
not ( n18491 , n18490 );
or ( n18492 , n18488 , n18491 );
not ( n18493 , n12186 );
not ( n18494 , n18493 );
not ( n18495 , n1947 );
or ( n18496 , n18494 , n18495 );
nand ( n18497 , n18496 , n2004 );
nand ( n18498 , n18492 , n18497 );
or ( n18499 , n18487 , n18498 );
nand ( n18500 , n12832 , n154 );
not ( n18501 , n18500 );
not ( n18502 , n13269 );
or ( n18503 , n18501 , n18502 );
not ( n18504 , n2142 );
and ( n18505 , n18504 , n2067 );
nand ( n18506 , n12873 , n1905 );
nor ( n18507 , n18505 , n18506 );
nand ( n18508 , n18503 , n18507 );
not ( n18509 , n18508 );
not ( n18510 , n1906 );
nand ( n18511 , n18510 , n13331 , n10834 );
not ( n18512 , n18511 );
or ( n18513 , n18509 , n18512 );
nand ( n18514 , n13331 , n2210 , n11718 , n1868 );
and ( n18515 , n1988 , n2000 );
and ( n18516 , n12828 , n1841 );
nor ( n18517 , n18515 , n18516 );
nand ( n18518 , n18517 , n13275 );
or ( n18519 , n18514 , n18518 );
not ( n18520 , n1918 );
not ( n18521 , n10882 );
or ( n18522 , n18520 , n18521 );
nand ( n18523 , n1866 , n10876 );
nand ( n18524 , n18522 , n18523 );
nand ( n18525 , n18524 , n12136 , n160 );
nand ( n18526 , n18519 , n18525 );
nand ( n18527 , n18513 , n18526 );
nand ( n18528 , n18499 , n18527 );
nand ( n18529 , n1985 , n1921 );
nand ( n18530 , n1916 , n18529 , n10865 , n12872 );
nand ( n18531 , n18530 , n2004 );
nand ( n18532 , n2147 , n1864 , n160 );
nor ( n18533 , n1876 , n10867 );
or ( n18534 , n12839 , n18533 );
nand ( n18535 , n18534 , n2006 );
nand ( n18536 , n18531 , n1951 , n18532 , n18535 );
not ( n18537 , n1954 );
not ( n18538 , n10794 );
nand ( n18539 , n18538 , n156 );
nand ( n18540 , n18537 , n18539 );
or ( n18541 , n18540 , n10878 );
nand ( n18542 , n18541 , n11722 );
not ( n18543 , n2018 );
not ( n18544 , n12873 );
and ( n18545 , n18543 , n18544 );
not ( n18546 , n11782 );
nor ( n18547 , n18545 , n18546 );
nand ( n18548 , n18542 , n18547 );
nor ( n18549 , n18536 , n18548 );
nand ( n18550 , n18528 , n18549 );
and ( n18551 , n12122 , n18550 );
not ( n18552 , n12122 );
not ( n18553 , n18550 );
and ( n18554 , n18552 , n18553 );
nor ( n18555 , n18551 , n18554 );
not ( n18556 , n18351 );
not ( n18557 , n1200 );
not ( n18558 , n1114 );
or ( n18559 , n18557 , n18558 );
nand ( n18560 , n18559 , n167 );
and ( n18561 , n17019 , n778 );
nand ( n18562 , n869 , n805 );
and ( n18563 , n18560 , n18561 , n18562 );
not ( n18564 , n10546 );
not ( n18565 , n1007 );
or ( n18566 , n18564 , n18565 );
not ( n18567 , n167 );
nand ( n18568 , n18566 , n18567 );
nand ( n18569 , n18563 , n18568 );
not ( n18570 , n10622 );
not ( n18571 , n902 );
not ( n18572 , n948 );
or ( n18573 , n18571 , n18572 );
nand ( n18574 , n18573 , n957 );
nor ( n18575 , n18570 , n18574 );
not ( n18576 , n18575 );
not ( n18577 , n1246 );
or ( n18578 , n18576 , n18577 );
nand ( n18579 , n18578 , n920 );
nand ( n18580 , n18579 , n17101 );
or ( n18581 , n18569 , n18580 );
not ( n18582 , n1066 );
and ( n18583 , n18582 , n10622 , n169 );
nor ( n18584 , n18583 , n10609 );
nand ( n18585 , n18581 , n18584 );
not ( n18586 , n18585 );
not ( n18587 , n830 );
not ( n18588 , n952 );
and ( n18589 , n18587 , n18588 );
nand ( n18590 , n835 , n812 );
and ( n18591 , n18590 , n995 );
nor ( n18592 , n18589 , n18591 );
not ( n18593 , n10566 );
not ( n18594 , n1037 );
or ( n18595 , n18593 , n18594 );
nand ( n18596 , n18595 , n169 );
and ( n18597 , n756 , n974 , n801 );
nor ( n18598 , n18597 , n1050 );
and ( n18599 , n18592 , n18596 , n18598 );
not ( n18600 , n1041 );
not ( n18601 , n919 );
or ( n18602 , n18600 , n18601 );
nand ( n18603 , n18602 , n167 );
not ( n18604 , n1057 );
nand ( n18605 , n18604 , n857 );
not ( n18606 , n10544 );
or ( n18607 , n18605 , n18606 );
nand ( n18608 , n18607 , n10609 );
and ( n18609 , n18599 , n18603 , n18608 );
not ( n18610 , n18609 );
or ( n18611 , n18586 , n18610 );
not ( n18612 , n10534 );
or ( n18613 , n18612 , n797 );
nand ( n18614 , n18613 , n847 );
nand ( n18615 , n18614 , n1013 , n10754 , n1230 );
nor ( n18616 , n18569 , n18615 );
or ( n18617 , n18616 , n169 );
nor ( n18618 , n935 , n766 );
not ( n18619 , n1235 );
not ( n18620 , n972 );
or ( n18621 , n18619 , n18620 );
nand ( n18622 , n18621 , n1186 );
nand ( n18623 , n18618 , n18622 );
and ( n18624 , n18623 , n920 );
nand ( n18625 , n904 , n169 );
and ( n18626 , n18625 , n10667 , n10536 );
buf ( n18627 , n1018 );
or ( n18628 , n18626 , n18627 );
not ( n18629 , n1001 );
not ( n18630 , n779 );
and ( n18631 , n18629 , n18630 );
not ( n18632 , n756 );
not ( n18633 , n10624 );
or ( n18634 , n18632 , n18633 );
nand ( n18635 , n18634 , n1050 );
nor ( n18636 , n18631 , n18635 );
nand ( n18637 , n18628 , n18636 );
nor ( n18638 , n18624 , n18637 );
nand ( n18639 , n18617 , n18638 );
nand ( n18640 , n18611 , n18639 );
not ( n18641 , n950 );
not ( n18642 , n10666 );
or ( n18643 , n18641 , n18642 );
nand ( n18644 , n18643 , n1178 );
or ( n18645 , n747 , n1205 );
nand ( n18646 , n18645 , n785 );
or ( n18647 , n18646 , n886 );
nand ( n18648 , n18647 , n10609 );
not ( n18649 , n1158 );
and ( n18650 , n18649 , n756 );
nor ( n18651 , n18650 , n874 );
and ( n18652 , n18644 , n18648 , n18651 );
nand ( n18653 , n18640 , n18652 );
not ( n18654 , n18653 );
and ( n18655 , n18556 , n18654 );
and ( n18656 , n18653 , n18351 );
nor ( n18657 , n18655 , n18656 );
not ( n18658 , n18657 );
and ( n18659 , n18555 , n18658 );
not ( n18660 , n18555 );
and ( n18661 , n18660 , n18657 );
nor ( n18662 , n18659 , n18661 );
xnor ( n18663 , n218 , n12244 );
not ( n18664 , n18663 );
and ( n18665 , n18662 , n18664 );
not ( n18666 , n18662 );
and ( n18667 , n18666 , n18663 );
nor ( n18668 , n18665 , n18667 );
or ( n18669 , n18668 , n1 );
xnor ( n18670 , n217 , n218 );
or ( n18671 , n2246 , n18670 );
nand ( n18672 , n18669 , n18671 );
not ( n18673 , n230 );
not ( n18674 , n18673 );
not ( n18675 , n18054 );
or ( n18676 , n18674 , n18675 );
or ( n18677 , n18058 , n18673 );
nand ( n18678 , n18676 , n18677 );
and ( n18679 , n18678 , n10336 );
not ( n18680 , n18678 );
buf ( n18681 , n10331 );
and ( n18682 , n18680 , n18681 );
or ( n18683 , n18679 , n18682 );
buf ( n18684 , n18232 );
and ( n18685 , n18684 , n17927 );
not ( n18686 , n18684 );
and ( n18687 , n18686 , n17917 );
nor ( n18688 , n18685 , n18687 );
not ( n18689 , n18688 );
and ( n18690 , n18683 , n18689 );
not ( n18691 , n18683 );
and ( n18692 , n18691 , n18688 );
nor ( n18693 , n18690 , n18692 );
or ( n18694 , n18693 , n1 );
and ( n18695 , n231 , n18673 );
not ( n18696 , n231 );
and ( n18697 , n18696 , n230 );
nor ( n18698 , n18695 , n18697 );
or ( n18699 , n2246 , n18698 );
nand ( n18700 , n18694 , n18699 );
nor ( n18701 , n3153 , n3042 , n3114 );
not ( n18702 , n18701 );
not ( n18703 , n10000 );
or ( n18704 , n18702 , n18703 );
nand ( n18705 , n10126 , n3235 );
nand ( n18706 , n18704 , n18705 );
and ( n18707 , n10061 , n3209 , n3094 );
nor ( n18708 , n18707 , n15214 );
nor ( n18709 , n15156 , n15260 );
nand ( n18710 , n3212 , n10091 );
nand ( n18711 , n18709 , n15459 , n3085 , n18710 );
nor ( n18712 , n18708 , n18711 );
or ( n18713 , n18706 , n18712 );
or ( n18714 , n17874 , n15467 );
nand ( n18715 , n18714 , n3199 );
and ( n18716 , n15146 , n15508 , n15172 , n119 );
and ( n18717 , n18715 , n18716 );
nand ( n18718 , n18713 , n18717 );
not ( n18719 , n15155 );
nand ( n18720 , n18719 , n3122 );
or ( n18721 , n18720 , n16009 );
nand ( n18722 , n18721 , n3164 );
and ( n18723 , n3230 , n118 );
not ( n18724 , n3226 );
not ( n18725 , n10009 );
or ( n18726 , n18724 , n18725 );
nand ( n18727 , n18726 , n117 );
nand ( n18728 , n18722 , n18723 , n18727 );
not ( n18729 , n3048 );
not ( n18730 , n3266 );
or ( n18731 , n18729 , n18730 );
nand ( n18732 , n18731 , n17905 );
and ( n18733 , n18728 , n18732 );
nor ( n18734 , n18733 , n10133 );
not ( n18735 , n3137 );
not ( n18736 , n3221 );
or ( n18737 , n18735 , n18736 );
nand ( n18738 , n15177 , n18014 );
nand ( n18739 , n18737 , n18738 );
nand ( n18740 , n18734 , n18739 );
nand ( n18741 , n18718 , n18740 );
nand ( n18742 , n15157 , n17904 , n10113 , n10037 );
not ( n18743 , n18742 );
not ( n18744 , n3086 );
not ( n18745 , n16033 );
nand ( n18746 , n18744 , n18745 , n17885 , n10035 );
not ( n18747 , n18746 );
or ( n18748 , n18743 , n18747 );
and ( n18749 , n3204 , n10030 );
nor ( n18750 , n18749 , n15171 );
nand ( n18751 , n18748 , n18750 );
and ( n18752 , n3191 , n115 );
nor ( n18753 , n18752 , n3106 );
not ( n18754 , n18753 );
not ( n18755 , n16038 );
not ( n18756 , n18755 );
or ( n18757 , n18754 , n18756 );
nand ( n18758 , n18757 , n3234 );
nand ( n18759 , n18758 , n10104 );
nand ( n18760 , n18751 , n18759 );
or ( n18761 , n15197 , n3071 );
or ( n18762 , n116 , n10110 );
nand ( n18763 , n18761 , n18762 , n3209 );
and ( n18764 , n18763 , n3235 );
not ( n18765 , n3194 );
not ( n18766 , n18765 );
not ( n18767 , n3082 );
or ( n18768 , n18766 , n18767 );
and ( n18769 , n3247 , n117 );
nand ( n18770 , n18768 , n18769 );
nand ( n18771 , n18770 , n18033 );
nor ( n18772 , n18764 , n18771 );
and ( n18773 , n18741 , n18760 , n18772 );
not ( n18774 , n18773 );
not ( n18775 , n238 );
and ( n18776 , n18774 , n18775 );
and ( n18777 , n18773 , n238 );
nor ( n18778 , n18776 , n18777 );
not ( n18779 , n18778 );
not ( n18780 , n17497 );
or ( n18781 , n18779 , n18780 );
or ( n18782 , n17497 , n18778 );
nand ( n18783 , n18781 , n18782 );
and ( n18784 , n18783 , n16106 );
not ( n18785 , n18783 );
and ( n18786 , n18785 , n16109 );
nor ( n18787 , n18784 , n18786 );
or ( n18788 , n18787 , n1 );
xnor ( n18789 , n238 , n239 );
or ( n18790 , n2246 , n18789 );
nand ( n18791 , n18788 , n18790 );
not ( n18792 , n11053 );
buf ( n18793 , n17806 );
not ( n18794 , n18793 );
or ( n18795 , n18792 , n18794 );
or ( n18796 , n18793 , n11053 );
nand ( n18797 , n18795 , n18796 );
xor ( n18798 , n240 , n17014 );
buf ( n18799 , n11828 );
xor ( n18800 , n18798 , n18799 );
not ( n18801 , n18800 );
and ( n18802 , n18797 , n18801 );
not ( n18803 , n18797 );
and ( n18804 , n18803 , n18800 );
nor ( n18805 , n18802 , n18804 );
or ( n18806 , n18805 , n1 );
xnor ( n18807 , n240 , n241 );
or ( n18808 , n2246 , n18807 );
nand ( n18809 , n18806 , n18808 );
not ( n18810 , n12986 );
not ( n18811 , n10654 );
and ( n18812 , n18810 , n18811 );
and ( n18813 , n12986 , n10654 );
nor ( n18814 , n18812 , n18813 );
not ( n18815 , n18814 );
not ( n18816 , n18815 );
not ( n18817 , n18793 );
not ( n18818 , n18817 );
or ( n18819 , n18816 , n18818 );
nand ( n18820 , n18814 , n18793 );
nand ( n18821 , n18819 , n18820 );
xor ( n18822 , n242 , n11828 );
not ( n18823 , n18822 );
and ( n18824 , n18821 , n18823 );
not ( n18825 , n18821 );
and ( n18826 , n18825 , n18822 );
nor ( n18827 , n18824 , n18826 );
or ( n18828 , n18827 , n1 );
xnor ( n18829 , n242 , n243 );
or ( n18830 , n2246 , n18829 );
nand ( n18831 , n18828 , n18830 );
not ( n18832 , n18657 );
not ( n18833 , n255 );
not ( n18834 , n13487 );
or ( n18835 , n18833 , n18834 );
or ( n18836 , n17955 , n255 );
nand ( n18837 , n18835 , n18836 );
not ( n18838 , n18837 );
or ( n18839 , n18832 , n18838 );
or ( n18840 , n18657 , n18837 );
nand ( n18841 , n18839 , n18840 );
and ( n18842 , n18841 , n18446 );
not ( n18843 , n18841 );
not ( n18844 , n18446 );
and ( n18845 , n18843 , n18844 );
nor ( n18846 , n18842 , n18845 );
or ( n18847 , n18846 , n1 );
xnor ( n18848 , n254 , n255 );
or ( n18849 , n2246 , n18848 );
nand ( n18850 , n18847 , n18849 );
not ( n18851 , n17199 );
not ( n18852 , n17168 );
or ( n18853 , n18851 , n18852 );
nand ( n18854 , n18853 , n17237 );
not ( n18855 , n250 );
xor ( n18856 , n18854 , n18855 );
xnor ( n18857 , n18856 , n15792 );
not ( n18858 , n15423 );
not ( n18859 , n3019 );
and ( n18860 , n18858 , n18859 );
and ( n18861 , n3019 , n15423 );
nor ( n18862 , n18860 , n18861 );
not ( n18863 , n18862 );
not ( n18864 , n18863 );
not ( n18865 , n16106 );
or ( n18866 , n18864 , n18865 );
or ( n18867 , n16106 , n18863 );
nand ( n18868 , n18866 , n18867 );
not ( n18869 , n18868 );
and ( n18870 , n18857 , n18869 );
not ( n18871 , n18857 );
and ( n18872 , n18871 , n18868 );
nor ( n18873 , n18870 , n18872 );
or ( n18874 , n18873 , n1 );
and ( n18875 , n251 , n18855 );
not ( n18876 , n251 );
and ( n18877 , n18876 , n250 );
nor ( n18878 , n18875 , n18877 );
or ( n18879 , n2246 , n18878 );
nand ( n18880 , n18874 , n18879 );
and ( n18881 , n1227 , n843 , n990 );
not ( n18882 , n18881 );
not ( n18883 , n10566 );
or ( n18884 , n18882 , n18883 );
nand ( n18885 , n18884 , n169 );
not ( n18886 , n18885 );
nand ( n18887 , n974 , n834 , n10703 );
and ( n18888 , n18887 , n961 );
nor ( n18889 , n18888 , n755 );
nor ( n18890 , n826 , n18889 );
nand ( n18891 , n10667 , n791 );
or ( n18892 , n10530 , n18891 );
nand ( n18893 , n18892 , n805 );
and ( n18894 , n18890 , n18893 );
nand ( n18895 , n793 , n798 );
not ( n18896 , n18895 );
not ( n18897 , n1244 );
or ( n18898 , n18896 , n18897 );
not ( n18899 , n914 );
nand ( n18900 , n18898 , n18899 );
nand ( n18901 , n18900 , n779 );
not ( n18902 , n987 );
not ( n18903 , n18899 );
or ( n18904 , n18902 , n18903 );
nand ( n18905 , n18904 , n167 );
not ( n18906 , n1073 );
not ( n18907 , n1170 );
or ( n18908 , n18906 , n18907 );
nand ( n18909 , n18908 , n995 );
nand ( n18910 , n18894 , n18901 , n18905 , n18909 );
or ( n18911 , n18886 , n18910 );
not ( n18912 , n1034 );
not ( n18913 , n1061 );
or ( n18914 , n18912 , n18913 );
nand ( n18915 , n770 , n783 );
nand ( n18916 , n920 , n18582 , n18915 , n832 );
nand ( n18917 , n18914 , n18916 );
or ( n18918 , n778 , n163 );
not ( n18919 , n1184 );
not ( n18920 , n760 );
not ( n18921 , n18920 );
and ( n18922 , n18919 , n18921 );
nor ( n18923 , n18922 , n10577 );
and ( n18924 , n10541 , n857 , n18918 , n18923 );
nand ( n18925 , n18917 , n18924 );
not ( n18926 , n18925 );
nand ( n18927 , n10663 , n834 );
not ( n18928 , n10536 );
not ( n18929 , n952 );
and ( n18930 , n18928 , n18929 );
and ( n18931 , n989 , n1019 );
nor ( n18932 , n18930 , n18931 );
nand ( n18933 , n18927 , n18932 , n1233 , n779 );
not ( n18934 , n18933 );
or ( n18935 , n18926 , n18934 );
nand ( n18936 , n10741 , n905 , n10632 );
and ( n18937 , n18936 , n167 );
not ( n18938 , n871 );
not ( n18939 , n18574 );
or ( n18940 , n18938 , n18939 );
and ( n18941 , n18562 , n1041 , n1050 );
nand ( n18942 , n18940 , n18941 );
nor ( n18943 , n18937 , n18942 );
nand ( n18944 , n18935 , n18943 );
nand ( n18945 , n18911 , n18944 );
not ( n18946 , n18899 );
not ( n18947 , n839 );
or ( n18948 , n18946 , n18947 );
not ( n18949 , n18627 );
nand ( n18950 , n18948 , n18949 );
nor ( n18951 , n17039 , n1166 );
nand ( n18952 , n784 , n779 );
nor ( n18953 , n18951 , n18952 );
not ( n18954 , n1001 );
not ( n18955 , n10667 );
or ( n18956 , n18954 , n18955 );
nand ( n18957 , n18956 , n805 );
nand ( n18958 , n17027 , n1010 );
and ( n18959 , n18953 , n18957 , n18958 );
nand ( n18960 , n18950 , n18959 );
not ( n18961 , n10700 );
or ( n18962 , n18961 , n10541 );
and ( n18963 , n935 , n167 );
not ( n18964 , n18562 );
nor ( n18965 , n18963 , n18964 );
nand ( n18966 , n18962 , n18965 );
and ( n18967 , n18960 , n18966 );
not ( n18968 , n806 );
nand ( n18969 , n18968 , n1158 );
and ( n18970 , n10567 , n18969 );
nor ( n18971 , n18967 , n18970 );
nand ( n18972 , n18945 , n18971 );
buf ( n18973 , n18972 );
xor ( n18974 , n18973 , n13369 );
xor ( n18975 , n260 , n12122 );
xnor ( n18976 , n18975 , n12244 );
xnor ( n18977 , n18974 , n18976 );
or ( n18978 , n18977 , n1 );
xnor ( n18979 , n260 , n261 );
or ( n18980 , n2246 , n18979 );
nand ( n18981 , n18978 , n18980 );
not ( n18982 , n9708 );
nand ( n18983 , n4172 , n203 );
not ( n18984 , n5217 );
not ( n18985 , n14614 );
or ( n18986 , n18984 , n18985 );
nand ( n18987 , n18986 , n5132 );
not ( n18988 , n14599 );
or ( n18989 , n4028 , n4035 , n18988 );
nand ( n18990 , n18989 , n4078 );
and ( n18991 , n18983 , n18987 , n18990 );
not ( n18992 , n18991 );
and ( n18993 , n5875 , n5090 , n202 );
nand ( n18994 , n18993 , n4182 , n4191 );
not ( n18995 , n14595 );
nand ( n18996 , n18995 , n4193 );
and ( n18997 , n18994 , n18996 );
nand ( n18998 , n4145 , n5158 );
not ( n18999 , n13161 );
nand ( n19000 , n3992 , n200 );
not ( n19001 , n19000 );
or ( n19002 , n18999 , n19001 );
nand ( n19003 , n19002 , n4068 );
nand ( n19004 , n4007 , n4121 , n4025 );
nand ( n19005 , n18998 , n19003 , n19004 , n204 );
nor ( n19006 , n18997 , n19005 );
not ( n19007 , n19006 );
or ( n19008 , n18992 , n19007 );
not ( n19009 , n5224 );
not ( n19010 , n5815 );
or ( n19011 , n19009 , n19010 );
nand ( n19012 , n19011 , n3986 );
nand ( n19013 , n4193 , n5132 );
nor ( n19014 , n5174 , n19013 );
nand ( n19015 , n19012 , n19014 );
nand ( n19016 , n4107 , n199 );
and ( n19017 , n19016 , n5829 );
nor ( n19018 , n19017 , n5179 );
or ( n19019 , n19015 , n19018 );
and ( n19020 , n13132 , n4051 );
nor ( n19021 , n5689 , n19020 );
not ( n19022 , n203 );
not ( n19023 , n4191 );
or ( n19024 , n19022 , n19023 );
nand ( n19025 , n19024 , n4077 );
nand ( n19026 , n19021 , n19025 );
nand ( n19027 , n19019 , n19026 );
and ( n19028 , n3975 , n199 );
nor ( n19029 , n19028 , n5183 );
nand ( n19030 , n5185 , n4058 );
nor ( n19031 , n19029 , n19030 );
not ( n19032 , n19031 );
and ( n19033 , n13178 , n3986 );
nor ( n19034 , n19033 , n13107 );
not ( n19035 , n19034 );
or ( n19036 , n19032 , n19035 );
not ( n19037 , n5691 );
nand ( n19038 , n19037 , n4151 , n5781 );
nand ( n19039 , n19036 , n19038 );
nand ( n19040 , n19027 , n19039 );
nand ( n19041 , n19008 , n19040 );
not ( n19042 , n14555 );
nand ( n19043 , n4136 , n3996 );
or ( n19044 , n19043 , n17732 );
or ( n19045 , n4049 , n3996 );
nand ( n19046 , n19044 , n19045 );
not ( n19047 , n19046 );
not ( n19048 , n203 );
or ( n19049 , n19047 , n19048 );
nand ( n19050 , n19049 , n4120 );
not ( n19051 , n19050 );
or ( n19052 , n19042 , n19051 );
nand ( n19053 , n4136 , n5158 );
or ( n19054 , n5675 , n19053 , n13101 );
or ( n19055 , n5190 , n5128 , n203 );
nand ( n19056 , n19054 , n19055 );
not ( n19057 , n5178 );
nor ( n19058 , n19057 , n17658 );
nand ( n19059 , n19056 , n19058 );
nand ( n19060 , n19052 , n19059 );
not ( n19061 , n13161 );
nand ( n19062 , n19061 , n4087 );
and ( n19063 , n5177 , n4052 , n19062 , n13102 );
and ( n19064 , n19041 , n19060 , n19063 );
not ( n19065 , n19064 );
and ( n19066 , n18982 , n19065 );
and ( n19067 , n9708 , n19064 );
nor ( n19068 , n19066 , n19067 );
not ( n19069 , n19068 );
not ( n19070 , n262 );
not ( n19071 , n4362 );
or ( n19072 , n19070 , n19071 );
or ( n19073 , n5395 , n262 );
nand ( n19074 , n19072 , n19073 );
not ( n19075 , n19074 );
and ( n19076 , n19069 , n19075 );
and ( n19077 , n19068 , n19074 );
nor ( n19078 , n19076 , n19077 );
not ( n19079 , n9819 );
and ( n19080 , n19078 , n19079 );
not ( n19081 , n19078 );
and ( n19082 , n19081 , n9819 );
nor ( n19083 , n19080 , n19082 );
or ( n19084 , n19083 , n1 );
xnor ( n19085 , n262 , n263 );
or ( n19086 , n2246 , n19085 );
nand ( n19087 , n19084 , n19086 );
xor ( n19088 , n15031 , n10172 );
not ( n19089 , n299 );
nor ( n19090 , n10194 , n2274 );
nor ( n19091 , n2325 , n10276 );
nor ( n19092 , n19091 , n2295 );
and ( n19093 , n19090 , n19092 , n2497 );
and ( n19094 , n15682 , n2395 , n16233 , n2265 );
or ( n19095 , n19093 , n19094 );
not ( n19096 , n2410 );
nor ( n19097 , n19096 , n2504 );
nand ( n19098 , n19095 , n19097 );
not ( n19099 , n14704 );
not ( n19100 , n10315 );
or ( n19101 , n19099 , n19100 );
nand ( n19102 , n19101 , n2424 );
nor ( n19103 , n10251 , n2316 );
nand ( n19104 , n15632 , n19103 );
nor ( n19105 , n19104 , n10274 );
nand ( n19106 , n19102 , n2299 , n19105 );
nand ( n19107 , n19098 , n19106 );
and ( n19108 , n14750 , n17352 );
not ( n19109 , n14732 );
not ( n19110 , n14674 );
or ( n19111 , n19109 , n19110 );
nand ( n19112 , n19111 , n134 );
nand ( n19113 , n19112 , n2506 );
and ( n19114 , n10309 , n19108 , n19113 );
not ( n19115 , n10240 );
not ( n19116 , n2270 );
or ( n19117 , n19115 , n19116 );
nand ( n19118 , n19117 , n16284 );
nand ( n19119 , n19118 , n2424 );
and ( n19120 , n14723 , n17347 , n19119 , n16248 );
or ( n19121 , n19114 , n19120 );
and ( n19122 , n2357 , n2389 );
and ( n19123 , n2293 , n2324 );
nor ( n19124 , n19122 , n19123 );
not ( n19125 , n19124 );
not ( n19126 , n10177 );
or ( n19127 , n19125 , n19126 );
nand ( n19128 , n14672 , n2424 );
nor ( n19129 , n14657 , n19128 );
nand ( n19130 , n19129 , n10315 );
nand ( n19131 , n19127 , n19130 );
and ( n19132 , n19131 , n10304 );
nand ( n19133 , n19121 , n19132 );
nand ( n19134 , n19133 , n135 );
not ( n19135 , n10250 );
not ( n19136 , n15594 );
or ( n19137 , n19135 , n19136 );
nand ( n19138 , n19137 , n2432 );
not ( n19139 , n14652 );
not ( n19140 , n2289 );
or ( n19141 , n19139 , n19140 );
nand ( n19142 , n19141 , n2470 );
not ( n19143 , n19142 );
or ( n19144 , n19138 , n19143 );
not ( n19145 , n2424 );
not ( n19146 , n15593 );
not ( n19147 , n10213 );
or ( n19148 , n19146 , n19147 );
nand ( n19149 , n19148 , n14720 );
not ( n19150 , n19149 );
or ( n19151 , n19145 , n19150 );
nand ( n19152 , n2394 , n14653 );
and ( n19153 , n15540 , n19152 , n10178 , n134 );
nand ( n19154 , n19151 , n19153 );
nand ( n19155 , n19144 , n19154 );
not ( n19156 , n19155 );
not ( n19157 , n131 );
not ( n19158 , n2499 );
nor ( n19159 , n19158 , n14735 );
not ( n19160 , n19159 );
or ( n19161 , n19157 , n19160 );
nor ( n19162 , n14675 , n2301 );
or ( n19163 , n19162 , n16288 );
nand ( n19164 , n19161 , n19163 );
nor ( n19165 , n2504 , n19164 );
not ( n19166 , n19165 );
or ( n19167 , n19156 , n19166 );
nand ( n19168 , n19167 , n2359 );
and ( n19169 , n15729 , n2461 );
and ( n19170 , n2377 , n2477 );
nor ( n19171 , n19169 , n19170 );
nand ( n19172 , n19107 , n19134 , n19168 , n19171 );
not ( n19173 , n19172 );
not ( n19174 , n19173 );
or ( n19175 , n19089 , n19174 );
not ( n19176 , n299 );
nand ( n19177 , n19176 , n19172 );
nand ( n19178 , n19175 , n19177 );
buf ( n19179 , n16340 );
not ( n19180 , n19179 );
and ( n19181 , n19178 , n19180 );
not ( n19182 , n19178 );
and ( n19183 , n19182 , n19179 );
nor ( n19184 , n19181 , n19183 );
xnor ( n19185 , n19088 , n19184 );
or ( n19186 , n19185 , n1 );
and ( n19187 , n300 , n19176 );
not ( n19188 , n300 );
and ( n19189 , n19188 , n299 );
nor ( n19190 , n19187 , n19189 );
or ( n19191 , n2246 , n19190 );
nand ( n19192 , n19186 , n19191 );
xor ( n19193 , n15140 , n10172 );
not ( n19194 , n305 );
not ( n19195 , n19173 );
or ( n19196 , n19194 , n19195 );
not ( n19197 , n305 );
nand ( n19198 , n19197 , n19172 );
nand ( n19199 , n19196 , n19198 );
buf ( n19200 , n16221 );
and ( n19201 , n19199 , n19200 );
not ( n19202 , n19199 );
not ( n19203 , n19200 );
and ( n19204 , n19202 , n19203 );
nor ( n19205 , n19201 , n19204 );
xnor ( n19206 , n19193 , n19205 );
or ( n19207 , n19206 , n1 );
and ( n19208 , n306 , n19197 );
not ( n19209 , n306 );
and ( n19210 , n19209 , n305 );
nor ( n19211 , n19208 , n19210 );
or ( n19212 , n2246 , n19211 );
nand ( n19213 , n19207 , n19212 );
xor ( n19214 , n17800 , n16970 );
not ( n19215 , n313 );
not ( n19216 , n10898 );
or ( n19217 , n19215 , n19216 );
or ( n19218 , n10898 , n313 );
nand ( n19219 , n19217 , n19218 );
xnor ( n19220 , n19214 , n19219 );
or ( n19221 , n19220 , n1 );
xnor ( n19222 , n313 , n314 );
or ( n19223 , n2246 , n19222 );
nand ( n19224 , n19221 , n19223 );
xnor ( n19225 , n15278 , n15030 );
not ( n19226 , n307 );
not ( n19227 , n19173 );
or ( n19228 , n19226 , n19227 );
or ( n19229 , n307 , n19173 );
nand ( n19230 , n19228 , n19229 );
xor ( n19231 , n19225 , n19230 );
not ( n19232 , n18041 );
nand ( n19233 , n17880 , n17835 , n17903 , n17912 );
not ( n19234 , n19233 );
or ( n19235 , n19232 , n19234 );
nand ( n19236 , n18240 , n18042 );
nand ( n19237 , n19235 , n19236 );
not ( n19238 , n19237 );
not ( n19239 , n14898 );
and ( n19240 , n19238 , n19239 );
and ( n19241 , n19237 , n14898 );
nor ( n19242 , n19240 , n19241 );
not ( n19243 , n19242 );
and ( n19244 , n19231 , n19243 );
not ( n19245 , n19231 );
and ( n19246 , n19245 , n19242 );
nor ( n19247 , n19244 , n19246 );
or ( n19248 , n19247 , n1 );
xnor ( n19249 , n307 , n308 );
or ( n19250 , n2246 , n19249 );
nand ( n19251 , n19248 , n19250 );
xor ( n19252 , n326 , n13358 );
not ( n19253 , n12244 );
xor ( n19254 , n19252 , n19253 );
not ( n19255 , n1803 );
not ( n19256 , n19255 );
not ( n19257 , n12000 );
not ( n19258 , n18972 );
not ( n19259 , n19258 );
or ( n19260 , n19257 , n19259 );
nand ( n19261 , n18972 , n11999 );
nand ( n19262 , n19260 , n19261 );
not ( n19263 , n19262 );
or ( n19264 , n19256 , n19263 );
or ( n19265 , n19255 , n19262 );
nand ( n19266 , n19264 , n19265 );
and ( n19267 , n19254 , n19266 );
not ( n19268 , n19254 );
not ( n19269 , n19266 );
and ( n19270 , n19268 , n19269 );
nor ( n19271 , n19267 , n19270 );
or ( n19272 , n19271 , n1 );
xnor ( n19273 , n326 , n327 );
or ( n19274 , n2246 , n19273 );
nand ( n19275 , n19272 , n19274 );
not ( n19276 , n5393 );
not ( n19277 , n5087 );
or ( n19278 , n19276 , n19277 );
nand ( n19279 , n5248 , n5392 );
nand ( n19280 , n19278 , n19279 );
and ( n19281 , n11288 , n340 );
not ( n19282 , n11288 );
not ( n19283 , n340 );
and ( n19284 , n19282 , n19283 );
nor ( n19285 , n19281 , n19284 );
and ( n19286 , n19280 , n19285 );
not ( n19287 , n19280 );
not ( n19288 , n19285 );
and ( n19289 , n19287 , n19288 );
nor ( n19290 , n19286 , n19289 );
nand ( n19291 , n19290 , n2246 );
not ( n19292 , n17756 );
not ( n19293 , n19292 );
not ( n19294 , n16838 );
not ( n19295 , n19294 );
or ( n19296 , n19293 , n19295 );
nand ( n19297 , n16838 , n17756 );
nand ( n19298 , n19296 , n19297 );
not ( n19299 , n19298 );
not ( n19300 , n5893 );
not ( n19301 , n4362 );
or ( n19302 , n19300 , n19301 );
not ( n19303 , n4362 );
nand ( n19304 , n5779 , n19303 );
nand ( n19305 , n19302 , n19304 );
not ( n19306 , n19305 );
or ( n19307 , n19299 , n19306 );
or ( n19308 , n19305 , n19298 );
nand ( n19309 , n19307 , n19308 );
or ( n19310 , n19291 , n19309 );
and ( n19311 , n341 , n19283 );
not ( n19312 , n341 );
and ( n19313 , n19312 , n340 );
nor ( n19314 , n19311 , n19313 );
or ( n19315 , n19314 , n2246 );
not ( n19316 , n19290 );
nand ( n19317 , n19309 , n19316 , n2246 );
nand ( n19318 , n19310 , n19315 , n19317 );
not ( n19319 , n349 );
xnor ( n19320 , n2512 , n19319 );
and ( n19321 , n19320 , n18681 );
not ( n19322 , n19320 );
and ( n19323 , n19322 , n10336 );
nor ( n19324 , n19321 , n19323 );
buf ( n19325 , n3430 );
and ( n19326 , n19325 , n17927 );
not ( n19327 , n19325 );
and ( n19328 , n19327 , n17917 );
nor ( n19329 , n19326 , n19328 );
not ( n19330 , n19329 );
and ( n19331 , n19324 , n19330 );
not ( n19332 , n19324 );
and ( n19333 , n19332 , n19329 );
nor ( n19334 , n19331 , n19333 );
or ( n19335 , n19334 , n1 );
and ( n19336 , n350 , n19319 );
not ( n19337 , n350 );
and ( n19338 , n19337 , n349 );
nor ( n19339 , n19336 , n19338 );
or ( n19340 , n2246 , n19339 );
nand ( n19341 , n19335 , n19340 );
xor ( n19342 , n355 , n12987 );
xnor ( n19343 , n19342 , n17014 );
not ( n19344 , n17107 );
not ( n19345 , n17641 );
or ( n19346 , n19344 , n19345 );
or ( n19347 , n17641 , n17107 );
nand ( n19348 , n19346 , n19347 );
not ( n19349 , n19348 );
and ( n19350 , n19343 , n19349 );
not ( n19351 , n19343 );
and ( n19352 , n19351 , n19348 );
nor ( n19353 , n19350 , n19352 );
or ( n19354 , n19353 , n1 );
xnor ( n19355 , n355 , n356 );
or ( n19356 , n2246 , n19355 );
nand ( n19357 , n19354 , n19356 );
buf ( n19358 , n14619 );
xor ( n19359 , n19358 , n13222 );
xor ( n19360 , n359 , n12662 );
xnor ( n19361 , n19360 , n12770 );
xnor ( n19362 , n19359 , n19361 );
or ( n19363 , n19362 , n1 );
xnor ( n19364 , n359 , n360 );
or ( n19365 , n2246 , n19364 );
nand ( n19366 , n19363 , n19365 );
nand ( n19367 , n15881 , n14974 );
and ( n19368 , n19367 , n2609 );
nor ( n19369 , n19368 , n144 );
not ( n19370 , n19369 );
not ( n19371 , n17221 );
or ( n19372 , n14995 , n19371 );
nand ( n19373 , n3321 , n2539 , n2580 );
nand ( n19374 , n19372 , n19373 );
and ( n19375 , n14984 , n2615 , n3352 );
nand ( n19376 , n19374 , n19375 );
nand ( n19377 , n2614 , n2686 );
or ( n19378 , n19377 , n14982 );
and ( n19379 , n138 , n142 );
nand ( n19380 , n2575 , n19379 );
or ( n19381 , n19380 , n141 );
nand ( n19382 , n19378 , n19381 );
not ( n19383 , n2547 );
and ( n19384 , n140 , n143 );
and ( n19385 , n19383 , n2583 , n19384 );
nor ( n19386 , n19382 , n19385 );
and ( n19387 , n19386 , n16207 , n16126 );
not ( n19388 , n19387 );
or ( n19389 , n19376 , n19388 );
not ( n19390 , n3384 );
nand ( n19391 , n19390 , n3381 , n143 );
and ( n19392 , n2717 , n2680 , n19391 , n16135 );
nand ( n19393 , n3391 , n19392 );
not ( n19394 , n142 );
nand ( n19395 , n19394 , n2590 , n2720 );
and ( n19396 , n3323 , n19395 , n16181 );
nor ( n19397 , n14950 , n15021 , n3425 );
or ( n19398 , n19396 , n19397 );
nand ( n19399 , n19398 , n15881 );
or ( n19400 , n19393 , n19399 );
nand ( n19401 , n19389 , n19400 );
not ( n19402 , n19401 );
or ( n19403 , n19370 , n19402 );
not ( n19404 , n2517 );
not ( n19405 , n19383 );
or ( n19406 , n19404 , n19405 );
nand ( n19407 , n19406 , n2626 );
or ( n19408 , n19407 , n14903 );
nand ( n19409 , n19408 , n141 );
not ( n19410 , n2755 );
not ( n19411 , n2618 );
not ( n19412 , n3384 );
or ( n19413 , n19411 , n19412 );
nand ( n19414 , n19413 , n14939 );
nor ( n19415 , n19410 , n19414 , n15871 );
nand ( n19416 , n19409 , n19415 );
nor ( n19417 , n19416 , n3347 );
not ( n19418 , n19417 );
not ( n19419 , n19387 );
or ( n19420 , n19418 , n19419 );
not ( n19421 , n19399 );
not ( n19422 , n3411 );
not ( n19423 , n3361 );
or ( n19424 , n19422 , n19423 );
nand ( n19425 , n19424 , n141 );
not ( n19426 , n19383 );
not ( n19427 , n2568 );
or ( n19428 , n19426 , n19427 );
nand ( n19429 , n19428 , n3319 );
nor ( n19430 , n19429 , n15009 , n17138 );
nand ( n19431 , n19421 , n19425 , n19430 );
nand ( n19432 , n19420 , n19431 );
not ( n19433 , n17158 );
not ( n19434 , n14969 );
or ( n19435 , n19433 , n19434 , n3370 );
nand ( n19436 , n19435 , n2585 );
nor ( n19437 , n2672 , n2604 );
or ( n19438 , n19437 , n17177 , n2564 );
nand ( n19439 , n19438 , n3284 );
and ( n19440 , n14955 , n19436 , n17433 , n19439 );
nand ( n19441 , n19432 , n19440 );
nand ( n19442 , n19403 , n19441 );
not ( n19443 , n3305 );
nand ( n19444 , n19443 , n17211 );
and ( n19445 , n19444 , n2639 );
or ( n19446 , n14964 , n2669 );
nand ( n19447 , n19446 , n17170 );
nor ( n19448 , n19445 , n19447 );
nand ( n19449 , n19442 , n19448 );
not ( n19450 , n19449 );
and ( n19451 , n19450 , n15140 );
not ( n19452 , n19450 );
and ( n19453 , n19452 , n15141 );
nor ( n19454 , n19451 , n19453 );
xnor ( n19455 , n19454 , n19237 );
not ( n19456 , n19173 );
not ( n19457 , n15030 );
or ( n19458 , n19456 , n19457 );
nand ( n19459 , n15031 , n19172 );
nand ( n19460 , n19458 , n19459 );
not ( n19461 , n361 );
buf ( n19462 , n18054 );
not ( n19463 , n19462 );
xor ( n19464 , n19461 , n19463 );
not ( n19465 , n19464 );
and ( n19466 , n19460 , n19465 );
not ( n19467 , n19460 );
and ( n19468 , n19467 , n19464 );
nor ( n19469 , n19466 , n19468 );
xor ( n19470 , n19455 , n19469 );
or ( n19471 , n19470 , n1 );
and ( n19472 , n362 , n19461 );
not ( n19473 , n362 );
and ( n19474 , n19473 , n361 );
nor ( n19475 , n19472 , n19474 );
or ( n19476 , n2246 , n19475 );
nand ( n19477 , n19471 , n19476 );
xor ( n19478 , n5491 , n13212 );
xnor ( n19479 , n19478 , n11422 );
not ( n19480 , n11293 );
not ( n19481 , n376 );
and ( n19482 , n19480 , n19481 );
and ( n19483 , n11293 , n376 );
nor ( n19484 , n19482 , n19483 );
nand ( n19485 , n19484 , n2246 );
or ( n19486 , n19479 , n19485 );
nor ( n19487 , n19484 , n1 );
nand ( n19488 , n19479 , n19487 );
xor ( n19489 , n376 , n377 );
nand ( n19490 , n19489 , n1 );
nand ( n19491 , n19486 , n19488 , n19490 );
buf ( n19492 , n9118 );
not ( n19493 , n7225 );
not ( n19494 , n18 );
and ( n19495 , n19493 , n19494 );
and ( n19496 , n7225 , n18 );
nor ( n19497 , n19495 , n19496 );
xnor ( n19498 , n19492 , n19497 );
not ( n19499 , n16537 );
not ( n19500 , n6555 );
or ( n19501 , n19499 , n19500 );
or ( n19502 , n6555 , n16537 );
nand ( n19503 , n19501 , n19502 );
nor ( n19504 , n19498 , n19503 );
or ( n19505 , n19504 , n1 );
not ( n19506 , n18 );
and ( n19507 , n35 , n19506 );
not ( n19508 , n35 );
and ( n19509 , n19508 , n18 );
nor ( n19510 , n19507 , n19509 );
or ( n19511 , n2246 , n19510 );
nand ( n19512 , n19505 , n19511 );
not ( n19513 , n7224 );
xor ( n19514 , n37 , n19513 );
xnor ( n19515 , n19514 , n16435 );
buf ( n19516 , n18077 );
not ( n19517 , n19516 );
and ( n19518 , n18106 , n19517 );
not ( n19519 , n18106 );
and ( n19520 , n19519 , n19516 );
nor ( n19521 , n19518 , n19520 );
and ( n19522 , n19515 , n19521 );
not ( n19523 , n19515 );
not ( n19524 , n19521 );
and ( n19525 , n19523 , n19524 );
nor ( n19526 , n19522 , n19525 );
or ( n19527 , n19526 , n1 );
xnor ( n19528 , n36 , n37 );
or ( n19529 , n2246 , n19528 );
nand ( n19530 , n19527 , n19529 );
not ( n19531 , n19492 );
not ( n19532 , n6962 );
or ( n19533 , n19531 , n19532 );
or ( n19534 , n19492 , n6962 );
nand ( n19535 , n19533 , n19534 );
not ( n19536 , n9216 );
xor ( n19537 , n45 , n19536 );
xnor ( n19538 , n19537 , n7225 );
not ( n19539 , n19538 );
and ( n19540 , n19535 , n19539 );
not ( n19541 , n19535 );
and ( n19542 , n19541 , n19538 );
nor ( n19543 , n19540 , n19542 );
or ( n19544 , n19543 , n1 );
xnor ( n19545 , n45 , n46 );
or ( n19546 , n2246 , n19545 );
nand ( n19547 , n19544 , n19546 );
not ( n19548 , n13818 );
xor ( n19549 , n19548 , n8006 );
xor ( n19550 , n51 , n18077 );
not ( n19551 , n16435 );
xnor ( n19552 , n19550 , n19551 );
xnor ( n19553 , n19549 , n19552 );
or ( n19554 , n19553 , n1 );
xnor ( n19555 , n51 , n52 );
or ( n19556 , n2246 , n19555 );
nand ( n19557 , n19554 , n19556 );
xor ( n19558 , n14035 , n8899 );
xor ( n19559 , n59 , n14390 );
buf ( n19560 , n13937 );
not ( n19561 , n19560 );
xor ( n19562 , n19559 , n19561 );
xnor ( n19563 , n19558 , n19562 );
or ( n19564 , n19563 , n1 );
xnor ( n19565 , n59 , n60 );
or ( n19566 , n2246 , n19565 );
nand ( n19567 , n19564 , n19566 );
not ( n19568 , n14141 );
xor ( n19569 , n11073 , n19568 );
xor ( n19570 , n63 , n14410 );
not ( n19571 , n8633 );
xnor ( n19572 , n19570 , n19571 );
xnor ( n19573 , n19569 , n19572 );
or ( n19574 , n19573 , n1 );
xnor ( n19575 , n63 , n64 );
or ( n19576 , n2246 , n19575 );
nand ( n19577 , n19574 , n19576 );
not ( n19578 , n7834 );
xor ( n19579 , n19578 , n13823 );
xor ( n19580 , n48 , n16435 );
xnor ( n19581 , n19580 , n7668 );
xnor ( n19582 , n19579 , n19581 );
or ( n19583 , n19582 , n1 );
xnor ( n19584 , n48 , n57 );
or ( n19585 , n2246 , n19584 );
nand ( n19586 , n19583 , n19585 );
xor ( n19587 , n8897 , n19568 );
xor ( n19588 , n61 , n19560 );
xnor ( n19589 , n19588 , n8633 );
xnor ( n19590 , n19587 , n19589 );
or ( n19591 , n19590 , n1 );
xnor ( n19592 , n61 , n62 );
or ( n19593 , n2246 , n19592 );
nand ( n19594 , n19591 , n19593 );
not ( n19595 , n14395 );
and ( n19596 , n58 , n19560 );
not ( n19597 , n58 );
and ( n19598 , n19597 , n13938 );
or ( n19599 , n19596 , n19598 );
not ( n19600 , n19599 );
or ( n19601 , n19595 , n19600 );
or ( n19602 , n19599 , n14395 );
nand ( n19603 , n19601 , n19602 );
and ( n19604 , n19603 , n9579 );
not ( n19605 , n19603 );
and ( n19606 , n19605 , n9578 );
nor ( n19607 , n19604 , n19606 );
or ( n19608 , n19607 , n1 );
xnor ( n19609 , n58 , n70 );
or ( n19610 , n2246 , n19609 );
nand ( n19611 , n19608 , n19610 );
not ( n19612 , n8505 );
not ( n19613 , n19612 );
not ( n19614 , n8400 );
not ( n19615 , n19614 );
or ( n19616 , n19613 , n19615 );
nand ( n19617 , n8505 , n8400 );
nand ( n19618 , n19616 , n19617 );
not ( n19619 , n19618 );
not ( n19620 , n9352 );
not ( n19621 , n80 );
not ( n19622 , n19621 );
and ( n19623 , n19620 , n19622 );
and ( n19624 , n9352 , n19621 );
nor ( n19625 , n19623 , n19624 );
not ( n19626 , n19625 );
or ( n19627 , n19619 , n19626 );
or ( n19628 , n19625 , n19618 );
nand ( n19629 , n19627 , n19628 );
and ( n19630 , n19629 , n9223 );
not ( n19631 , n19629 );
and ( n19632 , n19631 , n9224 );
nor ( n19633 , n19630 , n19632 );
or ( n19634 , n19633 , n1 );
and ( n19635 , n83 , n19621 );
not ( n19636 , n83 );
and ( n19637 , n19636 , n80 );
nor ( n19638 , n19635 , n19637 );
or ( n19639 , n2246 , n19638 );
nand ( n19640 , n19634 , n19639 );
not ( n19641 , n93 );
xor ( n19642 , n19641 , n9216 );
not ( n19643 , n19642 );
not ( n19644 , n8510 );
or ( n19645 , n19643 , n19644 );
or ( n19646 , n8510 , n19642 );
nand ( n19647 , n19645 , n19646 );
xnor ( n19648 , n19614 , n11076 );
and ( n19649 , n19647 , n19648 );
not ( n19650 , n19647 );
not ( n19651 , n19648 );
and ( n19652 , n19650 , n19651 );
nor ( n19653 , n19649 , n19652 );
or ( n19654 , n19653 , n1 );
and ( n19655 , n94 , n19641 );
not ( n19656 , n94 );
and ( n19657 , n19656 , n93 );
nor ( n19658 , n19655 , n19657 );
or ( n19659 , n2246 , n19658 );
nand ( n19660 , n19654 , n19659 );
xor ( n19661 , n9804 , n19305 );
not ( n19662 , n6155 );
not ( n19663 , n102 );
and ( n19664 , n19662 , n19663 );
and ( n19665 , n6271 , n102 );
nor ( n19666 , n19664 , n19665 );
buf ( n19667 , n14526 );
and ( n19668 , n19666 , n19667 );
not ( n19669 , n19666 );
not ( n19670 , n19667 );
and ( n19671 , n19669 , n19670 );
nor ( n19672 , n19668 , n19671 );
xnor ( n19673 , n19661 , n19672 );
or ( n19674 , n19673 , n1 );
not ( n19675 , n102 );
and ( n19676 , n222 , n19675 );
not ( n19677 , n222 );
and ( n19678 , n19677 , n102 );
nor ( n19679 , n19676 , n19678 );
or ( n19680 , n2246 , n19679 );
nand ( n19681 , n19674 , n19680 );
not ( n19682 , n19064 );
xor ( n19683 , n19682 , n12666 );
not ( n19684 , n223 );
xor ( n19685 , n19684 , n14526 );
and ( n19686 , n19685 , n9804 );
not ( n19687 , n19685 );
and ( n19688 , n19687 , n9805 );
nor ( n19689 , n19686 , n19688 );
xnor ( n19690 , n19683 , n19689 );
or ( n19691 , n19690 , n1 );
and ( n19692 , n224 , n19684 );
not ( n19693 , n224 );
and ( n19694 , n19693 , n223 );
nor ( n19695 , n19692 , n19694 );
or ( n19696 , n2246 , n19695 );
nand ( n19697 , n19691 , n19696 );
not ( n19698 , n18553 );
not ( n19699 , n225 );
and ( n19700 , n19698 , n19699 );
and ( n19701 , n18553 , n225 );
nor ( n19702 , n19700 , n19701 );
xor ( n19703 , n19702 , n19262 );
xor ( n19704 , n19703 , n18440 );
or ( n19705 , n19704 , n1 );
xnor ( n19706 , n225 , n226 );
or ( n19707 , n2246 , n19706 );
nand ( n19708 , n19705 , n19707 );
xor ( n19709 , n19358 , n19068 );
xor ( n19710 , n244 , n9804 );
xnor ( n19711 , n19710 , n15309 );
xnor ( n19712 , n19709 , n19711 );
or ( n19713 , n19712 , n1 );
xnor ( n19714 , n244 , n245 );
or ( n19715 , n2246 , n19714 );
nand ( n19716 , n19713 , n19715 );
xor ( n19717 , n19200 , n18237 );
xor ( n19718 , n252 , n16340 );
xnor ( n19719 , n19718 , n10336 );
xnor ( n19720 , n19717 , n19719 );
or ( n19721 , n19720 , n1 );
xnor ( n19722 , n252 , n253 );
or ( n19723 , n2246 , n19722 );
nand ( n19724 , n19721 , n19723 );
not ( n19725 , n18438 );
xor ( n19726 , n17800 , n19725 );
xor ( n19727 , n257 , n18553 );
xnor ( n19728 , n19727 , n2232 );
not ( n19729 , n19728 );
and ( n19730 , n19726 , n19729 );
not ( n19731 , n19726 );
and ( n19732 , n19731 , n19728 );
nor ( n19733 , n19730 , n19732 );
or ( n19734 , n19733 , n1 );
xnor ( n19735 , n256 , n257 );
or ( n19736 , n2246 , n19735 );
nand ( n19737 , n19734 , n19736 );
not ( n19738 , n18047 );
not ( n19739 , n17320 );
not ( n19740 , n3018 );
not ( n19741 , n19740 );
and ( n19742 , n19739 , n19741 );
and ( n19743 , n17320 , n3019 );
nor ( n19744 , n19742 , n19743 );
buf ( n19745 , n19744 );
not ( n19746 , n19745 );
or ( n19747 , n19738 , n19746 );
or ( n19748 , n19745 , n18047 );
nand ( n19749 , n19747 , n19748 );
nand ( n19750 , n19749 , n2246 );
buf ( n19751 , n19450 );
xor ( n19752 , n17401 , n19751 );
not ( n19753 , n272 );
not ( n19754 , n2512 );
and ( n19755 , n19753 , n19754 );
not ( n19756 , n2513 );
and ( n19757 , n19756 , n272 );
nor ( n19758 , n19755 , n19757 );
xnor ( n19759 , n19752 , n19758 );
or ( n19760 , n19750 , n19759 );
xnor ( n19761 , n272 , n273 );
or ( n19762 , n19761 , n2246 );
not ( n19763 , n19749 );
nand ( n19764 , n19759 , n19763 , n2246 );
nand ( n19765 , n19760 , n19762 , n19764 );
xor ( n19766 , n9995 , n18237 );
xor ( n19767 , n282 , n3430 );
xnor ( n19768 , n19767 , n16340 );
xnor ( n19769 , n19766 , n19768 );
or ( n19770 , n19769 , n1 );
xnor ( n19771 , n282 , n283 );
or ( n19772 , n2246 , n19771 );
nand ( n19773 , n19770 , n19772 );
not ( n19774 , n10760 );
not ( n19775 , n16963 );
or ( n19776 , n19774 , n19775 );
or ( n19777 , n10760 , n17626 );
nand ( n19778 , n19776 , n19777 );
not ( n19779 , n19778 );
not ( n19780 , n10905 );
not ( n19781 , n284 );
and ( n19782 , n19780 , n19781 );
and ( n19783 , n10898 , n284 );
nor ( n19784 , n19782 , n19783 );
not ( n19785 , n19784 );
or ( n19786 , n19779 , n19785 );
or ( n19787 , n19784 , n19778 );
nand ( n19788 , n19786 , n19787 );
and ( n19789 , n19788 , n18844 );
not ( n19790 , n19788 );
and ( n19791 , n19790 , n18446 );
nor ( n19792 , n19789 , n19791 );
or ( n19793 , n19792 , n1 );
xnor ( n19794 , n284 , n285 );
or ( n19795 , n2246 , n19794 );
nand ( n19796 , n19793 , n19795 );
xor ( n19797 , n19682 , n19305 );
not ( n19798 , n292 );
xor ( n19799 , n19798 , n4954 );
xor ( n19800 , n19799 , n19667 );
xnor ( n19801 , n19797 , n19800 );
or ( n19802 , n19801 , n1 );
and ( n19803 , n293 , n19798 );
not ( n19804 , n293 );
and ( n19805 , n19804 , n292 );
nor ( n19806 , n19803 , n19805 );
or ( n19807 , n2246 , n19806 );
nand ( n19808 , n19802 , n19807 );
xor ( n19809 , n12661 , n19068 );
not ( n19810 , n14526 );
not ( n19811 , n101 );
and ( n19812 , n19810 , n19811 );
not ( n19813 , n19810 );
and ( n19814 , n19813 , n101 );
nor ( n19815 , n19812 , n19814 );
and ( n19816 , n19815 , n15305 );
not ( n19817 , n19815 );
and ( n19818 , n19817 , n15309 );
nor ( n19819 , n19816 , n19818 );
xnor ( n19820 , n19809 , n19819 );
or ( n19821 , n19820 , n1 );
and ( n19822 , n296 , n19811 );
not ( n19823 , n296 );
and ( n19824 , n19823 , n101 );
nor ( n19825 , n19822 , n19824 );
or ( n19826 , n2246 , n19825 );
nand ( n19827 , n19821 , n19826 );
not ( n19828 , n15990 );
not ( n19829 , n15903 );
or ( n19830 , n19828 , n19829 );
or ( n19831 , n15990 , n15903 );
nand ( n19832 , n19830 , n19831 );
not ( n19833 , n19233 );
not ( n19834 , n15517 );
and ( n19835 , n19833 , n19834 );
and ( n19836 , n18241 , n15517 );
nor ( n19837 , n19835 , n19836 );
xor ( n19838 , n19832 , n19837 );
not ( n19839 , n17238 );
not ( n19840 , n15779 );
or ( n19841 , n19839 , n19840 );
or ( n19842 , n18854 , n15784 );
nand ( n19843 , n19841 , n19842 );
not ( n19844 , n19843 );
not ( n19845 , n19462 );
not ( n19846 , n303 );
not ( n19847 , n19846 );
and ( n19848 , n19845 , n19847 );
and ( n19849 , n19462 , n19846 );
nor ( n19850 , n19848 , n19849 );
not ( n19851 , n19850 );
or ( n19852 , n19844 , n19851 );
or ( n19853 , n19850 , n19843 );
nand ( n19854 , n19852 , n19853 );
xnor ( n19855 , n19838 , n19854 );
or ( n19856 , n19855 , n1 );
and ( n19857 , n304 , n19846 );
not ( n19858 , n304 );
and ( n19859 , n19858 , n303 );
nor ( n19860 , n19857 , n19859 );
or ( n19861 , n2246 , n19860 );
nand ( n19862 , n19856 , n19861 );
not ( n19863 , n2767 );
not ( n19864 , n19450 );
or ( n19865 , n19863 , n19864 );
nand ( n19866 , n19449 , n18054 );
nand ( n19867 , n19865 , n19866 );
xor ( n19868 , n19172 , n19867 );
xnor ( n19869 , n19868 , n15283 );
not ( n19870 , n14764 );
not ( n19871 , n309 );
or ( n19872 , n19870 , n19871 );
or ( n19873 , n14764 , n309 );
nand ( n19874 , n19872 , n19873 );
nand ( n19875 , n2246 , n19874 );
or ( n19876 , n19869 , n19875 );
nor ( n19877 , n19874 , n1 );
nand ( n19878 , n19869 , n19877 );
xor ( n19879 , n309 , n310 );
nand ( n19880 , n19879 , n1 );
nand ( n19881 , n19876 , n19878 , n19880 );
not ( n19882 , n11685 );
not ( n19883 , n13487 );
not ( n19884 , n10760 );
and ( n19885 , n19883 , n19884 );
and ( n19886 , n13487 , n10760 );
nor ( n19887 , n19885 , n19886 );
not ( n19888 , n19887 );
or ( n19889 , n19882 , n19888 );
or ( n19890 , n11685 , n19887 );
nand ( n19891 , n19889 , n19890 );
not ( n19892 , n10898 );
not ( n19893 , n311 );
and ( n19894 , n19892 , n19893 );
and ( n19895 , n10898 , n311 );
nor ( n19896 , n19894 , n19895 );
not ( n19897 , n19896 );
and ( n19898 , n19891 , n19897 );
not ( n19899 , n19891 );
and ( n19900 , n19899 , n19896 );
nor ( n19901 , n19898 , n19900 );
or ( n19902 , n19901 , n1 );
xnor ( n19903 , n311 , n312 );
or ( n19904 , n2246 , n19903 );
nand ( n19905 , n19902 , n19904 );
and ( n19906 , n17923 , n18862 );
not ( n19907 , n17923 );
and ( n19908 , n19907 , n18863 );
nor ( n19909 , n19906 , n19908 );
xor ( n19910 , n332 , n19756 );
and ( n19911 , n19909 , n19910 );
not ( n19912 , n19909 );
not ( n19913 , n19910 );
and ( n19914 , n19912 , n19913 );
nor ( n19915 , n19911 , n19914 );
or ( n19916 , n19915 , n1 );
xnor ( n19917 , n332 , n333 );
or ( n19918 , n2246 , n19917 );
nand ( n19919 , n19916 , n19918 );
not ( n19920 , n10769 );
not ( n19921 , n16969 );
or ( n19922 , n19920 , n19921 );
or ( n19923 , n16969 , n10769 );
nand ( n19924 , n19922 , n19923 );
xor ( n19925 , n336 , n2232 );
not ( n19926 , n19925 );
and ( n19927 , n19924 , n19926 );
not ( n19928 , n19924 );
and ( n19929 , n19928 , n19925 );
nor ( n19930 , n19927 , n19929 );
or ( n19931 , n19930 , n1 );
xnor ( n19932 , n336 , n337 );
or ( n19933 , n2246 , n19932 );
nand ( n19934 , n19931 , n19933 );
xor ( n19935 , n18862 , n19837 );
not ( n19936 , n15780 );
not ( n19937 , n344 );
and ( n19938 , n19936 , n19937 );
not ( n19939 , n15779 );
and ( n19940 , n19939 , n344 );
nor ( n19941 , n19938 , n19940 );
xnor ( n19942 , n17243 , n19941 );
xor ( n19943 , n19935 , n19942 );
or ( n19944 , n19943 , n1 );
xnor ( n19945 , n344 , n345 );
or ( n19946 , n2246 , n19945 );
nand ( n19947 , n19944 , n19946 );
buf ( n19948 , n18653 );
xor ( n19949 , n17800 , n19948 );
and ( n19950 , n11577 , n351 );
not ( n19951 , n11577 );
not ( n19952 , n351 );
and ( n19953 , n19951 , n19952 );
or ( n19954 , n19950 , n19953 );
buf ( n19955 , n18550 );
not ( n19956 , n19955 );
and ( n19957 , n19954 , n19956 );
not ( n19958 , n19954 );
and ( n19959 , n19958 , n19955 );
nor ( n19960 , n19957 , n19959 );
not ( n19961 , n19960 );
and ( n19962 , n19949 , n19961 );
not ( n19963 , n19949 );
and ( n19964 , n19963 , n19960 );
nor ( n19965 , n19962 , n19964 );
or ( n19966 , n19965 , n1 );
and ( n19967 , n352 , n19952 );
not ( n19968 , n352 );
and ( n19969 , n19968 , n351 );
nor ( n19970 , n19967 , n19969 );
or ( n19971 , n2246 , n19970 );
nand ( n19972 , n19966 , n19971 );
and ( n19973 , n17491 , n14893 );
not ( n19974 , n17491 );
and ( n19975 , n19974 , n14894 );
nor ( n19976 , n19973 , n19975 );
not ( n19977 , n18773 );
not ( n19978 , n19977 );
not ( n19979 , n19233 );
or ( n19980 , n19978 , n19979 );
or ( n19981 , n19233 , n19977 );
nand ( n19982 , n19980 , n19981 );
xor ( n19983 , n19976 , n19982 );
not ( n19984 , n19867 );
not ( n19985 , n371 );
and ( n19986 , n14759 , n19985 );
not ( n19987 , n14759 );
and ( n19988 , n19987 , n371 );
nor ( n19989 , n19986 , n19988 );
not ( n19990 , n19989 );
or ( n19991 , n19984 , n19990 );
or ( n19992 , n19989 , n19867 );
nand ( n19993 , n19991 , n19992 );
xnor ( n19994 , n19983 , n19993 );
or ( n19995 , n19994 , n1 );
and ( n19996 , n372 , n19985 );
not ( n19997 , n372 );
and ( n19998 , n19997 , n371 );
nor ( n19999 , n19996 , n19998 );
or ( n20000 , n2246 , n19999 );
nand ( n20001 , n19995 , n20000 );
xor ( n20002 , n5244 , n14624 );
xor ( n20003 , n369 , n12662 );
xnor ( n20004 , n20003 , n13224 );
xnor ( n20005 , n20002 , n20004 );
or ( n20006 , n20005 , n1 );
xnor ( n20007 , n369 , n370 );
or ( n20008 , n2246 , n20007 );
nand ( n20009 , n20006 , n20008 );
not ( n20010 , n3709 );
not ( n20011 , n16990 );
or ( n20012 , n20010 , n20011 );
nand ( n20013 , n3708 , n5889 );
nand ( n20014 , n20012 , n20013 );
not ( n20015 , n6185 );
nand ( n20016 , n20015 , n6267 );
not ( n20017 , n105 );
and ( n20018 , n20016 , n20017 );
not ( n20019 , n20016 );
and ( n20020 , n20019 , n105 );
nor ( n20021 , n20018 , n20020 );
and ( n20022 , n20014 , n20021 );
not ( n20023 , n20014 );
not ( n20024 , n20021 );
and ( n20025 , n20023 , n20024 );
nor ( n20026 , n20022 , n20025 );
and ( n20027 , n20026 , n9819 );
not ( n20028 , n20026 );
and ( n20029 , n20028 , n19079 );
nor ( n20030 , n20027 , n20029 );
or ( n20031 , n20030 , n1 );
and ( n20032 , n375 , n20017 );
not ( n20033 , n375 );
and ( n20034 , n20033 , n105 );
nor ( n20035 , n20032 , n20034 );
or ( n20036 , n2246 , n20035 );
nand ( n20037 , n20031 , n20036 );
not ( n20038 , n103 );
not ( n20039 , n16720 );
or ( n20040 , n20038 , n20039 );
not ( n20041 , n103 );
nand ( n20042 , n16719 , n20041 );
nand ( n20043 , n20040 , n20042 );
and ( n20044 , n20043 , n4653 );
not ( n20045 , n20043 );
not ( n20046 , n4653 );
and ( n20047 , n20045 , n20046 );
nor ( n20048 , n20044 , n20047 );
xnor ( n20049 , n4830 , n19298 );
not ( n20050 , n20049 );
and ( n20051 , n20048 , n20050 );
not ( n20052 , n20048 );
and ( n20053 , n20052 , n20049 );
nor ( n20054 , n20051 , n20053 );
or ( n20055 , n20054 , n1 );
and ( n20056 , n264 , n20041 );
not ( n20057 , n264 );
and ( n20058 , n20057 , n103 );
nor ( n20059 , n20056 , n20058 );
or ( n20060 , n2246 , n20059 );
nand ( n20061 , n20055 , n20060 );
xor ( n20062 , n19744 , n19982 );
and ( n20063 , n19449 , n18042 );
not ( n20064 , n19449 );
and ( n20065 , n20064 , n18041 );
nor ( n20066 , n20063 , n20065 );
and ( n20067 , n14759 , n276 );
not ( n20068 , n14759 );
not ( n20069 , n276 );
and ( n20070 , n20068 , n20069 );
nor ( n20071 , n20067 , n20070 );
xor ( n20072 , n20066 , n20071 );
xnor ( n20073 , n20062 , n20072 );
or ( n20074 , n20073 , n1 );
and ( n20075 , n277 , n20069 );
not ( n20076 , n277 );
and ( n20077 , n20076 , n276 );
nor ( n20078 , n20075 , n20077 );
or ( n20079 , n2246 , n20078 );
nand ( n20080 , n20074 , n20079 );
xor ( n20081 , n19548 , n18106 );
xor ( n20082 , n40 , n9118 );
xnor ( n20083 , n20082 , n19551 );
xnor ( n20084 , n20081 , n20083 );
or ( n20085 , n20084 , n1 );
xnor ( n20086 , n40 , n47 );
or ( n20087 , n2246 , n20086 );
nand ( n20088 , n20085 , n20087 );
nand ( n20089 , n19648 , n2246 );
not ( n20090 , n77 );
xor ( n20091 , n9352 , n20090 );
xnor ( n20092 , n20091 , n6963 );
or ( n20093 , n20089 , n20092 );
nand ( n20094 , n20092 , n19651 , n2246 );
and ( n20095 , n88 , n77 );
not ( n20096 , n88 );
and ( n20097 , n20096 , n20090 );
nor ( n20098 , n20095 , n20097 );
nand ( n20099 , n20098 , n1 );
nand ( n20100 , n20093 , n20094 , n20099 );
xor ( n20101 , n19948 , n12124 );
xor ( n20102 , n110 , n18435 );
xor ( n20103 , n20102 , n18553 );
xnor ( n20104 , n20101 , n20103 );
or ( n20105 , n20104 , n1 );
xnor ( n20106 , n110 , n219 );
or ( n20107 , n2246 , n20106 );
nand ( n20108 , n20105 , n20107 );
not ( n20109 , n18773 );
not ( n20110 , n17321 );
or ( n20111 , n20109 , n20110 );
nand ( n20112 , n19977 , n17320 );
nand ( n20113 , n20111 , n20112 );
xor ( n20114 , n18854 , n20113 );
xor ( n20115 , n246 , n17401 );
xnor ( n20116 , n20115 , n15784 );
xnor ( n20117 , n20114 , n20116 );
or ( n20118 , n20117 , n1 );
xnor ( n20119 , n246 , n247 );
or ( n20120 , n2246 , n20119 );
nand ( n20121 , n20118 , n20120 );
xor ( n20122 , n15990 , n20113 );
xor ( n20123 , n248 , n19939 );
xor ( n20124 , n20123 , n17492 );
xnor ( n20125 , n20122 , n20124 );
or ( n20126 , n20125 , n1 );
xnor ( n20127 , n248 , n249 );
or ( n20128 , n2246 , n20127 );
nand ( n20129 , n20126 , n20128 );
buf ( n20130 , n4211 );
not ( n20131 , n20130 );
not ( n20132 , n19298 );
or ( n20133 , n20131 , n20132 );
or ( n20134 , n19298 , n20130 );
nand ( n20135 , n20133 , n20134 );
xor ( n20136 , n265 , n16637 );
xnor ( n20137 , n20136 , n4653 );
and ( n20138 , n20135 , n20137 );
not ( n20139 , n20135 );
not ( n20140 , n20137 );
and ( n20141 , n20139 , n20140 );
nor ( n20142 , n20138 , n20141 );
or ( n20143 , n20142 , n1 );
xnor ( n20144 , n265 , n266 );
or ( n20145 , n2246 , n20144 );
nand ( n20146 , n20143 , n20145 );
xor ( n20147 , n330 , n20016 );
and ( n20148 , n20147 , n4373 );
not ( n20149 , n20147 );
and ( n20150 , n20149 , n3962 );
nor ( n20151 , n20148 , n20150 );
not ( n20152 , n19305 );
and ( n20153 , n20151 , n20152 );
not ( n20154 , n20151 );
and ( n20155 , n20154 , n19305 );
nor ( n20156 , n20153 , n20155 );
or ( n20157 , n20156 , n1 );
xnor ( n20158 , n330 , n331 );
or ( n20159 , n2246 , n20158 );
nand ( n20160 , n20157 , n20159 );
xor ( n20161 , n365 , n16719 );
xnor ( n20162 , n20161 , n16843 );
and ( n20163 , n20162 , n6019 );
not ( n20164 , n20162 );
and ( n20165 , n20164 , n6022 );
nor ( n20166 , n20163 , n20165 );
or ( n20167 , n20166 , n1 );
xnor ( n20168 , n365 , n366 );
or ( n20169 , n2246 , n20168 );
nand ( n20170 , n20167 , n20169 );
xor ( n20171 , n9995 , n19225 );
xor ( n20172 , n363 , n16221 );
xnor ( n20173 , n20172 , n16340 );
xnor ( n20174 , n20171 , n20173 );
or ( n20175 , n20174 , n1 );
xnor ( n20176 , n363 , n364 );
or ( n20177 , n2246 , n20176 );
nand ( n20178 , n20175 , n20177 );
xor ( n20179 , n18973 , n18658 );
xor ( n20180 , n373 , n18435 );
xnor ( n20181 , n20180 , n12244 );
xnor ( n20182 , n20179 , n20181 );
or ( n20183 , n20182 , n1 );
xnor ( n20184 , n373 , n374 );
or ( n20185 , n2246 , n20184 );
nand ( n20186 , n20183 , n20185 );
xor ( n20187 , n1271 , n19262 );
xor ( n20188 , n320 , n12122 );
xnor ( n20189 , n20188 , n13359 );
xnor ( n20190 , n20187 , n20189 );
or ( n20191 , n20190 , n1 );
xnor ( n20192 , n320 , n321 );
or ( n20193 , n2246 , n20192 );
nand ( n20194 , n20191 , n20193 );
not ( n20195 , n17757 );
xor ( n20196 , n20195 , n11156 );
xor ( n20197 , n234 , n16637 );
xnor ( n20198 , n20197 , n16719 );
xnor ( n20199 , n20196 , n20198 );
or ( n20200 , n20199 , n1 );
xnor ( n20201 , n234 , n235 );
or ( n20202 , n2246 , n20201 );
nand ( n20203 , n20200 , n20202 );
xnor ( n20204 , n297 , n15661 );
xor ( n20205 , n15908 , n20204 );
not ( n20206 , n18242 );
not ( n20207 , n15424 );
and ( n20208 , n20206 , n20207 );
and ( n20209 , n18242 , n15424 );
nor ( n20210 , n20208 , n20209 );
xnor ( n20211 , n20205 , n20210 );
or ( n20212 , n20211 , n1 );
xnor ( n20213 , n297 , n298 );
or ( n20214 , n2246 , n20213 );
nand ( n20215 , n20212 , n20214 );
xor ( n20216 , n109 , n18 );
not ( n20217 , n19811 );
nor ( n20218 , n100 , n101 );
not ( n20219 , n20218 );
not ( n20220 , n20219 );
not ( n20221 , n102 );
nand ( n20222 , n20221 , n101 );
nor ( n20223 , n20222 , n15298 );
not ( n20224 , n20223 );
not ( n20225 , n20224 );
or ( n20226 , n20220 , n20225 );
not ( n20227 , n99 );
nor ( n20228 , n20227 , n98 );
nand ( n20229 , n20226 , n20228 );
nor ( n20230 , n16723 , n99 );
nand ( n20231 , n20230 , n15298 );
nor ( n20232 , n101 , n102 );
or ( n20233 , n20231 , n20232 );
nand ( n20234 , n20229 , n20233 );
nand ( n20235 , n20234 , n20041 );
not ( n20236 , n20235 );
nor ( n20237 , n100 , n102 );
nand ( n20238 , n20237 , n16723 );
or ( n20239 , n20236 , n20238 );
and ( n20240 , n11185 , n103 );
nand ( n20241 , n20240 , n19675 , n98 );
and ( n20242 , n99 , n98 , n102 );
not ( n20243 , n20242 );
nand ( n20244 , n20241 , n20243 );
and ( n20245 , n20244 , n11125 );
nor ( n20246 , n98 , n99 );
and ( n20247 , n20246 , n19675 );
and ( n20248 , n20237 , n99 );
nor ( n20249 , n20247 , n20248 );
nand ( n20250 , n100 , n102 );
not ( n20251 , n20250 );
nand ( n20252 , n20251 , n20230 );
and ( n20253 , n20249 , n20252 );
nand ( n20254 , n103 , n104 );
nor ( n20255 , n20253 , n20254 );
nor ( n20256 , n20245 , n20255 );
nand ( n20257 , n20239 , n20256 );
not ( n20258 , n20257 );
or ( n20259 , n20217 , n20258 );
nand ( n20260 , n20232 , n100 );
nor ( n20261 , n20260 , n16723 );
and ( n20262 , n20261 , n99 );
not ( n20263 , n100 );
nand ( n20264 , n20263 , n99 );
nand ( n20265 , n20219 , n20264 );
and ( n20266 , n20265 , n16723 , n20041 );
nand ( n20267 , n20252 , n104 );
nor ( n20268 , n20262 , n20266 , n20267 );
not ( n20269 , n20268 );
not ( n20270 , n16723 );
nand ( n20271 , n101 , n102 );
nor ( n20272 , n20271 , n100 );
not ( n20273 , n20272 );
or ( n20274 , n20270 , n20273 );
nand ( n20275 , n20251 , n19811 );
nand ( n20276 , n20274 , n20275 );
and ( n20277 , n20276 , n20240 );
not ( n20278 , n20222 );
nand ( n20279 , n20278 , n99 );
not ( n20280 , n20279 );
and ( n20281 , n20280 , n103 );
nor ( n20282 , n20277 , n20281 );
not ( n20283 , n20282 );
or ( n20284 , n20269 , n20283 );
nand ( n20285 , n20041 , n98 );
not ( n20286 , n20285 );
and ( n20287 , n20237 , n20286 );
not ( n20288 , n20275 );
nor ( n20289 , n20287 , n20288 );
or ( n20290 , n20289 , n11185 );
not ( n20291 , n11185 );
not ( n20292 , n20272 );
or ( n20293 , n20291 , n20292 );
not ( n20294 , n20041 );
not ( n20295 , n20260 );
or ( n20296 , n20294 , n20295 );
nand ( n20297 , n20296 , n20285 );
nand ( n20298 , n20293 , n20297 );
nand ( n20299 , n20237 , n101 );
nand ( n20300 , n20299 , n20243 , n103 );
nand ( n20301 , n20298 , n20300 );
nand ( n20302 , n20290 , n20301 , n11125 );
nand ( n20303 , n20284 , n20302 );
nand ( n20304 , n20218 , n102 );
not ( n20305 , n20304 );
not ( n20306 , n20279 );
or ( n20307 , n20305 , n20306 );
nand ( n20308 , n20307 , n98 );
and ( n20309 , n20228 , n20251 , n101 );
nor ( n20310 , n99 , n100 );
nand ( n20311 , n20232 , n20310 );
not ( n20312 , n20311 );
nor ( n20313 , n20309 , n20312 );
nand ( n20314 , n20308 , n20313 );
nand ( n20315 , n20314 , n103 );
not ( n20316 , n19811 );
not ( n20317 , n20228 );
or ( n20318 , n20316 , n20317 );
or ( n20319 , n99 , n20222 );
nand ( n20320 , n20318 , n20319 );
and ( n20321 , n20320 , n20041 , n100 );
nor ( n20322 , n20321 , n20017 );
nand ( n20323 , n20303 , n20315 , n20322 );
or ( n20324 , n20311 , n103 );
nor ( n20325 , n15298 , n16723 );
nand ( n20326 , n20280 , n20325 );
not ( n20327 , n20238 );
nand ( n20328 , n20327 , n20240 );
nand ( n20329 , n20324 , n20326 , n20328 );
nand ( n20330 , n20329 , n104 );
not ( n20331 , n20272 );
or ( n20332 , n20331 , n20041 );
or ( n20333 , n20250 , n20254 );
nand ( n20334 , n20332 , n20333 );
and ( n20335 , n20334 , n20228 );
not ( n20336 , n20246 );
nor ( n20337 , n20336 , n20219 , n20041 );
nor ( n20338 , n20335 , n20337 , n105 );
not ( n20339 , n20285 );
nand ( n20340 , n20339 , n20272 );
nand ( n20341 , n20330 , n20235 , n20338 , n20340 );
nand ( n20342 , n20323 , n20341 );
nand ( n20343 , n20259 , n20342 );
and ( n20344 , n20261 , n103 );
and ( n20345 , n20242 , n20041 );
nor ( n20346 , n20344 , n20345 );
and ( n20347 , n20228 , n20272 );
and ( n20348 , n20223 , n11185 );
nor ( n20349 , n20347 , n20348 );
nand ( n20350 , n20346 , n20349 );
nand ( n20351 , n20246 , n19811 );
and ( n20352 , n20231 , n20351 );
nor ( n20353 , n20352 , n19675 );
or ( n20354 , n20350 , n20353 );
nand ( n20355 , n20354 , n20017 );
not ( n20356 , n20355 );
not ( n20357 , n102 );
not ( n20358 , n20240 );
or ( n20359 , n20357 , n20358 );
nand ( n20360 , n20359 , n20336 );
nand ( n20361 , n20360 , n100 , n101 );
not ( n20362 , n20361 );
or ( n20363 , n20356 , n20362 );
nand ( n20364 , n20363 , n11125 );
or ( n20365 , n20242 , n11125 );
nand ( n20366 , n20365 , n20041 );
not ( n20367 , n20366 );
not ( n20368 , n20315 );
or ( n20369 , n20367 , n20368 );
or ( n20370 , n20275 , n20246 );
or ( n20371 , n20279 , n100 );
nand ( n20372 , n20370 , n20371 );
nand ( n20373 , n20369 , n20372 );
nand ( n20374 , n20268 , n20261 , n20041 );
nand ( n20375 , n20364 , n20373 , n20374 );
nor ( n20376 , n20343 , n20375 );
xnor ( n20377 , n20216 , n20376 );
not ( n20378 , n20377 );
and ( n20379 , n110 , n20378 );
not ( n20380 , n110 );
and ( n20381 , n20380 , n20377 );
nor ( n20382 , n20379 , n20381 );
or ( n20383 , n20382 , n106 );
not ( n20384 , n106 );
not ( n20385 , n111 );
or ( n20386 , n20384 , n20385 );
nand ( n20387 , n20383 , n20386 );
xor ( n20388 , n223 , n110 );
xnor ( n20389 , n20388 , n20377 );
or ( n20390 , n20389 , n106 );
not ( n20391 , n227 );
or ( n20392 , n20384 , n20391 );
nand ( n20393 , n20390 , n20392 );
and ( n20394 , n45 , n7485 );
not ( n20395 , n45 );
and ( n20396 , n20395 , n11088 );
nor ( n20397 , n20394 , n20396 );
or ( n20398 , n20378 , n106 );
not ( n20399 , n108 );
not ( n20400 , n106 );
or ( n20401 , n20399 , n20400 );
nand ( n20402 , n20398 , n20401 );
not ( n20403 , n107 );
not ( n20404 , n106 );
or ( n20405 , n20403 , n20404 );
not ( n20406 , n20376 );
not ( n20407 , n18 );
and ( n20408 , n20406 , n20407 );
and ( n20409 , n20376 , n18 );
nor ( n20410 , n20408 , n20409 );
or ( n20411 , n20410 , n106 );
nand ( n20412 , n20405 , n20411 );
and ( n20413 , n65 , n14421 );
not ( n20414 , n65 );
not ( n20415 , n14421 );
and ( n20416 , n20414 , n20415 );
nor ( n20417 , n20413 , n20416 );
not ( n20418 , n14258 );
not ( n20419 , n14305 );
or ( n20420 , n20418 , n20419 );
or ( n20421 , n14305 , n14258 );
nand ( n20422 , n20420 , n20421 );
and ( n20423 , n58 , n14035 );
not ( n20424 , n58 );
and ( n20425 , n20424 , n14038 );
nor ( n20426 , n20423 , n20425 );
and ( n20427 , n48 , n19516 );
not ( n20428 , n48 );
and ( n20429 , n20428 , n19517 );
nor ( n20430 , n20427 , n20429 );
not ( n20431 , n37 );
not ( n20432 , n19492 );
or ( n20433 , n20431 , n20432 );
or ( n20434 , n37 , n19492 );
nand ( n20435 , n20433 , n20434 );
not ( n20436 , n7225 );
and ( n20437 , n40 , n20436 );
not ( n20438 , n40 );
and ( n20439 , n20438 , n7225 );
nor ( n20440 , n20437 , n20439 );
and ( n20441 , n71 , n8633 );
not ( n20442 , n71 );
and ( n20443 , n20442 , n19571 );
nor ( n20444 , n20441 , n20443 );
not ( n20445 , n84 );
not ( n20446 , n8002 );
or ( n20447 , n20445 , n20446 );
or ( n20448 , n84 , n8002 );
nand ( n20449 , n20447 , n20448 );
not ( n20450 , n78 );
not ( n20451 , n12436 );
or ( n20452 , n20450 , n20451 );
or ( n20453 , n78 , n12436 );
nand ( n20454 , n20452 , n20453 );
not ( n20455 , n11076 );
not ( n20456 , n80 );
or ( n20457 , n20455 , n20456 );
or ( n20458 , n80 , n11076 );
nand ( n20459 , n20457 , n20458 );
not ( n20460 , n8918 );
not ( n20461 , n55 );
or ( n20462 , n20460 , n20461 );
or ( n20463 , n55 , n8918 );
nand ( n20464 , n20462 , n20463 );
and ( n20465 , n63 , n19560 );
not ( n20466 , n63 );
not ( n20467 , n19560 );
and ( n20468 , n20466 , n20467 );
nor ( n20469 , n20465 , n20468 );
not ( n20470 , n95 );
not ( n20471 , n13946 );
or ( n20472 , n20470 , n20471 );
or ( n20473 , n95 , n13946 );
nand ( n20474 , n20472 , n20473 );
not ( n20475 , n86 );
not ( n20476 , n7668 );
or ( n20477 , n20475 , n20476 );
or ( n20478 , n86 , n7668 );
nand ( n20479 , n20477 , n20478 );
not ( n20480 , n59 );
not ( n20481 , n14134 );
or ( n20482 , n20480 , n20481 );
or ( n20483 , n59 , n14134 );
nand ( n20484 , n20482 , n20483 );
not ( n20485 , n93 );
not ( n20486 , n9352 );
or ( n20487 , n20485 , n20486 );
or ( n20488 , n93 , n9352 );
nand ( n20489 , n20487 , n20488 );
not ( n20490 , n19578 );
and ( n20491 , n81 , n20490 );
not ( n20492 , n81 );
and ( n20493 , n20492 , n19578 );
nor ( n20494 , n20491 , n20493 );
and ( n20495 , n8897 , n73 );
not ( n20496 , n8897 );
and ( n20497 , n20496 , n9241 );
nor ( n20498 , n20495 , n20497 );
not ( n20499 , n11077 );
not ( n20500 , n69 );
or ( n20501 , n20499 , n20500 );
or ( n20502 , n69 , n11077 );
nand ( n20503 , n20501 , n20502 );
not ( n20504 , n51 );
not ( n20505 , n13731 );
or ( n20506 , n20504 , n20505 );
or ( n20507 , n51 , n13731 );
nand ( n20508 , n20506 , n20507 );
not ( n20509 , n14291 );
not ( n20510 , n8264 );
or ( n20511 , n20509 , n20510 );
or ( n20512 , n8264 , n14291 );
nand ( n20513 , n20511 , n20512 );
not ( n20514 , n61 );
not ( n20515 , n14414 );
or ( n20516 , n20514 , n20515 );
or ( n20517 , n14414 , n61 );
nand ( n20518 , n20516 , n20517 );
and ( n20519 , n75 , n8757 );
not ( n20520 , n75 );
and ( n20521 , n20520 , n8758 );
nor ( n20522 , n20519 , n20521 );
and ( n20523 , n18 , n9016 );
not ( n20524 , n18 );
and ( n20525 , n20524 , n9017 );
nor ( n20526 , n20523 , n20525 );
not ( n20527 , n49 );
not ( n20528 , n19551 );
or ( n20529 , n20527 , n20528 );
or ( n20530 , n49 , n19551 );
nand ( n20531 , n20529 , n20530 );
and ( n20532 , n20400 , n97 );
and ( n20533 , n106 , n443 );
nor ( n20534 , n20532 , n20533 );
not ( n20535 , n20534 );
and ( n20536 , n20400 , n216 );
and ( n20537 , n106 , n407 );
nor ( n20538 , n20536 , n20537 );
not ( n20539 , n20538 );
and ( n20540 , n20400 , n64 );
and ( n20541 , n106 , n414 );
nor ( n20542 , n20540 , n20541 );
not ( n20543 , n20542 );
and ( n20544 , n20400 , n310 );
and ( n20545 , n106 , n409 );
nor ( n20546 , n20544 , n20545 );
not ( n20547 , n20546 );
and ( n20548 , n20400 , n374 );
and ( n20549 , n106 , n396 );
nor ( n20550 , n20548 , n20549 );
not ( n20551 , n20550 );
and ( n20552 , n20400 , n379 );
and ( n20553 , n106 , n436 );
nor ( n20554 , n20552 , n20553 );
not ( n20555 , n20554 );
and ( n20556 , n20400 , n341 );
and ( n20557 , n106 , n404 );
nor ( n20558 , n20556 , n20557 );
not ( n20559 , n20558 );
and ( n20560 , n20400 , n88 );
and ( n20561 , n106 , n449 );
nor ( n20562 , n20560 , n20561 );
not ( n20563 , n20562 );
and ( n20564 , n20400 , n47 );
and ( n20565 , n106 , n410 );
nor ( n20566 , n20564 , n20565 );
not ( n20567 , n20566 );
and ( n20568 , n20384 , n50 );
and ( n20569 , n106 , n429 );
nor ( n20570 , n20568 , n20569 );
not ( n20571 , n20570 );
and ( n20572 , n20384 , n35 );
and ( n20573 , n106 , n348 );
nor ( n20574 , n20572 , n20573 );
not ( n20575 , n20574 );
and ( n20576 , n20384 , n226 );
and ( n20577 , n106 , n406 );
nor ( n20578 , n20576 , n20577 );
not ( n20579 , n20578 );
and ( n20580 , n20400 , n44 );
and ( n20581 , n106 , n411 );
nor ( n20582 , n20580 , n20581 );
not ( n20583 , n20582 );
and ( n20584 , n20400 , n275 );
and ( n20585 , n106 , n430 );
nor ( n20586 , n20584 , n20585 );
not ( n20587 , n20586 );
and ( n20588 , n20384 , n372 );
and ( n20589 , n106 , n397 );
nor ( n20590 , n20588 , n20589 );
not ( n20591 , n20590 );
and ( n20592 , n20384 , n391 );
and ( n20593 , n106 , n431 );
nor ( n20594 , n20592 , n20593 );
not ( n20595 , n20594 );
and ( n20596 , n20384 , n52 );
and ( n20597 , n106 , n402 );
nor ( n20598 , n20596 , n20597 );
not ( n20599 , n20598 );
and ( n20600 , n20400 , n263 );
and ( n20601 , n106 , n413 );
nor ( n20602 , n20600 , n20601 );
not ( n20603 , n20602 );
and ( n20604 , n20400 , n289 );
and ( n20605 , n106 , n442 );
nor ( n20606 , n20604 , n20605 );
not ( n20607 , n20606 );
and ( n20608 , n20384 , n233 );
and ( n20609 , n106 , n441 );
nor ( n20610 , n20608 , n20609 );
not ( n20611 , n20610 );
and ( n20612 , n20400 , n62 );
and ( n20613 , n106 , n428 );
nor ( n20614 , n20612 , n20613 );
not ( n20615 , n20614 );
and ( n20616 , n20400 , n57 );
and ( n20617 , n106 , n403 );
nor ( n20618 , n20616 , n20617 );
not ( n20619 , n20618 );
and ( n20620 , n20400 , n89 );
and ( n20621 , n106 , n415 );
nor ( n20622 , n20620 , n20621 );
not ( n20623 , n20622 );
and ( n20624 , n20384 , n145 );
and ( n20625 , n106 , n417 );
nor ( n20626 , n20624 , n20625 );
not ( n20627 , n20626 );
and ( n20628 , n20384 , n266 );
and ( n20629 , n106 , n432 );
nor ( n20630 , n20628 , n20629 );
not ( n20631 , n20630 );
and ( n20632 , n20384 , n302 );
and ( n20633 , n106 , n437 );
nor ( n20634 , n20632 , n20633 );
not ( n20635 , n20634 );
and ( n20636 , n20384 , n337 );
and ( n20637 , n106 , n438 );
nor ( n20638 , n20636 , n20637 );
not ( n20639 , n20638 );
and ( n20640 , n20384 , n279 );
and ( n20641 , n106 , n423 );
nor ( n20642 , n20640 , n20641 );
not ( n20643 , n20642 );
and ( n20644 , n20384 , n325 );
and ( n20645 , n106 , n440 );
nor ( n20646 , n20644 , n20645 );
not ( n20647 , n20646 );
and ( n20648 , n20384 , n360 );
and ( n20649 , n106 , n400 );
nor ( n20650 , n20648 , n20649 );
not ( n20651 , n20650 );
and ( n20652 , n20400 , n323 );
and ( n20653 , n106 , n419 );
nor ( n20654 , n20652 , n20653 );
not ( n20655 , n20654 );
and ( n20656 , n20400 , n92 );
and ( n20657 , n106 , n416 );
nor ( n20658 , n20656 , n20657 );
not ( n20659 , n20658 );
and ( n20660 , n20384 , n224 );
and ( n20661 , n106 , n398 );
nor ( n20662 , n20660 , n20661 );
not ( n20663 , n20662 );
and ( n20664 , n20400 , n281 );
and ( n20665 , n106 , n424 );
nor ( n20666 , n20664 , n20665 );
not ( n20667 , n20666 );
and ( n20668 , n20400 , n247 );
and ( n20669 , n106 , n447 );
nor ( n20670 , n20668 , n20669 );
not ( n20671 , n20670 );
and ( n20672 , n20400 , n335 );
and ( n20673 , n106 , n426 );
nor ( n20674 , n20672 , n20673 );
not ( n20675 , n20674 );
and ( n20676 , n20384 , n76 );
and ( n20677 , n106 , n408 );
nor ( n20678 , n20676 , n20677 );
not ( n20679 , n20678 );
and ( n20680 , n20400 , n329 );
and ( n20681 , n106 , n446 );
nor ( n20682 , n20680 , n20681 );
not ( n20683 , n20682 );
and ( n20684 , n20400 , n231 );
and ( n20685 , n106 , n395 );
nor ( n20686 , n20684 , n20685 );
not ( n20687 , n20686 );
and ( n20688 , n20384 , n345 );
and ( n20689 , n106 , n394 );
nor ( n20690 , n20688 , n20689 );
not ( n20691 , n20690 );
and ( n20692 , n20384 , n222 );
and ( n20693 , n106 , n444 );
nor ( n20694 , n20692 , n20693 );
not ( n20695 , n20694 );
and ( n20696 , n20400 , n54 );
and ( n20697 , n106 , n433 );
nor ( n20698 , n20696 , n20697 );
not ( n20699 , n20698 );
and ( n20700 , n20384 , n268 );
and ( n20701 , n106 , n450 );
nor ( n20702 , n20700 , n20701 );
not ( n20703 , n20702 );
and ( n20704 , n20384 , n370 );
and ( n20705 , n106 , n399 );
nor ( n20706 , n20704 , n20705 );
not ( n20707 , n20706 );
and ( n20708 , n20400 , n70 );
and ( n20709 , n106 , n412 );
nor ( n20710 , n20708 , n20709 );
not ( n20711 , n20710 );
and ( n20712 , n20384 , n356 );
and ( n20713 , n106 , n422 );
nor ( n20714 , n20712 , n20713 );
not ( n20715 , n20714 );
and ( n20716 , n20384 , n347 );
and ( n20717 , n106 , n418 );
nor ( n20718 , n20716 , n20717 );
not ( n20719 , n20718 );
and ( n20720 , n20384 , n285 );
and ( n20721 , n106 , n445 );
nor ( n20722 , n20720 , n20721 );
not ( n20723 , n20722 );
and ( n20724 , n20384 , n362 );
and ( n20725 , n106 , n448 );
nor ( n20726 , n20724 , n20725 );
not ( n20727 , n20726 );
and ( n20728 , n20400 , n312 );
and ( n20729 , n106 , n405 );
nor ( n20730 , n20728 , n20729 );
not ( n20731 , n20730 );
and ( n20732 , n20384 , n237 );
and ( n20733 , n106 , n393 );
nor ( n20734 , n20732 , n20733 );
not ( n20735 , n20734 );
and ( n20736 , n20400 , n259 );
and ( n20737 , n106 , n435 );
nor ( n20738 , n20736 , n20737 );
not ( n20739 , n20738 );
and ( n20740 , n20384 , n377 );
and ( n20741 , n106 , n427 );
nor ( n20742 , n20740 , n20741 );
not ( n20743 , n20742 );
and ( n20744 , n20400 , n91 );
and ( n20745 , n106 , n425 );
nor ( n20746 , n20744 , n20745 );
not ( n20747 , n20746 );
xnor ( n20748 , n401 , n434 );
nor ( n20749 , n20748 , n106 );
and ( n20750 , n20384 , n60 );
and ( n20751 , n106 , n420 );
nor ( n20752 , n20750 , n20751 );
not ( n20753 , n20752 );
and ( n20754 , n20384 , n87 );
and ( n20755 , n106 , n421 );
nor ( n20756 , n20754 , n20755 );
not ( n20757 , n20756 );
nor ( n20758 , n106 , n401 );
nand ( n20759 , n401 , n434 );
and ( n20760 , n19614 , n18141 );
not ( n20761 , n19614 );
and ( n20762 , n20761 , n90 );
nor ( n20763 , n20760 , n20762 );
xor ( n20764 , n43 , n8268 );
xor ( n20765 , n39 , n6554 );
xnor ( n20766 , n41 , n9216 );
xor ( n20767 , n20759 , n439 );
nor ( n20768 , n20767 , n106 );
and ( n20769 , n19548 , n16436 );
not ( n20770 , n19548 );
and ( n20771 , n20770 , n53 );
nor ( n20772 , n20769 , n20771 );
and ( n20773 , n19612 , n20090 );
not ( n20774 , n19612 );
and ( n20775 , n20774 , n77 );
nor ( n20776 , n20773 , n20775 );
endmodule

