//NOTE: no-implementation module stub

module Delaya (
    input wire RSack,
    output reg delRSack
);

endmodule
