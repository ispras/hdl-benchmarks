// IWLS benchmark module "i4" printed on Wed May 29 16:38:48 2002
module i4(\V56(0) , \V28(0) , \V56(1) , \V28(1) , \V56(2) , \V28(2) , \V56(6) , \V28(6) , \V56(10) , \V28(10) , \V56(14) , \V28(14) , \V56(18) , \V28(18) , \V56(22) , \V28(22) , \V56(26) , \V28(26) , \V120(2) , \V88(2) , \V120(6) , \V88(6) , \V120(10) , \V88(10) , \V120(14) , \V88(14) , \V120(18) , \V88(18) , \V120(22) , \V88(22) , \V120(26) , \V88(26) , \V120(30) , \V88(30) , \V132(2) , \V126(2) , \V144(0) , \V28(3) , \V56(3) , \V144(1) , \V56(4) , \V28(4) , \V144(2) , \V28(5) , \V56(5) , \V144(4) , \V28(7) , \V56(7) , \V144(5) , \V56(8) , \V28(8) , \V144(6) , \V28(9) , \V56(9) , \V144(8) , \V28(11) , \V56(11) , \V144(9) , \V56(12) , \V28(12) , \V144(10) , \V28(13) , \V56(13) , \V144(12) , \V28(15) , \V56(15) , \V144(13) , \V56(16) , \V28(16) , \V144(14) , \V28(17) , \V56(17) , \V156(0) , \V28(19) , \V56(19) , \V156(1) , \V56(20) , \V28(20) , \V156(2) , \V28(21) , \V56(21) , \V156(4) , \V28(23) , \V56(23) , \V156(5) , \V56(24) , \V28(24) , \V156(6) , \V28(25) , \V56(25) , \V156(8) , \V28(27) , \V56(27) , \V156(9) , \V120(0) , \V88(0) , \V156(10) , \V88(1) , \V120(1) , \V156(12) , \V88(3) , \V120(3) , \V156(13) , \V120(4) , \V88(4) , \V156(14) , \V88(5) , \V120(5) , \V168(0) , \V88(7) , \V120(7) , \V168(1) , \V120(8) , \V88(8) , \V168(2) , \V88(9) , \V120(9) , \V168(4) , \V88(11) , \V120(11) , \V168(5) , \V120(12) , \V88(12) , \V168(6) , \V88(13) , \V120(13) , \V168(8) , \V88(15) , \V120(15) , \V168(9) , \V120(16) , \V88(16) , \V168(10) , \V88(17) , \V120(17) , \V168(12) , \V88(19) , \V120(19) , \V168(13) , \V120(20) , \V88(20) , \V168(14) , \V88(21) , \V120(21) , \V180(0) , \V88(23) , \V120(23) , \V180(1) , \V120(24) , \V88(24) , \V180(2) , \V88(25) , \V120(25) , \V180(4) , \V88(27) , \V120(27) , \V180(5) , \V120(28) , \V88(28) , \V180(6) , \V88(29) , \V120(29) , \V180(8) , \V88(31) , \V120(31) , \V180(9) , \V132(0) , \V126(0) , \V180(10) , \V126(1) , \V132(1) , \V180(12) , \V126(3) , \V132(3) , \V180(13) , \V132(4) , \V126(4) , \V180(14) , \V126(5) , \V132(5) , \V183(0) , \V183(1) , \V183(2) , \V186(0) , \V186(1) , \V186(2) , \V189(0) , \V189(1) , \V189(2) , \V192(0) , \V192(1) , \V192(2) , \V194(0) , \V194(1) , \V198(0) , \V198(1) , \V198(2) , \V198(3) );
input
  \V186(2) ,
  \V88(11) ,
  \V88(10) ,
  \V186(1) ,
  \V144(10) ,
  \V186(0) ,
  \V144(13) ,
  \V88(17) ,
  \V144(12) ,
  \V88(16) ,
  \V88(19) ,
  \V144(14) ,
  \V180(10) ,
  \V88(18) ,
  \V180(13) ,
  \V88(23) ,
  \V126(3) ,
  \V180(12) ,
  \V56(0) ,
  \V88(22) ,
  \V126(2) ,
  \V56(13) ,
  \V56(1) ,
  \V88(25) ,
  \V126(5) ,
  \V56(12) ,
  \V180(14) ,
  \V56(2) ,
  \V88(24) ,
  \V126(4) ,
  \V56(15) ,
  \V56(3) ,
  \V56(14) ,
  \V56(4) ,
  \V56(5) ,
  \V88(21) ,
  \V126(1) ,
  \V56(6) ,
  \V88(20) ,
  \V126(0) ,
  \V56(11) ,
  \V56(7) ,
  \V189(2) ,
  \V56(10) ,
  \V56(8) ,
  \V56(9) ,
  \V88(27) ,
  \V88(26) ,
  \V189(1) ,
  \V56(17) ,
  \V88(29) ,
  \V189(0) ,
  \V56(16) ,
  \V88(28) ,
  \V56(19) ,
  \V56(18) ,
  \V56(23) ,
  \V56(22) ,
  \V56(25) ,
  \V56(24) ,
  \V88(31) ,
  \V88(30) ,
  \V56(21) ,
  \V56(20) ,
  \V56(27) ,
  \V56(26) ,
  \V120(27) ,
  \V120(26) ,
  \V120(29) ,
  \V120(28) ,
  \V168(10) ,
  \V168(2) ,
  \V168(13) ,
  \V168(5) ,
  \V168(12) ,
  \V168(4) ,
  \V120(21) ,
  \V120(20) ,
  \V168(14) ,
  \V120(23) ,
  \V28(13) ,
  \V168(1) ,
  \V120(22) ,
  \V28(12) ,
  \V168(0) ,
  \V120(25) ,
  \V28(15) ,
  \V120(24) ,
  \V28(14) ,
  \V120(17) ,
  \V120(16) ,
  \V156(2) ,
  \V120(19) ,
  \V28(11) ,
  \V156(5) ,
  \V120(18) ,
  \V28(10) ,
  \V168(6) ,
  \V156(4) ,
  \V168(9) ,
  \V168(8) ,
  \V156(1) ,
  \V156(0) ,
  \V28(17) ,
  \V28(16) ,
  \V192(2) ,
  \V120(11) ,
  \V28(19) ,
  \V120(10) ,
  \V28(18) ,
  \V144(2) ,
  \V120(13) ,
  \V28(23) ,
  \V144(5) ,
  \V120(12) ,
  \V28(22) ,
  \V156(6) ,
  \V144(4) ,
  \V120(15) ,
  \V88(0) ,
  \V28(25) ,
  \V156(9) ,
  \V192(1) ,
  \V120(14) ,
  \V88(1) ,
  \V28(24) ,
  \V156(8) ,
  \V192(0) ,
  \V88(2) ,
  \V144(1) ,
  \V88(3) ,
  \V144(0) ,
  \V88(4) ,
  \V28(21) ,
  \V88(5) ,
  \V28(20) ,
  \V180(2) ,
  \V88(6) ,
  \V132(3) ,
  \V180(5) ,
  \V88(7) ,
  \V132(2) ,
  \V180(4) ,
  \V88(8) ,
  \V132(5) ,
  \V88(9) ,
  \V144(6) ,
  \V132(4) ,
  \V28(27) ,
  \V144(9) ,
  \V180(1) ,
  \V28(26) ,
  \V144(8) ,
  \V180(0) ,
  \V28(0) ,
  \V132(1) ,
  \V156(10) ,
  \V28(1) ,
  \V132(0) ,
  \V156(13) ,
  \V28(2) ,
  \V156(12) ,
  \V28(3) ,
  \V28(4) ,
  \V120(3) ,
  \V156(14) ,
  \V28(5) ,
  \V180(6) ,
  \V120(2) ,
  \V28(6) ,
  \V180(9) ,
  \V120(5) ,
  \V28(7) ,
  \V180(8) ,
  \V120(4) ,
  \V28(8) ,
  \V28(9) ,
  \V120(1) ,
  \V120(0) ,
  \V183(2) ,
  \V120(31) ,
  \V120(7) ,
  \V120(30) ,
  \V120(6) ,
  \V183(1) ,
  \V120(9) ,
  \V183(0) ,
  \V120(8) ,
  \V88(13) ,
  \V88(12) ,
  \V88(15) ,
  \V88(14) ;
output
  \V194(1) ,
  \V194(0) ,
  \V198(3) ,
  \V198(2) ,
  \V198(1) ,
  \V198(0) ;
wire
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  V199,
  \V274(3) ,
  \V274(2) ,
  \V274(1) ,
  V200,
  V201,
  V202,
  V203,
  V204,
  V205,
  V206,
  V207,
  V208,
  V209,
  V210,
  V211,
  V212,
  V213,
  V214,
  V215,
  V216,
  V217,
  V218,
  V219,
  V220,
  V221,
  V222,
  V223,
  V224,
  V225,
  V226,
  V230,
  V231,
  V232,
  V233,
  V234,
  V235,
  V236,
  V237,
  V238,
  V239,
  V240,
  V241,
  V245,
  V246,
  V247,
  V248,
  V249,
  V250,
  V251,
  V252,
  V253,
  V254,
  V255,
  V256,
  V260,
  V261,
  V262,
  V263,
  V264,
  V265,
  V266,
  V267,
  V268,
  V269,
  V270,
  V271,
  V275,
  V276,
  V277,
  V278,
  V279,
  V280,
  V281,
  V282,
  V283,
  V284,
  V285,
  V286,
  \V229(3) ,
  \V229(2) ,
  \V229(1) ,
  \V244(3) ,
  \V244(2) ,
  \V244(1) ,
  \V259(3) ,
  \V259(2) ,
  \V259(1) ;
assign
  \[0]  = \V28(0)  & \V56(0) ,
  \[1]  = \V28(1)  & \V56(1) ,
  \[2]  = V276 | (V217 | (V215 | (V199 | (V216 | (V275 | V277))))),
  \[3]  = V279 | (V232 | (V230 | (V203 | (V231 | (V278 | V280))))),
  \[4]  = V282 | (V247 | (V245 | (V207 | (V246 | (V281 | V283))))),
  \[5]  = V285 | (V262 | (V260 | (V211 | (V261 | (V284 | V286))))),
  V199 = \V28(2)  & \V56(2) ,
  \V274(3)  = V270 | (V214 | (V269 | V271)),
  \V274(2)  = V267 | (V213 | (V266 | V268)),
  \V274(1)  = V264 | (V212 | (V263 | V265)),
  V200 = \V28(6)  & \V56(6) ,
  V201 = \V28(10)  & \V56(10) ,
  V202 = \V28(14)  & \V56(14) ,
  V203 = \V28(18)  & \V56(18) ,
  V204 = \V28(22)  & \V56(22) ,
  V205 = \V28(26)  & \V56(26) ,
  V206 = \V88(2)  & \V120(2) ,
  V207 = \V88(6)  & \V120(6) ,
  V208 = \V88(10)  & \V120(10) ,
  V209 = \V88(14)  & \V120(14) ,
  V210 = \V88(18)  & \V120(18) ,
  V211 = \V88(22)  & \V120(22) ,
  V212 = \V88(26)  & \V120(26) ,
  V213 = \V88(30)  & \V120(30) ,
  V214 = \V126(2)  & \V132(2) ,
  V215 = \V56(3)  & (\V28(3)  & \V144(0) ),
  V216 = \V144(0)  & (\V28(4)  & (\V56(4)  & \V144(1) )),
  V217 = \V144(1)  & (\V56(5)  & (\V28(5)  & (\V144(0)  & \V144(2) ))),
  V218 = \V56(7)  & (\V28(7)  & \V144(4) ),
  V219 = \V144(4)  & (\V28(8)  & (\V56(8)  & \V144(5) )),
  V220 = \V144(5)  & (\V56(9)  & (\V28(9)  & (\V144(4)  & \V144(6) ))),
  V221 = \V56(11)  & (\V28(11)  & \V144(8) ),
  V222 = \V144(8)  & (\V28(12)  & (\V56(12)  & \V144(9) )),
  V223 = \V144(9)  & (\V56(13)  & (\V28(13)  & (\V144(8)  & \V144(10) ))),
  V224 = \V56(15)  & (\V28(15)  & \V144(12) ),
  V225 = \V144(12)  & (\V28(16)  & (\V56(16)  & \V144(13) )),
  V226 = \V144(13)  & (\V56(17)  & (\V28(17)  & (\V144(12)  & \V144(14) ))),
  V230 = \V56(19)  & (\V28(19)  & \V156(0) ),
  V231 = \V156(0)  & (\V28(20)  & (\V56(20)  & \V156(1) )),
  V232 = \V156(1)  & (\V56(21)  & (\V28(21)  & (\V156(0)  & \V156(2) ))),
  V233 = \V56(23)  & (\V28(23)  & \V156(4) ),
  V234 = \V156(4)  & (\V28(24)  & (\V56(24)  & \V156(5) )),
  V235 = \V156(5)  & (\V56(25)  & (\V28(25)  & (\V156(4)  & \V156(6) ))),
  V236 = \V56(27)  & (\V28(27)  & \V156(8) ),
  V237 = \V156(8)  & (\V88(0)  & (\V120(0)  & \V156(9) )),
  V238 = \V156(9)  & (\V120(1)  & (\V88(1)  & (\V156(8)  & \V156(10) ))),
  V239 = \V120(3)  & (\V88(3)  & \V156(12) ),
  V240 = \V156(12)  & (\V88(4)  & (\V120(4)  & \V156(13) )),
  V241 = \V156(13)  & (\V120(5)  & (\V88(5)  & (\V156(12)  & \V156(14) ))),
  V245 = \V120(7)  & (\V88(7)  & \V168(0) ),
  V246 = \V168(0)  & (\V88(8)  & (\V120(8)  & \V168(1) )),
  V247 = \V168(1)  & (\V120(9)  & (\V88(9)  & (\V168(0)  & \V168(2) ))),
  V248 = \V120(11)  & (\V88(11)  & \V168(4) ),
  V249 = \V168(4)  & (\V88(12)  & (\V120(12)  & \V168(5) )),
  V250 = \V168(5)  & (\V120(13)  & (\V88(13)  & (\V168(4)  & \V168(6) ))),
  V251 = \V120(15)  & (\V88(15)  & \V168(8) ),
  V252 = \V168(8)  & (\V88(16)  & (\V120(16)  & \V168(9) )),
  V253 = \V168(9)  & (\V120(17)  & (\V88(17)  & (\V168(8)  & \V168(10) ))),
  V254 = \V120(19)  & (\V88(19)  & \V168(12) ),
  V255 = \V168(12)  & (\V88(20)  & (\V120(20)  & \V168(13) )),
  V256 = \V168(13)  & (\V120(21)  & (\V88(21)  & (\V168(12)  & \V168(14) ))),
  V260 = \V120(23)  & (\V88(23)  & \V180(0) ),
  V261 = \V180(0)  & (\V88(24)  & (\V120(24)  & \V180(1) )),
  V262 = \V180(1)  & (\V120(25)  & (\V88(25)  & (\V180(0)  & \V180(2) ))),
  V263 = \V120(27)  & (\V88(27)  & \V180(4) ),
  V264 = \V180(4)  & (\V88(28)  & (\V120(28)  & \V180(5) )),
  V265 = \V180(5)  & (\V120(29)  & (\V88(29)  & (\V180(4)  & \V180(6) ))),
  V266 = \V120(31)  & (\V88(31)  & \V180(8) ),
  V267 = \V180(8)  & (\V126(0)  & (\V132(0)  & \V180(9) )),
  V268 = \V180(9)  & (\V132(1)  & (\V126(1)  & (\V180(8)  & \V180(10) ))),
  V269 = \V132(3)  & (\V126(3)  & \V180(12) ),
  V270 = \V180(12)  & (\V126(4)  & (\V132(4)  & \V180(13) )),
  V271 = \V180(13)  & (\V132(5)  & (\V126(5)  & (\V180(12)  & \V180(14) ))),
  V275 = \V229(1)  & \V183(0) ,
  V276 = \V183(0)  & (\V229(2)  & \V183(1) ),
  V277 = \V183(1)  & (\V229(3)  & (\V183(0)  & \V183(2) )),
  V278 = \V244(1)  & \V186(0) ,
  V279 = \V186(0)  & (\V244(2)  & \V186(1) ),
  V280 = \V186(1)  & (\V244(3)  & (\V186(0)  & \V186(2) )),
  V281 = \V259(1)  & \V189(0) ,
  V282 = \V189(0)  & (\V259(2)  & \V189(1) ),
  V283 = \V189(1)  & (\V259(3)  & (\V189(0)  & \V189(2) )),
  V284 = \V274(1)  & \V192(0) ,
  V285 = \V192(0)  & (\V274(2)  & \V192(1) ),
  V286 = \V192(1)  & (\V274(3)  & (\V192(0)  & \V192(2) )),
  \V229(3)  = V225 | (V202 | (V224 | V226)),
  \V229(2)  = V222 | (V201 | (V221 | V223)),
  \V229(1)  = V219 | (V200 | (V218 | V220)),
  \V244(3)  = V240 | (V206 | (V239 | V241)),
  \V244(2)  = V237 | (V205 | (V236 | V238)),
  \V244(1)  = V234 | (V204 | (V233 | V235)),
  \V194(1)  = \[1] ,
  \V194(0)  = \[0] ,
  \V259(3)  = V255 | (V210 | (V254 | V256)),
  \V259(2)  = V252 | (V209 | (V251 | V253)),
  \V259(1)  = V249 | (V208 | (V248 | V250)),
  \V198(3)  = \[5] ,
  \V198(2)  = \[4] ,
  \V198(1)  = \[3] ,
  \V198(0)  = \[2] ;
endmodule

