// IWLS benchmark module "bigkey" printed on Wed May 29 21:51:13 2002
module bigkey(\key<255> , \key<254> , \key<253> , \key<252> , \key<251> , \key<250> , \key<249> , \key<248> , \key<247> , \key<246> , \key<245> , \key<244> , \key<243> , \key<242> , \key<241> , \key<240> , \key<239> , \key<238> , \key<237> , \key<236> , \key<235> , \key<234> , \key<233> , \key<232> , \key<231> , \key<230> , \key<229> , \key<228> , \key<227> , \key<226> , \key<225> , \key<224> , \key<223> , \key<222> , \key<221> , \key<220> , \key<219> , \key<218> , \key<217> , \key<216> , \key<215> , \key<214> , \key<213> , \key<212> , \key<211> , \key<210> , \key<209> , \key<208> , \key<207> , \key<206> , \key<205> , \key<204> , \key<203> , \key<202> , \key<201> , \key<200> , \key<199> , \key<198> , \key<197> , \key<196> , \key<195> , \key<194> , \key<193> , \key<192> , \key<191> , \key<190> , \key<189> , \key<188> , \key<187> , \key<186> , \key<185> , \key<184> , \key<183> , \key<182> , \key<181> , \key<180> , \key<179> , \key<178> , \key<177> , \key<176> , \key<175> , \key<174> , \key<173> , \key<172> , \key<171> , \key<170> , \key<169> , \key<168> , \key<167> , \key<166> , \key<165> , \key<164> , \key<163> , \key<162> , \key<161> , \key<160> , \key<159> , \key<158> , \key<157> , \key<156> , \key<155> , \key<154> , \key<153> , \key<152> , \key<151> , \key<150> , \key<149> , \key<148> , \key<147> , \key<146> , \key<145> , \key<144> , \key<143> , \key<142> , \key<141> , \key<140> , \key<139> , \key<138> , \key<137> , \key<136> , \key<135> , \key<134> , \key<133> , \key<132> , \key<131> , \key<130> , \key<129> , \key<128> , \key<127> , \key<126> , \key<125> , \key<124> , \key<123> , \key<122> , \key<121> , \key<120> , \key<119> , \key<118> , \key<117> , \key<116> , \key<115> , \key<114> , \key<113> , \key<112> , \key<111> , \key<110> , \key<109> , \key<108> , \key<107> , \key<106> , \key<105> , \key<104> , \key<103> , \key<102> , \key<101> , \key<100> , \key<99> , \key<98> , \key<97> , \key<96> , \key<95> , \key<94> , \key<93> , \key<92> , \key<91> , \key<90> , \key<89> , \key<88> , \key<87> , \key<86> , \key<85> , \key<84> , \key<83> , \key<82> , \key<81> , \key<80> , \key<79> , \key<78> , \key<77> , \key<76> , \key<75> , \key<74> , \key<73> , \key<72> , \key<71> , \key<70> , \key<69> , \key<68> , \key<67> , \key<66> , \key<65> , \key<64> , \key<63> , \key<62> , \key<61> , \key<60> , \key<59> , \key<58> , \key<57> , \key<56> , \key<55> , \key<54> , \key<53> , \key<52> , \key<51> , \key<50> , \key<49> , \key<48> , \key<47> , \key<46> , \key<45> , \key<44> , \key<43> , \key<42> , \key<41> , \key<40> , \key<39> , \key<38> , \key<37> , \key<36> , \key<35> , \key<34> , \key<33> , \key<32> , \key<31> , \key<30> , \key<29> , \key<28> , \key<27> , \key<26> , \key<25> , \key<24> , \key<23> , \key<22> , \key<21> , \key<20> , \key<19> , \key<18> , \key<17> , \key<16> , \key<15> , \key<14> , \key<13> , \key<12> , \key<11> , \key<10> , \key<9> , \key<8> , \key<7> , \key<6> , \key<5> , \key<4> , \key<3> , \key<2> , \key<1> , \key<0> , \encrypt<0> , \start<0> , \count<3> , \count<2> , \count<1> , \count<0> , \new_count<3> , \new_count<2> , \new_count<1> , \new_count<0> , \data_ready<0> , \KSi<191> , \KSi<190> , \KSi<189> , \KSi<188> , \KSi<187> , \KSi<186> , \KSi<185> , \KSi<184> , \KSi<183> , \KSi<182> , \KSi<181> , \KSi<180> , \KSi<179> , \KSi<178> , \KSi<177> , \KSi<176> , \KSi<175> , \KSi<174> , \KSi<173> , \KSi<172> , \KSi<171> , \KSi<170> , \KSi<169> , \KSi<168> , \KSi<167> , \KSi<166> , \KSi<165> , \KSi<164> , \KSi<163> , \KSi<162> , \KSi<161> , \KSi<160> , \KSi<159> , \KSi<158> , \KSi<157> , \KSi<156> , \KSi<155> , \KSi<154> , \KSi<153> , \KSi<152> , \KSi<151> , \KSi<150> , \KSi<149> , \KSi<148> , \KSi<147> , \KSi<146> , \KSi<145> , \KSi<144> , \KSi<143> , \KSi<142> , \KSi<141> , \KSi<140> , \KSi<139> , \KSi<138> , \KSi<137> , \KSi<136> , \KSi<135> , \KSi<134> , \KSi<133> , \KSi<132> , \KSi<131> , \KSi<130> , \KSi<129> , \KSi<128> , \KSi<127> , \KSi<126> , \KSi<125> , \KSi<124> , \KSi<123> , \KSi<122> , \KSi<121> , \KSi<120> , \KSi<119> , \KSi<118> , \KSi<117> , \KSi<116> , \KSi<115> , \KSi<114> , \KSi<113> , \KSi<112> , \KSi<111> , \KSi<110> , \KSi<109> , \KSi<108> , \KSi<107> , \KSi<106> , \KSi<105> , \KSi<104> , \KSi<103> , \KSi<102> , \KSi<101> , \KSi<100> , \KSi<99> , \KSi<98> , \KSi<97> , \KSi<96> , \KSi<95> , \KSi<94> , \KSi<93> , \KSi<92> , \KSi<91> , \KSi<90> , \KSi<89> , \KSi<88> , \KSi<87> , \KSi<86> , \KSi<85> , \KSi<84> , \KSi<83> , \KSi<82> , \KSi<81> , \KSi<80> , \KSi<79> , \KSi<78> , \KSi<77> , \KSi<76> , \KSi<75> , \KSi<74> , \KSi<73> , \KSi<72> , \KSi<71> , \KSi<70> , \KSi<69> , \KSi<68> , \KSi<67> , \KSi<66> , \KSi<65> , \KSi<64> , \KSi<63> , \KSi<62> , \KSi<61> , \KSi<60> , \KSi<59> , \KSi<58> , \KSi<57> , \KSi<56> , \KSi<55> , \KSi<54> , \KSi<53> , \KSi<52> , \KSi<51> , \KSi<50> , \KSi<49> , \KSi<48> , \KSi<47> , \KSi<46> , \KSi<45> , \KSi<44> , \KSi<43> , \KSi<42> , \KSi<41> , \KSi<40> , \KSi<39> , \KSi<38> , \KSi<37> , \KSi<36> , \KSi<35> , \KSi<34> , \KSi<33> , \KSi<32> , \KSi<31> , \KSi<30> , \KSi<29> , \KSi<28> , \KSi<27> , \KSi<26> , \KSi<25> , \KSi<24> , \KSi<23> , \KSi<22> , \KSi<21> , \KSi<20> , \KSi<19> , \KSi<18> , \KSi<17> , \KSi<16> , \KSi<15> , \KSi<14> , \KSi<13> , \KSi<12> , \KSi<11> , \KSi<10> , \KSi<9> , \KSi<8> , \KSi<7> , \KSi<6> , \KSi<5> , \KSi<4> , \KSi<3> , \KSi<2> , \KSi<1> , \KSi<0> );
input
  \key<156> ,
  \key<155> ,
  \key<158> ,
  \key<157> ,
  \key<159> ,
  \key<240> ,
  \key<14> ,
  \key<13> ,
  \key<242> ,
  \key<12> ,
  \key<241> ,
  \key<11> ,
  \key<244> ,
  \key<10> ,
  \key<243> ,
  \key<246> ,
  \key<245> ,
  \key<248> ,
  \key<247> ,
  \key<249> ,
  \key<19> ,
  \key<18> ,
  \key<17> ,
  \key<0> ,
  \key<16> ,
  \key<1> ,
  \key<15> ,
  \key<2> ,
  \key<230> ,
  \key<24> ,
  \key<3> ,
  \key<23> ,
  \key<4> ,
  \key<232> ,
  \key<22> ,
  \key<5> ,
  \key<231> ,
  \key<21> ,
  \key<6> ,
  \key<234> ,
  \key<20> ,
  \key<7> ,
  \key<233> ,
  \key<8> ,
  \key<236> ,
  \key<9> ,
  \key<235> ,
  \key<238> ,
  \key<237> ,
  \key<239> ,
  \key<29> ,
  \key<28> ,
  \key<27> ,
  \key<26> ,
  \key<25> ,
  \key<220> ,
  \key<34> ,
  \key<33> ,
  \key<222> ,
  \key<32> ,
  \key<221> ,
  \key<31> ,
  \key<224> ,
  \key<30> ,
  \key<223> ,
  \key<226> ,
  \key<225> ,
  \key<228> ,
  \key<227> ,
  \key<229> ,
  \key<39> ,
  \key<38> ,
  \key<37> ,
  \key<36> ,
  \key<35> ,
  \key<210> ,
  \key<44> ,
  \key<43> ,
  \key<212> ,
  \key<42> ,
  \key<211> ,
  \key<41> ,
  \key<214> ,
  \key<40> ,
  \key<213> ,
  \key<216> ,
  \key<215> ,
  \key<218> ,
  \key<217> ,
  \key<219> ,
  \key<49> ,
  \key<48> ,
  \key<47> ,
  \key<46> ,
  \key<45> ,
  \key<200> ,
  \key<54> ,
  \key<53> ,
  \key<202> ,
  \key<52> ,
  \key<201> ,
  \key<51> ,
  \key<204> ,
  \key<50> ,
  \key<203> ,
  \key<206> ,
  \key<205> ,
  \key<208> ,
  \key<207> ,
  \key<209> ,
  \key<59> ,
  \key<58> ,
  \key<57> ,
  \key<56> ,
  \key<55> ,
  \key<64> ,
  \key<63> ,
  \key<62> ,
  \key<61> ,
  \key<60> ,
  \key<69> ,
  \key<68> ,
  \key<67> ,
  \key<66> ,
  \key<65> ,
  \key<74> ,
  \key<73> ,
  \key<72> ,
  \key<71> ,
  \key<70> ,
  \key<79> ,
  \key<78> ,
  \key<77> ,
  \key<76> ,
  \key<75> ,
  \key<84> ,
  \key<83> ,
  \key<82> ,
  \key<81> ,
  \key<80> ,
  \key<89> ,
  \key<88> ,
  \key<87> ,
  \key<86> ,
  \key<85> ,
  \key<94> ,
  \key<93> ,
  \key<92> ,
  \key<91> ,
  \key<90> ,
  \key<99> ,
  \key<98> ,
  \key<97> ,
  \key<96> ,
  \key<95> ,
  \start<0> ,
  \key<140> ,
  \key<250> ,
  \key<142> ,
  \key<252> ,
  \key<141> ,
  \key<251> ,
  \key<144> ,
  \key<254> ,
  \key<143> ,
  \key<253> ,
  \key<146> ,
  \key<145> ,
  \key<255> ,
  \key<148> ,
  \key<147> ,
  \key<149> ,
  \key<130> ,
  \key<132> ,
  \key<131> ,
  \key<134> ,
  \key<133> ,
  \key<136> ,
  \key<135> ,
  \key<138> ,
  \key<137> ,
  \key<139> ,
  \count<0> ,
  \count<3> ,
  \key<120> ,
  \count<1> ,
  \key<122> ,
  \count<2> ,
  \key<121> ,
  \key<124> ,
  \key<123> ,
  \key<126> ,
  \key<125> ,
  \key<128> ,
  \key<127> ,
  \key<129> ,
  \key<110> ,
  \key<112> ,
  \key<111> ,
  \key<114> ,
  \key<113> ,
  \key<116> ,
  \key<115> ,
  \key<118> ,
  \key<117> ,
  \key<119> ,
  \key<100> ,
  \key<102> ,
  \key<101> ,
  \key<104> ,
  \key<103> ,
  \key<106> ,
  \key<105> ,
  \key<108> ,
  \key<107> ,
  \key<109> ,
  \key<190> ,
  \key<192> ,
  \key<191> ,
  \key<194> ,
  \key<193> ,
  \key<196> ,
  \key<195> ,
  \key<198> ,
  \key<197> ,
  \key<199> ,
  \key<180> ,
  \key<182> ,
  \key<181> ,
  \key<184> ,
  \key<183> ,
  \key<186> ,
  \key<185> ,
  \key<188> ,
  \key<187> ,
  \key<189> ,
  \key<170> ,
  \key<172> ,
  \key<171> ,
  \key<174> ,
  \key<173> ,
  \key<176> ,
  \key<175> ,
  \key<178> ,
  \key<177> ,
  \key<179> ,
  \encrypt<0> ,
  \key<160> ,
  \key<162> ,
  \key<161> ,
  \key<164> ,
  \key<163> ,
  \key<166> ,
  \key<165> ,
  \key<168> ,
  \key<167> ,
  \key<169> ,
  \key<150> ,
  \key<152> ,
  \key<151> ,
  \key<154> ,
  \key<153> ;
output
  \KSi<130> ,
  \KSi<131> ,
  \KSi<132> ,
  \KSi<133> ,
  \KSi<134> ,
  \KSi<135> ,
  \KSi<136> ,
  \KSi<137> ,
  \KSi<138> ,
  \KSi<139> ,
  \KSi<100> ,
  \KSi<101> ,
  \KSi<102> ,
  \KSi<103> ,
  \KSi<104> ,
  \KSi<105> ,
  \KSi<106> ,
  \KSi<107> ,
  \KSi<108> ,
  \KSi<109> ,
  \KSi<190> ,
  \KSi<191> ,
  \KSi<160> ,
  \KSi<161> ,
  \KSi<162> ,
  \KSi<163> ,
  \KSi<164> ,
  \KSi<165> ,
  \KSi<166> ,
  \KSi<167> ,
  \KSi<168> ,
  \KSi<169> ,
  \KSi<150> ,
  \KSi<151> ,
  \KSi<152> ,
  \KSi<153> ,
  \KSi<154> ,
  \KSi<155> ,
  \KSi<156> ,
  \KSi<157> ,
  \KSi<158> ,
  \KSi<159> ,
  \KSi<0> ,
  \KSi<1> ,
  \KSi<2> ,
  \KSi<3> ,
  \KSi<4> ,
  \KSi<180> ,
  \KSi<5> ,
  \KSi<181> ,
  \KSi<6> ,
  \KSi<182> ,
  \KSi<7> ,
  \KSi<183> ,
  \KSi<8> ,
  \KSi<184> ,
  \KSi<9> ,
  \KSi<185> ,
  \KSi<186> ,
  \KSi<187> ,
  \KSi<188> ,
  \KSi<189> ,
  \KSi<170> ,
  \KSi<171> ,
  \KSi<172> ,
  \KSi<173> ,
  \KSi<174> ,
  \KSi<175> ,
  \KSi<176> ,
  \KSi<177> ,
  \KSi<178> ,
  \KSi<179> ,
  \new_count<0> ,
  \new_count<3> ,
  \new_count<1> ,
  \new_count<2> ,
  \KSi<12> ,
  \KSi<11> ,
  \KSi<14> ,
  \KSi<13> ,
  \KSi<10> ,
  \KSi<19> ,
  \KSi<16> ,
  \KSi<15> ,
  \KSi<18> ,
  \KSi<17> ,
  \KSi<22> ,
  \KSi<21> ,
  \KSi<24> ,
  \KSi<23> ,
  \KSi<20> ,
  \KSi<29> ,
  \KSi<26> ,
  \KSi<25> ,
  \KSi<28> ,
  \KSi<27> ,
  \KSi<32> ,
  \KSi<31> ,
  \KSi<34> ,
  \KSi<33> ,
  \KSi<30> ,
  \KSi<39> ,
  \KSi<36> ,
  \KSi<35> ,
  \KSi<38> ,
  \KSi<37> ,
  \KSi<42> ,
  \KSi<41> ,
  \KSi<44> ,
  \KSi<43> ,
  \KSi<40> ,
  \KSi<49> ,
  \KSi<46> ,
  \KSi<45> ,
  \KSi<48> ,
  \KSi<47> ,
  \KSi<52> ,
  \KSi<51> ,
  \KSi<54> ,
  \KSi<53> ,
  \KSi<50> ,
  \KSi<59> ,
  \KSi<56> ,
  \KSi<55> ,
  \KSi<58> ,
  \KSi<57> ,
  \KSi<62> ,
  \KSi<61> ,
  \KSi<64> ,
  \KSi<63> ,
  \KSi<60> ,
  \KSi<69> ,
  \KSi<66> ,
  \data_ready<0> ,
  \KSi<65> ,
  \KSi<68> ,
  \KSi<67> ,
  \KSi<72> ,
  \KSi<71> ,
  \KSi<74> ,
  \KSi<73> ,
  \KSi<70> ,
  \KSi<79> ,
  \KSi<76> ,
  \KSi<75> ,
  \KSi<78> ,
  \KSi<77> ,
  \KSi<82> ,
  \KSi<81> ,
  \KSi<84> ,
  \KSi<83> ,
  \KSi<80> ,
  \KSi<89> ,
  \KSi<86> ,
  \KSi<85> ,
  \KSi<88> ,
  \KSi<87> ,
  \KSi<92> ,
  \KSi<91> ,
  \KSi<94> ,
  \KSi<93> ,
  \KSi<90> ,
  \KSi<99> ,
  \KSi<96> ,
  \KSi<95> ,
  \KSi<98> ,
  \KSi<97> ,
  \KSi<120> ,
  \KSi<121> ,
  \KSi<122> ,
  \KSi<123> ,
  \KSi<124> ,
  \KSi<125> ,
  \KSi<126> ,
  \KSi<127> ,
  \KSi<128> ,
  \KSi<129> ,
  \KSi<110> ,
  \KSi<111> ,
  \KSi<112> ,
  \KSi<113> ,
  \KSi<114> ,
  \KSi<115> ,
  \KSi<116> ,
  \KSi<117> ,
  \KSi<118> ,
  \KSi<119> ,
  \KSi<140> ,
  \KSi<141> ,
  \KSi<142> ,
  \KSi<143> ,
  \KSi<144> ,
  \KSi<145> ,
  \KSi<146> ,
  \KSi<147> ,
  \KSi<148> ,
  \KSi<149> ;
reg
  \D<0> ,
  \D<1> ,
  \D<2> ,
  \D<3> ,
  \D<4> ,
  \D<5> ,
  \D<6> ,
  \C<10> ,
  \D<7> ,
  \C<11> ,
  \D<8> ,
  \C<12> ,
  \D<9> ,
  \C<13> ,
  \C<14> ,
  \C<15> ,
  \C<16> ,
  \C<17> ,
  \C<18> ,
  \C<19> ,
  \C<20> ,
  \C<21> ,
  \C<22> ,
  \C<23> ,
  \C<24> ,
  \C<25> ,
  \C<26> ,
  \C<27> ,
  \C<28> ,
  \C<29> ,
  \C<30> ,
  \C<31> ,
  \C<32> ,
  \C<33> ,
  \C<34> ,
  \C<35> ,
  \C<36> ,
  \C<37> ,
  \C<38> ,
  \C<39> ,
  \C<40> ,
  \C<41> ,
  \C<42> ,
  \C<43> ,
  \C<44> ,
  \C<45> ,
  \C<46> ,
  \C<47> ,
  \C<48> ,
  \C<49> ,
  \C<50> ,
  \C<51> ,
  \C<52> ,
  \C<53> ,
  \C<54> ,
  \C<55> ,
  \C<56> ,
  \C<57> ,
  \C<58> ,
  \C<59> ,
  \C<60> ,
  \C<61> ,
  \C<62> ,
  \C<63> ,
  \C<64> ,
  \C<65> ,
  \C<66> ,
  \C<67> ,
  \C<68> ,
  \C<69> ,
  \C<70> ,
  \C<71> ,
  \C<72> ,
  \C<73> ,
  \C<74> ,
  \C<75> ,
  \C<76> ,
  \C<77> ,
  \C<78> ,
  \C<79> ,
  \C<80> ,
  \C<81> ,
  \C<82> ,
  \C<83> ,
  \C<84> ,
  \C<85> ,
  \C<86> ,
  \C<87> ,
  \C<88> ,
  \C<89> ,
  \C<90> ,
  \C<91> ,
  \D<10> ,
  \C<92> ,
  \D<11> ,
  \C<93> ,
  \D<12> ,
  \C<94> ,
  \D<13> ,
  \C<95> ,
  \D<14> ,
  \C<96> ,
  \D<15> ,
  \C<97> ,
  \D<16> ,
  \C<98> ,
  \D<17> ,
  \C<99> ,
  \D<18> ,
  \D<19> ,
  \D<20> ,
  \D<21> ,
  \D<22> ,
  \D<23> ,
  \D<24> ,
  \D<25> ,
  \D<26> ,
  \D<27> ,
  \D<28> ,
  \D<29> ,
  \D<30> ,
  \D<31> ,
  \D<32> ,
  \D<33> ,
  \D<34> ,
  \D<35> ,
  \D<36> ,
  \D<37> ,
  \D<38> ,
  \D<39> ,
  \D<40> ,
  \D<41> ,
  \D<42> ,
  \D<43> ,
  \D<44> ,
  \D<45> ,
  \D<46> ,
  \D<47> ,
  \D<48> ,
  \D<49> ,
  \D<50> ,
  \D<51> ,
  \D<52> ,
  \D<53> ,
  \D<54> ,
  \D<55> ,
  \D<56> ,
  \D<57> ,
  \D<58> ,
  \D<59> ,
  \D<60> ,
  \D<61> ,
  \D<62> ,
  \D<63> ,
  \D<64> ,
  \D<65> ,
  \D<66> ,
  \D<67> ,
  \D<68> ,
  \D<69> ,
  \C<100> ,
  \D<70> ,
  \C<101> ,
  \D<71> ,
  \C<102> ,
  \D<72> ,
  \C<103> ,
  \D<73> ,
  \C<104> ,
  \D<74> ,
  \C<105> ,
  \D<75> ,
  \C<106> ,
  \D<76> ,
  \C<107> ,
  \D<77> ,
  \C<108> ,
  \C<0> ,
  \D<78> ,
  \C<109> ,
  \C<1> ,
  \D<79> ,
  \C<2> ,
  \C<3> ,
  \C<4> ,
  \C<5> ,
  \C<6> ,
  \C<7> ,
  \C<110> ,
  \C<8> ,
  \D<80> ,
  \C<111> ,
  \C<9> ,
  \D<81> ,
  \D<82> ,
  \D<83> ,
  \D<84> ,
  \D<85> ,
  \D<86> ,
  \D<87> ,
  \D<88> ,
  \D<89> ,
  \D<90> ,
  \D<91> ,
  \D<92> ,
  \D<93> ,
  \D<94> ,
  \D<95> ,
  \D<96> ,
  \D<97> ,
  \D<98> ,
  \D<99> ,
  \D<100> ,
  \D<101> ,
  \D<102> ,
  \D<103> ,
  \D<104> ,
  \D<105> ,
  \D<106> ,
  \D<107> ,
  \D<108> ,
  \D<109> ,
  \D<110> ,
  \D<111> ;
wire
  \[378] ,
  \[568] ,
  \new_D<98> ,
  \[379] ,
  \[569] ,
  \new_D<91> ,
  \new_D<92> ,
  \new_D<93> ,
  \new_D<94> ,
  \[380] ,
  \[570] ,
  \new_D<90> ,
  \[381] ,
  \[571] ,
  \[382] ,
  \[572] ,
  \[383] ,
  \[573] ,
  \[384] ,
  \[574] ,
  \[385] ,
  \[575] ,
  \[386] ,
  \[576] ,
  \[387] ,
  \[577] ,
  \main/$MINUS_4_1/sum<3>8.1 ,
  \[388] ,
  \[578] ,
  \new_C<111> ,
  \[389] ,
  \[579] ,
  \new_C<110> ,
  \[390] ,
  \[580] ,
  \[391] ,
  \[581] ,
  \[392] ,
  \[582] ,
  \[393] ,
  \[583] ,
  \[394] ,
  \[584] ,
  \[395] ,
  \[585] ,
  \[396] ,
  \[586] ,
  \[397] ,
  \[587] ,
  \[398] ,
  \[588] ,
  \[399] ,
  \[589] ,
  \[590] ,
  \[591] ,
  \[592] ,
  \[593] ,
  \[594] ,
  \[595] ,
  \[596] ,
  \[597] ,
  \[598] ,
  \[599] ,
  \new_D<59> ,
  \main/$PLUS_5_1/sum<2>5.1 ,
  \new_D<55> ,
  \new_D<56> ,
  \new_D<57> ,
  \new_D<58> ,
  \new_D<51> ,
  \new_D<52> ,
  \new_D<53> ,
  \new_D<54> ,
  \new_D<50> ,
  \new_D<69> ,
  \new_D<65> ,
  \new_D<66> ,
  \new_D<67> ,
  \new_D<68> ,
  \new_D<61> ,
  \new_D<62> ,
  \new_D<63> ,
  \new_D<64> ,
  \new_D<60> ,
  \new_D<79> ,
  \new_D<75> ,
  \new_D<76> ,
  \new_D<77> ,
  \new_D<78> ,
  \new_D<71> ,
  \new_D<72> ,
  \new_D<73> ,
  \new_D<74> ,
  \new_D<70> ,
  \new_D<111> ,
  \new_D<89> ,
  \new_D<85> ,
  \new_D<110> ,
  \new_D<86> ,
  \new_D<87> ,
  \new_D<88> ,
  \new_D<81> ,
  \new_D<82> ,
  \new_D<83> ,
  \new_D<84> ,
  \new_C<109> ,
  \new_D<80> ,
  \main/$MINUS_4_1/sum<2>8.1 ,
  \new_C<106> ,
  \new_C<105> ,
  \new_C<108> ,
  \new_C<107> ,
  \new_C<102> ,
  \new_C<101> ,
  \new_C<104> ,
  \new_C<103> ,
  \new_C<100> ,
  \[400] ,
  \[401] ,
  \[402] ,
  \[403] ,
  \[404] ,
  \[405] ,
  \[406] ,
  \[407] ,
  \[408] ,
  \[409] ,
  \[410] ,
  \[600] ,
  \[411] ,
  \[601] ,
  \[412] ,
  \[602] ,
  \[413] ,
  \[603] ,
  \[224] ,
  \[414] ,
  \[604] ,
  \[225] ,
  \[415] ,
  \[605] ,
  \[226] ,
  \[416] ,
  \[606] ,
  \[227] ,
  \[417] ,
  \[607] ,
  \[228] ,
  \[418] ,
  \[608] ,
  \[229] ,
  \[419] ,
  \[609] ,
  \[230] ,
  \[420] ,
  \[610] ,
  \[231] ,
  \[421] ,
  \[611] ,
  \[232] ,
  \[422] ,
  \[612] ,
  \[233] ,
  \[423] ,
  \[613] ,
  \[234] ,
  \[424] ,
  \[614] ,
  \[235] ,
  \[425] ,
  \[615] ,
  \[236] ,
  \[426] ,
  \[616] ,
  \new_D<1> ,
  \[237] ,
  \[427] ,
  \[617] ,
  \new_D<2> ,
  \[238] ,
  \[428] ,
  \[618] ,
  \new_D<3> ,
  \[239] ,
  \[429] ,
  \[619] ,
  \new_D<4> ,
  \new_D<0> ,
  \new_D<9> ,
  \[240] ,
  \[430] ,
  \[620] ,
  \[241] ,
  \[431] ,
  \[621] ,
  \[242] ,
  \[432] ,
  \[622] ,
  \new_D<5> ,
  \[243] ,
  \[433] ,
  \[623] ,
  \new_D<6> ,
  \[244] ,
  \[434] ,
  \[624] ,
  \main/$PLUS_5_1/sum<1>5.1 ,
  \new_D<7> ,
  \[245] ,
  \[435] ,
  \[625] ,
  \new_D<8> ,
  \[246] ,
  \[436] ,
  \[626] ,
  \[247] ,
  \[437] ,
  \[627] ,
  \[248] ,
  \[438] ,
  \[628] ,
  \[249] ,
  \[439] ,
  \[629] ,
  \[250] ,
  \[440] ,
  \[630] ,
  \[251] ,
  \[441] ,
  \[631] ,
  \[252] ,
  \[442] ,
  \[632] ,
  \[253] ,
  \[443] ,
  \[633] ,
  \[254] ,
  \[444] ,
  \[634] ,
  \[255] ,
  \[445] ,
  \[635] ,
  \[256] ,
  \[446] ,
  \[636] ,
  \[257] ,
  \[447] ,
  \[637] ,
  \[258] ,
  \[448] ,
  \[638] ,
  \[259] ,
  \[449] ,
  \[639] ,
  \new_D<109> ,
  \new_D<106> ,
  \new_D<105> ,
  \new_D<108> ,
  \new_D<107> ,
  \[260] ,
  \[450] ,
  \[640] ,
  \new_D<102> ,
  \[261] ,
  \[451] ,
  \[641] ,
  \new_D<101> ,
  \[262] ,
  \[452] ,
  \[642] ,
  \new_D<104> ,
  \[263] ,
  \[453] ,
  \[643] ,
  \new_D<103> ,
  \[264] ,
  \[454] ,
  \[644] ,
  \[265] ,
  \[455] ,
  \[266] ,
  \[456] ,
  \new_D<100> ,
  \[267] ,
  \[457] ,
  \[268] ,
  \[458] ,
  \[269] ,
  \[459] ,
  \[270] ,
  \[460] ,
  \new_C<19> ,
  \[271] ,
  \[461] ,
  \[272] ,
  \main/$PLUS_5_1/c<0>5.3 ,
  \main/$PLUS_5_1/c<0>5.4 ,
  \[462] ,
  \[273] ,
  \[463] ,
  \[274] ,
  \[464] ,
  \new_C<15> ,
  \[275] ,
  \[465] ,
  \new_C<16> ,
  \[276] ,
  \[466] ,
  \new_C<17> ,
  \[277] ,
  \[467] ,
  \new_C<18> ,
  \[278] ,
  \[468] ,
  \new_C<11> ,
  \[279] ,
  \[469] ,
  \new_C<12> ,
  \new_C<13> ,
  \new_C<14> ,
  \$$COND0<0>5.1 ,
  \new_C<10> ,
  \[280] ,
  \[470] ,
  \new_C<29> ,
  \[281] ,
  \[471] ,
  \[282] ,
  \[472] ,
  \[283] ,
  \[473] ,
  \[284] ,
  \[474] ,
  \new_C<25> ,
  \main/$MINUS_4_1/sum<1>8.1 ,
  \[285] ,
  \[475] ,
  \new_C<26> ,
  \[286] ,
  \[476] ,
  \new_C<27> ,
  \[287] ,
  \[477] ,
  \new_C<28> ,
  \[288] ,
  \[478] ,
  \new_C<21> ,
  \[289] ,
  \[479] ,
  \new_C<22> ,
  \new_C<23> ,
  \new_C<24> ,
  \new_C<20> ,
  \[290] ,
  \[480] ,
  \new_C<39> ,
  \[291] ,
  \[481] ,
  \[292] ,
  \[482] ,
  \[293] ,
  \[483] ,
  \[294] ,
  \[484] ,
  \new_C<35> ,
  \[295] ,
  \[485] ,
  \new_C<36> ,
  \[296] ,
  \[486] ,
  \new_C<37> ,
  \[297] ,
  \[487] ,
  \new_C<38> ,
  \[298] ,
  \[488] ,
  \new_C<31> ,
  \[299] ,
  \[489] ,
  \new_C<32> ,
  \main/$PLUS_5_1/sum<0>5.1 ,
  \new_C<33> ,
  \new_C<34> ,
  \new_C<30> ,
  \[490] ,
  \new_C<49> ,
  \[491] ,
  \[492] ,
  \[493] ,
  \[494] ,
  \new_C<45> ,
  \[495] ,
  \new_C<46> ,
  \[496] ,
  \new_C<47> ,
  \[497] ,
  \new_C<48> ,
  \[498] ,
  \new_C<41> ,
  \[499] ,
  \new_C<42> ,
  \new_C<43> ,
  \new_C<44> ,
  \new_C<40> ,
  \main/$MINUS_4_1/sum<0>8.1 ,
  \new_C<99> ,
  \new_D<19> ,
  \new_C<95> ,
  \new_C<96> ,
  \main/$MINUS_4_1/c<0>8.3 ,
  \main/$MINUS_4_1/c<0>8.4 ,
  \new_D<15> ,
  \new_C<97> ,
  \new_D<16> ,
  \new_C<98> ,
  \new_D<17> ,
  \new_C<91> ,
  \new_D<18> ,
  \new_C<92> ,
  \new_D<11> ,
  \new_C<93> ,
  \new_D<12> ,
  \new_C<94> ,
  \new_D<13> ,
  \new_D<14> ,
  \new_C<90> ,
  \[300] ,
  \new_D<10> ,
  \[301] ,
  \new_D<29> ,
  \[302] ,
  \[303] ,
  \[304] ,
  \[305] ,
  \new_D<25> ,
  \[306] ,
  \new_D<26> ,
  \[307] ,
  \new_D<27> ,
  \[308] ,
  \new_D<28> ,
  \[309] ,
  \new_D<21> ,
  \new_D<22> ,
  \new_D<23> ,
  \new_D<24> ,
  \[310] ,
  \[500] ,
  \new_D<20> ,
  \[311] ,
  \[501] ,
  \new_D<39> ,
  \[312] ,
  \[502] ,
  \[313] ,
  \[503] ,
  \[314] ,
  \[504] ,
  \[315] ,
  \[505] ,
  \new_D<35> ,
  \[316] ,
  \[506] ,
  \new_D<36> ,
  \[317] ,
  \[507] ,
  \new_D<37> ,
  \[318] ,
  \[508] ,
  \new_D<38> ,
  \[319] ,
  \[509] ,
  \new_D<31> ,
  \new_D<32> ,
  \new_D<33> ,
  \new_D<34> ,
  \[320] ,
  \[510] ,
  \new_D<30> ,
  \[321] ,
  \[511] ,
  \new_D<49> ,
  \[322] ,
  \[512] ,
  \[323] ,
  \[513] ,
  \[324] ,
  \[514] ,
  \[325] ,
  \[515] ,
  \new_D<45> ,
  \[326] ,
  \[516] ,
  \new_C<1> ,
  \new_D<46> ,
  \[327] ,
  \[517] ,
  \new_C<2> ,
  \new_D<47> ,
  \[328] ,
  \[518] ,
  \new_C<3> ,
  \new_D<48> ,
  \[329] ,
  \[519] ,
  \new_C<4> ,
  \new_D<41> ,
  \new_D<42> ,
  \new_D<43> ,
  \new_D<44> ,
  \new_C<0> ,
  \new_C<9> ,
  \[330] ,
  \[520] ,
  \new_C<59> ,
  \new_D<40> ,
  \[331] ,
  \[521] ,
  \main/$PLUS_5_1/sum<3>5.1 ,
  \[332] ,
  \[522] ,
  \new_C<5> ,
  \[333] ,
  \[523] ,
  \new_C<6> ,
  \[334] ,
  \[524] ,
  \new_C<55> ,
  \new_C<7> ,
  \[335] ,
  \[525] ,
  \new_C<56> ,
  \new_C<8> ,
  \[336] ,
  \[526] ,
  \new_C<57> ,
  \[337] ,
  \[527] ,
  \new_C<58> ,
  \[338] ,
  \[528] ,
  \new_C<51> ,
  \[339] ,
  \[529] ,
  \new_C<52> ,
  \new_C<53> ,
  \new_C<54> ,
  \new_C<50> ,
  \[340] ,
  \[530] ,
  \new_C<69> ,
  \[341] ,
  \[531] ,
  \[342] ,
  \[532] ,
  \[343] ,
  \[533] ,
  \[344] ,
  \[534] ,
  \new_C<65> ,
  \[345] ,
  \[535] ,
  \new_C<66> ,
  \[346] ,
  \[536] ,
  \new_C<67> ,
  \[347] ,
  \[537] ,
  \new_C<68> ,
  \[348] ,
  \[538] ,
  \new_C<61> ,
  \[349] ,
  \[539] ,
  \new_C<62> ,
  \new_C<63> ,
  \new_C<64> ,
  \new_C<60> ,
  \[350] ,
  \[540] ,
  \new_C<79> ,
  \[351] ,
  \[541] ,
  \[352] ,
  \[542] ,
  \[353] ,
  \[543] ,
  \[354] ,
  \[544] ,
  \new_C<75> ,
  \[355] ,
  \[545] ,
  \new_C<76> ,
  \[356] ,
  \[546] ,
  \new_C<77> ,
  \[357] ,
  \[547] ,
  \new_C<78> ,
  \[358] ,
  \[548] ,
  \new_C<71> ,
  \[359] ,
  \[549] ,
  \new_C<72> ,
  \new_C<73> ,
  \new_C<74> ,
  \new_C<70> ,
  \[360] ,
  \[550] ,
  \new_C<89> ,
  \[361] ,
  \[551] ,
  \[362] ,
  \[552] ,
  \[363] ,
  \[553] ,
  \[364] ,
  \[554] ,
  \new_C<85> ,
  \[365] ,
  \[555] ,
  \new_C<86> ,
  \[366] ,
  \[556] ,
  \new_C<87> ,
  \[367] ,
  \[557] ,
  \new_C<88> ,
  \[368] ,
  \[558] ,
  \new_C<81> ,
  \[369] ,
  \[559] ,
  \new_C<82> ,
  \new_C<83> ,
  \new_C<84> ,
  \new_C<80> ,
  \[370] ,
  \[560] ,
  \[371] ,
  \[561] ,
  \new_D<99> ,
  \[372] ,
  \[562] ,
  \[373] ,
  \[563] ,
  \[374] ,
  \[564] ,
  \[375] ,
  \[565] ,
  \$$COND1<0>8.1 ,
  \new_D<95> ,
  \[376] ,
  \[566] ,
  \new_D<96> ,
  \[377] ,
  \[567] ,
  \new_D<97> ;
assign
  \[378]  = \C<43> ,
  \[568]  = \new_D<76> ,
  \new_D<98>  = (~\$$COND0<0>5.1  & (\C<98>  & (\D<98>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<98>  & (\D<98>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<98>  & (~\D<98>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<98>  & (~\D<98>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<98>  & (\D<98>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<98>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<98>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<197>  & (\encrypt<0>  & \start<0> )) | (\key<205>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[379]  = \C<35> ,
  \[569]  = \new_D<75> ,
  \new_D<91>  = (~\$$COND0<0>5.1  & (\C<91>  & (\D<91>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<91>  & (\D<91>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<91>  & (~\D<91>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<91>  & (~\D<91>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<91>  & (\D<91>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<91>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<91>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<253>  & (\encrypt<0>  & \start<0> )) | (\key<198>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<92>  = (~\$$COND0<0>5.1  & (\C<92>  & (\D<92>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<92>  & (\D<92>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<92>  & (~\D<92>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<92>  & (~\D<92>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<92>  & (\D<92>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<92>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<92>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<245>  & (\encrypt<0>  & \start<0> )) | (\key<253>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<93>  = (~\$$COND0<0>5.1  & (\C<93>  & (\D<93>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<93>  & (\D<93>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<93>  & (~\D<93>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<93>  & (~\D<93>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<93>  & (\D<93>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<93>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<93>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<237>  & (\encrypt<0>  & \start<0> )) | (\key<245>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<94>  = (~\$$COND0<0>5.1  & (\C<94>  & (\D<94>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<94>  & (\D<94>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<94>  & (~\D<94>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<94>  & (~\D<94>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<94>  & (\D<94>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<94>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<94>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<229>  & (\encrypt<0>  & \start<0> )) | (\key<237>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<130>  = \[290] ,
  \KSi<131>  = \[289] ,
  \KSi<132>  = \[288] ,
  \[380]  = \C<53> ,
  \[570]  = \new_D<74> ,
  \KSi<133>  = \[287] ,
  \new_D<90>  = (~\$$COND0<0>5.1  & (\C<90>  & (\D<90>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<90>  & (\D<90>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<90>  & (~\D<90>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<90>  & (~\D<90>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<90>  & (\D<90>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<90>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<90>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<198>  & (\encrypt<0>  & \start<0> )) | (\key<206>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[381]  = \C<31> ,
  \[571]  = \new_D<73> ,
  \KSi<134>  = \[286] ,
  \[382]  = \C<39> ,
  \[572]  = \new_D<72> ,
  \KSi<135>  = \[285] ,
  \[383]  = \C<46> ,
  \[573]  = \new_D<71> ,
  \KSi<136>  = \[284] ,
  \[384]  = \C<50> ,
  \[574]  = \new_D<70> ,
  \KSi<137>  = \[283] ,
  \[385]  = \C<37> ,
  \[575]  = \new_D<69> ,
  \KSi<138>  = \[282] ,
  \[386]  = \C<48> ,
  \[576]  = \new_D<68> ,
  \KSi<139>  = \[281] ,
  \[387]  = \C<33> ,
  \[577]  = \new_D<67> ,
  \main/$MINUS_4_1/sum<3>8.1  = (~\main/$MINUS_4_1/c<0>8.4  & ~\count<3> ) | (\main/$MINUS_4_1/c<0>8.4  & \count<3> ),
  \[388]  = \C<42> ,
  \[578]  = \new_D<66> ,
  \new_C<111>  = (~\$$COND0<0>5.1  & (~\D<111>  & (\C<111>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<111>  & (~\C<111>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<111>  & (\C<111>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<111>  & (~\C<111>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<111>  & (\C<111>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<111>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<111>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<56>  & (\encrypt<0>  & \start<0> )) | (\key<227>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[389]  = \C<55> ,
  \[579]  = \new_D<65> ,
  \new_C<110>  = (~\$$COND0<0>5.1  & (~\D<110>  & (\C<110>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<110>  & (~\C<110>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<110>  & (\C<110>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<110>  & (~\C<110>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<110>  & (\C<110>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<110>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<110>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<227>  & (\encrypt<0>  & \start<0> )) | (\key<235>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[390]  = \C<30> ,
  \[580]  = \new_D<64> ,
  \[391]  = \C<32> ,
  \[581]  = \new_D<63> ,
  \[392]  = \C<28> ,
  \[582]  = \new_D<62> ,
  \[393]  = \C<51> ,
  \[583]  = \new_D<61> ,
  \[394]  = \C<38> ,
  \[584]  = \new_D<60> ,
  \[395]  = \C<44> ,
  \[585]  = \new_D<59> ,
  \[396]  = \C<41> ,
  \[586]  = \new_D<58> ,
  \[397]  = \C<1> ,
  \[587]  = \new_D<57> ,
  \[398]  = \C<12> ,
  \[588]  = \new_D<56> ,
  \[399]  = \C<19> ,
  \[589]  = \new_D<55> ,
  \[590]  = \new_D<54> ,
  \[591]  = \new_D<53> ,
  \[592]  = \new_D<52> ,
  \[593]  = \new_D<51> ,
  \[594]  = \new_D<50> ,
  \[595]  = \new_D<49> ,
  \[596]  = \new_D<48> ,
  \[597]  = \new_D<47> ,
  \[598]  = \new_D<46> ,
  \[599]  = \new_D<45> ,
  \KSi<100>  = \[320] ,
  \KSi<101>  = \[319] ,
  \KSi<102>  = \[318] ,
  \KSi<103>  = \[317] ,
  \KSi<104>  = \[316] ,
  \new_D<59>  = (~\$$COND0<0>5.1  & (\C<59>  & (\D<59>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<59>  & (\D<59>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<59>  & (~\D<59>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<59>  & (~\D<59>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<59>  & (\D<59>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<59>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<59>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<158>  & (\encrypt<0>  & \start<0> )) | (\key<166>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<105>  = \[315] ,
  \main/$PLUS_5_1/sum<2>5.1  = (~\main/$PLUS_5_1/c<0>5.3  & \count<2> ) | (\main/$PLUS_5_1/c<0>5.3  & ~\count<2> ),
  \KSi<106>  = \[314] ,
  \KSi<107>  = \[313] ,
  \KSi<108>  = \[312] ,
  \new_D<55>  = (~\$$COND0<0>5.1  & (\C<55>  & (\D<55>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<55>  & (\D<55>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<55>  & (~\D<55>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<55>  & (~\D<55>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<55>  & (\D<55>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<55>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<55>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<190>  & (\encrypt<0>  & \start<0> )) | (\key<67>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<109>  = \[311] ,
  \new_D<56>  = (~\$$COND0<0>5.1  & (\C<56>  & (\D<56>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<56>  & (\D<56>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<56>  & (~\D<56>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<56>  & (~\D<56>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<56>  & (\D<56>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<56>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<56>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<182>  & (\encrypt<0>  & \start<0> )) | (\key<190>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<57>  = (~\$$COND0<0>5.1  & (\C<57>  & (\D<57>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<57>  & (\D<57>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<57>  & (~\D<57>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<57>  & (~\D<57>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<57>  & (\D<57>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<57>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<57>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<174>  & (\encrypt<0>  & \start<0> )) | (\key<182>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<58>  = (~\$$COND0<0>5.1  & (\C<58>  & (\D<58>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<58>  & (\D<58>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<58>  & (~\D<58>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<58>  & (~\D<58>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<58>  & (\D<58>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<58>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<58>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<166>  & (\encrypt<0>  & \start<0> )) | (\key<174>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<51>  = (~\$$COND0<0>5.1  & (\C<51>  & (\D<51>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<51>  & (\D<51>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<51>  & (~\D<51>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<51>  & (~\D<51>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<51>  & (\D<51>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<51>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<51>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<91>  & (\encrypt<0>  & \start<0> )) | (\key<68>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<52>  = (~\$$COND0<0>5.1  & (\C<52>  & (\D<52>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<52>  & (\D<52>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<52>  & (~\D<52>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<52>  & (~\D<52>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<52>  & (\D<52>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<52>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<52>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<83>  & (\encrypt<0>  & \start<0> )) | (\key<91>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<53>  = (~\$$COND0<0>5.1  & (\C<53>  & (\D<53>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<53>  & (\D<53>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<53>  & (~\D<53>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<53>  & (~\D<53>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<53>  & (\D<53>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<53>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<53>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<75>  & (\encrypt<0>  & \start<0> )) | (\key<83>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<54>  = (~\$$COND0<0>5.1  & (\C<54>  & (\D<54>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<54>  & (\D<54>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<54>  & (~\D<54>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<54>  & (~\D<54>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<54>  & (\D<54>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<54>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<54>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<67>  & (\encrypt<0>  & \start<0> )) | (\key<75>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<50>  = (~\$$COND0<0>5.1  & (\C<50>  & (\D<50>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<50>  & (\D<50>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<50>  & (~\D<50>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<50>  & (~\D<50>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<50>  & (\D<50>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<50>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<50>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<68>  & (\encrypt<0>  & \start<0> )) | (\key<76>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<69>  = (~\$$COND0<0>5.1  & (\C<69>  & (\D<69>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<69>  & (\D<69>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<69>  & (~\D<69>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<69>  & (~\D<69>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<69>  & (\D<69>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<69>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<69>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<141>  & (\encrypt<0>  & \start<0> )) | (\key<149>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<65>  = (~\$$COND0<0>5.1  & (\C<65>  & (\D<65>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<65>  & (\D<65>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<65>  & (~\D<65>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<65>  & (~\D<65>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<65>  & (\D<65>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<65>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<65>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<173>  & (\encrypt<0>  & \start<0> )) | (\key<181>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<66>  = (~\$$COND0<0>5.1  & (\C<66>  & (\D<66>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<66>  & (\D<66>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<66>  & (~\D<66>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<66>  & (~\D<66>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<66>  & (\D<66>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<66>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<66>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<165>  & (\encrypt<0>  & \start<0> )) | (\key<173>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<67>  = (~\$$COND0<0>5.1  & (\C<67>  & (\D<67>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<67>  & (\D<67>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<67>  & (~\D<67>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<67>  & (~\D<67>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<67>  & (\D<67>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<67>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<67>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<157>  & (\encrypt<0>  & \start<0> )) | (\key<165>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<68>  = (~\$$COND0<0>5.1  & (\C<68>  & (\D<68>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<68>  & (\D<68>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<68>  & (~\D<68>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<68>  & (~\D<68>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<68>  & (\D<68>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<68>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<68>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<149>  & (\encrypt<0>  & \start<0> )) | (\key<157>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<61>  = (~\$$COND0<0>5.1  & (\C<61>  & (\D<61>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<61>  & (\D<61>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<61>  & (~\D<61>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<61>  & (~\D<61>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<61>  & (\D<61>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<61>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<61>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<142>  & (\encrypt<0>  & \start<0> )) | (\key<150>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<62>  = (~\$$COND0<0>5.1  & (\C<62>  & (\D<62>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<62>  & (\D<62>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<62>  & (~\D<62>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<62>  & (~\D<62>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<62>  & (\D<62>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<62>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<62>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<134>  & (\encrypt<0>  & \start<0> )) | (\key<142>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<63>  = (~\$$COND0<0>5.1  & (\C<63>  & (\D<63>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<63>  & (\D<63>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<63>  & (~\D<63>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<63>  & (~\D<63>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<63>  & (\D<63>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<63>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<63>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<189>  & (\encrypt<0>  & \start<0> )) | (\key<134>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<64>  = (~\$$COND0<0>5.1  & (\C<64>  & (\D<64>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<64>  & (\D<64>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<64>  & (~\D<64>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<64>  & (~\D<64>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<64>  & (\D<64>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<64>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<64>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<181>  & (\encrypt<0>  & \start<0> )) | (\key<189>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<60>  = (~\$$COND0<0>5.1  & (\C<60>  & (\D<60>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<60>  & (\D<60>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<60>  & (~\D<60>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<60>  & (~\D<60>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<60>  & (\D<60>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<60>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<60>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<150>  & (\encrypt<0>  & \start<0> )) | (\key<158>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<79>  = (~\$$COND0<0>5.1  & (\C<79>  & (\D<79>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<79>  & (\D<79>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<79>  & (~\D<79>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<79>  & (~\D<79>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<79>  & (\D<79>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<79>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<79>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<155>  & (\encrypt<0>  & \start<0> )) | (\key<132>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<75>  = (~\$$COND0<0>5.1  & (\C<75>  & (\D<75>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<75>  & (\D<75>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<75>  & (~\D<75>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<75>  & (~\D<75>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<75>  & (\D<75>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<75>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<75>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<156>  & (\encrypt<0>  & \start<0> )) | (\key<164>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<76>  = (~\$$COND0<0>5.1  & (\C<76>  & (\D<76>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<76>  & (\D<76>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<76>  & (~\D<76>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<76>  & (~\D<76>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<76>  & (\D<76>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<76>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<76>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<148>  & (\encrypt<0>  & \start<0> )) | (\key<156>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<77>  = (~\$$COND0<0>5.1  & (\C<77>  & (\D<77>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<77>  & (\D<77>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<77>  & (~\D<77>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<77>  & (~\D<77>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<77>  & (\D<77>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<77>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<77>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<140>  & (\encrypt<0>  & \start<0> )) | (\key<148>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<78>  = (~\$$COND0<0>5.1  & (\C<78>  & (\D<78>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<78>  & (\D<78>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<78>  & (~\D<78>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<78>  & (~\D<78>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<78>  & (\D<78>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<78>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<78>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<132>  & (\encrypt<0>  & \start<0> )) | (\key<140>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<71>  = (~\$$COND0<0>5.1  & (\C<71>  & (\D<71>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<71>  & (\D<71>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<71>  & (~\D<71>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<71>  & (~\D<71>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<71>  & (\D<71>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<71>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<71>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<188>  & (\encrypt<0>  & \start<0> )) | (\key<133>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<72>  = (~\$$COND0<0>5.1  & (\C<72>  & (\D<72>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<72>  & (\D<72>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<72>  & (~\D<72>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<72>  & (~\D<72>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<72>  & (\D<72>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<72>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<72>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<180>  & (\encrypt<0>  & \start<0> )) | (\key<188>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<73>  = (~\$$COND0<0>5.1  & (\C<73>  & (\D<73>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<73>  & (\D<73>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<73>  & (~\D<73>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<73>  & (~\D<73>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<73>  & (\D<73>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<73>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<73>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<172>  & (\encrypt<0>  & \start<0> )) | (\key<180>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<74>  = (~\$$COND0<0>5.1  & (\C<74>  & (\D<74>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<74>  & (\D<74>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<74>  & (~\D<74>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<74>  & (~\D<74>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<74>  & (\D<74>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<74>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<74>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<164>  & (\encrypt<0>  & \start<0> )) | (\key<172>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<190>  = \[230] ,
  \KSi<191>  = \[229] ,
  \new_D<70>  = (~\$$COND0<0>5.1  & (\C<70>  & (\D<70>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<70>  & (\D<70>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<70>  & (~\D<70>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<70>  & (~\D<70>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<70>  & (\D<70>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<70>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<70>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<133>  & (\encrypt<0>  & \start<0> )) | (\key<141>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<111>  = (~\$$COND0<0>5.1  & (\C<111>  & (\D<111>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<111>  & (\D<111>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<111>  & (~\D<111>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<111>  & (~\D<111>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<111>  & (\D<111>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<111>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<111>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<62>  & (\encrypt<0>  & \start<0> )) | (\key<195>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<89>  = (~\$$COND0<0>5.1  & (\C<89>  & (\D<89>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<89>  & (\D<89>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<89>  & (~\D<89>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<89>  & (~\D<89>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<89>  & (\D<89>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<89>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<89>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<206>  & (\encrypt<0>  & \start<0> )) | (\key<214>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<85>  = (~\$$COND0<0>5.1  & (\C<85>  & (\D<85>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<85>  & (\D<85>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<85>  & (~\D<85>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<85>  & (~\D<85>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<85>  & (\D<85>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<85>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<85>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<238>  & (\encrypt<0>  & \start<0> )) | (\key<246>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<110>  = (~\$$COND0<0>5.1  & (\C<110>  & (\D<110>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<110>  & (\D<110>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<110>  & (~\D<110>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<110>  & (~\D<110>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<110>  & (\D<110>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<110>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<110>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<195>  & (\encrypt<0>  & \start<0> )) | (\key<203>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<86>  = (~\$$COND0<0>5.1  & (\C<86>  & (\D<86>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<86>  & (\D<86>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<86>  & (~\D<86>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<86>  & (~\D<86>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<86>  & (\D<86>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<86>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<86>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<230>  & (\encrypt<0>  & \start<0> )) | (\key<238>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<87>  = (~\$$COND0<0>5.1  & (\C<87>  & (\D<87>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<87>  & (\D<87>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<87>  & (~\D<87>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<87>  & (~\D<87>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<87>  & (\D<87>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<87>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<87>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<222>  & (\encrypt<0>  & \start<0> )) | (\key<230>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<88>  = (~\$$COND0<0>5.1  & (\C<88>  & (\D<88>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<88>  & (\D<88>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<88>  & (~\D<88>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<88>  & (~\D<88>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<88>  & (\D<88>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<88>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<88>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<214>  & (\encrypt<0>  & \start<0> )) | (\key<222>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<81>  = (~\$$COND0<0>5.1  & (\C<81>  & (\D<81>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<81>  & (\D<81>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<81>  & (~\D<81>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<81>  & (~\D<81>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<81>  & (\D<81>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<81>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<81>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<139>  & (\encrypt<0>  & \start<0> )) | (\key<147>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<82>  = (~\$$COND0<0>5.1  & (\C<82>  & (\D<82>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<82>  & (\D<82>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<82>  & (~\D<82>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<82>  & (~\D<82>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<82>  & (\D<82>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<82>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<82>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<131>  & (\encrypt<0>  & \start<0> )) | (\key<139>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<83>  = (~\$$COND0<0>5.1  & (\C<83>  & (\D<83>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<83>  & (\D<83>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<83>  & (~\D<83>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<83>  & (~\D<83>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<83>  & (\D<83>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<83>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<83>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<254>  & (\encrypt<0>  & \start<0> )) | (\key<131>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<84>  = (~\$$COND0<0>5.1  & (\C<84>  & (\D<84>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<84>  & (\D<84>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<84>  & (~\D<84>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<84>  & (~\D<84>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<84>  & (\D<84>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<84>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<84>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<246>  & (\encrypt<0>  & \start<0> )) | (\key<254>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<109>  = (~\$$COND0<0>5.1  & (~\D<109>  & (\C<109>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<109>  & (~\C<109>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<109>  & (\C<109>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<109>  & (~\C<109>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<109>  & (\C<109>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<109>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<109>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<235>  & (\encrypt<0>  & \start<0> )) | (\key<243>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<80>  = (~\$$COND0<0>5.1  & (\C<80>  & (\D<80>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<80>  & (\D<80>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<80>  & (~\D<80>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<80>  & (~\D<80>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<80>  & (\D<80>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<80>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<80>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<147>  & (\encrypt<0>  & \start<0> )) | (\key<155>  & (~\encrypt<0>  & \start<0> ))))))))),
  \main/$MINUS_4_1/sum<2>8.1  = (~\main/$MINUS_4_1/c<0>8.3  & ~\count<2> ) | (\main/$MINUS_4_1/c<0>8.3  & \count<2> ),
  \new_C<106>  = (~\$$COND0<0>5.1  & (~\D<106>  & (\C<106>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<106>  & (~\C<106>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<106>  & (\C<106>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<106>  & (~\C<106>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<106>  & (\C<106>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<106>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<106>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<194>  & (\encrypt<0>  & \start<0> )) | (\key<202>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<105>  = (~\$$COND0<0>5.1  & (~\D<105>  & (\C<105>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<105>  & (~\C<105>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<105>  & (\C<105>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<105>  & (~\C<105>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<105>  & (\C<105>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<105>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<105>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<202>  & (\encrypt<0>  & \start<0> )) | (\key<210>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<108>  = (~\$$COND0<0>5.1  & (~\D<108>  & (\C<108>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<108>  & (~\C<108>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<108>  & (\C<108>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<108>  & (~\C<108>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<108>  & (\C<108>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<108>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<108>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<243>  & (\encrypt<0>  & \start<0> )) | (\key<251>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<107>  = (~\$$COND0<0>5.1  & (~\D<107>  & (\C<107>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<107>  & (~\C<107>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<107>  & (\C<107>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<107>  & (~\C<107>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<107>  & (\C<107>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<107>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<107>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<251>  & (\encrypt<0>  & \start<0> )) | (\key<194>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<102>  = (~\$$COND0<0>5.1  & (~\D<102>  & (\C<102>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<102>  & (~\C<102>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<102>  & (\C<102>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<102>  & (~\C<102>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<102>  & (\C<102>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<102>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<102>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<226>  & (\encrypt<0>  & \start<0> )) | (\key<234>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<101>  = (~\$$COND0<0>5.1  & (~\D<101>  & (\C<101>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<101>  & (~\C<101>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<101>  & (\C<101>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<101>  & (~\C<101>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<101>  & (\C<101>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<101>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<101>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<234>  & (\encrypt<0>  & \start<0> )) | (\key<242>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<104>  = (~\$$COND0<0>5.1  & (~\D<104>  & (\C<104>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<104>  & (~\C<104>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<104>  & (\C<104>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<104>  & (~\C<104>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<104>  & (\C<104>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<104>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<104>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<210>  & (\encrypt<0>  & \start<0> )) | (\key<218>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<103>  = (~\$$COND0<0>5.1  & (~\D<103>  & (\C<103>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<103>  & (~\C<103>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<103>  & (\C<103>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<103>  & (~\C<103>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<103>  & (\C<103>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<103>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<103>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<218>  & (\encrypt<0>  & \start<0> )) | (\key<226>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<100>  = (~\$$COND0<0>5.1  & (~\D<100>  & (\C<100>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<100>  & (~\C<100>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<100>  & (\C<100>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<100>  & (~\C<100>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<100>  & (\C<100>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<100>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<100>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<242>  & (\encrypt<0>  & \start<0> )) | (\key<250>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[400]  = \C<26> ,
  \[401]  = \C<6> ,
  \[402]  = \C<15> ,
  \[403]  = \C<7> ,
  \[404]  = \C<25> ,
  \[405]  = \C<3> ,
  \[406]  = \C<11> ,
  \[407]  = \C<18> ,
  \[408]  = \C<22> ,
  \[409]  = \C<9> ,
  \KSi<160>  = \[260] ,
  \KSi<161>  = \[259] ,
  \KSi<162>  = \[258] ,
  \[410]  = \C<20> ,
  \[600]  = \new_D<44> ,
  \KSi<163>  = \[257] ,
  \[411]  = \C<5> ,
  \[601]  = \new_D<43> ,
  \KSi<164>  = \[256] ,
  \[412]  = \C<14> ,
  \[602]  = \new_D<42> ,
  \KSi<165>  = \[255] ,
  \[413]  = \C<27> ,
  \[603]  = \new_D<41> ,
  \KSi<166>  = \[254] ,
  \[224]  = (\main/$PLUS_5_1/sum<3>5.1  & (\encrypt<0>  & ~\start<0> )) | ((\main/$MINUS_4_1/sum<3>8.1  & (~\encrypt<0>  & ~\start<0> )) | (~\encrypt<0>  & \start<0> )),
  \[414]  = \C<2> ,
  \[604]  = \new_D<40> ,
  \KSi<167>  = \[253] ,
  \[225]  = (\main/$PLUS_5_1/sum<2>5.1  & (\encrypt<0>  & ~\start<0> )) | ((\main/$MINUS_4_1/sum<2>8.1  & (~\encrypt<0>  & ~\start<0> )) | (~\encrypt<0>  & \start<0> )),
  \[415]  = \C<4> ,
  \[605]  = \new_D<39> ,
  \KSi<168>  = \[252] ,
  \[226]  = (\main/$PLUS_5_1/sum<1>5.1  & (\encrypt<0>  & ~\start<0> )) | ((\main/$MINUS_4_1/sum<1>8.1  & (~\encrypt<0>  & ~\start<0> )) | (~\encrypt<0>  & \start<0> )),
  \[416]  = \C<0> ,
  \[606]  = \new_D<38> ,
  \KSi<169>  = \[251] ,
  \[227]  = (\main/$PLUS_5_1/sum<0>5.1  & (\encrypt<0>  & ~\start<0> )) | ((\main/$MINUS_4_1/sum<0>8.1  & (~\encrypt<0>  & ~\start<0> )) | (~\encrypt<0>  & \start<0> )),
  \[417]  = \C<23> ,
  \[607]  = \new_D<37> ,
  \[228]  = (~\count<3>  & (~\count<2>  & (~\count<1>  & (~\count<0>  & (~\encrypt<0>  & ~\start<0> ))))) | (\count<3>  & (\count<2>  & (\count<1>  & (\count<0>  & (\encrypt<0>  & ~\start<0> ))))),
  \[418]  = \C<10> ,
  \[608]  = \new_D<36> ,
  \[229]  = \D<87> ,
  \[419]  = \C<16> ,
  \[609]  = \new_D<35> ,
  \KSi<150>  = \[270] ,
  \KSi<151>  = \[269] ,
  \KSi<152>  = \[268] ,
  \[230]  = \D<84> ,
  \[420]  = \C<13> ,
  \[610]  = \new_D<34> ,
  \KSi<153>  = \[267] ,
  \[231]  = \D<91> ,
  \[421]  = \new_C<111> ,
  \[611]  = \new_D<33> ,
  \KSi<154>  = \[266] ,
  \[232]  = \D<105> ,
  \[422]  = \new_C<110> ,
  \[612]  = \new_D<32> ,
  \KSi<155>  = \[265] ,
  \[233]  = \D<87> ,
  \[423]  = \new_C<109> ,
  \[613]  = \new_D<31> ,
  \KSi<156>  = \[264] ,
  \[234]  = \D<101> ,
  \[424]  = \new_C<108> ,
  \[614]  = \new_D<30> ,
  \KSi<157>  = \[263] ,
  \[235]  = \D<108> ,
  \[425]  = \new_C<107> ,
  \[615]  = \new_D<29> ,
  \KSi<158>  = \[262] ,
  \[236]  = \D<89> ,
  \[426]  = \new_C<106> ,
  \[616]  = \new_D<28> ,
  \KSi<159>  = \[261] ,
  \new_D<1>  = (~\$$COND0<0>5.1  & (\C<1>  & (\D<1>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<1>  & (\D<1>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<1>  & (~\D<1>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<1>  & (~\D<1>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<1>  & (\D<1>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<1>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<1>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<46>  & (\encrypt<0>  & \start<0> )) | (\key<54>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[237]  = \D<111> ,
  \[427]  = \new_C<105> ,
  \[617]  = \new_D<27> ,
  \new_D<2>  = (~\$$COND0<0>5.1  & (\C<2>  & (\D<2>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<2>  & (\D<2>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<2>  & (~\D<2>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<2>  & (~\D<2>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<2>  & (\D<2>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<2>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<2>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<38>  & (\encrypt<0>  & \start<0> )) | (\key<46>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[238]  = \D<94> ,
  \[428]  = \new_C<104> ,
  \[618]  = \new_D<26> ,
  \new_D<3>  = (~\$$COND0<0>5.1  & (\C<3>  & (\D<3>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<3>  & (\D<3>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<3>  & (~\D<3>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<3>  & (~\D<3>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<3>  & (\D<3>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<3>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<3>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<30>  & (\encrypt<0>  & \start<0> )) | (\key<38>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[239]  = \D<104> ,
  \[429]  = \new_C<103> ,
  \[619]  = \new_D<25> ,
  \KSi<0>  = \[420] ,
  \new_D<4>  = (~\$$COND0<0>5.1  & (\C<4>  & (\D<4>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<4>  & (\D<4>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<4>  & (~\D<4>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<4>  & (~\D<4>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<4>  & (\D<4>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<4>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<4>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<22>  & (\encrypt<0>  & \start<0> )) | (\key<30>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<1>  = \[419] ,
  \KSi<2>  = \[418] ,
  \KSi<3>  = \[417] ,
  \KSi<4>  = \[416] ,
  \KSi<180>  = \[240] ,
  \new_D<0>  = (~\$$COND0<0>5.1  & (\C<0>  & (\D<0>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<0>  & (\D<0>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<0>  & (~\D<0>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<0>  & (~\D<0>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<0>  & (\D<0>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<0>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<0>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<54>  & (\encrypt<0>  & \start<0> )) | (\key<62>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<5>  = \[415] ,
  \KSi<181>  = \[239] ,
  \new_D<9>  = (~\$$COND0<0>5.1  & (\C<9>  & (\D<9>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<9>  & (\D<9>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<9>  & (~\D<9>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<9>  & (~\D<9>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<9>  & (\D<9>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<9>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<9>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<45>  & (\encrypt<0>  & \start<0> )) | (\key<53>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<6>  = \[414] ,
  \KSi<182>  = \[238] ,
  \[240]  = \D<99> ,
  \[430]  = \new_C<102> ,
  \[620]  = \new_D<24> ,
  \KSi<7>  = \[413] ,
  \KSi<183>  = \[237] ,
  \[241]  = \D<103> ,
  \[431]  = \new_C<101> ,
  \[621]  = \new_D<23> ,
  \KSi<8>  = \[412] ,
  \KSi<184>  = \[236] ,
  \[242]  = \D<88> ,
  \[432]  = \new_C<100> ,
  \[622]  = \new_D<22> ,
  \KSi<9>  = \[411] ,
  \KSi<185>  = \[235] ,
  \new_D<5>  = (~\$$COND0<0>5.1  & (\C<5>  & (\D<5>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<5>  & (\D<5>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<5>  & (~\D<5>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<5>  & (~\D<5>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<5>  & (\D<5>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<5>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<5>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<14>  & (\encrypt<0>  & \start<0> )) | (\key<22>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[243]  = \D<100> ,
  \[433]  = \new_C<99> ,
  \[623]  = \new_D<21> ,
  \KSi<186>  = \[234] ,
  \new_D<6>  = (~\$$COND0<0>5.1  & (\C<6>  & (\D<6>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<6>  & (\D<6>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<6>  & (~\D<6>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<6>  & (~\D<6>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<6>  & (\D<6>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<6>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<6>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<6>  & (\encrypt<0>  & \start<0> )) | (\key<14>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[244]  = \D<106> ,
  \[434]  = \new_C<98> ,
  \[624]  = \new_D<20> ,
  \main/$PLUS_5_1/sum<1>5.1  = (~\count<0>  & \count<1> ) | (\count<0>  & ~\count<1> ),
  \KSi<187>  = \[233] ,
  \new_D<7>  = (~\$$COND0<0>5.1  & (\C<7>  & (\D<7>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<7>  & (\D<7>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<7>  & (~\D<7>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<7>  & (~\D<7>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<7>  & (\D<7>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<7>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<7>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<61>  & (\encrypt<0>  & \start<0> )) | (\key<6>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[245]  = \D<95> ,
  \[435]  = \new_C<97> ,
  \[625]  = \new_D<19> ,
  \KSi<188>  = \[232] ,
  \new_D<8>  = (~\$$COND0<0>5.1  & (\C<8>  & (\D<8>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<8>  & (\D<8>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<8>  & (~\D<8>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<8>  & (~\D<8>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<8>  & (\D<8>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<8>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<8>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<53>  & (\encrypt<0>  & \start<0> )) | (\key<61>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[246]  = \D<85> ,
  \[436]  = \new_C<96> ,
  \[626]  = \new_D<18> ,
  \KSi<189>  = \[231] ,
  \[247]  = \D<110> ,
  \[437]  = \new_C<95> ,
  \[627]  = \new_D<17> ,
  \[248]  = \D<102> ,
  \[438]  = \new_C<94> ,
  \[628]  = \new_D<16> ,
  \[249]  = \D<92> ,
  \[439]  = \new_C<93> ,
  \[629]  = \new_D<15> ,
  \KSi<170>  = \[250] ,
  \KSi<171>  = \[249] ,
  \KSi<172>  = \[248] ,
  \[250]  = \D<86> ,
  \[440]  = \new_C<92> ,
  \[630]  = \new_D<14> ,
  \KSi<173>  = \[247] ,
  \[251]  = \D<107> ,
  \[441]  = \new_C<91> ,
  \[631]  = \new_D<13> ,
  \KSi<174>  = \[246] ,
  \[252]  = \D<104> ,
  \[442]  = \new_C<90> ,
  \[632]  = \new_D<12> ,
  \KSi<175>  = \[245] ,
  \[253]  = \D<59> ,
  \[443]  = \new_C<89> ,
  \[633]  = \new_D<11> ,
  \KSi<176>  = \[244] ,
  \[254]  = \D<56> ,
  \[444]  = \new_C<88> ,
  \[634]  = \new_D<10> ,
  \KSi<177>  = \[243] ,
  \[255]  = \D<63> ,
  \[445]  = \new_C<87> ,
  \[635]  = \new_D<9> ,
  \KSi<178>  = \[242] ,
  \[256]  = \D<77> ,
  \[446]  = \new_C<86> ,
  \[636]  = \new_D<8> ,
  \KSi<179>  = \[241] ,
  \[257]  = \D<69> ,
  \[447]  = \new_C<85> ,
  \[637]  = \new_D<7> ,
  \[258]  = \D<73> ,
  \[448]  = \new_C<84> ,
  \[638]  = \new_D<6> ,
  \[259]  = \D<80> ,
  \[449]  = \new_C<83> ,
  \[639]  = \new_D<5> ,
  \new_D<109>  = (~\$$COND0<0>5.1  & (\C<109>  & (\D<109>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<109>  & (\D<109>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<109>  & (~\D<109>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<109>  & (~\D<109>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<109>  & (\D<109>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<109>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<109>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<203>  & (\encrypt<0>  & \start<0> )) | (\key<211>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<106>  = (~\$$COND0<0>5.1  & (\C<106>  & (\D<106>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<106>  & (\D<106>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<106>  & (~\D<106>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<106>  & (~\D<106>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<106>  & (\D<106>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<106>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<106>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<196>  & (\encrypt<0>  & \start<0> )) | (\key<204>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<105>  = (~\$$COND0<0>5.1  & (\C<105>  & (\D<105>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<105>  & (\D<105>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<105>  & (~\D<105>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<105>  & (~\D<105>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<105>  & (\D<105>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<105>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<105>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<204>  & (\encrypt<0>  & \start<0> )) | (\key<212>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<108>  = (~\$$COND0<0>5.1  & (\C<108>  & (\D<108>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<108>  & (\D<108>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<108>  & (~\D<108>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<108>  & (~\D<108>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<108>  & (\D<108>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<108>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<108>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<211>  & (\encrypt<0>  & \start<0> )) | (\key<219>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<107>  = (~\$$COND0<0>5.1  & (\C<107>  & (\D<107>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<107>  & (\D<107>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<107>  & (~\D<107>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<107>  & (~\D<107>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<107>  & (\D<107>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<107>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<107>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<219>  & (\encrypt<0>  & \start<0> )) | (\key<196>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[260]  = \D<61> ,
  \[450]  = \new_C<82> ,
  \[640]  = \new_D<4> ,
  \new_D<102>  = (~\$$COND0<0>5.1  & (\C<102>  & (\D<102>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<102>  & (\D<102>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<102>  & (~\D<102>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<102>  & (~\D<102>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<102>  & (\D<102>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<102>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<102>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<228>  & (\encrypt<0>  & \start<0> )) | (\key<172>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[261]  = \D<83> ,
  \[451]  = \new_C<81> ,
  \[641]  = \new_D<3> ,
  \new_D<101>  = (~\$$COND0<0>5.1  & (\C<101>  & (\D<101>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<101>  & (\D<101>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<101>  & (~\D<101>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<101>  & (~\D<101>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<101>  & (\D<101>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<101>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<101>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<172>  & (\encrypt<0>  & \start<0> )) | (\key<244>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[262]  = \D<66> ,
  \[452]  = \new_C<80> ,
  \[642]  = \new_D<2> ,
  \new_D<104>  = (~\$$COND0<0>5.1  & (\C<104>  & (\D<104>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<104>  & (\D<104>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<104>  & (~\D<104>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<104>  & (~\D<104>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<104>  & (\D<104>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<104>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<104>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<212>  & (\encrypt<0>  & \start<0> )) | (\key<220>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[263]  = \D<76> ,
  \[453]  = \new_C<79> ,
  \[643]  = \new_D<1> ,
  \new_D<103>  = (~\$$COND0<0>5.1  & (\C<103>  & (\D<103>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<103>  & (\D<103>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<103>  & (~\D<103>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<103>  & (~\D<103>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<103>  & (\D<103>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<103>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<103>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<220>  & (\encrypt<0>  & \start<0> )) | (\key<228>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[264]  = \D<71> ,
  \[454]  = \new_C<78> ,
  \[644]  = \new_D<0> ,
  \[265]  = \D<75> ,
  \[455]  = \new_C<77> ,
  \[266]  = \D<60> ,
  \[456]  = \new_C<76> ,
  \new_D<100>  = (~\$$COND0<0>5.1  & (\C<100>  & (\D<100>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<100>  & (\D<100>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<100>  & (~\D<100>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<100>  & (~\D<100>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<100>  & (\D<100>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<100>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<100>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<244>  & (\encrypt<0>  & \start<0> )) | (\key<252>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[267]  = \D<70> ,
  \[457]  = \new_C<75> ,
  \[268]  = \D<78> ,
  \[458]  = \new_C<74> ,
  \[269]  = \D<67> ,
  \[459]  = \new_C<73> ,
  \[270]  = \D<57> ,
  \[460]  = \new_C<72> ,
  \new_C<19>  = (~\$$COND0<0>5.1  & (~\D<19>  & (\C<19>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<19>  & (~\C<19>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<19>  & (\C<19>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<19>  & (~\C<19>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<19>  & (\C<19>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<19>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<19>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<26>  & (\encrypt<0>  & \start<0> )) | (\key<34>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[271]  = \D<82> ,
  \[461]  = \new_C<71> ,
  \[272]  = \D<74> ,
  \main/$PLUS_5_1/c<0>5.3  = \count<0>  & \count<1> ,
  \main/$PLUS_5_1/c<0>5.4  = \main/$PLUS_5_1/c<0>5.3  & \count<2> ,
  \[462]  = \new_C<70> ,
  \[273]  = \D<64> ,
  \[463]  = \new_C<69> ,
  \[274]  = \D<58> ,
  \[464]  = \new_C<68> ,
  \new_C<15>  = (~\$$COND0<0>5.1  & (~\D<15>  & (\C<15>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<15>  & (~\C<15>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<15>  & (\C<15>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<15>  & (~\C<15>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<15>  & (\C<15>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<15>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<15>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<58>  & (\encrypt<0>  & \start<0> )) | (\key<1>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[275]  = \D<79> ,
  \[465]  = \new_C<67> ,
  \new_C<16>  = (~\$$COND0<0>5.1  & (~\D<16>  & (\C<16>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<16>  & (~\C<16>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<16>  & (\C<16>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<16>  & (~\C<16>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<16>  & (\C<16>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<16>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<16>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<50>  & (\encrypt<0>  & \start<0> )) | (\key<58>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[276]  = \D<68> ,
  \[466]  = \new_C<66> ,
  \new_C<17>  = (~\$$COND0<0>5.1  & (~\D<17>  & (\C<17>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<17>  & (~\C<17>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<17>  & (\C<17>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<17>  & (~\C<17>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<17>  & (\C<17>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<17>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<17>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<42>  & (\encrypt<0>  & \start<0> )) | (\key<50>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[277]  = \D<31> ,
  \[467]  = \new_C<65> ,
  \new_C<18>  = (~\$$COND0<0>5.1  & (~\D<18>  & (\C<18>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<18>  & (~\C<18>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<18>  & (\C<18>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<18>  & (~\C<18>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<18>  & (\C<18>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<18>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<18>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<34>  & (\encrypt<0>  & \start<0> )) | (\key<42>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[278]  = \D<28> ,
  \[468]  = \new_C<64> ,
  \new_C<11>  = (~\$$COND0<0>5.1  & (~\D<11>  & (\C<11>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<11>  & (~\C<11>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<11>  & (\C<11>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<11>  & (~\C<11>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<11>  & (\C<11>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<11>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<11>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<25>  & (\encrypt<0>  & \start<0> )) | (\key<33>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[279]  = \D<35> ,
  \[469]  = \new_C<63> ,
  \new_C<12>  = (~\$$COND0<0>5.1  & (~\D<12>  & (\C<12>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<12>  & (~\C<12>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<12>  & (\C<12>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<12>  & (~\C<12>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<12>  & (\C<12>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<12>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<12>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<17>  & (\encrypt<0>  & \start<0> )) | (\key<25>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<13>  = (~\$$COND0<0>5.1  & (~\D<13>  & (\C<13>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<13>  & (~\C<13>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<13>  & (\C<13>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<13>  & (~\C<13>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<13>  & (\C<13>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<13>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<13>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<9>  & (\encrypt<0>  & \start<0> )) | (\key<17>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<14>  = (~\$$COND0<0>5.1  & (~\D<14>  & (\C<14>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<14>  & (~\C<14>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<14>  & (\C<14>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<14>  & (~\C<14>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<14>  & (\C<14>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<14>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<14>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<1>  & (\encrypt<0>  & \start<0> )) | (\key<9>  & (~\encrypt<0>  & \start<0> ))))))))),
  \$$COND0<0>5.1  = (~\count<3>  & (~\count<2>  & (~\count<1>  & ~\count<0> ))) | ((~\count<3>  & (\count<2>  & (\count<1>  & \count<0> ))) | (\count<3>  & (\count<2>  & (\count<1>  & ~\count<0> )))),
  \new_C<10>  = (~\$$COND0<0>5.1  & (~\D<10>  & (\C<10>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<10>  & (~\C<10>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<10>  & (\C<10>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<10>  & (~\C<10>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<10>  & (\C<10>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<10>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<10>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<33>  & (\encrypt<0>  & \start<0> )) | (\key<41>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[280]  = \D<49> ,
  \[470]  = \new_C<62> ,
  \new_C<29>  = (~\$$COND0<0>5.1  & (~\D<29>  & (\C<29>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<29>  & (~\C<29>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<29>  & (\C<29>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<29>  & (~\C<29>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<29>  & (\C<29>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<29>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<29>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<104>  & (\encrypt<0>  & \start<0> )) | (\key<112>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[281]  = \D<31> ,
  \[471]  = \new_C<61> ,
  \[282]  = \D<45> ,
  \[472]  = \new_C<60> ,
  \[283]  = \D<52> ,
  \[473]  = \new_C<59> ,
  \[284]  = \D<33> ,
  \[474]  = \new_C<58> ,
  \new_C<25>  = (~\$$COND0<0>5.1  & (~\D<25>  & (\C<25>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<25>  & (~\C<25>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<25>  & (\C<25>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<25>  & (~\C<25>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<25>  & (\C<25>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<25>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<25>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<43>  & (\encrypt<0>  & \start<0> )) | (\key<51>  & (~\encrypt<0>  & \start<0> ))))))))),
  \main/$MINUS_4_1/sum<1>8.1  = (~\count<0>  & ~\count<1> ) | (\count<0>  & \count<1> ),
  \[285]  = \D<55> ,
  \[475]  = \new_C<57> ,
  \new_C<26>  = (~\$$COND0<0>5.1  & (~\D<26>  & (\C<26>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<26>  & (~\C<26>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<26>  & (\C<26>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<26>  & (~\C<26>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<26>  & (\C<26>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<26>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<26>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<35>  & (\encrypt<0>  & \start<0> )) | (\key<43>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[286]  = \D<38> ,
  \[476]  = \new_C<56> ,
  \new_C<27>  = (~\$$COND0<0>5.1  & (~\D<27>  & (\C<27>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<27>  & (~\C<27>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<27>  & (\C<27>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<27>  & (~\C<27>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<27>  & (\C<27>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<27>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<27>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<120>  & (\encrypt<0>  & \start<0> )) | (\key<35>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[287]  = \D<48> ,
  \[477]  = \new_C<55> ,
  \new_C<28>  = (~\$$COND0<0>5.1  & (~\D<28>  & (\C<28>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<28>  & (~\C<28>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<28>  & (\C<28>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<28>  & (~\C<28>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<28>  & (\C<28>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<28>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<28>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<112>  & (\encrypt<0>  & \start<0> )) | (\key<120>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[288]  = \D<43> ,
  \[478]  = \new_C<54> ,
  \new_C<21>  = (~\$$COND0<0>5.1  & (~\D<21>  & (\C<21>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<21>  & (~\C<21>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<21>  & (\C<21>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<21>  & (~\C<21>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<21>  & (\C<21>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<21>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<21>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<10>  & (\encrypt<0>  & \start<0> )) | (\key<18>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[289]  = \D<47> ,
  \[479]  = \new_C<53> ,
  \new_C<22>  = (~\$$COND0<0>5.1  & (~\D<22>  & (\C<22>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<22>  & (~\C<22>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<22>  & (\C<22>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<22>  & (~\C<22>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<22>  & (\C<22>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<22>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<22>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<2>  & (\encrypt<0>  & \start<0> )) | (\key<10>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<23>  = (~\$$COND0<0>5.1  & (~\D<23>  & (\C<23>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<23>  & (~\C<23>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<23>  & (\C<23>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<23>  & (~\C<23>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<23>  & (\C<23>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<23>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<23>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<59>  & (\encrypt<0>  & \start<0> )) | (\key<2>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<24>  = (~\$$COND0<0>5.1  & (~\D<24>  & (\C<24>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<24>  & (~\C<24>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<24>  & (\C<24>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<24>  & (~\C<24>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<24>  & (\C<24>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<24>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<24>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<51>  & (\encrypt<0>  & \start<0> )) | (\key<59>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<20>  = (~\$$COND0<0>5.1  & (~\D<20>  & (\C<20>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<20>  & (~\C<20>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<20>  & (\C<20>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<20>  & (~\C<20>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<20>  & (\C<20>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<20>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<20>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<18>  & (\encrypt<0>  & \start<0> )) | (\key<26>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[290]  = \D<32> ,
  \[480]  = \new_C<52> ,
  \new_C<39>  = (~\$$COND0<0>5.1  & (~\D<39>  & (\C<39>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<39>  & (~\C<39>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<39>  & (\C<39>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<39>  & (~\C<39>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<39>  & (\C<39>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<39>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<39>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<89>  & (\encrypt<0>  & \start<0> )) | (\key<97>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[291]  = \D<44> ,
  \[481]  = \new_C<51> ,
  \[292]  = \D<50> ,
  \[482]  = \new_C<50> ,
  \[293]  = \D<39> ,
  \[483]  = \new_C<49> ,
  \[294]  = \D<29> ,
  \[484]  = \new_C<48> ,
  \new_C<35>  = (~\$$COND0<0>5.1  & (~\D<35>  & (\C<35>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<35>  & (~\C<35>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<35>  & (\C<35>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<35>  & (~\C<35>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<35>  & (\C<35>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<35>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<35>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<121>  & (\encrypt<0>  & \start<0> )) | (\key<64>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[295]  = \D<54> ,
  \[485]  = \new_C<47> ,
  \new_C<36>  = (~\$$COND0<0>5.1  & (~\D<36>  & (\C<36>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<36>  & (~\C<36>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<36>  & (\C<36>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<36>  & (~\C<36>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<36>  & (\C<36>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<36>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<36>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<113>  & (\encrypt<0>  & \start<0> )) | (\key<121>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[296]  = \D<46> ,
  \[486]  = \new_C<46> ,
  \new_C<37>  = (~\$$COND0<0>5.1  & (~\D<37>  & (\C<37>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<37>  & (~\C<37>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<37>  & (\C<37>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<37>  & (~\C<37>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<37>  & (\C<37>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<37>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<37>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<105>  & (\encrypt<0>  & \start<0> )) | (\key<113>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[297]  = \D<36> ,
  \[487]  = \new_C<45> ,
  \new_C<38>  = (~\$$COND0<0>5.1  & (~\D<38>  & (\C<38>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<38>  & (~\C<38>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<38>  & (\C<38>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<38>  & (~\C<38>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<38>  & (\C<38>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<38>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<38>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<97>  & (\encrypt<0>  & \start<0> )) | (\key<105>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[298]  = \D<30> ,
  \[488]  = \new_C<44> ,
  \new_C<31>  = (~\$$COND0<0>5.1  & (~\D<31>  & (\C<31>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<31>  & (~\C<31>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<31>  & (\C<31>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<31>  & (~\C<31>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<31>  & (\C<31>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<31>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<31>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<88>  & (\encrypt<0>  & \start<0> )) | (\key<96>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[299]  = \D<51> ,
  \[489]  = \new_C<43> ,
  \new_C<32>  = (~\$$COND0<0>5.1  & (~\D<32>  & (\C<32>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<32>  & (~\C<32>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<32>  & (\C<32>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<32>  & (~\C<32>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<32>  & (\C<32>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<32>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<32>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<80>  & (\encrypt<0>  & \start<0> )) | (\key<88>  & (~\encrypt<0>  & \start<0> ))))))))),
  \main/$PLUS_5_1/sum<0>5.1  = ~\count<0> ,
  \new_C<33>  = (~\$$COND0<0>5.1  & (~\D<33>  & (\C<33>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<33>  & (~\C<33>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<33>  & (\C<33>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<33>  & (~\C<33>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<33>  & (\C<33>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<33>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<33>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<72>  & (\encrypt<0>  & \start<0> )) | (\key<80>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<34>  = (~\$$COND0<0>5.1  & (~\D<34>  & (\C<34>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<34>  & (~\C<34>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<34>  & (\C<34>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<34>  & (~\C<34>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<34>  & (\C<34>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<34>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<34>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<64>  & (\encrypt<0>  & \start<0> )) | (\key<72>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<30>  = (~\$$COND0<0>5.1  & (~\D<30>  & (\C<30>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<30>  & (~\C<30>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<30>  & (\C<30>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<30>  & (~\C<30>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<30>  & (\C<30>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<30>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<30>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<96>  & (\encrypt<0>  & \start<0> )) | (\key<104>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[490]  = \new_C<42> ,
  \new_C<49>  = (~\$$COND0<0>5.1  & (~\D<49>  & (\C<49>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<49>  & (~\C<49>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<49>  & (\C<49>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<49>  & (~\C<49>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<49>  & (\C<49>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<49>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<49>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<74>  & (\encrypt<0>  & \start<0> )) | (\key<82>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[491]  = \new_C<41> ,
  \[492]  = \new_C<40> ,
  \[493]  = \new_C<39> ,
  \[494]  = \new_C<38> ,
  \new_C<45>  = (~\$$COND0<0>5.1  & (~\D<45>  & (\C<45>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<45>  & (~\C<45>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<45>  & (\C<45>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<45>  & (~\C<45>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<45>  & (\C<45>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<45>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<45>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<106>  & (\encrypt<0>  & \start<0> )) | (\key<114>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[495]  = \new_C<37> ,
  \new_C<46>  = (~\$$COND0<0>5.1  & (~\D<46>  & (\C<46>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<46>  & (~\C<46>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<46>  & (\C<46>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<46>  & (~\C<46>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<46>  & (\C<46>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<46>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<46>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<98>  & (\encrypt<0>  & \start<0> )) | (\key<106>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[496]  = \new_C<36> ,
  \new_C<47>  = (~\$$COND0<0>5.1  & (~\D<47>  & (\C<47>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<47>  & (~\C<47>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<47>  & (\C<47>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<47>  & (~\C<47>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<47>  & (\C<47>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<47>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<47>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<90>  & (\encrypt<0>  & \start<0> )) | (\key<98>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[497]  = \new_C<35> ,
  \new_C<48>  = (~\$$COND0<0>5.1  & (~\D<48>  & (\C<48>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<48>  & (~\C<48>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<48>  & (\C<48>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<48>  & (~\C<48>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<48>  & (\C<48>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<48>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<48>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<82>  & (\encrypt<0>  & \start<0> )) | (\key<90>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[498]  = \new_C<34> ,
  \new_C<41>  = (~\$$COND0<0>5.1  & (~\D<41>  & (\C<41>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<41>  & (~\C<41>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<41>  & (\C<41>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<41>  & (~\C<41>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<41>  & (\C<41>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<41>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<41>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<73>  & (\encrypt<0>  & \start<0> )) | (\key<81>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[499]  = \new_C<33> ,
  \new_C<42>  = (~\$$COND0<0>5.1  & (~\D<42>  & (\C<42>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<42>  & (~\C<42>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<42>  & (\C<42>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<42>  & (~\C<42>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<42>  & (\C<42>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<42>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<42>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<65>  & (\encrypt<0>  & \start<0> )) | (\key<73>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_count<0>  = \[227] ,
  \new_C<43>  = (~\$$COND0<0>5.1  & (~\D<43>  & (\C<43>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<43>  & (~\C<43>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<43>  & (\C<43>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<43>  & (~\C<43>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<43>  & (\C<43>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<43>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<43>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<122>  & (\encrypt<0>  & \start<0> )) | (\key<65>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<44>  = (~\$$COND0<0>5.1  & (~\D<44>  & (\C<44>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<44>  & (~\C<44>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<44>  & (\C<44>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<44>  & (~\C<44>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<44>  & (\C<44>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<44>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<44>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<114>  & (\encrypt<0>  & \start<0> )) | (\key<122>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_count<3>  = \[224] ,
  \new_count<1>  = \[226] ,
  \new_C<40>  = (~\$$COND0<0>5.1  & (~\D<40>  & (\C<40>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<40>  & (~\C<40>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<40>  & (\C<40>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<40>  & (~\C<40>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<40>  & (\C<40>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<40>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<40>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<81>  & (\encrypt<0>  & \start<0> )) | (\key<89>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_count<2>  = \[225] ,
  \KSi<12>  = \[408] ,
  \KSi<11>  = \[409] ,
  \KSi<14>  = \[406] ,
  \KSi<13>  = \[407] ,
  \KSi<10>  = \[410] ,
  \KSi<19>  = \[401] ,
  \KSi<16>  = \[404] ,
  \KSi<15>  = \[405] ,
  \KSi<18>  = \[402] ,
  \KSi<17>  = \[403] ,
  \KSi<22>  = \[398] ,
  \KSi<21>  = \[399] ,
  \KSi<24>  = \[396] ,
  \KSi<23>  = \[397] ,
  \KSi<20>  = \[400] ,
  \KSi<29>  = \[391] ,
  \KSi<26>  = \[394] ,
  \KSi<25>  = \[395] ,
  \KSi<28>  = \[392] ,
  \KSi<27>  = \[393] ,
  \KSi<32>  = \[388] ,
  \KSi<31>  = \[389] ,
  \KSi<34>  = \[386] ,
  \KSi<33>  = \[387] ,
  \KSi<30>  = \[390] ,
  \KSi<39>  = \[381] ,
  \KSi<36>  = \[384] ,
  \KSi<35>  = \[385] ,
  \KSi<38>  = \[382] ,
  \KSi<37>  = \[383] ,
  \KSi<42>  = \[378] ,
  \KSi<41>  = \[379] ,
  \KSi<44>  = \[376] ,
  \KSi<43>  = \[377] ,
  \main/$MINUS_4_1/sum<0>8.1  = ~\count<0> ,
  \new_C<99>  = (~\$$COND0<0>5.1  & (~\D<99>  & (\C<99>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<99>  & (~\C<99>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<99>  & (\C<99>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<99>  & (~\C<99>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<99>  & (\C<99>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<99>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<99>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<250>  & (\encrypt<0>  & \start<0> )) | (\key<193>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<19>  = (~\$$COND0<0>5.1  & (\C<19>  & (\D<19>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<19>  & (\D<19>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<19>  & (~\D<19>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<19>  & (~\D<19>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<19>  & (\D<19>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<19>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<19>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<28>  & (\encrypt<0>  & \start<0> )) | (\key<36>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<40>  = \[380] ,
  \new_C<95>  = (~\$$COND0<0>5.1  & (~\D<95>  & (\C<95>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<95>  & (~\C<95>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<95>  & (\C<95>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<95>  & (~\C<95>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<95>  & (\C<95>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<95>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<95>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<217>  & (\encrypt<0>  & \start<0> )) | (\key<225>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<49>  = \[371] ,
  \new_C<96>  = (~\$$COND0<0>5.1  & (~\D<96>  & (\C<96>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<96>  & (~\C<96>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<96>  & (\C<96>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<96>  & (~\C<96>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<96>  & (\C<96>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<96>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<96>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<209>  & (\encrypt<0>  & \start<0> )) | (\key<217>  & (~\encrypt<0>  & \start<0> ))))))))),
  \main/$MINUS_4_1/c<0>8.3  = \count<0>  | \count<1> ,
  \main/$MINUS_4_1/c<0>8.4  = \main/$MINUS_4_1/c<0>8.3  | \count<2> ,
  \new_D<15>  = (~\$$COND0<0>5.1  & (\C<15>  & (\D<15>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<15>  & (\D<15>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<15>  & (~\D<15>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<15>  & (~\D<15>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<15>  & (\D<15>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<15>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<15>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<60>  & (\encrypt<0>  & \start<0> )) | (\key<5>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<97>  = (~\$$COND0<0>5.1  & (~\D<97>  & (\C<97>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<97>  & (~\C<97>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<97>  & (\C<97>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<97>  & (~\C<97>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<97>  & (\C<97>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<97>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<97>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<201>  & (\encrypt<0>  & \start<0> )) | (\key<209>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<16>  = (~\$$COND0<0>5.1  & (\C<16>  & (\D<16>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<16>  & (\D<16>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<16>  & (~\D<16>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<16>  & (~\D<16>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<16>  & (\D<16>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<16>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<16>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<52>  & (\encrypt<0>  & \start<0> )) | (\key<60>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<98>  = (~\$$COND0<0>5.1  & (~\D<98>  & (\C<98>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<98>  & (~\C<98>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<98>  & (\C<98>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<98>  & (~\C<98>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<98>  & (\C<98>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<98>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<98>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<193>  & (\encrypt<0>  & \start<0> )) | (\key<201>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<17>  = (~\$$COND0<0>5.1  & (\C<17>  & (\D<17>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<17>  & (\D<17>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<17>  & (~\D<17>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<17>  & (~\D<17>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<17>  & (\D<17>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<17>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<17>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<44>  & (\encrypt<0>  & \start<0> )) | (\key<52>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<46>  = \[374] ,
  \new_C<91>  = (~\$$COND0<0>5.1  & (~\D<91>  & (\C<91>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<91>  & (~\C<91>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<91>  & (\C<91>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<91>  & (~\C<91>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<91>  & (\C<91>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<91>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<91>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<249>  & (\encrypt<0>  & \start<0> )) | (\key<192>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<18>  = (~\$$COND0<0>5.1  & (\C<18>  & (\D<18>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<18>  & (\D<18>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<18>  & (~\D<18>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<18>  & (~\D<18>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<18>  & (\D<18>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<18>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<18>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<36>  & (\encrypt<0>  & \start<0> )) | (\key<44>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<45>  = \[375] ,
  \new_C<92>  = (~\$$COND0<0>5.1  & (~\D<92>  & (\C<92>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<92>  & (~\C<92>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<92>  & (\C<92>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<92>  & (~\C<92>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<92>  & (\C<92>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<92>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<92>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<241>  & (\encrypt<0>  & \start<0> )) | (\key<249>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<11>  = (~\$$COND0<0>5.1  & (\C<11>  & (\D<11>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<11>  & (\D<11>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<11>  & (~\D<11>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<11>  & (~\D<11>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<11>  & (\D<11>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<11>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<11>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<29>  & (\encrypt<0>  & \start<0> )) | (\key<37>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<48>  = \[372] ,
  \new_C<93>  = (~\$$COND0<0>5.1  & (~\D<93>  & (\C<93>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<93>  & (~\C<93>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<93>  & (\C<93>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<93>  & (~\C<93>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<93>  & (\C<93>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<93>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<93>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<233>  & (\encrypt<0>  & \start<0> )) | (\key<241>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<12>  = (~\$$COND0<0>5.1  & (\C<12>  & (\D<12>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<12>  & (\D<12>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<12>  & (~\D<12>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<12>  & (~\D<12>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<12>  & (\D<12>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<12>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<12>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<21>  & (\encrypt<0>  & \start<0> )) | (\key<29>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<47>  = \[373] ,
  \new_C<94>  = (~\$$COND0<0>5.1  & (~\D<94>  & (\C<94>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<94>  & (~\C<94>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<94>  & (\C<94>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<94>  & (~\C<94>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<94>  & (\C<94>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<94>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<94>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<225>  & (\encrypt<0>  & \start<0> )) | (\key<233>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<13>  = (~\$$COND0<0>5.1  & (\C<13>  & (\D<13>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<13>  & (\D<13>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<13>  & (~\D<13>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<13>  & (~\D<13>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<13>  & (\D<13>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<13>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<13>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<13>  & (\encrypt<0>  & \start<0> )) | (\key<21>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<52>  = \[368] ,
  \new_D<14>  = (~\$$COND0<0>5.1  & (\C<14>  & (\D<14>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<14>  & (\D<14>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<14>  & (~\D<14>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<14>  & (~\D<14>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<14>  & (\D<14>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<14>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<14>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<5>  & (\encrypt<0>  & \start<0> )) | (\key<13>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<51>  = \[369] ,
  \KSi<54>  = \[366] ,
  \KSi<53>  = \[367] ,
  \new_C<90>  = (~\$$COND0<0>5.1  & (~\D<90>  & (\C<90>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<90>  & (~\C<90>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<90>  & (\C<90>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<90>  & (~\C<90>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<90>  & (\C<90>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<90>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<90>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<192>  & (\encrypt<0>  & \start<0> )) | (\key<200>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[300]  = \D<40> ,
  \new_D<10>  = (~\$$COND0<0>5.1  & (\C<10>  & (\D<10>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<10>  & (\D<10>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<10>  & (~\D<10>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<10>  & (~\D<10>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<10>  & (\D<10>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<10>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<10>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<37>  & (\encrypt<0>  & \start<0> )) | (\key<45>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[301]  = \D<3> ,
  \new_D<29>  = (~\$$COND0<0>5.1  & (\C<29>  & (\D<29>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<29>  & (\D<29>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<29>  & (~\D<29>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<29>  & (~\D<29>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<29>  & (\D<29>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<29>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<29>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<110>  & (\encrypt<0>  & \start<0> )) | (\key<118>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[302]  = \D<0> ,
  \KSi<50>  = \[370] ,
  \[303]  = \D<7> ,
  \[304]  = \D<21> ,
  \[305]  = \D<13> ,
  \KSi<59>  = \[361] ,
  \new_D<25>  = (~\$$COND0<0>5.1  & (\C<25>  & (\D<25>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<25>  & (\D<25>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<25>  & (~\D<25>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<25>  & (~\D<25>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<25>  & (\D<25>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<25>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<25>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<11>  & (\encrypt<0>  & \start<0> )) | (\key<19>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[306]  = \D<17> ,
  \new_D<26>  = (~\$$COND0<0>5.1  & (\C<26>  & (\D<26>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<26>  & (\D<26>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<26>  & (~\D<26>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<26>  & (~\D<26>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<26>  & (\D<26>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<26>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<26>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<3>  & (\encrypt<0>  & \start<0> )) | (\key<11>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[307]  = \D<24> ,
  \new_D<27>  = (~\$$COND0<0>5.1  & (\C<27>  & (\D<27>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<27>  & (\D<27>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<27>  & (~\D<27>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<27>  & (~\D<27>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<27>  & (\D<27>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<27>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<27>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<126>  & (\encrypt<0>  & \start<0> )) | (\key<3>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[308]  = \D<5> ,
  \KSi<56>  = \[364] ,
  \new_D<28>  = (~\$$COND0<0>5.1  & (\C<28>  & (\D<28>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<28>  & (\D<28>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<28>  & (~\D<28>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<28>  & (~\D<28>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<28>  & (\D<28>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<28>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<28>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<118>  & (\encrypt<0>  & \start<0> )) | (\key<126>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[309]  = \D<27> ,
  \KSi<55>  = \[365] ,
  \new_D<21>  = (~\$$COND0<0>5.1  & (\C<21>  & (\D<21>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<21>  & (\D<21>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<21>  & (~\D<21>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<21>  & (~\D<21>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<21>  & (\D<21>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<21>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<21>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<12>  & (\encrypt<0>  & \start<0> )) | (\key<20>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<58>  = \[362] ,
  \new_D<22>  = (~\$$COND0<0>5.1  & (\C<22>  & (\D<22>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<22>  & (\D<22>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<22>  & (~\D<22>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<22>  & (~\D<22>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<22>  & (\D<22>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<22>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<22>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<4>  & (\encrypt<0>  & \start<0> )) | (\key<12>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<57>  = \[363] ,
  \new_D<23>  = (~\$$COND0<0>5.1  & (\C<23>  & (\D<23>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<23>  & (\D<23>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<23>  & (~\D<23>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<23>  & (~\D<23>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<23>  & (\D<23>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<23>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<23>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<27>  & (\encrypt<0>  & \start<0> )) | (\key<4>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<62>  = \[358] ,
  \new_D<24>  = (~\$$COND0<0>5.1  & (\C<24>  & (\D<24>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<24>  & (\D<24>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<24>  & (~\D<24>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<24>  & (~\D<24>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<24>  & (\D<24>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<24>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<24>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<19>  & (\encrypt<0>  & \start<0> )) | (\key<27>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<61>  = \[359] ,
  \KSi<64>  = \[356] ,
  \KSi<63>  = \[357] ,
  \[310]  = \D<10> ,
  \[500]  = \new_C<32> ,
  \new_D<20>  = (~\$$COND0<0>5.1  & (\C<20>  & (\D<20>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<20>  & (\D<20>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<20>  & (~\D<20>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<20>  & (~\D<20>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<20>  & (\D<20>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<20>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<20>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<20>  & (\encrypt<0>  & \start<0> )) | (\key<28>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[311]  = \D<20> ,
  \[501]  = \new_C<31> ,
  \new_D<39>  = (~\$$COND0<0>5.1  & (\C<39>  & (\D<39>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<39>  & (\D<39>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<39>  & (~\D<39>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<39>  & (~\D<39>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<39>  & (\D<39>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<39>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<39>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<93>  & (\encrypt<0>  & \start<0> )) | (\key<101>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[312]  = \D<15> ,
  \KSi<60>  = \[360] ,
  \[502]  = \new_C<30> ,
  \[313]  = \D<19> ,
  \[503]  = \new_C<29> ,
  \[314]  = \D<4> ,
  \[504]  = \new_C<28> ,
  \[315]  = \D<16> ,
  \KSi<69>  = \[351] ,
  \[505]  = \new_C<27> ,
  \new_D<35>  = (~\$$COND0<0>5.1  & (\C<35>  & (\D<35>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<35>  & (\D<35>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<35>  & (~\D<35>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<35>  & (~\D<35>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<35>  & (\D<35>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<35>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<35>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<125>  & (\encrypt<0>  & \start<0> )) | (\key<70>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[316]  = \D<22> ,
  \[506]  = \new_C<26> ,
  \new_D<36>  = (~\$$COND0<0>5.1  & (\C<36>  & (\D<36>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<36>  & (\D<36>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<36>  & (~\D<36>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<36>  & (~\D<36>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<36>  & (\D<36>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<36>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<36>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<117>  & (\encrypt<0>  & \start<0> )) | (\key<125>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[317]  = \D<11> ,
  \[507]  = \new_C<25> ,
  \new_D<37>  = (~\$$COND0<0>5.1  & (\C<37>  & (\D<37>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<37>  & (\D<37>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<37>  & (~\D<37>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<37>  & (~\D<37>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<37>  & (\D<37>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<37>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<37>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<109>  & (\encrypt<0>  & \start<0> )) | (\key<117>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[318]  = \D<1> ,
  \KSi<66>  = \[354] ,
  \[508]  = \new_C<24> ,
  \data_ready<0>  = \[228] ,
  \new_D<38>  = (~\$$COND0<0>5.1  & (\C<38>  & (\D<38>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<38>  & (\D<38>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<38>  & (~\D<38>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<38>  & (~\D<38>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<38>  & (\D<38>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<38>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<38>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<101>  & (\encrypt<0>  & \start<0> )) | (\key<109>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[319]  = \D<26> ,
  \KSi<65>  = \[355] ,
  \[509]  = \new_C<23> ,
  \new_D<31>  = (~\$$COND0<0>5.1  & (\C<31>  & (\D<31>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<31>  & (\D<31>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<31>  & (~\D<31>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<31>  & (~\D<31>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<31>  & (\D<31>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<31>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<31>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<94>  & (\encrypt<0>  & \start<0> )) | (\key<102>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<68>  = \[352] ,
  \new_D<32>  = (~\$$COND0<0>5.1  & (\C<32>  & (\D<32>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<32>  & (\D<32>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<32>  & (~\D<32>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<32>  & (~\D<32>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<32>  & (\D<32>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<32>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<32>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<86>  & (\encrypt<0>  & \start<0> )) | (\key<94>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<67>  = \[353] ,
  \new_D<33>  = (~\$$COND0<0>5.1  & (\C<33>  & (\D<33>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<33>  & (\D<33>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<33>  & (~\D<33>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<33>  & (~\D<33>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<33>  & (\D<33>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<33>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<33>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<78>  & (\encrypt<0>  & \start<0> )) | (\key<86>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<72>  = \[348] ,
  \new_D<34>  = (~\$$COND0<0>5.1  & (\C<34>  & (\D<34>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<34>  & (\D<34>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<34>  & (~\D<34>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<34>  & (~\D<34>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<34>  & (\D<34>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<34>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<34>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<70>  & (\encrypt<0>  & \start<0> )) | (\key<78>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<71>  = \[349] ,
  \KSi<74>  = \[346] ,
  \KSi<73>  = \[347] ,
  \[320]  = \D<18> ,
  \[510]  = \new_C<22> ,
  \new_D<30>  = (~\$$COND0<0>5.1  & (\C<30>  & (\D<30>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<30>  & (\D<30>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<30>  & (~\D<30>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<30>  & (~\D<30>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<30>  & (\D<30>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<30>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<30>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<102>  & (\encrypt<0>  & \start<0> )) | (\key<110>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[321]  = \D<8> ,
  \[511]  = \new_C<21> ,
  \new_D<49>  = (~\$$COND0<0>5.1  & (\C<49>  & (\D<49>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<49>  & (\D<49>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<49>  & (~\D<49>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<49>  & (~\D<49>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<49>  & (\D<49>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<49>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<49>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<76>  & (\encrypt<0>  & \start<0> )) | (\key<84>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[322]  = \D<2> ,
  \KSi<70>  = \[350] ,
  \[512]  = \new_C<20> ,
  \[323]  = \D<23> ,
  \[513]  = \new_C<19> ,
  \[324]  = \D<12> ,
  \[514]  = \new_C<18> ,
  \[325]  = \C<85> ,
  \KSi<79>  = \[341] ,
  \[515]  = \new_C<17> ,
  \new_D<45>  = (~\$$COND0<0>5.1  & (\C<45>  & (\D<45>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<45>  & (\D<45>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<45>  & (~\D<45>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<45>  & (~\D<45>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<45>  & (\D<45>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<45>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<45>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<44>  & (\encrypt<0>  & \start<0> )) | (\key<116>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[326]  = \C<96> ,
  \[516]  = \new_C<16> ,
  \new_C<1>  = (~\$$COND0<0>5.1  & (~\D<1>  & (\C<1>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<1>  & (~\C<1>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<1>  & (\C<1>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<1>  & (~\C<1>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<1>  & (\C<1>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<1>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<1>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<40>  & (\encrypt<0>  & \start<0> )) | (\key<48>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<46>  = (~\$$COND0<0>5.1  & (\C<46>  & (\D<46>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<46>  & (\D<46>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<46>  & (~\D<46>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<46>  & (~\D<46>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<46>  & (\D<46>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<46>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<46>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<100>  & (\encrypt<0>  & \start<0> )) | (\key<44>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[327]  = \C<103> ,
  \[517]  = \new_C<15> ,
  \new_C<2>  = (~\$$COND0<0>5.1  & (~\D<2>  & (\C<2>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<2>  & (~\C<2>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<2>  & (\C<2>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<2>  & (~\C<2>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<2>  & (\C<2>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<2>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<2>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<32>  & (\encrypt<0>  & \start<0> )) | (\key<40>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<47>  = (~\$$COND0<0>5.1  & (\C<47>  & (\D<47>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<47>  & (\D<47>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<47>  & (~\D<47>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<47>  & (~\D<47>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<47>  & (\D<47>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<47>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<47>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<92>  & (\encrypt<0>  & \start<0> )) | (\key<100>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[328]  = \C<110> ,
  \KSi<76>  = \[344] ,
  \[518]  = \new_C<14> ,
  \new_C<3>  = (~\$$COND0<0>5.1  & (~\D<3>  & (\C<3>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<3>  & (~\C<3>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<3>  & (\C<3>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<3>  & (~\C<3>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<3>  & (\C<3>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<3>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<3>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<24>  & (\encrypt<0>  & \start<0> )) | (\key<32>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<48>  = (~\$$COND0<0>5.1  & (\C<48>  & (\D<48>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<48>  & (\D<48>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<48>  & (~\D<48>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<48>  & (~\D<48>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<48>  & (\D<48>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<48>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<48>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<84>  & (\encrypt<0>  & \start<0> )) | (\key<92>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[329]  = \C<90> ,
  \KSi<75>  = \[345] ,
  \[519]  = \new_C<13> ,
  \new_C<4>  = (~\$$COND0<0>5.1  & (~\D<4>  & (\C<4>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<4>  & (~\C<4>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<4>  & (\C<4>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<4>  & (~\C<4>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<4>  & (\C<4>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<4>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<4>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<16>  & (\encrypt<0>  & \start<0> )) | (\key<24>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<41>  = (~\$$COND0<0>5.1  & (\C<41>  & (\D<41>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<41>  & (\D<41>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<41>  & (~\D<41>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<41>  & (~\D<41>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<41>  & (\D<41>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<41>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<41>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<77>  & (\encrypt<0>  & \start<0> )) | (\key<85>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<78>  = \[342] ,
  \new_D<42>  = (~\$$COND0<0>5.1  & (\C<42>  & (\D<42>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<42>  & (\D<42>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<42>  & (~\D<42>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<42>  & (~\D<42>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<42>  & (\D<42>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<42>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<42>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<69>  & (\encrypt<0>  & \start<0> )) | (\key<77>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<77>  = \[343] ,
  \new_D<43>  = (~\$$COND0<0>5.1  & (\C<43>  & (\D<43>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<43>  & (\D<43>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<43>  & (~\D<43>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<43>  & (~\D<43>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<43>  & (\D<43>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<43>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<43>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<124>  & (\encrypt<0>  & \start<0> )) | (\key<69>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<82>  = \[338] ,
  \new_D<44>  = (~\$$COND0<0>5.1  & (\C<44>  & (\D<44>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<44>  & (\D<44>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<44>  & (~\D<44>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<44>  & (~\D<44>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<44>  & (\D<44>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<44>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<44>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<116>  & (\encrypt<0>  & \start<0> )) | (\key<124>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<81>  = \[339] ,
  \new_C<0>  = (~\$$COND0<0>5.1  & (~\D<0>  & (\C<0>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<0>  & (~\C<0>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<0>  & (\C<0>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<0>  & (~\C<0>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<0>  & (\C<0>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<0>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<0>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<48>  & (\encrypt<0>  & \start<0> )) | (\key<56>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<84>  = \[336] ,
  \new_C<9>  = (~\$$COND0<0>5.1  & (~\D<9>  & (\C<9>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<9>  & (~\C<9>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<9>  & (\C<9>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<9>  & (~\C<9>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<9>  & (\C<9>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<9>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<9>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<41>  & (\encrypt<0>  & \start<0> )) | (\key<49>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<83>  = \[337] ,
  \[330]  = \C<109> ,
  \[520]  = \new_C<12> ,
  \new_C<59>  = (~\$$COND0<0>5.1  & (~\D<59>  & (\C<59>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<59>  & (~\C<59>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<59>  & (\C<59>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<59>  & (~\C<59>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<59>  & (\C<59>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<59>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<59>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<152>  & (\encrypt<0>  & \start<0> )) | (\key<160>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_D<40>  = (~\$$COND0<0>5.1  & (\C<40>  & (\D<40>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<40>  & (\D<40>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<40>  & (~\D<40>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<40>  & (~\D<40>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<40>  & (\D<40>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<40>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<40>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<85>  & (\encrypt<0>  & \start<0> )) | (\key<93>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[331]  = \C<91> ,
  \[521]  = \new_C<11> ,
  \main/$PLUS_5_1/sum<3>5.1  = (~\main/$PLUS_5_1/c<0>5.4  & \count<3> ) | (\main/$PLUS_5_1/c<0>5.4  & ~\count<3> ),
  \[332]  = \C<109> ,
  \KSi<80>  = \[340] ,
  \[522]  = \new_C<10> ,
  \new_C<5>  = (~\$$COND0<0>5.1  & (~\D<5>  & (\C<5>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<5>  & (~\C<5>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<5>  & (\C<5>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<5>  & (~\C<5>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<5>  & (\C<5>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<5>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<5>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<8>  & (\encrypt<0>  & \start<0> )) | (\key<16>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[333]  = \C<87> ,
  \[523]  = \new_C<9> ,
  \new_C<6>  = (~\$$COND0<0>5.1  & (~\D<6>  & (\C<6>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<6>  & (~\C<6>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<6>  & (\C<6>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<6>  & (~\C<6>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<6>  & (\C<6>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<6>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<6>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<0>  & (\encrypt<0>  & \start<0> )) | (\key<8>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[334]  = \C<95> ,
  \[524]  = \new_C<8> ,
  \new_C<55>  = (~\$$COND0<0>5.1  & (~\D<55>  & (\C<55>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<55>  & (~\C<55>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<55>  & (\C<55>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<55>  & (~\C<55>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<55>  & (\C<55>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<55>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<55>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<184>  & (\encrypt<0>  & \start<0> )) | (\key<99>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<7>  = (~\$$COND0<0>5.1  & (~\D<7>  & (\C<7>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<7>  & (~\C<7>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<7>  & (\C<7>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<7>  & (~\C<7>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<7>  & (\C<7>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<7>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<7>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<57>  & (\encrypt<0>  & \start<0> )) | (\key<0>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[335]  = \C<102> ,
  \KSi<89>  = \[331] ,
  \[525]  = \new_C<7> ,
  \new_C<56>  = (~\$$COND0<0>5.1  & (~\D<56>  & (\C<56>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<56>  & (~\C<56>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<56>  & (\C<56>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<56>  & (~\C<56>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<56>  & (\C<56>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<56>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<56>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<176>  & (\encrypt<0>  & \start<0> )) | (\key<184>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<8>  = (~\$$COND0<0>5.1  & (~\D<8>  & (\C<8>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<8>  & (~\C<8>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<8>  & (\C<8>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<8>  & (~\C<8>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<8>  & (\C<8>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<8>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<8>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<49>  & (\encrypt<0>  & \start<0> )) | (\key<57>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[336]  = \C<106> ,
  \[526]  = \new_C<6> ,
  \new_C<57>  = (~\$$COND0<0>5.1  & (~\D<57>  & (\C<57>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<57>  & (~\C<57>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<57>  & (\C<57>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<57>  & (~\C<57>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<57>  & (\C<57>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<57>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<57>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<168>  & (\encrypt<0>  & \start<0> )) | (\key<176>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[337]  = \C<93> ,
  \[527]  = \new_C<5> ,
  \new_C<58>  = (~\$$COND0<0>5.1  & (~\D<58>  & (\C<58>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<58>  & (~\C<58>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<58>  & (\C<58>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<58>  & (~\C<58>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<58>  & (\C<58>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<58>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<58>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<160>  & (\encrypt<0>  & \start<0> )) | (\key<168>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[338]  = \C<104> ,
  \KSi<86>  = \[334] ,
  \[528]  = \new_C<4> ,
  \new_C<51>  = (~\$$COND0<0>5.1  & (~\D<51>  & (\C<51>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<51>  & (~\C<51>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<51>  & (\C<51>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<51>  & (~\C<51>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<51>  & (\C<51>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<51>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<51>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<123>  & (\encrypt<0>  & \start<0> )) | (\key<66>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[339]  = \C<89> ,
  \KSi<85>  = \[335] ,
  \[529]  = \new_C<3> ,
  \new_C<52>  = (~\$$COND0<0>5.1  & (~\D<52>  & (\C<52>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<52>  & (~\C<52>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<52>  & (\C<52>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<52>  & (~\C<52>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<52>  & (\C<52>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<52>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<52>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<115>  & (\encrypt<0>  & \start<0> )) | (\key<123>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<88>  = \[332] ,
  \new_C<53>  = (~\$$COND0<0>5.1  & (~\D<53>  & (\C<53>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<53>  & (~\C<53>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<53>  & (\C<53>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<53>  & (~\C<53>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<53>  & (\C<53>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<53>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<53>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<107>  & (\encrypt<0>  & \start<0> )) | (\key<115>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<87>  = \[333] ,
  \new_C<54>  = (~\$$COND0<0>5.1  & (~\D<54>  & (\C<54>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<54>  & (~\C<54>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<54>  & (\C<54>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<54>  & (~\C<54>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<54>  & (\C<54>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<54>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<54>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<99>  & (\encrypt<0>  & \start<0> )) | (\key<107>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<92>  = \[328] ,
  \KSi<91>  = \[329] ,
  \KSi<94>  = \[326] ,
  \KSi<93>  = \[327] ,
  \new_C<50>  = (~\$$COND0<0>5.1  & (~\D<50>  & (\C<50>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<50>  & (~\C<50>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<50>  & (\C<50>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<50>  & (~\C<50>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<50>  & (\C<50>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<50>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<50>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<66>  & (\encrypt<0>  & \start<0> )) | (\key<74>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[340]  = \C<98> ,
  \[530]  = \new_C<2> ,
  \new_C<69>  = (~\$$COND0<0>5.1  & (~\D<69>  & (\C<69>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<69>  & (~\C<69>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<69>  & (\C<69>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<69>  & (~\C<69>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<69>  & (\C<69>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<69>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<69>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<137>  & (\encrypt<0>  & \start<0> )) | (\key<145>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[341]  = \C<111> ,
  \[531]  = \new_C<1> ,
  \[342]  = \C<86> ,
  \KSi<90>  = \[330] ,
  \[532]  = \new_C<0> ,
  \[343]  = \C<88> ,
  \[533]  = \new_D<111> ,
  \[344]  = \C<84> ,
  \[534]  = \new_D<110> ,
  \new_C<65>  = (~\$$COND0<0>5.1  & (~\D<65>  & (\C<65>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<65>  & (~\C<65>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<65>  & (\C<65>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<65>  & (~\C<65>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<65>  & (\C<65>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<65>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<65>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<169>  & (\encrypt<0>  & \start<0> )) | (\key<177>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[345]  = \C<107> ,
  \KSi<99>  = \[321] ,
  \[535]  = \new_D<109> ,
  \new_C<66>  = (~\$$COND0<0>5.1  & (~\D<66>  & (\C<66>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<66>  & (~\C<66>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<66>  & (\C<66>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<66>  & (~\C<66>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<66>  & (\C<66>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<66>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<66>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<161>  & (\encrypt<0>  & \start<0> )) | (\key<169>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[346]  = \C<94> ,
  \[536]  = \new_D<108> ,
  \new_C<67>  = (~\$$COND0<0>5.1  & (~\D<67>  & (\C<67>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<67>  & (~\C<67>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<67>  & (\C<67>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<67>  & (~\C<67>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<67>  & (\C<67>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<67>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<67>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<153>  & (\encrypt<0>  & \start<0> )) | (\key<161>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[347]  = \C<100> ,
  \[537]  = \new_D<107> ,
  \new_C<68>  = (~\$$COND0<0>5.1  & (~\D<68>  & (\C<68>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<68>  & (~\C<68>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<68>  & (\C<68>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<68>  & (~\C<68>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<68>  & (\C<68>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<68>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<68>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<145>  & (\encrypt<0>  & \start<0> )) | (\key<153>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[348]  = \C<97> ,
  \KSi<96>  = \[324] ,
  \[538]  = \new_D<106> ,
  \new_C<61>  = (~\$$COND0<0>5.1  & (~\D<61>  & (\C<61>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<61>  & (~\C<61>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<61>  & (\C<61>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<61>  & (~\C<61>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<61>  & (\C<61>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<61>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<61>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<136>  & (\encrypt<0>  & \start<0> )) | (\key<144>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[349]  = \C<57> ,
  \KSi<95>  = \[325] ,
  \[539]  = \new_D<105> ,
  \new_C<62>  = (~\$$COND0<0>5.1  & (~\D<62>  & (\C<62>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<62>  & (~\C<62>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<62>  & (\C<62>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<62>  & (~\C<62>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<62>  & (\C<62>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<62>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<62>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<128>  & (\encrypt<0>  & \start<0> )) | (\key<136>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<98>  = \[322] ,
  \new_C<63>  = (~\$$COND0<0>5.1  & (~\D<63>  & (\C<63>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<63>  & (~\C<63>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<63>  & (\C<63>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<63>  & (~\C<63>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<63>  & (\C<63>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<63>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<63>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<185>  & (\encrypt<0>  & \start<0> )) | (\key<128>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<97>  = \[323] ,
  \new_C<64>  = (~\$$COND0<0>5.1  & (~\D<64>  & (\C<64>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<64>  & (~\C<64>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<64>  & (\C<64>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<64>  & (~\C<64>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<64>  & (\C<64>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<64>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<64>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<177>  & (\encrypt<0>  & \start<0> )) | (\key<185>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<120>  = \[300] ,
  \KSi<121>  = \[299] ,
  \new_C<60>  = (~\$$COND0<0>5.1  & (~\D<60>  & (\C<60>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<60>  & (~\C<60>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<60>  & (\C<60>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<60>  & (~\C<60>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<60>  & (\C<60>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<60>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<60>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<144>  & (\encrypt<0>  & \start<0> )) | (\key<152>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<122>  = \[298] ,
  \[350]  = \C<68> ,
  \[540]  = \new_D<104> ,
  \new_C<79>  = (~\$$COND0<0>5.1  & (~\D<79>  & (\C<79>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<79>  & (~\C<79>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<79>  & (\C<79>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<79>  & (~\C<79>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<79>  & (\C<79>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<79>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<79>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<187>  & (\encrypt<0>  & \start<0> )) | (\key<130>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<123>  = \[297] ,
  \[351]  = \C<75> ,
  \[541]  = \new_D<103> ,
  \KSi<124>  = \[296] ,
  \[352]  = \C<82> ,
  \[542]  = \new_D<102> ,
  \KSi<125>  = \[295] ,
  \[353]  = \C<62> ,
  \[543]  = \new_D<101> ,
  \KSi<126>  = \[294] ,
  \[354]  = \C<71> ,
  \[544]  = \new_D<100> ,
  \new_C<75>  = (~\$$COND0<0>5.1  & (~\D<75>  & (\C<75>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<75>  & (~\C<75>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<75>  & (\C<75>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<75>  & (~\C<75>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<75>  & (\C<75>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<75>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<75>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<154>  & (\encrypt<0>  & \start<0> )) | (\key<162>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<127>  = \[293] ,
  \[355]  = \C<63> ,
  \[545]  = \new_D<99> ,
  \new_C<76>  = (~\$$COND0<0>5.1  & (~\D<76>  & (\C<76>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<76>  & (~\C<76>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<76>  & (\C<76>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<76>  & (~\C<76>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<76>  & (\C<76>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<76>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<76>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<146>  & (\encrypt<0>  & \start<0> )) | (\key<154>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<128>  = \[292] ,
  \[356]  = \C<81> ,
  \[546]  = \new_D<98> ,
  \new_C<77>  = (~\$$COND0<0>5.1  & (~\D<77>  & (\C<77>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<77>  & (~\C<77>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<77>  & (\C<77>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<77>  & (~\C<77>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<77>  & (\C<77>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<77>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<77>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<138>  & (\encrypt<0>  & \start<0> )) | (\key<146>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<129>  = \[291] ,
  \[357]  = \C<59> ,
  \[547]  = \new_D<97> ,
  \new_C<78>  = (~\$$COND0<0>5.1  & (~\D<78>  & (\C<78>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<78>  & (~\C<78>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<78>  & (\C<78>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<78>  & (~\C<78>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<78>  & (\C<78>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<78>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<78>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<130>  & (\encrypt<0>  & \start<0> )) | (\key<138>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[358]  = \C<67> ,
  \[548]  = \new_D<96> ,
  \new_C<71>  = (~\$$COND0<0>5.1  & (~\D<71>  & (\C<71>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<71>  & (~\C<71>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<71>  & (\C<71>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<71>  & (~\C<71>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<71>  & (\C<71>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<71>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<71>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<186>  & (\encrypt<0>  & \start<0> )) | (\key<129>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[359]  = \C<74> ,
  \[549]  = \new_D<95> ,
  \new_C<72>  = (~\$$COND0<0>5.1  & (~\D<72>  & (\C<72>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<72>  & (~\C<72>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<72>  & (\C<72>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<72>  & (~\C<72>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<72>  & (\C<72>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<72>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<72>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<178>  & (\encrypt<0>  & \start<0> )) | (\key<186>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<73>  = (~\$$COND0<0>5.1  & (~\D<73>  & (\C<73>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<73>  & (~\C<73>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<73>  & (\C<73>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<73>  & (~\C<73>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<73>  & (\C<73>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<73>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<73>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<170>  & (\encrypt<0>  & \start<0> )) | (\key<178>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<74>  = (~\$$COND0<0>5.1  & (~\D<74>  & (\C<74>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<74>  & (~\C<74>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<74>  & (\C<74>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<74>  & (~\C<74>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<74>  & (\C<74>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<74>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<74>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<162>  & (\encrypt<0>  & \start<0> )) | (\key<170>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<110>  = \[310] ,
  \KSi<111>  = \[309] ,
  \new_C<70>  = (~\$$COND0<0>5.1  & (~\D<70>  & (\C<70>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<70>  & (~\C<70>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<70>  & (\C<70>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<70>  & (~\C<70>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<70>  & (\C<70>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<70>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<70>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<129>  & (\encrypt<0>  & \start<0> )) | (\key<137>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<112>  = \[308] ,
  \[360]  = \C<78> ,
  \[550]  = \new_D<94> ,
  \new_C<89>  = (~\$$COND0<0>5.1  & (~\D<89>  & (\C<89>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<89>  & (~\C<89>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<89>  & (\C<89>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<89>  & (~\C<89>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<89>  & (\C<89>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<89>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<89>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<200>  & (\encrypt<0>  & \start<0> )) | (\key<208>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<113>  = \[307] ,
  \[361]  = \C<65> ,
  \[551]  = \new_D<93> ,
  \KSi<114>  = \[306] ,
  \[362]  = \C<76> ,
  \[552]  = \new_D<92> ,
  \KSi<115>  = \[305] ,
  \[363]  = \C<61> ,
  \[553]  = \new_D<91> ,
  \KSi<116>  = \[304] ,
  \[364]  = \C<70> ,
  \[554]  = \new_D<90> ,
  \new_C<85>  = (~\$$COND0<0>5.1  & (~\D<85>  & (\C<85>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<85>  & (~\C<85>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<85>  & (\C<85>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<85>  & (~\C<85>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<85>  & (\C<85>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<85>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<85>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<232>  & (\encrypt<0>  & \start<0> )) | (\key<240>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<117>  = \[303] ,
  \[365]  = \C<83> ,
  \[555]  = \new_D<89> ,
  \new_C<86>  = (~\$$COND0<0>5.1  & (~\D<86>  & (\C<86>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<86>  & (~\C<86>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<86>  & (\C<86>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<86>  & (~\C<86>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<86>  & (\C<86>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<86>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<86>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<224>  & (\encrypt<0>  & \start<0> )) | (\key<232>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<118>  = \[302] ,
  \[366]  = \C<58> ,
  \[556]  = \new_D<88> ,
  \new_C<87>  = (~\$$COND0<0>5.1  & (~\D<87>  & (\C<87>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<87>  & (~\C<87>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<87>  & (\C<87>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<87>  & (~\C<87>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<87>  & (\C<87>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<87>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<87>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<216>  & (\encrypt<0>  & \start<0> )) | (\key<224>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<119>  = \[301] ,
  \[367]  = \C<60> ,
  \[557]  = \new_D<87> ,
  \new_C<88>  = (~\$$COND0<0>5.1  & (~\D<88>  & (\C<88>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<88>  & (~\C<88>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<88>  & (\C<88>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<88>  & (~\C<88>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<88>  & (\C<88>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<88>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<88>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<208>  & (\encrypt<0>  & \start<0> )) | (\key<216>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[368]  = \C<56> ,
  \[558]  = \new_D<86> ,
  \new_C<81>  = (~\$$COND0<0>5.1  & (~\D<81>  & (\C<81>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<81>  & (~\C<81>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<81>  & (\C<81>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<81>  & (~\C<81>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<81>  & (\C<81>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<81>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<81>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<171>  & (\encrypt<0>  & \start<0> )) | (\key<179>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[369]  = \C<79> ,
  \[559]  = \new_D<85> ,
  \new_C<82>  = (~\$$COND0<0>5.1  & (~\D<82>  & (\C<82>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<82>  & (~\C<82>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<82>  & (\C<82>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<82>  & (~\C<82>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<82>  & (\C<82>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<82>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<82>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<163>  & (\encrypt<0>  & \start<0> )) | (\key<171>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<83>  = (~\$$COND0<0>5.1  & (~\D<83>  & (\C<83>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<83>  & (~\C<83>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<83>  & (\C<83>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<83>  & (~\C<83>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<83>  & (\C<83>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<83>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<83>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<248>  & (\encrypt<0>  & \start<0> )) | (\key<163>  & (~\encrypt<0>  & \start<0> ))))))))),
  \new_C<84>  = (~\$$COND0<0>5.1  & (~\D<84>  & (\C<84>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<84>  & (~\C<84>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<84>  & (\C<84>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<84>  & (~\C<84>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<84>  & (\C<84>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<84>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<84>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<240>  & (\encrypt<0>  & \start<0> )) | (\key<248>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<140>  = \[280] ,
  \KSi<141>  = \[279] ,
  \new_C<80>  = (~\$$COND0<0>5.1  & (~\D<80>  & (\C<80>  & (\encrypt<0>  & ~\start<0> )))) | ((~\$$COND0<0>5.1  & (\D<80>  & (~\C<80>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\D<80>  & (\C<80>  & (\encrypt<0>  & ~\start<0> )))) | ((~\D<80>  & (~\C<80>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<80>  & (\C<80>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\D<80>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\C<80>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<179>  & (\encrypt<0>  & \start<0> )) | (\key<187>  & (~\encrypt<0>  & \start<0> ))))))))),
  \KSi<142>  = \[278] ,
  \[370]  = \C<66> ,
  \[560]  = \new_D<84> ,
  \KSi<143>  = \[277] ,
  \[371]  = \C<72> ,
  \[561]  = \new_D<83> ,
  \KSi<144>  = \[276] ,
  \new_D<99>  = (~\$$COND0<0>5.1  & (\C<99>  & (\D<99>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<99>  & (\D<99>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<99>  & (~\D<99>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<99>  & (~\D<99>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<99>  & (\D<99>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<99>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<99>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<252>  & (\encrypt<0>  & \start<0> )) | (\key<197>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[372]  = \C<69> ,
  \[562]  = \new_D<82> ,
  \KSi<145>  = \[275] ,
  \[373]  = \C<29> ,
  \[563]  = \new_D<81> ,
  \KSi<146>  = \[274] ,
  \[374]  = \C<40> ,
  \[564]  = \new_D<80> ,
  \KSi<147>  = \[273] ,
  \[375]  = \C<47> ,
  \[565]  = \new_D<79> ,
  \$$COND1<0>8.1  = (~\count<3>  & (~\count<2>  & (~\count<1>  & ~\count<0> ))) | ((~\count<3>  & (~\count<2>  & (~\count<1>  & \count<0> ))) | ((\count<3>  & (~\count<2>  & (~\count<1>  & ~\count<0> ))) | (\count<3>  & (\count<2>  & (\count<1>  & \count<0> ))))),
  \KSi<148>  = \[272] ,
  \new_D<95>  = (~\$$COND0<0>5.1  & (\C<95>  & (\D<95>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<95>  & (\D<95>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<95>  & (~\D<95>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<95>  & (~\D<95>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<95>  & (\D<95>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<95>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<95>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<221>  & (\encrypt<0>  & \start<0> )) | (\key<229>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[376]  = \C<54> ,
  \[566]  = \new_D<78> ,
  \KSi<149>  = \[271] ,
  \new_D<96>  = (~\$$COND0<0>5.1  & (\C<96>  & (\D<96>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<96>  & (\D<96>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<96>  & (~\D<96>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<96>  & (~\D<96>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<96>  & (\D<96>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<96>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<96>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<213>  & (\encrypt<0>  & \start<0> )) | (\key<221>  & (~\encrypt<0>  & \start<0> ))))))))),
  \[377]  = \C<34> ,
  \[567]  = \new_D<77> ,
  \new_D<97>  = (~\$$COND0<0>5.1  & (\C<97>  & (\D<97>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (~\C<97>  & (\D<97>  & (\encrypt<0>  & ~\start<0> )))) | ((\$$COND0<0>5.1  & (\C<97>  & (~\D<97>  & (\encrypt<0>  & ~\start<0> )))) | ((~\C<97>  & (~\D<97>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<97>  & (\D<97>  & (~\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> )))) | ((\C<97>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\D<97>  & (\$$COND1<0>8.1  & (~\encrypt<0>  & ~\start<0> ))) | ((\key<205>  & (\encrypt<0>  & \start<0> )) | (\key<213>  & (~\encrypt<0>  & \start<0> )))))))));
always begin
  \D<0>  = \[644] ;
  \D<1>  = \[643] ;
  \D<2>  = \[642] ;
  \D<3>  = \[641] ;
  \D<4>  = \[640] ;
  \D<5>  = \[639] ;
  \D<6>  = \[638] ;
  \C<10>  = \[522] ;
  \D<7>  = \[637] ;
  \C<11>  = \[521] ;
  \D<8>  = \[636] ;
  \C<12>  = \[520] ;
  \D<9>  = \[635] ;
  \C<13>  = \[519] ;
  \C<14>  = \[518] ;
  \C<15>  = \[517] ;
  \C<16>  = \[516] ;
  \C<17>  = \[515] ;
  \C<18>  = \[514] ;
  \C<19>  = \[513] ;
  \C<20>  = \[512] ;
  \C<21>  = \[511] ;
  \C<22>  = \[510] ;
  \C<23>  = \[509] ;
  \C<24>  = \[508] ;
  \C<25>  = \[507] ;
  \C<26>  = \[506] ;
  \C<27>  = \[505] ;
  \C<28>  = \[504] ;
  \C<29>  = \[503] ;
  \C<30>  = \[502] ;
  \C<31>  = \[501] ;
  \C<32>  = \[500] ;
  \C<33>  = \[499] ;
  \C<34>  = \[498] ;
  \C<35>  = \[497] ;
  \C<36>  = \[496] ;
  \C<37>  = \[495] ;
  \C<38>  = \[494] ;
  \C<39>  = \[493] ;
  \C<40>  = \[492] ;
  \C<41>  = \[491] ;
  \C<42>  = \[490] ;
  \C<43>  = \[489] ;
  \C<44>  = \[488] ;
  \C<45>  = \[487] ;
  \C<46>  = \[486] ;
  \C<47>  = \[485] ;
  \C<48>  = \[484] ;
  \C<49>  = \[483] ;
  \C<50>  = \[482] ;
  \C<51>  = \[481] ;
  \C<52>  = \[480] ;
  \C<53>  = \[479] ;
  \C<54>  = \[478] ;
  \C<55>  = \[477] ;
  \C<56>  = \[476] ;
  \C<57>  = \[475] ;
  \C<58>  = \[474] ;
  \C<59>  = \[473] ;
  \C<60>  = \[472] ;
  \C<61>  = \[471] ;
  \C<62>  = \[470] ;
  \C<63>  = \[469] ;
  \C<64>  = \[468] ;
  \C<65>  = \[467] ;
  \C<66>  = \[466] ;
  \C<67>  = \[465] ;
  \C<68>  = \[464] ;
  \C<69>  = \[463] ;
  \C<70>  = \[462] ;
  \C<71>  = \[461] ;
  \C<72>  = \[460] ;
  \C<73>  = \[459] ;
  \C<74>  = \[458] ;
  \C<75>  = \[457] ;
  \C<76>  = \[456] ;
  \C<77>  = \[455] ;
  \C<78>  = \[454] ;
  \C<79>  = \[453] ;
  \C<80>  = \[452] ;
  \C<81>  = \[451] ;
  \C<82>  = \[450] ;
  \C<83>  = \[449] ;
  \C<84>  = \[448] ;
  \C<85>  = \[447] ;
  \C<86>  = \[446] ;
  \C<87>  = \[445] ;
  \C<88>  = \[444] ;
  \C<89>  = \[443] ;
  \C<90>  = \[442] ;
  \C<91>  = \[441] ;
  \D<10>  = \[634] ;
  \C<92>  = \[440] ;
  \D<11>  = \[633] ;
  \C<93>  = \[439] ;
  \D<12>  = \[632] ;
  \C<94>  = \[438] ;
  \D<13>  = \[631] ;
  \C<95>  = \[437] ;
  \D<14>  = \[630] ;
  \C<96>  = \[436] ;
  \D<15>  = \[629] ;
  \C<97>  = \[435] ;
  \D<16>  = \[628] ;
  \C<98>  = \[434] ;
  \D<17>  = \[627] ;
  \C<99>  = \[433] ;
  \D<18>  = \[626] ;
  \D<19>  = \[625] ;
  \D<20>  = \[624] ;
  \D<21>  = \[623] ;
  \D<22>  = \[622] ;
  \D<23>  = \[621] ;
  \D<24>  = \[620] ;
  \D<25>  = \[619] ;
  \D<26>  = \[618] ;
  \D<27>  = \[617] ;
  \D<28>  = \[616] ;
  \D<29>  = \[615] ;
  \D<30>  = \[614] ;
  \D<31>  = \[613] ;
  \D<32>  = \[612] ;
  \D<33>  = \[611] ;
  \D<34>  = \[610] ;
  \D<35>  = \[609] ;
  \D<36>  = \[608] ;
  \D<37>  = \[607] ;
  \D<38>  = \[606] ;
  \D<39>  = \[605] ;
  \D<40>  = \[604] ;
  \D<41>  = \[603] ;
  \D<42>  = \[602] ;
  \D<43>  = \[601] ;
  \D<44>  = \[600] ;
  \D<45>  = \[599] ;
  \D<46>  = \[598] ;
  \D<47>  = \[597] ;
  \D<48>  = \[596] ;
  \D<49>  = \[595] ;
  \D<50>  = \[594] ;
  \D<51>  = \[593] ;
  \D<52>  = \[592] ;
  \D<53>  = \[591] ;
  \D<54>  = \[590] ;
  \D<55>  = \[589] ;
  \D<56>  = \[588] ;
  \D<57>  = \[587] ;
  \D<58>  = \[586] ;
  \D<59>  = \[585] ;
  \D<60>  = \[584] ;
  \D<61>  = \[583] ;
  \D<62>  = \[582] ;
  \D<63>  = \[581] ;
  \D<64>  = \[580] ;
  \D<65>  = \[579] ;
  \D<66>  = \[578] ;
  \D<67>  = \[577] ;
  \D<68>  = \[576] ;
  \D<69>  = \[575] ;
  \C<100>  = \[432] ;
  \D<70>  = \[574] ;
  \C<101>  = \[431] ;
  \D<71>  = \[573] ;
  \C<102>  = \[430] ;
  \D<72>  = \[572] ;
  \C<103>  = \[429] ;
  \D<73>  = \[571] ;
  \C<104>  = \[428] ;
  \D<74>  = \[570] ;
  \C<105>  = \[427] ;
  \D<75>  = \[569] ;
  \C<106>  = \[426] ;
  \D<76>  = \[568] ;
  \C<107>  = \[425] ;
  \D<77>  = \[567] ;
  \C<108>  = \[424] ;
  \C<0>  = \[532] ;
  \D<78>  = \[566] ;
  \C<109>  = \[423] ;
  \C<1>  = \[531] ;
  \D<79>  = \[565] ;
  \C<2>  = \[530] ;
  \C<3>  = \[529] ;
  \C<4>  = \[528] ;
  \C<5>  = \[527] ;
  \C<6>  = \[526] ;
  \C<7>  = \[525] ;
  \C<110>  = \[422] ;
  \C<8>  = \[524] ;
  \D<80>  = \[564] ;
  \C<111>  = \[421] ;
  \C<9>  = \[523] ;
  \D<81>  = \[563] ;
  \D<82>  = \[562] ;
  \D<83>  = \[561] ;
  \D<84>  = \[560] ;
  \D<85>  = \[559] ;
  \D<86>  = \[558] ;
  \D<87>  = \[557] ;
  \D<88>  = \[556] ;
  \D<89>  = \[555] ;
  \D<90>  = \[554] ;
  \D<91>  = \[553] ;
  \D<92>  = \[552] ;
  \D<93>  = \[551] ;
  \D<94>  = \[550] ;
  \D<95>  = \[549] ;
  \D<96>  = \[548] ;
  \D<97>  = \[547] ;
  \D<98>  = \[546] ;
  \D<99>  = \[545] ;
  \D<100>  = \[544] ;
  \D<101>  = \[543] ;
  \D<102>  = \[542] ;
  \D<103>  = \[541] ;
  \D<104>  = \[540] ;
  \D<105>  = \[539] ;
  \D<106>  = \[538] ;
  \D<107>  = \[537] ;
  \D<108>  = \[536] ;
  \D<109>  = \[535] ;
  \D<110>  = \[534] ;
  \D<111>  = \[533] ;
end
initial begin
  \D<0>  = 0;
  \D<1>  = 0;
  \D<2>  = 0;
  \D<3>  = 0;
  \D<4>  = 0;
  \D<5>  = 0;
  \D<6>  = 0;
  \C<10>  = 0;
  \D<7>  = 0;
  \C<11>  = 0;
  \D<8>  = 0;
  \C<12>  = 0;
  \D<9>  = 0;
  \C<13>  = 0;
  \C<14>  = 0;
  \C<15>  = 0;
  \C<16>  = 0;
  \C<17>  = 0;
  \C<18>  = 0;
  \C<19>  = 0;
  \C<20>  = 0;
  \C<21>  = 0;
  \C<22>  = 0;
  \C<23>  = 0;
  \C<24>  = 0;
  \C<25>  = 0;
  \C<26>  = 0;
  \C<27>  = 0;
  \C<28>  = 0;
  \C<29>  = 0;
  \C<30>  = 0;
  \C<31>  = 0;
  \C<32>  = 0;
  \C<33>  = 0;
  \C<34>  = 0;
  \C<35>  = 0;
  \C<36>  = 0;
  \C<37>  = 0;
  \C<38>  = 0;
  \C<39>  = 0;
  \C<40>  = 0;
  \C<41>  = 0;
  \C<42>  = 0;
  \C<43>  = 0;
  \C<44>  = 0;
  \C<45>  = 0;
  \C<46>  = 0;
  \C<47>  = 0;
  \C<48>  = 0;
  \C<49>  = 0;
  \C<50>  = 0;
  \C<51>  = 0;
  \C<52>  = 0;
  \C<53>  = 0;
  \C<54>  = 0;
  \C<55>  = 0;
  \C<56>  = 0;
  \C<57>  = 0;
  \C<58>  = 0;
  \C<59>  = 0;
  \C<60>  = 0;
  \C<61>  = 0;
  \C<62>  = 0;
  \C<63>  = 0;
  \C<64>  = 0;
  \C<65>  = 0;
  \C<66>  = 0;
  \C<67>  = 0;
  \C<68>  = 0;
  \C<69>  = 0;
  \C<70>  = 0;
  \C<71>  = 0;
  \C<72>  = 0;
  \C<73>  = 0;
  \C<74>  = 0;
  \C<75>  = 0;
  \C<76>  = 0;
  \C<77>  = 0;
  \C<78>  = 0;
  \C<79>  = 0;
  \C<80>  = 0;
  \C<81>  = 0;
  \C<82>  = 0;
  \C<83>  = 0;
  \C<84>  = 0;
  \C<85>  = 0;
  \C<86>  = 0;
  \C<87>  = 0;
  \C<88>  = 0;
  \C<89>  = 0;
  \C<90>  = 0;
  \C<91>  = 0;
  \D<10>  = 0;
  \C<92>  = 0;
  \D<11>  = 0;
  \C<93>  = 0;
  \D<12>  = 0;
  \C<94>  = 0;
  \D<13>  = 0;
  \C<95>  = 0;
  \D<14>  = 0;
  \C<96>  = 0;
  \D<15>  = 0;
  \C<97>  = 0;
  \D<16>  = 0;
  \C<98>  = 0;
  \D<17>  = 0;
  \C<99>  = 0;
  \D<18>  = 0;
  \D<19>  = 0;
  \D<20>  = 0;
  \D<21>  = 0;
  \D<22>  = 0;
  \D<23>  = 0;
  \D<24>  = 0;
  \D<25>  = 0;
  \D<26>  = 0;
  \D<27>  = 0;
  \D<28>  = 0;
  \D<29>  = 0;
  \D<30>  = 0;
  \D<31>  = 0;
  \D<32>  = 0;
  \D<33>  = 0;
  \D<34>  = 0;
  \D<35>  = 0;
  \D<36>  = 0;
  \D<37>  = 0;
  \D<38>  = 0;
  \D<39>  = 0;
  \D<40>  = 0;
  \D<41>  = 0;
  \D<42>  = 0;
  \D<43>  = 0;
  \D<44>  = 0;
  \D<45>  = 0;
  \D<46>  = 0;
  \D<47>  = 0;
  \D<48>  = 0;
  \D<49>  = 0;
  \D<50>  = 0;
  \D<51>  = 0;
  \D<52>  = 0;
  \D<53>  = 0;
  \D<54>  = 0;
  \D<55>  = 0;
  \D<56>  = 0;
  \D<57>  = 0;
  \D<58>  = 0;
  \D<59>  = 0;
  \D<60>  = 0;
  \D<61>  = 0;
  \D<62>  = 0;
  \D<63>  = 0;
  \D<64>  = 0;
  \D<65>  = 0;
  \D<66>  = 0;
  \D<67>  = 0;
  \D<68>  = 0;
  \D<69>  = 0;
  \C<100>  = 0;
  \D<70>  = 0;
  \C<101>  = 0;
  \D<71>  = 0;
  \C<102>  = 0;
  \D<72>  = 0;
  \C<103>  = 0;
  \D<73>  = 0;
  \C<104>  = 0;
  \D<74>  = 0;
  \C<105>  = 0;
  \D<75>  = 0;
  \C<106>  = 0;
  \D<76>  = 0;
  \C<107>  = 0;
  \D<77>  = 0;
  \C<108>  = 0;
  \C<0>  = 0;
  \D<78>  = 0;
  \C<109>  = 0;
  \C<1>  = 0;
  \D<79>  = 0;
  \C<2>  = 0;
  \C<3>  = 0;
  \C<4>  = 0;
  \C<5>  = 0;
  \C<6>  = 0;
  \C<7>  = 0;
  \C<110>  = 0;
  \C<8>  = 0;
  \D<80>  = 0;
  \C<111>  = 0;
  \C<9>  = 0;
  \D<81>  = 0;
  \D<82>  = 0;
  \D<83>  = 0;
  \D<84>  = 0;
  \D<85>  = 0;
  \D<86>  = 0;
  \D<87>  = 0;
  \D<88>  = 0;
  \D<89>  = 0;
  \D<90>  = 0;
  \D<91>  = 0;
  \D<92>  = 0;
  \D<93>  = 0;
  \D<94>  = 0;
  \D<95>  = 0;
  \D<96>  = 0;
  \D<97>  = 0;
  \D<98>  = 0;
  \D<99>  = 0;
  \D<100>  = 0;
  \D<101>  = 0;
  \D<102>  = 0;
  \D<103>  = 0;
  \D<104>  = 0;
  \D<105>  = 0;
  \D<106>  = 0;
  \D<107>  = 0;
  \D<108>  = 0;
  \D<109>  = 0;
  \D<110>  = 0;
  \D<111>  = 0;
end
endmodule

