module s1488_bench(
  blif_clk_net,
  blif_reset_net,
  CLR,
  v6,
  v5,
  v4,
  v3,
  v2,
  v1,
  v0,
  v13_D_20,
  v13_D_21,
  v13_D_16,
  v13_D_22,
  v13_D_19,
  v13_D_18,
  v13_D_11,
  v13_D_23,
  v13_D_6,
  v13_D_15,
  v13_D_9,
  v13_D_10,
  v13_D_8,
  v13_D_24,
  v13_D_14,
  v13_D_7,
  v13_D_17,
  v13_D_12,
  v13_D_13);
input blif_clk_net;
input blif_reset_net;
input CLR;
input v6;
input v5;
input v4;
input v3;
input v2;
input v1;
input v0;
output v13_D_20;
output v13_D_21;
output v13_D_16;
output v13_D_22;
output v13_D_19;
output v13_D_18;
output v13_D_11;
output v13_D_23;
output v13_D_6;
output v13_D_15;
output v13_D_9;
output v13_D_10;
output v13_D_8;
output v13_D_24;
output v13_D_14;
output v13_D_7;
output v13_D_17;
output v13_D_12;
output v13_D_13;
reg v12;
reg v11;
reg v10;
reg v9;
reg v8;
reg v7;
wire IIII88;
wire IIII108;
wire IIII267;
wire Av13_D_23B;
wire C199D;
wire IIII365;
wire C131DE;
wire C26D;
wire IIII188;
wire C172D;
wire C185D;
wire C119D;
wire IIII134;
wire IIII27;
wire IIII547;
wire IIII534;
wire IIII177;
wire IIII197;
wire IIII28;
wire IIII226;
wire IIII253;
wire C161D;
wire IIII300;
wire IIII468;
wire C76D;
wire IIII145;
wire IIII203;
wire IIII93;
wire II659;
wire II686;
wire IIII263;
wire C168D;
wire II689;
wire C27D;
wire C110D;
wire IIII69;
wire IIII288;
wire IIII83;
wire C160D;
wire IIII405;
wire IIII41;
wire C90D;
wire v13_D_1;
wire IIII387;
wire Av13_D_13B;
wire C29D;
wire IIII34;
wire IIII429;
wire IIII236;
wire II704;
wire C123D;
wire C153D;
wire C124DE;
wire IIII500;
wire IIII409;
wire IIII321;
wire IIII489;
wire IIII498;
wire C99D;
wire v3E;
wire IIII296;
wire IIII518;
wire IIII129;
wire C82D;
wire v4E;
wire IIII442;
wire IIII318;
wire C104DE;
wire C38D;
wire IIII161;
wire IIII506;
wire v13_D_2C;
wire IIII98;
wire C86D;
wire IIII533;
wire C105D;
wire IIII151;
wire IIII35;
wire Av13_D_9B;
wire Av13_D_0B;
wire II692;
wire C118D;
wire IIII415;
wire C144DE;
wire IIII475;
wire IIII278;
wire C88D;
wire IIII368;
wire C83D;
wire IIII105;
wire IIII444;
wire II716;
wire IIII359;
wire C138D;
wire IIII482;
wire C67D;
wire IIII554;
wire Av13_D_3B;
wire IIII72;
wire C215D;
wire IIII210;
wire IIII68;
wire IIII452;
wire Av13_D_11B;
wire IIII406;
wire IIII227;
wire IIII82;
wire IIII213;
wire v12E;
wire II114;
wire C202D;
wire II329;
wire IIII464;
wire IIII245;
wire C78D;
wire IIII157;
wire II142;
wire C109D;
wire IIII269;
wire C104D;
wire C167D;
wire IIII310;
wire IIII317;
wire C194DE;
wire C184D;
wire Av13_D_14B;
wire IIII297;
wire II650;
wire C169D;
wire IIII435;
wire C44D;
wire IIII91;
wire IIII329;
wire II707;
wire IIII123;
wire C180D;
wire IIII449;
wire II294;
wire IIII342;
wire IIII360;
wire II246;
wire IIII114;
wire C42D;
wire IIII302;
wire C126D;
wire IIII282;
wire IIII40;
wire Av13_D_24B;
wire C59D;
wire C45D;
wire IIII79;
wire v13_D_4C;
wire IIII212;
wire C117D;
wire IIII386;
wire II368;
wire v2E;
wire IIII222;
wire IIII501;
wire IIII71;
wire IIII483;
wire IIII260;
wire IIII86;
wire IIII92;
wire C120D;
wire IIII470;
wire IIII117;
wire C48D;
wire C188D;
wire C146D;
wire IIII58;
wire IIII39;
wire IIII55;
wire IIII128;
wire Av13_D_20B;
wire IIII95;
wire IIII516;
wire IIII281;
wire IIII513;
wire C81DE;
wire II722;
wire C189D;
wire IIII375;
wire IIII106;
wire IIII73;
wire C63D;
wire IIII243;
wire IIII299;
wire C100D;
wire IIII311;
wire IIII148;
wire IIII31;
wire C139D;
wire IIII399;
wire C115D;
wire C186D;
wire C191DE;
wire C134D;
wire IIII287;
wire IIII43;
wire C102D;
wire C97D;
wire IIII341;
wire IIII393;
wire IIII420;
wire IIII48;
wire IIII390;
wire C54D;
wire C30D;
wire II491;
wire IIII520;
wire C207D;
wire IIII127;
wire C98D;
wire IIII170;
wire C150D;
wire II683;
wire II642;
wire IIII196;
wire IIII167;
wire C74D;
wire IIII433;
wire IIII133;
wire IIII339;
wire C55D;
wire C133D;
wire v13_D_1C;
wire v13_D_0;
wire IIII275;
wire IIII205;
wire IIII186;
wire IIII200;
wire IIII471;
wire C141D;
wire IIII116;
wire Av13_D_10B;
wire IIII280;
wire IIII308;
wire IIII54;
wire IIII555;
wire IIII389;
wire C35D;
wire v10E;
wire v7E;
wire IIII350;
wire II653;
wire C220DE;
wire C53D;
wire C166D;
wire IIII199;
wire IIII59;
wire IIII146;
wire IIII262;
wire IIII323;
wire C201D;
wire IIII89;
wire II159;
wire IIII362;
wire IIII36;
wire IIII333;
wire Av13_D_8B;
wire IIII332;
wire IIII276;
wire C77D;
wire IIII242;
wire IIII237;
wire C43D;
wire IIII378;
wire C200D;
wire C177D;
wire C57D;
wire C56D;
wire II101;
wire IIII326;
wire IIII560;
wire IIII476;
wire IIII414;
wire C220D;
wire IIII169;
wire IIII450;
wire C129DE;
wire IIII438;
wire C218DE;
wire C148D;
wire IIII514;
wire IIII247;
wire IIII119;
wire Av13_D_2B;
wire C179D;
wire IIII49;
wire IIII495;
wire C140D;
wire IIII140;
wire C31D;
wire IIII432;
wire C49D;
wire IIII171;
wire IIII430;
wire C187D;
wire IIII80;
wire IIII223;
wire IIII546;
wire C164D;
wire C221D;
wire IIII441;
wire C180DE;
wire v5E;
wire IIII160;
wire v9E;
wire IIII402;
wire C70D;
wire C196D;
wire IIII220;
wire IIII478;
wire IIII272;
wire IIII137;
wire Av13_D_17B;
wire C116D;
wire IIII384;
wire C124D;
wire C166DE;
wire C176D;
wire C137D;
wire IIII97;
wire C142D;
wire C46D;
wire IIII352;
wire IIII369;
wire II497;
wire C165D;
wire C73D;
wire IIII372;
wire II674;
wire C181D;
wire C72D;
wire IIII473;
wire IIII131;
wire IIII446;
wire C91D;
wire IIII62;
wire IIII216;
wire IIII126;
wire IIII45;
wire IIII392;
wire C217D;
wire IIII395;
wire IIII423;
wire v13_D_4;
wire IIII234;
wire IIII508;
wire IIII494;
wire IIII377;
wire C39D;
wire C144D;
wire Av13_D_6B;
wire IIII64;
wire IIII233;
wire IIII84;
wire C89D;
wire Av13_D_22B;
wire IIII439;
wire IIII215;
wire IIII285;
wire IIII503;
wire C128D;
wire IIII130;
wire C130D;
wire C175D;
wire IIII38;
wire IIII320;
wire Av13_D_7B;
wire C37D;
wire C47D;
wire C28D;
wire IIII305;
wire IIII528;
wire IIII456;
wire II671;
wire C191D;
wire IIII485;
wire C113D;
wire C135D;
wire C118DE;
wire C70DE;
wire C112D;
wire II695;
wire Av13_D_21B;
wire v0E;
wire IIII96;
wire IIII396;
wire IIII180;
wire Av13_D_1B;
wire C147D;
wire C195D;
wire IIII153;
wire C87D;
wire IIII256;
wire IIII229;
wire IIII293;
wire IIII447;
wire IIII87;
wire IIII463;
wire IIII291;
wire IIII174;
wire C223D;
wire C90DE;
wire IIII76;
wire Av13_D_16B;
wire Av13_D_5B;
wire v13_D_3C;
wire IIII191;
wire IIII240;
wire IIII425;
wire v11E;
wire IIII347;
wire II542;
wire IIII273;
wire II668;
wire IIII154;
wire IIII189;
wire II548;
wire IIII325;
wire IIII479;
wire IIII538;
wire IIII173;
wire v8E;
wire C157D;
wire IIII111;
wire IIII284;
wire IIII419;
wire Av13_D_18B;
wire IIII239;
wire IIII75;
wire IIII403;
wire C214D;
wire IIII166;
wire C114D;
wire II677;
wire IIII103;
wire IIII52;
wire IIII354;
wire IIII44;
wire IIII336;
wire Av13_D_12B;
wire IIII412;
wire IIII109;
wire IIII104;
wire C85D;
wire C71D;
wire C173D;
wire IIII270;
wire C209D;
wire C162D;
wire C117DE;
wire IIII346;
wire IIII60;
wire C156D;
wire C75D;
wire C108D;
wire II373;
wire II680;
wire IIII457;
wire C79D;
wire C93D;
wire C81D;
wire C145D;
wire C84D;
wire IIII232;
wire Av13_D_15B;
wire IIII306;
wire II254;
wire IIII383;
wire C111D;
wire C163D;
wire C108DE;
wire IIII32;
wire IIII315;
wire IIII380;
wire IIII192;
wire C80D;
wire II665;
wire C203D;
wire C36D;
wire C129D;
wire C151D;
wire C95D;
wire v1E;
wire IIII163;
wire IIII100;
wire C125D;
wire IIII179;
wire IIII208;
wire C40D;
wire C183D;
wire Av13_D_4B;
wire C143D;
wire IIII136;
wire IIII492;
wire IIII363;
wire IIII250;
wire v13_D_0C;
wire C155D;
wire IIII524;
wire C58D;
wire IIII453;
wire IIII328;
wire IIII224;
wire IIII338;
wire C30DE;
wire C165DE;
wire IIII460;
wire IIII113;
wire IIII142;
wire C218D;
wire C193D;
wire C178D;
wire IIII63;
wire C65D;
wire IIII259;
wire v13_D_2;
wire C174D;
wire IIII66;
wire IIII185;
wire C216D;
wire IIII202;
wire C222D;
wire II710;
wire IIII510;
wire C131D;
wire IIII164;
wire IIII124;
wire IIII505;
wire C225D;
wire C157DE;
wire C92D;
wire IIII251;
wire C106D;
wire IIII182;
wire IIII152;
wire IIII537;
wire II143;
wire II701;
wire C206D;
wire IIII218;
wire IIII158;
wire C83DE;
wire C50D;
wire IIII294;
wire IIII335;
wire IIII51;
wire C170D;
wire IIII398;
wire IIII175;
wire IIII149;
wire IIII436;
wire II656;
wire IIII29;
wire C205D;
wire IIII417;
wire IIII156;
wire C195DE;
wire C122D;
wire C96D;
wire C52D;
wire IIII257;
wire C51D;
wire IIII101;
wire C211D;
wire IIII374;
wire II698;
wire IIII176;
wire II610;
wire C194D;
wire C69D;
wire C141DE;
wire IIII461;
wire IIII486;
wire IIII266;
wire v6E;
wire IIII357;
wire C224D;
wire C158D;
wire IIII248;
wire C213D;
wire IIII371;
wire IIII219;
wire IIII314;
wire C132D;
wire IIII194;
wire v13_D_5C;
wire C107D;
wire C152D;
wire IIII356;
wire C34D;
wire IIII344;
wire IIII78;
wire C159D;
wire IIII366;
wire IIII427;
wire C138DE;
wire C103D;
wire IIII381;
wire C49DE;
wire C190D;
wire IIII497;
wire IIII46;
wire IIII120;
wire v13_D_3;
wire C219D;
wire IIII254;
wire II719;
wire C60D;
wire IIII183;
wire IIII65;
wire C192D;
wire IIII559;
wire IIII141;
wire IIII491;
wire II713;
wire II662;
wire IIII206;
wire C210D;
wire IIII349;
wire C208D;
wire C208DE;
wire IIII230;
wire C33D;
wire C127D;
wire C41D;
wire IIII209;
wire IIII466;
wire v13_D_5;
wire IIII303;
wire Av13_D_19B;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    v12 <= 0;
  else
    v12 <= v13_D_5C;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    v11 <= 0;
  else
    v11 <= v13_D_4C;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    v10 <= 0;
  else
    v10 <= v13_D_3C;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    v9 <= 0;
  else
    v9 <= v13_D_2C;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    v8 <= 0;
  else
    v8 <= v13_D_1C;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    v7 <= 0;
  else
    v7 <= v13_D_0C;
assign IIII88 = (v2E&C43D);
assign IIII108 = (C181D&C83DE);
assign IIII267 = (C214D&v7E&v10E);
assign Av13_D_23B = (C216D&v7E&v8E);
assign C199D = (IIII191)|(IIII192);
assign IIII365 = (C56D&v8&v11);
assign C131DE = ((~C131D));
assign C26D = (IIII414)|(IIII415);
assign IIII188 = (C175D&v11);
assign C172D = (IIII478)|(IIII479);
assign v13_D_19 = ((~II665));
assign IIII27 = (C184D&v7);
assign C185D = (IIII491)|(IIII492);
assign C119D = (IIII349)|(IIII350);
assign IIII134 = (v7E&v10&C151D);
assign IIII547 = (v10&v11E);
assign IIII534 = (v8E&v10E);
assign IIII177 = (C137D&C127D);
assign IIII197 = (C158D&v7&v11E);
assign IIII28 = (v7E&C188D);
assign IIII226 = (v8E&v10E&C144DE);
assign IIII253 = (v1E&v10E&C138DE);
assign C161D = (IIII314)|(IIII315);
assign IIII300 = (v0E&C105D);
assign IIII468 = (v9&C83DE);
assign C76D = (C131DE)|(IIII427);
assign IIII145 = (C49DE&C166DE&C220DE);
assign IIII93 = (v7E&C147D);
assign IIII203 = (C34D&v9);
assign II659 = ((~Av13_D_21B));
assign II686 = ((~Av13_D_12B));
assign IIII263 = (v7E&v11&C41D);
assign C168D = (C159D)|(v9);
assign II689 = ((~Av13_D_11B));
assign C27D = (IIII500)|(IIII501);
assign C110D = (IIII229)|(IIII230);
assign IIII69 = (v7&C202D);
assign IIII288 = (v7E&C203D);
assign IIII83 = (C225D&v11);
assign C160D = (IIII341)|(IIII342);
assign IIII405 = (v8E&v9E&C194DE);
assign IIII41 = (v7&v12E&C96D);
assign v13_D_1 = ((~II719));
assign C90D = (v9)|(v12E);
assign IIII387 = (v8E&v9E&C124DE);
assign Av13_D_13B = (IIII27)|(IIII28)|(IIII29);
assign C29D = (C138DE)|(IIII466);
assign IIII34 = (C91D&C165DE);
assign IIII429 = (v9E&C30DE);
assign IIII236 = (v2E&v8&C219D);
assign v13_D_20 = ((~II662));
assign II704 = ((~Av13_D_6B));
assign C123D = (C157DE)|(IIII208)|(IIII209)|(IIII210);
assign C153D = (IIII133)|(IIII134);
assign C124DE = ((~C124D));
assign IIII500 = (v8&v11&C83DE);
assign IIII409 = (v9&v11E);
assign IIII321 = (C33D&v11E&v12E);
assign IIII489 = (v8E&v11);
assign IIII498 = (v8&C117DE);
assign C99D = (IIII111)|(IIII113)|(IIII114);
assign v3E = ((~v3));
assign IIII296 = (v8E&v9E&C124DE&C83DE);
assign IIII518 = ((~II101));
assign IIII129 = (v8E&C72D);
assign C82D = (IIII392)|(IIII393);
assign v4E = ((~v4));
assign IIII442 = (v7E&v8E&v9E);
assign IIII318 = (v11&C118D);
assign C104DE = ((~C104D));
assign C38D = (IIII116)|(IIII117);
assign IIII161 = (C144DE&C191D);
assign IIII506 = (v7E&v9&v10E&v12E);
assign v13_D_2C = (v13_D_2&CLR);
assign IIII98 = (v8E&v12&C87D);
assign C86D = (v9)|(IIII524);
assign IIII533 = (v9&v10);
assign C105D = (IIII449)|(IIII450);
assign v13_D_23 = ((~II653));
assign IIII151 = (v9&C138DE);
assign IIII35 = (C79D&v7&v9&v12E);
assign Av13_D_9B = (C153D&v12E);
assign Av13_D_0B = (IIII71)|(IIII72)|(IIII73);
assign II692 = ((~Av13_D_10B));
assign C118D = (v2E)|(v10E);
assign IIII415 = (v8E&v11E&v12E);
assign C144DE = ((~C144D));
assign IIII475 = (v2E&v8&C138DE);
assign IIII278 = (v10E&C138DE);
assign C88D = (IIII259)|(IIII260);
assign IIII368 = (C30D&C90DE);
assign C83D = (v4E)|(v5E);
assign IIII105 = (v8&C113D);
assign IIII444 = (v3E&v9E);
assign II716 = ((~Av13_D_2B));
assign IIII359 = (v12E&C165DE);
assign C138D = (v11E)|(v12E);
assign IIII482 = (v2&C220DE);
assign C67D = (IIII160)|(IIII161);
assign IIII554 = (v2E&v8&v9E);
assign Av13_D_3B = (IIII34)|(IIII35)|(IIII36);
assign IIII72 = (C38D&v7E);
assign C215D = (IIII438)|(IIII439);
assign IIII210 = (v9&C120D);
assign IIII68 = (C206D&v12E);
assign IIII452 = (v12E&C220DE);
assign Av13_D_11B = (IIII140)|(IIII141)|(IIII142);
assign IIII406 = (v8&v11&C117DE);
assign IIII82 = (v0E&C217D&C108DE);
assign IIII227 = (C139D&v8&v10);
assign IIII213 = (C57D&v10E);
assign v13_D_10 = ((~II692));
assign v12E = ((~v12));
assign II114 = ((~v2));
assign C202D = (IIII272)|(IIII273);
assign II329 = (v3&v7E&v10);
assign IIII464 = (v8E&v10E&v11);
assign IIII245 = (C185D&v8E);
assign C78D = (IIII452)|(IIII453);
assign IIII157 = (C82D&v9E);
assign II142 = (v7E&v9&v11E);
assign C109D = (IIII338)|(IIII339);
assign IIII269 = (v11E&C108DE&C83DE);
assign C104D = (v1)|(v6E);
assign C167D = (IIII380)|(IIII381);
assign IIII310 = (v6E&v9&v12E&C124DE);
assign IIII317 = (v10&v11E);
assign C194DE = ((~C194D));
assign C184D = (IIII182)|(IIII183);
assign Av13_D_14B = (IIII78)|(IIII79)|(IIII80);
assign IIII297 = (C209D&C208D&v11);
assign II650 = ((~Av13_D_24B));
assign C169D = (IIII232)|(IIII233)|(v12)|(IIII234);
assign IIII435 = (v12&C165DE);
assign v13_D_24 = ((~II650));
assign C44D = (IIII473)|(C124DE);
assign IIII91 = (C148D&C131DE);
assign IIII329 = (v9&v12&C30D);
assign II707 = ((~Av13_D_5B));
assign IIII123 = (v8&C162D);
assign C180D = (C194DE)|(v11E);
assign IIII449 = (C108DE&C83DE);
assign II294 = ((~IIII352));
assign IIII342 = (C159D&v8E);
assign IIII360 = (v3E&C59D);
assign II246 = ((~v11));
assign IIII114 = (v9&C97D);
assign C42D = (IIII432)|(IIII433);
assign IIII302 = (v11E&C157DE);
assign C126D = (IIII239)|(IIII240);
assign IIII40 = (v2&C92D);
assign IIII282 = (C36D&v12);
assign Av13_D_24B = (IIII82)|(IIII83)|(IIII84);
assign C59D = (IIII537)|(IIII538);
assign C45D = (C90DE)|(v11E);
assign IIII79 = (v8&C170D);
assign v13_D_4C = (v13_D_4&CLR);
assign IIII212 = (v9E&C49DE);
assign C117D = (v9E)|(v2);
assign IIII386 = (v0&C104D&v8&C30DE);
assign II368 = (v7&v8&v9E);
assign v13_D_7 = ((~II701));
assign v2E = ((~v2));
assign IIII222 = (C156D&C83DE);
assign IIII501 = (v8E&v11E);
assign IIII71 = (v2E&C28D);
assign IIII483 = (v8E&v9E&v11E&C83DE);
assign IIII260 = (v3E&C78D);
assign IIII86 = (C54D&C165DE);
assign IIII92 = (v7&C140D);
assign C120D = (C144D)|(IIII425);
assign IIII470 = (v8&v12E&C83DE);
assign IIII117 = (v8E&C35D);
assign C48D = (IIII136)|(IIII137);
assign C188D = (IIII54)|(IIII55);
assign IIII58 = (C75D&C129DE);
assign C146D = (IIII398)|(IIII399);
assign IIII39 = (C103D&v10E);
assign IIII55 = (C187D&v12E);
assign IIII128 = (v8&C69D);
assign Av13_D_20B = (C138DE&C220DE&C104D&II329);
assign IIII95 = (C76D&C81DE);
assign IIII516 = (v1&v12);
assign IIII281 = (v3E&C29D);
assign IIII513 = (v12E&C166DE&II142);
assign C81DE = ((~C81D));
assign II722 = ((~Av13_D_0B));
assign C189D = (IIII362)|(IIII363);
assign IIII375 = (C86D&v10E);
assign IIII73 = (v7&C31D&v8);
assign IIII106 = (v8E&C114D);
assign C63D = (IIII317)|(IIII318);
assign IIII243 = (C131D&v9&C144DE);
assign IIII299 = (v11E&C108DE);
assign C100D = (IIII429)|(IIII430);
assign IIII311 = (C71D&v9E);
assign IIII148 = (v9&v10E&C144DE);
assign IIII31 = (C108DE&C83DE&II642);
assign C139D = (IIII332)|(IIII333);
assign IIII399 = (v8&C141D);
assign C115D = (IIII299)|(IIII300);
assign C186D = (C49DE)|(IIII245);
assign C191DE = ((~C191D));
assign C134D = (IIII163)|(IIII164);
assign IIII287 = (v9&v11);
assign IIII43 = (v8&v10&C108DE);
assign C102D = (IIII65)|(IIII66)|(II610);
assign C97D = ((~II373));
assign IIII341 = (v11E&C118DE);
assign IIII393 = ((~II143));
assign IIII420 = (v2E&v7&C131DE);
assign IIII48 = (C177D&v8E);
assign IIII390 = (C220D&v10E);
assign C54D = (C90DE)|(IIII412);
assign C30D = (v10E)|(v11E);
assign II491 = (IIII173)|(IIII174)|(IIII175);
assign IIII520 = (v3E&v6E);
assign C207D = (IIII68)|(IIII69);
assign IIII127 = (C73D&v10E);
assign C98D = (C144D)|(IIII444);
assign IIII170 = (v10&v11E);
assign C150D = ((~II294));
assign II683 = ((~Av13_D_13B));
assign II642 = (v7E&v8E&C124DE);
assign IIII196 = (C161D&v11);
assign IIII167 = (v8&v11&C129D);
assign C74D = (IIII129)|(IIII130)|(IIII131)|(II542);
assign IIII433 = (v10&C144DE);
assign IIII133 = (C152D&v9);
assign IIII339 = (v8E&C144DE);
assign C55D = (IIII475)|(IIII476);
assign C133D = (C49DE)|(IIII278);
assign v13_D_14 = ((~II680));
assign v13_D_1C = (v13_D_1&CLR);
assign v13_D_0 = ((~II722));
assign IIII275 = (v7&v8&C90DE);
assign IIII205 = (v8E&C30DE);
assign IIII186 = (v8&v11&C117DE);
assign IIII200 = (v12E&C124D);
assign IIII471 = (v1&v10E&v12);
assign C141D = (v10E)|(v12);
assign IIII116 = (C37D&v9);
assign Av13_D_10B = (IIII123)|(IIII124);
assign IIII280 = (v1E&C26D);
assign IIII308 = (C111D&C144DE);
assign IIII54 = (C186D&v9E);
assign IIII555 = (v0&v8E&v11);
assign v13_D_8 = ((~II698));
assign IIII389 = (v8&v9&v10);
assign C35D = (IIII202)|(IIII203);
assign v10E = ((~v10));
assign v7E = ((~v7));
assign v13_D_13 = ((~II683));
assign II653 = ((~Av13_D_23B));
assign IIII350 = (v11&C117D);
assign C220DE = ((~C220D));
assign C53D = (IIII151)|(IIII152)|(IIII153)|(IIII154);
assign C166D = (v3E)|(v6E);
assign IIII199 = (v9E&C63D);
assign IIII59 = (v7&C67D);
assign IIII146 = (C223D&v8E&v9E);
assign IIII262 = (C42D&v8);
assign IIII323 = (v10E&C127D);
assign IIII89 = (v7&C48D);
assign C201D = (IIII503)|(v12E);
assign II159 = ((~C83D));
assign IIII36 = (v7E&C89D);
assign IIII362 = (v8&C138DE);
assign Av13_D_8B = (IIII91)|(IIII92)|(IIII93);
assign IIII333 = (v11E&v12E);
assign IIII332 = (C138D&v9E);
assign IIII276 = (C27D&v7E&v9&v12E);
assign C77D = (C104D)|(v0E);
assign IIII242 = (C130D&C165DE);
assign IIII237 = (v7&v12E&C221D);
assign C43D = (IIII262)|(IIII263);
assign C200D = (IIII513)|(IIII514);
assign IIII378 = (C218D&v5E&v9&v12E);
assign C177D = (IIII75)|(IIII76);
assign C57D = (IIII365)|(IIII366);
assign II101 = ((~v9));
assign C56D = (v9)|(IIII516);
assign IIII326 = (C81DE&C129D);
assign IIII560 = (v7E&v12E);
assign IIII476 = (v8E&v9&v11E&v12E);
assign IIII414 = (v6&C138DE);
assign C220D = (v8E)|(v9E);
assign IIII169 = (C195D&v8E);
assign IIII450 = (v3&v8&C138DE&C104DE);
assign C129DE = ((~C129D));
assign IIII438 = (v0&v10&C144DE);
assign C218DE = ((~C218D));
assign C148D = (C90DE)|(IIII409);
assign IIII514 = (v2&v7&v9E&C138DE);
assign IIII247 = (v10&C144DE);
assign IIII119 = (C126D&v8);
assign Av13_D_2B = (IIII58)|(IIII59)|(IIII60);
assign IIII49 = (v8&C176D);
assign C179D = (v10)|(IIII518);
assign IIII495 = (v9&v11&C131DE);
assign C140D = (IIII226)|(IIII227);
assign IIII140 = (v8E&v10E&C144DE);
assign C31D = (IIII368)|(IIII369);
assign IIII432 = (v7&C90DE);
assign C49D = (C141D)|(v11);
assign IIII430 = (v1E&v9&v10E);
assign IIII171 = (v8&C193D);
assign v13_D_9 = ((~II695));
assign C187D = (IIII108)|(IIII109);
assign IIII80 = (v7&v12E&C192D);
assign IIII223 = (v7E&C160D&v9E);
assign IIII546 = (v0&v11);
assign C164D = (IIII222)|(IIII223)|(IIII224);
assign C221D = (IIII389)|(IIII390);
assign IIII441 = (v11&C220DE);
assign C180DE = ((~C180D));
assign v5E = ((~v5));
assign IIII160 = (v8&C65D);
assign v9E = ((~v9));
assign IIII402 = (v8&v9E&C30DE);
assign C70D = (v0)|(v11E);
assign C196D = (IIII170)|(v12)|(IIII171)|(II497);
assign IIII220 = (C51D&v12);
assign IIII478 = (v10E&C83DE);
assign IIII272 = (v10E&C144DE);
assign IIII137 = (v8&C46D);
assign Av13_D_17B = (IIII31)|(IIII32);
assign C116D = (IIII103)|(IIII104)|(IIII105)|(IIII106);
assign IIII384 = (v10E&C138DE);
assign C124D = (v10)|(v11);
assign C166DE = ((~C166D));
assign C176D = (IIII188)|(IIII189);
assign C137D = (C117DE)|(IIII489);
assign IIII97 = (C88D&v11E);
assign C142D = (v0)|(v12);
assign C46D = (IIII247)|(IIII248);
assign v13_D_16 = ((~II674));
assign IIII352 = (v8&C124D);
assign IIII369 = (v9&C124DE);
assign II497 = (C208DE)|(C83DE)|(IIII169);
assign C165D = (v8E)|(v11);
assign C73D = (IIII269)|(IIII270);
assign IIII372 = (C129D&v12E);
assign II674 = ((~Av13_D_16B));
assign C181D = (IIII185)|(IIII186);
assign C72D = (IIII310)|(IIII311);
assign IIII473 = (v0E&C30DE);
assign IIII131 = (v9&v11E&C157DE);
assign IIII446 = (v11E&C90DE);
assign C91D = (IIII346)|(IIII347);
assign IIII62 = (v6E&C95D);
assign IIII216 = (C189D&v9E);
assign IIII126 = (v2&C58D);
assign IIII45 = (C116D&v7E);
assign IIII392 = (C81D&v11E);
assign C217D = (IIII419)|(IIII420);
assign IIII395 = (C157D&v9E);
assign IIII423 = (v3E&C157DE);
assign v13_D_4 = ((~II710));
assign IIII234 = (v8&C167D);
assign IIII508 = (v9E&v11E);
assign IIII494 = (v8E&v10&C108DE);
assign IIII377 = (v7&v10&C90DE);
assign C39D = (IIII423)|(v9);
assign C144D = (v11E)|(v12);
assign Av13_D_6B = (IIII119)|(IIII120);
assign IIII64 = (v11E&C157DE);
assign IIII233 = (C168D&v8E);
assign IIII84 = (v7E&C224D);
assign C89D = (IIII95)|(IIII96)|(IIII97)|(IIII98);
assign Av13_D_22B = (IIII266)|(IIII267);
assign IIII439 = (v6&v12&C124DE);
assign IIII215 = (v1&v9&C144DE);
assign IIII285 = (C222D&v10E);
assign IIII503 = (v9E&C30DE);
assign C128D = (IIII405)|(IIII406);
assign IIII130 = (C60D&C83D);
assign C130D = (IIII371)|(IIII372);
assign C175D = (IIII325)|(IIII326);
assign IIII38 = (C102D&v7E);
assign IIII320 = (v11&C141D);
assign Av13_D_7B = (IIII51)|(IIII52);
assign C37D = (IIII280)|(IIII281)|(IIII282);
assign C47D = (IIII533)|(IIII534);
assign C28D = (IIII275)|(IIII276);
assign IIII305 = (v9&C49DE);
assign IIII528 = (v9E&v11);
assign IIII456 = (v9&C30DE);
assign II671 = ((~Av13_D_17B));
assign C191D = (v10E)|(v9);
assign IIII485 = (v6&C141DE&C220DE);
assign C113D = (IIII148)|(IIII149);
assign C135D = (IIII100)|(IIII101);
assign C118DE = ((~C118D));
assign C70DE = ((~C70D));
assign C112D = (IIII308)|(v9E);
assign Av13_D_21B = (C213D&v7E&v10E&v12E);
assign II695 = ((~Av13_D_9B));
assign v0E = ((~v0));
assign IIII96 = (v8&C85D);
assign v13_D_6 = ((~II704));
assign IIII396 = (v10E&v12E);
assign IIII180 = (C173D&v9E);
assign Av13_D_1B = (IIII86)|(IIII87)|(IIII88)|(IIII89);
assign C147D = (IIII176)|(IIII177)|(II491);
assign C195D = (C180DE)|(v9);
assign IIII153 = (C52D&v8E);
assign C87D = (IIII374)|(IIII375);
assign IIII256 = (v9&v10&C138DE);
assign IIII229 = (v9&v10&C144DE);
assign IIII447 = (v8E&v9&v10E&v12E);
assign IIII293 = (C138DE&C118DE&II368);
assign IIII87 = (C53D&v7E);
assign IIII463 = (C165DE&C191DE);
assign IIII291 = (C142D&v11);
assign IIII174 = (v8E&C143D);
assign C223D = (IIII284)|(IIII285);
assign C90DE = ((~C90D));
assign IIII76 = (v7E&C174D);
assign Av13_D_16B = (C200D&v8&v10);
assign Av13_D_5B = (IIII43)|(IIII44)|(IIII45)|(IIII46);
assign v13_D_3C = (v13_D_3&CLR);
assign IIII191 = (v8&v11&C117DE);
assign IIII240 = (C125D&v9E);
assign IIII425 = (v8E&v10E);
assign v11E = ((~v11));
assign IIII347 = (C90D&v10E);
assign II542 = (IIII126)|(IIII127)|(IIII128);
assign II668 = ((~Av13_D_18B));
assign IIII273 = (C201D&v8);
assign IIII154 = (v2&C40D);
assign IIII189 = (v7&v12E);
assign II548 = (C199D&v4&v5E);
assign IIII325 = (v10&C90DE);
assign IIII479 = (v0&v11);
assign IIII538 = (v8&v12E);
assign IIII173 = (C146D&v11E);
assign C157D = (v10E)|(v12E);
assign v8E = ((~v8));
assign IIII111 = (C98D&v10E);
assign IIII284 = (v11E&C157DE);
assign IIII419 = (v5E&v7E&v8E&C30DE);
assign Av13_D_18B = (C210D&v7E&v12E);
assign IIII239 = (v9&v12&C124DE);
assign IIII75 = (C129DE&C144DE);
assign IIII403 = (v9&v12E&C124DE&II254);
assign C214D = (IIII460)|(IIII461);
assign IIII166 = (C205D&v10);
assign C114D = (IIII456)|(IIII457);
assign II677 = ((~Av13_D_15B));
assign IIII52 = (C135D&v7E);
assign IIII103 = (C115D&v10);
assign IIII354 = (C191D&v11);
assign IIII44 = (v2E&C106D);
assign v13_D_15 = ((~II677));
assign IIII336 = (C124D&v12);
assign Av13_D_12B = (IIII48)|(IIII49);
assign IIII412 = (v3&v10E&v12E);
assign IIII109 = (C179D&v2&v8&v11);
assign IIII104 = (v3&C107D&v12);
assign C85D = (IIII156)|(IIII157)|(IIII158);
assign C71D = (IIII383)|(IIII384);
assign C173D = (IIII302)|(IIII303);
assign C209D = (IIII497)|(IIII498);
assign IIII270 = (v1E&C55D);
assign C162D = (IIII196)|(IIII197);
assign C117DE = ((~C117D));
assign IIII346 = (v12&C191DE);
assign IIII60 = (v7E&C74D);
assign C156D = (IIII441)|(IIII442);
assign C108D = (v9)|(v12);
assign C75D = (IIII359)|(IIII360);
assign II373 = ((~IIII194));
assign II680 = ((~Av13_D_14B));
assign IIII457 = (v6&C124DE&C90DE);
assign C79D = ((~II246));
assign C93D = (C191DE)|(IIII468);
assign C81D = (v2E)|(v12);
assign C145D = (IIII528)|(v12);
assign C84D = (C138DE)|(IIII344);
assign IIII232 = (C165D&C83DE);
assign Av13_D_15B = (v7E&v12E&II548);
assign IIII306 = (C129DE&C138D);
assign II254 = (v1&v6&v7E&v8E);
assign IIII383 = (C70D&C141DE);
assign C111D = (C83DE)|(v2);
assign C163D = (C129DE)|(IIII510);
assign C108DE = ((~C108D));
assign IIII32 = (C207D&v2);
assign IIII315 = (C155D&v12E&C129D);
assign IIII380 = (v2&v11);
assign IIII192 = (v8E&v9E&C44D);
assign II665 = ((~Av13_D_19B));
assign C80D = (IIII250)|(IIII251);
assign C203D = (C70DE)|(IIII508);
assign C36D = (C165DE)|(v10E);
assign C129D = (v9)|(v10);
assign C151D = (IIII554)|(IIII555);
assign C95D = (IIII446)|(IIII447);
assign v1E = ((~v1));
assign IIII163 = (v11E&v12E&C118DE);
assign v13_D_12 = ((~II686));
assign IIII100 = (C134D&v9E);
assign C125D = (IIII335)|(IIII336);
assign IIII179 = (v9&v10&C144DE);
assign IIII208 = (C122D&v11E);
assign C40D = (IIII253)|(IIII254);
assign C183D = (IIII305)|(IIII306);
assign Av13_D_4B = (IIII38)|(IIII39)|(IIII40)|(IIII41);
assign C143D = (C49DE)|(v9)|(IIII291);
assign IIII136 = (C47D&C144DE);
assign IIII492 = (v10&v11E);
assign IIII363 = (v1E&C178D);
assign IIII250 = (C77D&v3&C138DE);
assign v13_D_0C = (v13_D_0&CLR);
assign C155D = (v2)|(v7);
assign IIII524 = (v6&v11E);
assign C58D = (IIII212)|(IIII213);
assign IIII453 = (v10E&v12);
assign IIII328 = (v3&v12E&C124DE);
assign IIII224 = (C163D&v8E&v11);
assign IIII338 = (C108D&C165DE);
assign C30DE = ((~C30D));
assign C165DE = ((~C165D));
assign IIII460 = (v2E&v12E&C165DE);
assign IIII113 = (v2E&v12E&C93D);
assign IIII142 = (v7E&C169D);
assign C193D = ((~II114));
assign C218D = (v7E)|(v10);
assign C178D = (IIII559)|(IIII560);
assign IIII63 = (v8&C99D);
assign C65D = (IIII199)|(IIII200);
assign IIII259 = (v12E&C129DE&C83DE);
assign v13_D_2 = ((~II716));
assign v13_D_11 = ((~II689));
assign C174D = (IIII179)|(IIII180);
assign IIII66 = (v8E&v12E&C100D);
assign IIII185 = (v8E&C195DE);
assign C216D = (IIII256)|(IIII257);
assign IIII202 = (v9E&C144DE&C83DE&C194DE);
assign C222D = (C138DE)|(IIII417);
assign II710 = ((~Av13_D_4B));
assign IIII510 = (v9&v10);
assign C131D = (v8E)|(v10);
assign IIII124 = (C164D&v12E);
assign IIII164 = (C133D&v8E);
assign IIII505 = (v7&v8&C138DE&C191DE);
assign C225D = (IIII236)|(IIII237);
assign C157DE = ((~C157D));
assign IIII251 = (v6E&v11E&v12E);
assign C92D = (IIII505)|(IIII506);
assign IIII182 = (v8E&v10E&C144DE);
assign C106D = (IIII402)|(IIII403);
assign IIII152 = (v8&v12E&C129DE);
assign IIII537 = (v6E&v7E&v8E&v12);
assign II143 = ((~v10E));
assign II701 = ((~Av13_D_7B));
assign C206D = (IIII166)|(IIII167);
assign IIII218 = (v12E&C44D&C83DE);
assign IIII158 = (C84D&v10E);
assign C83DE = ((~C83D));
assign C50D = (IIII520)|(v11);
assign IIII335 = (v12E&C218DE);
assign IIII294 = (C211D&v3&v7E&v11E);
assign IIII51 = (C132D&v7);
assign C170D = (C124DE)|(v9E);
assign IIII398 = (v12E&C118DE);
assign v13_D_22 = ((~II656));
assign IIII175 = (v9&C144D);
assign v13_D_18 = ((~II668));
assign IIII149 = (C112D&v10);
assign IIII436 = (v8E&v9&C144DE);
assign II656 = ((~Av13_D_22B));
assign IIII29 = (C190D&v10);
assign C205D = (IIII287)|(IIII288);
assign IIII417 = (v5E&v11E&v12E);
assign IIII156 = (C80D&v9);
assign C195DE = ((~C195D));
assign C122D = (v12)|(IIII323);
assign C96D = (IIII463)|(IIII464);
assign C52D = (IIII218)|(IIII219)|(IIII220);
assign IIII257 = (C215D&v9E);
assign C51D = (IIII356)|(IIII357);
assign IIII101 = (C127D&C128D&v12E);
assign C211D = (IIII485)|(IIII486);
assign IIII374 = (v9E&C30DE);
assign II698 = ((~Av13_D_8B));
assign IIII176 = (v10E&C145D);
assign II610 = (IIII62)|(IIII63)|(IIII64);
assign C194D = (v0)|(v10E);
assign C69D = (IIII328)|(IIII329);
assign C141DE = ((~C141D));
assign IIII461 = (v8E&v9&v12);
assign IIII486 = (v6E&v8E&v12&C129DE);
assign IIII357 = (v10&v11E);
assign v6E = ((~v6));
assign IIII266 = (v7&C49DE&C220DE);
assign C224D = (IIII145)|(IIII146);
assign C158D = (IIII395)|(IIII396);
assign IIII248 = (C45D&v10E);
assign IIII371 = (v10E&C90DE);
assign C213D = (IIII482)|(IIII483);
assign IIII219 = (C49D&v9);
assign IIII314 = (v10&C90DE);
assign C132D = (IIII242)|(IIII243);
assign IIII194 = (v3&v12&C77D);
assign v13_D_5C = (v13_D_5&CLR);
assign C107D = (IIII386)|(IIII387);
assign C152D = (IIII205)|(IIII206);
assign IIII356 = (C50D&v10E);
assign C34D = (IIII320)|(IIII321);
assign IIII344 = ((~II159));
assign IIII78 = (v7E&C196D);
assign C159D = (IIII546)|(IIII547);
assign IIII366 = (v8E&v9&v11E&v12E);
assign IIII427 = (v8E&v9&v10);
assign C138DE = ((~C138D));
assign C103D = (IIII435)|(IIII436);
assign IIII381 = (C166D&v11E);
assign C49DE = ((~C49D));
assign C190D = (IIII215)|(IIII216);
assign IIII497 = (v8E&v9E&C194DE);
assign IIII46 = (v7&C110D);
assign IIII120 = (v7E&C123D);
assign v13_D_17 = ((~II671));
assign v13_D_3 = ((~II713));
assign C219D = (IIII377)|(IIII378);
assign II719 = ((~Av13_D_1B));
assign IIII254 = (C39D&v8E);
assign C60D = (IIII494)|(IIII495);
assign IIII183 = (C183D&v8);
assign IIII65 = (v9&C185D);
assign v13_D_21 = ((~II659));
assign C192D = (v8)|(IIII354);
assign IIII559 = (v8&v11);
assign IIII141 = (C170D&v8);
assign IIII491 = (v10E&C138DE);
assign II713 = ((~Av13_D_3B));
assign II662 = ((~Av13_D_20B));
assign IIII206 = (v7&C150D);
assign C210D = (IIII296)|(IIII297);
assign IIII349 = (C118D&v11E);
assign C208DE = ((~C208D));
assign C208D = (v5)|(v4);
assign IIII230 = (C109D&v10E);
assign C33D = (v6E)|(v10);
assign C127D = (v5E)|(v4);
assign C41D = (IIII470)|(IIII471);
assign IIII209 = (v8&C119D);
assign IIII466 = (v8E&v11E&v12E);
assign v13_D_5 = ((~II707));
assign IIII303 = (C172D&v12E);
assign Av13_D_19B = (IIII293)|(IIII294);
endmodule
