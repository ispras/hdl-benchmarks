module test ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , 
 n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , 
 n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , 
 n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , 
 n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , 
 n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , 
 n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , 
 n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , 
 n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , 
 n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , 
 n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , 
 n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , 
 n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , 
 n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , 
 n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , 
 n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , 
 n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , 
 n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , 
 n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , 
 n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , 
 n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , 
 n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , 
 n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , 
 n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , 
 n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , 
 n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , 
 n381 , n382 , n383 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , 
 n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , 
 n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , 
 n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , 
 n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , 
 n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , 
 n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , 
 n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , 
 n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , 
 n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , 
 n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , 
 n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , 
 n121 , n122 , n123 , n124 , n125 , n126 , n127 ;
output n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , 
 n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , 
 n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , 
 n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , 
 n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , 
 n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , 
 n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , 
 n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , 
 n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , 
 n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , 
 n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , 
 n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , 
 n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , 
 n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , 
 n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , 
 n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , 
 n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , 
 n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , 
 n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , 
 n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , 
 n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , 
 n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , 
 n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , 
 n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , 
 n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , 
 n379 , n380 , n381 , n382 , n383 ;
wire n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , 
 n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , 
 n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , 
 n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , 
 n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , 
 n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , 
 n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , 
 n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , 
 n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , 
 n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , 
 n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , 
 n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , 
 n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , 
 n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , 
 n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , 
 n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , 
 n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , 
 n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , 
 n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , 
 n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , 
 n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , 
 n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , 
 n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , 
 n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , 
 n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , 
 n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , 
 n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , 
 n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , 
 n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , 
 n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , 
 n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , 
 n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , 
 n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , 
 n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , 
 n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , 
 n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , 
 n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , 
 n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , 
 n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , 
 n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , 
 n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , 
 n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , 
 n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , 
 n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , 
 n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , 
 n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , 
 n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , 
 n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , 
 n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , 
 n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , 
 n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , 
 n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , 
 n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , 
 n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , 
 n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , 
 n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , 
 n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , 
 n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , 
 n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , 
 n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , 
 n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , 
 n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , 
 n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , 
 n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , 
 n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , 
 n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , 
 n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , 
 n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , 
 n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , 
 n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , 
 n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , 
 n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , 
 n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , 
 n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , 
 n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , 
 n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , 
 n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , 
 n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , 
 n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , 
 n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , 
 n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , 
 n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , 
 n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , 
 n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , 
 n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , 
 n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , 
 n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , 
 n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , 
 n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , 
 n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , 
 n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , 
 n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , 
 n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , 
 n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , 
 n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , 
 n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , 
 n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , 
 n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , 
 n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , 
 n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , 
 n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , 
 n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , 
 n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , 
 n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , 
 n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , 
 n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , 
 n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , 
 n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , 
 n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , 
 n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , 
 n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , 
 n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , 
 n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , 
 n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , 
 n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , 
 n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , 
 n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , 
 n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , 
 n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , 
 n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , 
 n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , 
 n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , 
 n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , 
 n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , 
 n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , 
 n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , 
 n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , 
 n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , 
 n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , 
 n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , 
 n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , 
 n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , 
 n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , 
 n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , 
 n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , 
 n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , 
 n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , 
 n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , 
 n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , 
 n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , 
 n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , 
 n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , 
 n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , 
 n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , 
 n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , 
 n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , 
 n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , 
 n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , 
 n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , 
 n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , 
 n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , 
 n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , 
 n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , 
 n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , 
 n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , 
 n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , 
 n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , 
 n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , 
 n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , 
 n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , 
 n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , 
 n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , 
 n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , 
 n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , 
 n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , 
 n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , 
 n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , 
 n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , 
 n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , 
 n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , 
 n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , 
 n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , 
 n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , 
 n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , 
 n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , 
 n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , 
 n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , 
 n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , 
 n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , 
 n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , 
 n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , 
 n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , 
 n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , 
 n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , 
 n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , 
 n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , 
 n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , 
 n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , 
 n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , 
 n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , 
 n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , 
 n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , 
 n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , 
 n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , 
 n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , 
 n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , 
 n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , 
 n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , 
 n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , 
 n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , 
 n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , 
 n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , 
 n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , 
 n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , 
 n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , 
 n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , 
 n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , 
 n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , 
 n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , 
 n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , 
 n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , 
 n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , 
 n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , 
 n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , 
 n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , 
 n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , 
 n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , 
 n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , 
 n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , 
 n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , 
 n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , 
 n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , 
 n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , 
 n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , 
 n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , 
 n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , 
 n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , 
 n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , 
 n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , 
 n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , 
 n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , 
 n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , 
 n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , 
 n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , 
 n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , 
 n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , 
 n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , 
 n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , 
 n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , 
 n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , 
 n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , 
 n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , 
 n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , 
 n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , 
 n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , 
 n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , 
 n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , 
 n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , 
 n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , 
 n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , 
 n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , 
 n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , 
 n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , 
 n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , 
 n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , 
 n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , 
 n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , 
 n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , 
 n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , 
 n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , 
 n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , 
 n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , 
 n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , 
 n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , 
 n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , 
 n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , 
 n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , 
 n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , 
 n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , 
 n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , 
 n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , 
 n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , 
 n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , 
 n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , 
 n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , 
 n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , 
 n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , 
 n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , 
 n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , 
 n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , 
 n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , 
 n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , 
 n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , 
 n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , 
 n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , 
 n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , 
 n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , 
 n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , 
 n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , 
 n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , 
 n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , 
 n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , 
 n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , 
 n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , 
 n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , 
 n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , 
 n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , 
 n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , 
 n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , 
 n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , 
 n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , 
 n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , 
 n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , 
 n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , 
 n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , 
 n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , 
 n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , 
 n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , 
 n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , 
 n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , 
 n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , 
 n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , 
 n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , 
 n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , 
 n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , 
 n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , 
 n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , 
 n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , 
 n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , 
 n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , 
 n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , 
 n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , 
 n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , 
 n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , 
 n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , 
 n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , 
 n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , 
 n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , 
 n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , 
 n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , 
 n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , 
 n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , 
 n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , 
 n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , 
 n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , 
 n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , 
 n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , 
 n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , 
 n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , 
 n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , 
 n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , 
 n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , 
 n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , 
 n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , 
 n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , 
 n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , 
 n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , 
 n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , 
 n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , 
 n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , 
 n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , 
 n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , 
 n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , 
 n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , 
 n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , 
 n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , 
 n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , 
 n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , 
 n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , 
 n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , 
 n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , 
 n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , 
 n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , 
 n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , 
 n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , 
 n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , 
 n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , 
 n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , 
 n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , 
 n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , 
 n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , 
 n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , 
 n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , 
 n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , 
 n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , 
 n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , 
 n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , 
 n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , 
 n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , 
 n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , 
 n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , 
 n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , 
 n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , 
 n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , 
 n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , 
 n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , 
 n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , 
 n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , 
 n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , 
 n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , 
 n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , 
 n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , 
 n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , 
 n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , 
 n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , 
 n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , 
 n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , 
 n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , 
 n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , 
 n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , 
 n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , 
 n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , 
 n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , 
 n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , 
 n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , 
 n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , 
 n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , 
 n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , 
 n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , 
 n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , 
 n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , 
 n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , 
 n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , 
 n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , 
 n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , 
 n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , 
 n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , 
 n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , 
 n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , 
 n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , 
 n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , 
 n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , 
 n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , 
 n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , 
 n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , 
 n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , 
 n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , 
 n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , 
 n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , 
 n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , 
 n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , 
 n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , 
 n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , 
 n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , 
 n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , 
 n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , 
 n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , 
 n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , 
 n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , 
 n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , 
 n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , 
 n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , 
 n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , 
 n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , 
 n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , 
 n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , 
 n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , 
 n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , 
 n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , 
 n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , 
 n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , 
 n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , 
 n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , 
 n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , 
 n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , 
 n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , 
 n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , 
 n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , 
 n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , 
 n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , 
 n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , 
 n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , 
 n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , 
 n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , 
 n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , 
 n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , 
 n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , 
 n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , 
 n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , 
 n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , 
 n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , 
 n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , 
 n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , 
 n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , 
 n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , 
 n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , 
 n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , 
 n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , 
 n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , 
 n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , 
 n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , 
 n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , 
 n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , 
 n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , 
 n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , 
 n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , 
 n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , 
 n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , 
 n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , 
 n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , 
 n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , 
 n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , 
 n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , 
 n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , 
 n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , 
 n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , 
 n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , 
 n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , 
 n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , 
 n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , 
 n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , 
 n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , 
 n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , 
 n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , 
 n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , 
 n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , 
 n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , 
 n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , 
 n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , 
 n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , 
 n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , 
 n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , 
 n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , 
 n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , 
 n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , 
 n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , 
 n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , 
 n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , 
 n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , 
 n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , 
 n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , 
 n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , 
 n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , 
 n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , 
 n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , 
 n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , 
 n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , 
 n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , 
 n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , 
 n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , 
 n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , 
 n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , 
 n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , 
 n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , 
 n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , 
 n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , 
 n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , 
 n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , 
 n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , 
 n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , 
 n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , 
 n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , 
 n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , 
 n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , 
 n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , 
 n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , 
 n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , 
 n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , 
 n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , 
 n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , 
 n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , 
 n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , 
 n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , 
 n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , 
 n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , 
 n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , 
 n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , 
 n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , 
 n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , 
 n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , 
 n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , 
 n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , 
 n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , 
 n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , 
 n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , 
 n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , 
 n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , 
 n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , 
 n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , 
 n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , 
 n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , 
 n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , 
 n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , 
 n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , 
 n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , 
 n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , 
 n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , 
 n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , 
 n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , 
 n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , 
 n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , 
 n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , 
 n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , 
 n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , 
 n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , 
 n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , 
 n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , 
 n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , 
 n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , 
 n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , 
 n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , 
 n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , 
 n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , 
 n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , 
 n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , 
 n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , 
 n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , 
 n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , 
 n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , 
 n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , 
 n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , 
 n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , 
 n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , 
 n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , 
 n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , 
 n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , 
 n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , 
 n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , 
 n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , 
 n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , 
 n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , 
 n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , 
 n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , 
 n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , 
 n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , 
 n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , 
 n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , 
 n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , 
 n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , 
 n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , 
 n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , 
 n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , 
 n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , 
 n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , 
 n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , 
 n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , 
 n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , 
 n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , 
 n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , 
 n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , 
 n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , 
 n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , 
 n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , 
 n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , 
 n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , 
 n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , 
 n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , 
 n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , 
 n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , 
 n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , 
 n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , 
 n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , 
 n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , 
 n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , 
 n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , 
 n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , 
 n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , 
 n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , 
 n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , 
 n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , 
 n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , 
 n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , 
 n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , 
 n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , 
 n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , 
 n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , 
 n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , 
 n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , 
 n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , 
 n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , 
 n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , 
 n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , 
 n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , 
 n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , 
 n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , 
 n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , 
 n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , 
 n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , 
 n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , 
 n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , 
 n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , 
 n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , 
 n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , 
 n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , 
 n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , 
 n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , 
 n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , 
 n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , 
 n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , 
 n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , 
 n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , 
 n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , 
 n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , 
 n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , 
 n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , 
 n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , 
 n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , 
 n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , 
 n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , 
 n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , 
 n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , 
 n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , 
 n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , 
 n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , 
 n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , 
 n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , 
 n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , 
 n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , 
 n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , 
 n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , 
 n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , 
 n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , 
 n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , 
 n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , 
 n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , 
 n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , 
 n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , 
 n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , 
 n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , 
 n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , 
 n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , 
 n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , 
 n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , 
 n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , 
 n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , 
 n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , 
 n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , 
 n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , 
 n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , 
 n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , 
 n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , 
 n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , 
 n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , 
 n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , 
 n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , 
 n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , 
 n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , 
 n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , 
 n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , 
 n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , 
 n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , 
 n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , 
 n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , 
 n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , 
 n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , 
 n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , 
 n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , 
 n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , 
 n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , 
 n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , 
 n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , 
 n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , 
 n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , 
 n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , 
 n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , 
 n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , 
 n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , 
 n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , 
 n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , 
 n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , 
 n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , 
 n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , 
 n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , 
 n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , 
 n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , 
 n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , 
 n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , 
 n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , 
 n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , 
 n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , 
 n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , 
 n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , 
 n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , 
 n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , 
 n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , 
 n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , 
 n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , 
 n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , 
 n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , 
 n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , 
 n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , 
 n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , 
 n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , 
 n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , 
 n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , 
 n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , 
 n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , 
 n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , 
 n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , 
 n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , 
 n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , 
 n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , 
 n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , 
 n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , 
 n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , 
 n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , 
 n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , 
 n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , 
 n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , 
 n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , 
 n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , 
 n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , 
 n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , 
 n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , 
 n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , 
 n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , 
 n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , 
 n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , 
 n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , 
 n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , 
 n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , 
 n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , 
 n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , 
 n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , 
 n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , 
 n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , 
 n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , 
 n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , 
 n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , 
 n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , 
 n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , 
 n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , 
 n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , 
 n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , 
 n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , 
 n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , 
 n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , 
 n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , 
 n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , 
 n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , 
 n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , 
 n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , 
 n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , 
 n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , 
 n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , 
 n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , 
 n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , 
 n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , 
 n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , 
 n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , 
 n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , 
 n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , 
 n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , 
 n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , 
 n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , 
 n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , 
 n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , 
 n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , 
 n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , 
 n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , 
 n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , 
 n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , 
 n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , 
 n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , 
 n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , 
 n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , 
 n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , 
 n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , 
 n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , 
 n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , 
 n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , 
 n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , 
 n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , 
 n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , 
 n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , 
 n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , 
 n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , 
 n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , 
 n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , 
 n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , 
 n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , 
 n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , 
 n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , 
 n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , 
 n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , 
 n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , 
 n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , 
 n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , 
 n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , 
 n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , 
 n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , 
 n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , 
 n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , 
 n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , 
 n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , 
 n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , 
 n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , 
 n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , 
 n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , 
 n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , 
 n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , 
 n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , 
 n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , 
 n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , 
 n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , 
 n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , 
 n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , 
 n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , 
 n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , 
 n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , 
 n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , 
 n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , 
 n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , 
 n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , 
 n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , 
 n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , 
 n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , 
 n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , 
 n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , 
 n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , 
 n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , 
 n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , 
 n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , 
 n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , 
 n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , 
 n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , 
 n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , 
 n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , 
 n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , 
 n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , 
 n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , 
 n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , 
 n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , 
 n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , 
 n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , 
 n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , 
 n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , 
 n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , 
 n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , 
 n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , 
 n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , 
 n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , 
 n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , 
 n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , 
 n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , 
 n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , 
 n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , 
 n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , 
 n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , 
 n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , 
 n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , 
 n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , 
 n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , 
 n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , 
 n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , 
 n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , 
 n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , 
 n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , 
 n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , 
 n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , 
 n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , 
 n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , 
 n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , 
 n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , 
 n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , 
 n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , 
 n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , 
 n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , 
 n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , 
 n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , 
 n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , 
 n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , 
 n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , 
 n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , 
 n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , 
 n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , 
 n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , 
 n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , 
 n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , 
 n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , 
 n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , 
 n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , 
 n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , 
 n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , 
 n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , 
 n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , 
 n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , 
 n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , 
 n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , 
 n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , 
 n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , 
 n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , 
 n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , 
 n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , 
 n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , 
 n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , 
 n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , 
 n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , 
 n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , 
 n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , 
 n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , 
 n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , 
 n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , 
 n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , 
 n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , 
 n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , 
 n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , 
 n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , 
 n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , 
 n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , 
 n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , 
 n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , 
 n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , 
 n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , 
 n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , 
 n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , 
 n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , 
 n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , 
 n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , 
 n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , 
 n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , 
 n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , 
 n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , 
 n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , 
 n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , 
 n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , 
 n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , 
 n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , 
 n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , 
 n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , 
 n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , 
 n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , 
 n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , 
 n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , 
 n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , 
 n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , 
 n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , 
 n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , 
 n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , 
 n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , 
 n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , 
 n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , 
 n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , 
 n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , 
 n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , 
 n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , 
 n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , 
 n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , 
 n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , 
 n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , 
 n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , 
 n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , 
 n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , 
 n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , 
 n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , 
 n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , 
 n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , 
 n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , 
 n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , 
 n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , 
 n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , 
 n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , 
 n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , 
 n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , 
 n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , 
 n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , 
 n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , 
 n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , 
 n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , 
 n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , 
 n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , 
 n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , 
 n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , 
 n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , 
 n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , 
 n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , 
 n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , 
 n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , 
 n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , 
 n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , 
 n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , 
 n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , 
 n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , 
 n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , 
 n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , 
 n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , 
 n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , 
 n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , 
 n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , 
 n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , 
 n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , 
 n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , 
 n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , 
 n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , 
 n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , 
 n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , 
 n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , 
 n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , 
 n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , 
 n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , 
 n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , 
 n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , 
 n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , 
 n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , 
 n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , 
 n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , 
 n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , 
 n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , 
 n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , 
 n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , 
 n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , 
 n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , 
 n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , 
 n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , 
 n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , 
 n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , 
 n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , 
 n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , 
 n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , 
 n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , 
 n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , 
 n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , 
 n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , 
 n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , 
 n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , 
 n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , 
 n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , 
 n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , 
 n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , 
 n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , 
 n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , 
 n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , 
 n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , 
 n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , 
 n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , 
 n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , 
 n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , 
 n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , 
 n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , 
 n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , 
 n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , 
 n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , 
 n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , 
 n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , 
 n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , 
 n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , 
 n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , 
 n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , 
 n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , 
 n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , 
 n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , 
 n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , 
 n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , 
 n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , 
 n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , 
 n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , 
 n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , 
 n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , 
 n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , 
 n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , 
 n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , 
 n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , 
 n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , 
 n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , 
 n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , 
 n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , 
 n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , 
 n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , 
 n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , 
 n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , 
 n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , 
 n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , 
 n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , 
 n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , 
 n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , 
 n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , 
 n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , 
 n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , 
 n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , 
 n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , 
 n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , 
 n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , 
 n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , 
 n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , 
 n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , 
 n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , 
 n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , 
 n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , 
 n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , 
 n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , 
 n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , 
 n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , 
 n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , 
 n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , 
 n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , 
 n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , 
 n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , 
 n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , 
 n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , 
 n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , 
 n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , 
 n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , 
 n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , 
 n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , 
 n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , 
 n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , 
 n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , 
 n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , 
 n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , 
 n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , 
 n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , 
 n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , 
 n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , 
 n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , 
 n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , 
 n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , 
 n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , 
 n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , 
 n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , 
 n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , 
 n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , 
 n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , 
 n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , 
 n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , 
 n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , 
 n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , 
 n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , 
 n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , 
 n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , 
 n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , 
 n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , 
 n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , 
 n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , 
 n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , 
 n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , 
 n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , 
 n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , 
 n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , 
 n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , 
 n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , 
 n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , 
 n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , 
 n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , 
 n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , 
 n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , 
 n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , 
 n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , 
 n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , 
 n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , 
 n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , 
 n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , 
 n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , 
 n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , 
 n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , 
 n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , 
 n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , 
 n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , 
 n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , 
 n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , 
 n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , 
 n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , 
 n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , 
 n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , 
 n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , 
 n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , 
 n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , 
 n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , 
 n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , 
 n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , 
 n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , 
 n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , 
 n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , 
 n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , 
 n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , 
 n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , 
 n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , 
 n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , 
 n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , 
 n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , 
 n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , 
 n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , 
 n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , 
 n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , 
 n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , 
 n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , 
 n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , 
 n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , 
 n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , 
 n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , 
 n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , 
 n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , 
 n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , 
 n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , 
 n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , 
 n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , 
 n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , 
 n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , 
 n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , 
 n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , 
 n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , 
 n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , 
 n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , 
 n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , 
 n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , 
 n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , 
 n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , 
 n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , 
 n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , 
 n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , 
 n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , 
 n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , 
 n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , 
 n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , 
 n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , 
 n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , 
 n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , 
 n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , 
 n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , 
 n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , 
 n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , 
 n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , 
 n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , 
 n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , 
 n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , 
 n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , 
 n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , 
 n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , 
 n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , 
 n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , 
 n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , 
 n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , 
 n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , 
 n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , 
 n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , 
 n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , 
 n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , 
 n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , 
 n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , 
 n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , 
 n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , 
 n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , 
 n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , 
 n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , 
 n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , 
 n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , 
 n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , 
 n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , 
 n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , 
 n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , 
 n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , 
 n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , 
 n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , 
 n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , 
 n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , 
 n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , 
 n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , 
 n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , 
 n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , 
 n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , 
 n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , 
 n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , 
 n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , 
 n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , 
 n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , 
 n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , 
 n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , 
 n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , 
 n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , 
 n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , 
 n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , 
 n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , 
 n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , 
 n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , 
 n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , 
 n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , 
 n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , 
 n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , 
 n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , 
 n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , 
 n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , 
 n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , 
 n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , 
 n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , 
 n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , 
 n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , 
 n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , 
 n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , 
 n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , 
 n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , 
 n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , 
 n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , 
 n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , 
 n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , 
 n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , 
 n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , 
 n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , 
 n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , 
 n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , 
 n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , 
 n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , 
 n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , 
 n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , 
 n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , 
 n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , 
 n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , 
 n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , 
 n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , 
 n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , 
 n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , 
 n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , 
 n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , 
 n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , 
 n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , 
 n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , 
 n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , 
 n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , 
 n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , 
 n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , 
 n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , 
 n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , 
 n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , 
 n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , 
 n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , 
 n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , 
 n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , 
 n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , 
 n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , 
 n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , 
 n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , 
 n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , 
 n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , 
 n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , 
 n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , 
 n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , 
 n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , 
 n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , 
 n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , 
 n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , 
 n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , 
 n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , 
 n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , 
 n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , 
 n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , 
 n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , 
 n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , 
 n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , 
 n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , 
 n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , 
 n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , 
 n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , 
 n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , 
 n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , 
 n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , 
 n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , 
 n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , 
 n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , 
 n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , 
 n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , 
 n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , 
 n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , 
 n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , 
 n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , 
 n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , 
 n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , 
 n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , 
 n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , 
 n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , 
 n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , 
 n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , 
 n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , 
 n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , 
 n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , 
 n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , 
 n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , 
 n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , 
 n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , 
 n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , 
 n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , 
 n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , 
 n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , 
 n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , 
 n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , 
 n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , 
 n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , 
 n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , 
 n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , 
 n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , 
 n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , 
 n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , 
 n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , 
 n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , 
 n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , 
 n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , 
 n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , 
 n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , 
 n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , 
 n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , 
 n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , 
 n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , 
 n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , 
 n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , 
 n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , 
 n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , 
 n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , 
 n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , 
 n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , 
 n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , 
 n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , 
 n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , 
 n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , 
 n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , 
 n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , 
 n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , 
 n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , 
 n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , 
 n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , 
 n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , 
 n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , 
 n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , 
 n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , 
 n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , 
 n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , 
 n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , 
 n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , 
 n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , 
 n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , 
 n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , 
 n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , 
 n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , 
 n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , 
 n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , 
 n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , 
 n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , 
 n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , 
 n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , 
 n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , 
 n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , 
 n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , 
 n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , 
 n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , 
 n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , 
 n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , 
 n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , 
 n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , 
 n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , 
 n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , 
 n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , 
 n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , 
 n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , 
 n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , 
 n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , 
 n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , 
 n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , 
 n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , 
 n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , 
 n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , 
 n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , 
 n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , 
 n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , 
 n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , 
 n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , 
 n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , 
 n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , 
 n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , 
 n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , 
 n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , 
 n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , 
 n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , 
 n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , 
 n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , 
 n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , 
 n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , 
 n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , 
 n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , 
 n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , 
 n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , 
 n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , 
 n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , 
 n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , 
 n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , 
 n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , 
 n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , 
 n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , 
 n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , 
 n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , 
 n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , 
 n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , 
 n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , 
 n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , 
 n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , 
 n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , 
 n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , 
 n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , 
 n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , 
 n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , 
 n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , 
 n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , 
 n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , 
 n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , 
 n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , 
 n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , 
 n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , 
 n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , 
 n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , 
 n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , 
 n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , 
 n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , 
 n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , 
 n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , 
 n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , 
 n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , 
 n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , 
 n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , 
 n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , 
 n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , 
 n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , 
 n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , 
 n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , 
 n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , 
 n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , 
 n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , 
 n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , 
 n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , 
 n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , 
 n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , 
 n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , 
 n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , 
 n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , 
 n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , 
 n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , 
 n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , 
 n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , 
 n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , 
 n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , 
 n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , 
 n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , 
 n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , 
 n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , 
 n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , 
 n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , 
 n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , 
 n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , 
 n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , 
 n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , 
 n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , 
 n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , 
 n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , 
 n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , 
 n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , 
 n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , 
 n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , 
 n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , 
 n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , 
 n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , 
 n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , 
 n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , 
 n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , 
 n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , 
 n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , 
 n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , 
 n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , 
 n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , 
 n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , 
 n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , 
 n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , 
 n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , 
 n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , 
 n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , 
 n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , 
 n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , 
 n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , 
 n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , 
 n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , 
 n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , 
 n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , 
 n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , 
 n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , 
 n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , 
 n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , 
 n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , 
 n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , 
 n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , 
 n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , 
 n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , 
 n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , 
 n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , 
 n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , 
 n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , 
 n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , 
 n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , 
 n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , 
 n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , 
 n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , 
 n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , 
 n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , 
 n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , 
 n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , 
 n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , 
 n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , 
 n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , 
 n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , 
 n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , 
 n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , 
 n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , 
 n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , 
 n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , 
 n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , 
 n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , 
 n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , 
 n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , 
 n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , 
 n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , 
 n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , 
 n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , 
 n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , 
 n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , 
 n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , 
 n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , 
 n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , 
 n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , 
 n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , 
 n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , 
 n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , 
 n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , 
 n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , 
 n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , 
 n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , 
 n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , 
 n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , 
 n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , 
 n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , 
 n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , 
 n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , 
 n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , 
 n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , 
 n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , 
 n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , 
 n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , 
 n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , 
 n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , 
 n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , 
 n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , 
 n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , 
 n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , 
 n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , 
 n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , 
 n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , 
 n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , 
 n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , 
 n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , 
 n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , 
 n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , 
 n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , 
 n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , 
 n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , 
 n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , 
 n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , 
 n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , 
 n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , 
 n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , 
 n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , 
 n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , 
 n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , 
 n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , 
 n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , 
 n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , 
 n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , 
 n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , 
 n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , 
 n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , 
 n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , 
 n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , 
 n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , 
 n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , 
 n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , 
 n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , 
 n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , 
 n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , 
 n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , 
 n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , 
 n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , 
 n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , 
 n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , 
 n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , 
 n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , 
 n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , 
 n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , 
 n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , 
 n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , 
 n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , 
 n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , 
 n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , 
 n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , 
 n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , 
 n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , 
 n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , 
 n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , 
 n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , 
 n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , 
 n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , 
 n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , 
 n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , 
 n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , 
 n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , 
 n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , 
 n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , 
 n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , 
 n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , 
 n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , 
 n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , 
 n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , 
 n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , 
 n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , 
 n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , 
 n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , 
 n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , 
 n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , 
 n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , 
 n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , 
 n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , 
 n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , 
 n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , 
 n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , 
 n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , 
 n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , 
 n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , 
 n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , 
 n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , 
 n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , 
 n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , 
 n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , 
 n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , 
 n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , 
 n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , 
 n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , 
 n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , 
 n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , 
 n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , 
 n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , 
 n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , 
 n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , 
 n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , 
 n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , 
 n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , 
 n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , 
 n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , 
 n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , 
 n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , 
 n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , 
 n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , 
 n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , 
 n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , 
 n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , 
 n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , 
 n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , 
 n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , 
 n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , 
 n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , 
 n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , 
 n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , 
 n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , 
 n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , 
 n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , 
 n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , 
 n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , 
 n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , 
 n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , 
 n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , 
 n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , 
 n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , 
 n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , 
 n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , 
 n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , 
 n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , 
 n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , 
 n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , 
 n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , 
 n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , 
 n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , 
 n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , 
 n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , 
 n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , 
 n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , 
 n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , 
 n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , 
 n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , 
 n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , 
 n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , 
 n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , 
 n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , 
 n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , 
 n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , 
 n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , 
 n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , 
 n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , 
 n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , 
 n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , 
 n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , 
 n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , 
 n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , 
 n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , 
 n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , 
 n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , 
 n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , 
 n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , 
 n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , 
 n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , 
 n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , 
 n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , 
 n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , 
 n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , 
 n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , 
 n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , 
 n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , 
 n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , 
 n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , 
 n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , 
 n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , 
 n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , 
 n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , 
 n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , 
 n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , 
 n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , 
 n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , 
 n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , 
 n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , 
 n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , 
 n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , 
 n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , 
 n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , 
 n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , 
 n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , 
 n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , 
 n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , 
 n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , 
 n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , 
 n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , 
 n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , 
 n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , 
 n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , 
 n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , 
 n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , 
 n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , 
 n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , 
 n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , 
 n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , 
 n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , 
 n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , 
 n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , 
 n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , 
 n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , 
 n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , 
 n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , 
 n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , 
 n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , 
 n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , 
 n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , 
 n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , 
 n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , 
 n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , 
 n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , 
 n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , 
 n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , 
 n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , 
 n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , 
 n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , 
 n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , 
 n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , 
 n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , 
 n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , 
 n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , 
 n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , 
 n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , 
 n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , 
 n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , 
 n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , 
 n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , 
 n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , 
 n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , 
 n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , 
 n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , 
 n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , 
 n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , 
 n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , 
 n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , 
 n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , 
 n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , 
 n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , 
 n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , 
 n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , 
 n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , 
 n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , 
 n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , 
 n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , 
 n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , 
 n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , 
 n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , 
 n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , 
 n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , 
 n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , 
 n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , 
 n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , 
 n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , 
 n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , 
 n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , 
 n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , 
 n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , 
 n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , 
 n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , 
 n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , 
 n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , 
 n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , 
 n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , 
 n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , 
 n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , 
 n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , 
 n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , 
 n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , 
 n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , 
 n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , 
 n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , 
 n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , 
 n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , 
 n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , 
 n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , 
 n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , 
 n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , 
 n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , 
 n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , 
 n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , 
 n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , 
 n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , 
 n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , 
 n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , 
 n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , 
 n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , 
 n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , 
 n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , 
 n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , 
 n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , 
 n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , 
 n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , 
 n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , 
 n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , 
 n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , 
 n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , 
 n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , 
 n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , 
 n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , 
 n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , 
 n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , 
 n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , 
 n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , 
 n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , 
 n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , 
 n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , 
 n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , 
 n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , 
 n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , 
 n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , 
 n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , 
 n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , 
 n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , 
 n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , 
 n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , 
 n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , 
 n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , 
 n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , 
 n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , 
 n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , 
 n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , 
 n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , 
 n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , 
 n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , 
 n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , 
 n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , 
 n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , 
 n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , 
 n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , 
 n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , 
 n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , 
 n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , 
 n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , 
 n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , 
 n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , 
 n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , 
 n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , 
 n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , 
 n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , 
 n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , 
 n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , 
 n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , 
 n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , 
 n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , 
 n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , 
 n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , 
 n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , 
 n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , 
 n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , 
 n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , 
 n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , 
 n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , 
 n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , 
 n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , 
 n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , 
 n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , 
 n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , 
 n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , 
 n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , 
 n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , 
 n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , 
 n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , 
 n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , 
 n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , 
 n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , 
 n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , 
 n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , 
 n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , 
 n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , 
 n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , 
 n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , 
 n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , 
 n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , 
 n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , 
 n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , 
 n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , 
 n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , 
 n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , 
 n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , 
 n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , 
 n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , 
 n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , 
 n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , 
 n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , 
 n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , 
 n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , 
 n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , 
 n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , 
 n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , 
 n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , 
 n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , 
 n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , 
 n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , 
 n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , 
 n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , 
 n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , 
 n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , 
 n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , 
 n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , 
 n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , 
 n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , 
 n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , 
 n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , 
 n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , 
 n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , 
 n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , 
 n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , 
 n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , 
 n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , 
 n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , 
 n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , 
 n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , 
 n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , 
 n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , 
 n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , 
 n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , 
 n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , 
 n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , 
 n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , 
 n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , 
 n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , 
 n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , 
 n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , 
 n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , 
 n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , 
 n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , 
 n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , 
 n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , 
 n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , 
 n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , 
 n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , 
 n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , 
 n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , 
 n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , 
 n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , 
 n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , 
 n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , 
 n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , 
 n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , 
 n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , 
 n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , 
 n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , 
 n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , 
 n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , 
 n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , 
 n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , 
 n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , 
 n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , 
 n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , 
 n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , 
 n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , 
 n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , 
 n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , 
 n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , 
 n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , 
 n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , 
 n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , 
 n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , 
 n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , 
 n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , 
 n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , 
 n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , 
 n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , 
 n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , 
 n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , 
 n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , 
 n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , 
 n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , 
 n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , 
 n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , 
 n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , 
 n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , 
 n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , 
 n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , 
 n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , 
 n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , 
 n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , 
 n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , 
 n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , 
 n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , 
 n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , 
 n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , 
 n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , 
 n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , 
 n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , 
 n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , 
 n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , 
 n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , 
 n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , 
 n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , 
 n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , 
 n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , 
 n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , 
 n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , 
 n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , 
 n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , 
 n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , 
 n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , 
 n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , 
 n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , 
 n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , 
 n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , 
 n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , 
 n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , 
 n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , 
 n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , 
 n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , 
 n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , 
 n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , 
 n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , 
 n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , 
 n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , 
 n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , 
 n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , 
 n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , 
 n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , 
 n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , 
 n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , 
 n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , 
 n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , 
 n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , 
 n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , 
 n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , 
 n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , 
 n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , 
 n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , 
 n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , 
 n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , 
 n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , 
 n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , 
 n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , 
 n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , 
 n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , 
 n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , 
 n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , 
 n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , 
 n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , 
 n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , 
 n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , 
 n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , 
 n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , 
 n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , 
 n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , 
 n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , 
 n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , 
 n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , 
 n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , 
 n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , 
 n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , 
 n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , 
 n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , 
 n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , 
 n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , 
 n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , 
 n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , 
 n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , 
 n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , 
 n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , 
 n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , 
 n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , 
 n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , 
 n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , 
 n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , 
 n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , 
 n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , 
 n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , 
 n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , 
 n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , 
 n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , 
 n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , 
 n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , 
 n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , 
 n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , 
 n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , 
 n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , 
 n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , 
 n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , 
 n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , 
 n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , 
 n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , 
 n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , 
 n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , 
 n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , 
 n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , 
 n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , 
 n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , 
 n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , 
 n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , 
 n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , 
 n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , 
 n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , 
 n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , 
 n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , 
 n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , 
 n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , 
 n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , 
 n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , 
 n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , 
 n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , 
 n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , 
 n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , 
 n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , 
 n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , 
 n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , 
 n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , 
 n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , 
 n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , 
 n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , 
 n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , 
 n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , 
 n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , 
 n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , 
 n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , 
 n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , 
 n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , 
 n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , 
 n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , 
 n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , 
 n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , 
 n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , 
 n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , 
 n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , 
 n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , 
 n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , 
 n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , 
 n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , 
 n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , 
 n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , 
 n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , 
 n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , 
 n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , 
 n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , 
 n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , 
 n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , 
 n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , 
 n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , 
 n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , 
 n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , 
 n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , 
 n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , 
 n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , 
 n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , 
 n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , 
 n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , 
 n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , 
 n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , 
 n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , 
 n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , 
 n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , 
 n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , 
 n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , 
 n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , 
 n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , 
 n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , 
 n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , 
 n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , 
 n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , 
 n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , 
 n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , 
 n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , 
 n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , 
 n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , 
 n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , 
 n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , 
 n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , 
 n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , 
 n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , 
 n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , 
 n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , 
 n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , 
 n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , 
 n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , 
 n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , 
 n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , 
 n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , 
 n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , 
 n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , 
 n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , 
 n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , 
 n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , 
 n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , 
 n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , 
 n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , 
 n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , 
 n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , 
 n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , 
 n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , 
 n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , 
 n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , 
 n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , 
 n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , 
 n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , 
 n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , 
 n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , 
 n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , 
 n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , 
 n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , 
 n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , 
 n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , 
 n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , 
 n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , 
 n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , 
 n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , 
 n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , 
 n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , 
 n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , 
 n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , 
 n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , 
 n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , 
 n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , 
 n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , 
 n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , 
 n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , 
 n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , 
 n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , 
 n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , 
 n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , 
 n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , 
 n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , 
 n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , 
 n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , 
 n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , 
 n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , 
 n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , 
 n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , 
 n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , 
 n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , 
 n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , 
 n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , 
 n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , 
 n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , 
 n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , 
 n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , 
 n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , 
 n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , 
 n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , 
 n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , 
 n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , 
 n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , 
 n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , 
 n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , 
 n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , 
 n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , 
 n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , 
 n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , 
 n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , 
 n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , 
 n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , 
 n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , 
 n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , 
 n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , 
 n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , 
 n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , 
 n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , 
 n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , 
 n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , 
 n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , 
 n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , 
 n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , 
 n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , 
 n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , 
 n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , 
 n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , 
 n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , 
 n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , 
 n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , 
 n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , 
 n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , 
 n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , 
 n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , 
 n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , 
 n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , 
 n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , 
 n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , 
 n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , 
 n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , 
 n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , 
 n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , 
 n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , 
 n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , 
 n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , 
 n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , 
 n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , 
 n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , 
 n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , 
 n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , 
 n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , 
 n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , 
 n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , 
 n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , 
 n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , 
 n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , 
 n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , 
 n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , 
 n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , 
 n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , 
 n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , 
 n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , 
 n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , 
 n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , 
 n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , 
 n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , 
 n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , 
 n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , 
 n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , 
 n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , 
 n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , 
 n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , 
 n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , 
 n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , 
 n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , 
 n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , 
 n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , 
 n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , 
 n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , 
 n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , 
 n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , 
 n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , 
 n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , 
 n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , 
 n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , 
 n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , 
 n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , 
 n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , 
 n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , 
 n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , 
 n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , 
 n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , 
 n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , 
 n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , 
 n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , 
 n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , 
 n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , 
 n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , 
 n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , 
 n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , 
 n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , 
 n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , 
 n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , 
 n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , 
 n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , 
 n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , 
 n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , 
 n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , 
 n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , 
 n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , 
 n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , 
 n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , 
 n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , 
 n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , 
 n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , 
 n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , 
 n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , 
 n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , 
 n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , 
 n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , 
 n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , 
 n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , 
 n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , 
 n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , 
 n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , 
 n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , 
 n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , 
 n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , 
 n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , 
 n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , 
 n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , 
 n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , 
 n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , 
 n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , 
 n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , 
 n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , 
 n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , 
 n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , 
 n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , 
 n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , 
 n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , 
 n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , 
 n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , 
 n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , 
 n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , 
 n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , 
 n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , 
 n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , 
 n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , 
 n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , 
 n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , 
 n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , 
 n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , 
 n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , 
 n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , 
 n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , 
 n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , 
 n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , 
 n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , 
 n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , 
 n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , 
 n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , 
 n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , 
 n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , 
 n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , 
 n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , 
 n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , 
 n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , 
 n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , 
 n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , 
 n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , 
 n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , 
 n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , 
 n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , 
 n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , 
 n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , 
 n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , 
 n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , 
 n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , 
 n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , 
 n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , 
 n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , 
 n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , 
 n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , 
 n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , 
 n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , 
 n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , 
 n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , 
 n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , 
 n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , 
 n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , 
 n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , 
 n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , 
 n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , 
 n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , 
 n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , 
 n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , 
 n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , 
 n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , 
 n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , 
 n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , 
 n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , 
 n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , 
 n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , 
 n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , 
 n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , 
 n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , 
 n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , 
 n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , 
 n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , 
 n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , 
 n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , 
 n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , 
 n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , 
 n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , 
 n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , 
 n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , 
 n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , 
 n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , 
 n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , 
 n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , 
 n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , 
 n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , 
 n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , 
 n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , 
 n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , 
 n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , 
 n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , 
 n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , 
 n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , 
 n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , 
 n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , 
 n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , 
 n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , 
 n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , 
 n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , 
 n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , 
 n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , 
 n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , 
 n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , 
 n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , 
 n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , 
 n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , 
 n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , 
 n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , 
 n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , 
 n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , 
 n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , 
 n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , 
 n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , 
 n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , 
 n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , 
 n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , 
 n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , 
 n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , 
 n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , 
 n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , 
 n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , 
 n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , 
 n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , 
 n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , 
 n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , 
 n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , 
 n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , 
 n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , 
 n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , 
 n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , 
 n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , 
 n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , 
 n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , 
 n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , 
 n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , 
 n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , 
 n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , 
 n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , 
 n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , 
 n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , 
 n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , 
 n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , 
 n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , 
 n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , 
 n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , 
 n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , 
 n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , 
 n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , 
 n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , 
 n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , 
 n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , 
 n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , 
 n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , 
 n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , 
 n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , 
 n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , 
 n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , 
 n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , 
 n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , 
 n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , 
 n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , 
 n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , 
 n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , 
 n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , 
 n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , 
 n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , 
 n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , 
 n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , 
 n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , 
 n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , 
 n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , 
 n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , 
 n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , 
 n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , 
 n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , 
 n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , 
 n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , 
 n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , 
 n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , 
 n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , 
 n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , 
 n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , 
 n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , 
 n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , 
 n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , 
 n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , 
 n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , 
 n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , 
 n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , 
 n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , 
 n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , 
 n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , 
 n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , 
 n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , 
 n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , 
 n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , 
 n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , 
 n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , 
 n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , 
 n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , 
 n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , 
 n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , 
 n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , 
 n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , 
 n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , 
 n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , 
 n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , 
 n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , 
 n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , 
 n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , 
 n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , 
 n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , 
 n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , 
 n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , 
 n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , 
 n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , 
 n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , 
 n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , 
 n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , 
 n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , 
 n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , 
 n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , 
 n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , 
 n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , 
 n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , 
 n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , 
 n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , 
 n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , 
 n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , 
 n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , 
 n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , 
 n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , 
 n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , 
 n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , 
 n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , 
 n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , 
 n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , 
 n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , 
 n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , 
 n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , 
 n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , 
 n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , 
 n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , 
 n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , 
 n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , 
 n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , 
 n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , 
 n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , 
 n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , 
 n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , 
 n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , 
 n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , 
 n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , 
 n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , 
 n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , 
 n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , 
 n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , 
 n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , 
 n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , 
 n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , 
 n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , 
 n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , 
 n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , 
 n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , 
 n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , 
 n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , 
 n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , 
 n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , 
 n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , 
 n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , 
 n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , 
 n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , 
 n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , 
 n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , 
 n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , 
 n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , 
 n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , 
 n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , 
 n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , 
 n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , 
 n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , 
 n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , 
 n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , 
 n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , 
 n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , 
 n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , 
 n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , 
 n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , 
 n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , 
 n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , 
 n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , 
 n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , 
 n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , 
 n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , 
 n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , 
 n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , 
 n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , 
 n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , 
 n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , 
 n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , 
 n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , 
 n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , 
 n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , 
 n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , 
 n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , 
 n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , 
 n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , 
 n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , 
 n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , 
 n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , 
 n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , 
 n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , 
 n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , 
 n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , 
 n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , 
 n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , 
 n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , 
 n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , 
 n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , 
 n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , 
 n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , 
 n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , 
 n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , 
 n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , 
 n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , 
 n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , 
 n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , 
 n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , 
 n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , 
 n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , 
 n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , 
 n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , 
 n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , 
 n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , 
 n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , 
 n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , 
 n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , 
 n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , 
 n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , 
 n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , 
 n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , 
 n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , 
 n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , 
 n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , 
 n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , 
 n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , 
 n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , 
 n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , 
 n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , 
 n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , 
 n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , 
 n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , 
 n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , 
 n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , 
 n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , 
 n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , 
 n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , 
 n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , 
 n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , 
 n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , 
 n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , 
 n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , 
 n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , 
 n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , 
 n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , 
 n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , 
 n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , 
 n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , 
 n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , 
 n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , 
 n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , 
 n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , 
 n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , 
 n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , 
 n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , 
 n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , 
 n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , 
 n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , 
 n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , 
 n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , 
 n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , 
 n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , 
 n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , 
 n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , 
 n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , 
 n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , 
 n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , 
 n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , 
 n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , 
 n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , 
 n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , 
 n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , 
 n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , 
 n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , 
 n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , 
 n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , 
 n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , 
 n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , 
 n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , 
 n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , 
 n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , 
 n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , 
 n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , 
 n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , 
 n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , 
 n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , 
 n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , 
 n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , 
 n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , 
 n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , 
 n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , 
 n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , 
 n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , 
 n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , 
 n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , 
 n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , 
 n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , 
 n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , 
 n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , 
 n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , 
 n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , 
 n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , 
 n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , 
 n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , 
 n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , 
 n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , 
 n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , 
 n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , 
 n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , 
 n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , 
 n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , 
 n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , 
 n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , 
 n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , 
 n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , 
 n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , 
 n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , 
 n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , 
 n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , 
 n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , 
 n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , 
 n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , 
 n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , 
 n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , 
 n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , 
 n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , 
 n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , 
 n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , 
 n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , 
 n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , 
 n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , 
 n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , 
 n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , 
 n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , 
 n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , 
 n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , 
 n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , 
 n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , 
 n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , 
 n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , 
 n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , 
 n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , 
 n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , 
 n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , 
 n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , 
 n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , 
 n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , 
 n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , 
 n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , 
 n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , 
 n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , 
 n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , 
 n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , 
 n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , 
 n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , 
 n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , 
 n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , 
 n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , 
 n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , 
 n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , 
 n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , 
 n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , 
 n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , 
 n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , 
 n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , 
 n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , 
 n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , 
 n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , 
 n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , 
 n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , 
 n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , 
 n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , 
 n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , 
 n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , 
 n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , 
 n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , 
 n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , 
 n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , 
 n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , 
 n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , 
 n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , 
 n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , 
 n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , 
 n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , 
 n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , 
 n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , 
 n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , 
 n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , 
 n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , 
 n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , 
 n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , 
 n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , 
 n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , 
 n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , 
 n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , 
 n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , 
 n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , 
 n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , 
 n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , 
 n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , 
 n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , 
 n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , 
 n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , 
 n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , 
 n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , 
 n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , 
 n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , 
 n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , 
 n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , 
 n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , 
 n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , 
 n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , 
 n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , 
 n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , 
 n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , 
 n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , 
 n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , 
 n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , 
 n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , 
 n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , 
 n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , 
 n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , 
 n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , 
 n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , 
 n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , 
 n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , 
 n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , 
 n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , 
 n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , 
 n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , 
 n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , 
 n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , 
 n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , 
 n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , 
 n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , 
 n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , 
 n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , 
 n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , 
 n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , 
 n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , 
 n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , 
 n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , 
 n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , 
 n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , 
 n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , 
 n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , 
 n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , 
 n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , 
 n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , 
 n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , 
 n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , 
 n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , 
 n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , 
 n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , 
 n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , 
 n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , 
 n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , 
 n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , 
 n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , 
 n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , 
 n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , 
 n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , 
 n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , 
 n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , 
 n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , 
 n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , 
 n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , 
 n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , 
 n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , 
 n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , 
 n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , 
 n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , 
 n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , 
 n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , 
 n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , 
 n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , 
 n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , 
 n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , 
 n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , 
 n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , 
 n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , 
 n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , 
 n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , 
 n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , 
 n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , 
 n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , 
 n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , 
 n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , 
 n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , 
 n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , 
 n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , 
 n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , 
 n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , 
 n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , 
 n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , 
 n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , 
 n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , 
 n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , 
 n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , 
 n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , 
 n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , 
 n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , 
 n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , 
 n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , 
 n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , 
 n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , 
 n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , 
 n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , 
 n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , 
 n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , 
 n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , 
 n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , 
 n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , 
 n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , 
 n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , 
 n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , 
 n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , 
 n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , 
 n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , 
 n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , 
 n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , 
 n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , 
 n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , 
 n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , 
 n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , 
 n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , 
 n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , 
 n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , 
 n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , 
 n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , 
 n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , 
 n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , 
 n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , 
 n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , 
 n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , 
 n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , 
 n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , 
 n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , 
 n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , 
 n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , 
 n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , 
 n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , 
 n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , 
 n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , 
 n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , 
 n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , 
 n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , 
 n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , 
 n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , 
 n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , 
 n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , 
 n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , 
 n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , 
 n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , 
 n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , 
 n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , 
 n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , 
 n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , 
 n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , 
 n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , 
 n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , 
 n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , 
 n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , 
 n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , 
 n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , 
 n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , 
 n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , 
 n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , 
 n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , 
 n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , 
 n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , 
 n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , 
 n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , 
 n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , 
 n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , 
 n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , 
 n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , 
 n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , 
 n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , 
 n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , 
 n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , 
 n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , 
 n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , 
 n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , 
 n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , 
 n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , 
 n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , 
 n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , 
 n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , 
 n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , 
 n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , 
 n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , 
 n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , 
 n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , 
 n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , 
 n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , 
 n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , 
 n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , 
 n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , 
 n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , 
 n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , 
 n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , 
 n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , 
 n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , 
 n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , 
 n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , 
 n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , 
 n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , 
 n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , 
 n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , 
 n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , 
 n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , 
 n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , 
 n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , 
 n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , 
 n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , 
 n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , 
 n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , 
 n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , 
 n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , 
 n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , 
 n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , 
 n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , 
 n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , 
 n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , 
 n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , 
 n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , 
 n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , 
 n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , 
 n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , 
 n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , 
 n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , 
 n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , 
 n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , 
 n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , 
 n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , 
 n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , 
 n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , 
 n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , 
 n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , 
 n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , 
 n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , 
 n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , 
 n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , 
 n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , 
 n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , 
 n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , 
 n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , 
 n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , 
 n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , 
 n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , 
 n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , 
 n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , 
 n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , 
 n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , 
 n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , 
 n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , 
 n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , 
 n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , 
 n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , 
 n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , 
 n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , 
 n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , 
 n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , 
 n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , 
 n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , 
 n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , 
 n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , 
 n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , 
 n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , 
 n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , 
 n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , 
 n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , 
 n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , 
 n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , 
 n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , 
 n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , 
 n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , 
 n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , 
 n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , 
 n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , 
 n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , 
 n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , 
 n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , 
 n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , 
 n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , 
 n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , 
 n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , 
 n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , 
 n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , 
 n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , 
 n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , 
 n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , 
 n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , 
 n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , 
 n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , 
 n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , 
 n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , 
 n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , 
 n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , 
 n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , 
 n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , 
 n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , 
 n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , 
 n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , 
 n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , 
 n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , 
 n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , 
 n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , 
 n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , 
 n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , 
 n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , 
 n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , 
 n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , 
 n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , 
 n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , 
 n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , 
 n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , 
 n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , 
 n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , 
 n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , 
 n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , 
 n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , 
 n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , 
 n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , 
 n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , 
 n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , 
 n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , 
 n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , 
 n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , 
 n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , 
 n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , 
 n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , 
 n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , 
 n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , 
 n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , 
 n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , 
 n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , 
 n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , 
 n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , 
 n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , 
 n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , 
 n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , 
 n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , 
 n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , 
 n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , 
 n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , 
 n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , 
 n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , 
 n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , 
 n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , 
 n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , 
 n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , 
 n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , 
 n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , 
 n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , 
 n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , 
 n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , 
 n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , 
 n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , 
 n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , 
 n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , 
 n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , 
 n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , 
 n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , 
 n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , 
 n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , 
 n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , 
 n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , 
 n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , 
 n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , 
 n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , 
 n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , 
 n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , 
 n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , 
 n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , 
 n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , 
 n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , 
 n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , 
 n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , 
 n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , 
 n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , 
 n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , 
 n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , 
 n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , 
 n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , 
 n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , 
 n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , 
 n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , 
 n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , 
 n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , 
 n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , 
 n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , 
 n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , 
 n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , 
 n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , 
 n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , 
 n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , 
 n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , 
 n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , 
 n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , 
 n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , 
 n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , 
 n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , 
 n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , 
 n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , 
 n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , 
 n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , 
 n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , 
 n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , 
 n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , 
 n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , 
 n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , 
 n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , 
 n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , 
 n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , 
 n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , 
 n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , 
 n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , 
 n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , 
 n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , 
 n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , 
 n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , 
 n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , 
 n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , 
 n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , 
 n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , 
 n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , 
 n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , 
 n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , 
 n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , 
 n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , 
 n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , 
 n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , 
 n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , 
 n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , 
 n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , 
 n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , 
 n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , 
 n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , 
 n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , 
 n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , 
 n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , 
 n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , 
 n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , 
 n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , 
 n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , 
 n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , 
 n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , 
 n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , 
 n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , 
 n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , 
 n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , 
 n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , 
 n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , 
 n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , 
 n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , 
 n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , 
 n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , 
 n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , 
 n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , 
 n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , 
 n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , 
 n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , 
 n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , 
 n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , 
 n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , 
 n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , 
 n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , 
 n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , 
 n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , 
 n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , 
 n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , 
 n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , 
 n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , 
 n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , 
 n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , 
 n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , 
 n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , 
 n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , 
 n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , 
 n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , 
 n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , 
 n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , 
 n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , 
 n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , 
 n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , 
 n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , 
 n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , 
 n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , 
 n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , 
 n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , 
 n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , 
 n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , 
 n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , 
 n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , 
 n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , 
 n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , 
 n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , 
 n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , 
 n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , 
 n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , 
 n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , 
 n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , 
 n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , 
 n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , 
 n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , 
 n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , 
 n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , 
 n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , 
 n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , 
 n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , 
 n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , 
 n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , 
 n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , 
 n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , 
 n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , 
 n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , 
 n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , 
 n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , 
 n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , 
 n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , 
 n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , 
 n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , 
 n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , 
 n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , 
 n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , 
 n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , 
 n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , 
 n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , 
 n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , 
 n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , 
 n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , 
 n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , 
 n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , 
 n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , 
 n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , 
 n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , 
 n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , 
 n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , 
 n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , 
 n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , 
 n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , 
 n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , 
 n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , 
 n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , 
 n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , 
 n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , 
 n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , 
 n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , 
 n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , 
 n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , 
 n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , 
 n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , 
 n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , 
 n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , 
 n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , 
 n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , 
 n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , 
 n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , 
 n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , 
 n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , 
 n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , 
 n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , 
 n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , 
 n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , 
 n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , 
 n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , 
 n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , 
 n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , 
 n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , 
 n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , 
 n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , 
 n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , 
 n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , 
 n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , 
 n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , 
 n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , 
 n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , 
 n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , 
 n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , 
 n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , 
 n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , 
 n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , 
 n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , 
 n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , 
 n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , 
 n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , 
 n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , 
 n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , 
 n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , 
 n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , 
 n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , 
 n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , 
 n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , 
 n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , 
 n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , 
 n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , 
 n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , 
 n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , 
 n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , 
 n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , 
 n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , 
 n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , 
 n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , 
 n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , 
 n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , 
 n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , 
 n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , 
 n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , 
 n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , 
 n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , 
 n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , 
 n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , 
 n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , 
 n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , 
 n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , 
 n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , 
 n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , 
 n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , 
 n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , 
 n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , 
 n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , 
 n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , 
 n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , 
 n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , 
 n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , 
 n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , 
 n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , 
 n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , 
 n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , 
 n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , 
 n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , 
 n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , 
 n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , 
 n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , 
 n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , 
 n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , 
 n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , 
 n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , 
 n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , 
 n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , 
 n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , 
 n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , 
 n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , 
 n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , 
 n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , 
 n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , 
 n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , 
 n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , 
 n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , 
 n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , 
 n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , 
 n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , 
 n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , 
 n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , 
 n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , 
 n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , 
 n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , 
 n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , 
 n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , 
 n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , 
 n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , 
 n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , 
 n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , 
 n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , 
 n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , 
 n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , 
 n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , 
 n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , 
 n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , 
 n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , 
 n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , 
 n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , 
 n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , 
 n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , 
 n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , 
 n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , 
 n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , 
 n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , 
 n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , 
 n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , 
 n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , 
 n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , 
 n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , 
 n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , 
 n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , 
 n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , 
 n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , 
 n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , 
 n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , 
 n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , 
 n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , 
 n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , 
 n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , 
 n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , 
 n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , 
 n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , 
 n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , 
 n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , 
 n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , 
 n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , 
 n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , 
 n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , 
 n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , 
 n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , 
 n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , 
 n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , 
 n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , 
 n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , 
 n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , 
 n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , 
 n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , 
 n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , 
 n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , 
 n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , 
 n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , 
 n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , 
 n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , 
 n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , 
 n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , 
 n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , 
 n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , 
 n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , 
 n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , 
 n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , 
 n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , 
 n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , 
 n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , 
 n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , 
 n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , 
 n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , 
 n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , 
 n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , 
 n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , 
 n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , 
 n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , 
 n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , 
 n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , 
 n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , 
 n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , 
 n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , 
 n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , 
 n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , 
 n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , 
 n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , 
 n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , 
 n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , 
 n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , 
 n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , 
 n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , 
 n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , 
 n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , 
 n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , 
 n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , 
 n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , 
 n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , 
 n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , 
 n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , 
 n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , 
 n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , 
 n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , 
 n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , 
 n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , 
 n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , 
 n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , 
 n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , 
 n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , 
 n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , 
 n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , 
 n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , 
 n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , 
 n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , 
 n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , 
 n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , 
 n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , 
 n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , 
 n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , 
 n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , 
 n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , 
 n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , 
 n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , 
 n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , 
 n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , 
 n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , 
 n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , 
 n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , 
 n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , 
 n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , 
 n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , 
 n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , 
 n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , 
 n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , 
 n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , 
 n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , 
 n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , 
 n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , 
 n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , 
 n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , 
 n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , 
 n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , 
 n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , 
 n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , 
 n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , 
 n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , 
 n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , 
 n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , 
 n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , 
 n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , 
 n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , 
 n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , 
 n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , 
 n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , 
 n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , 
 n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , 
 n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , 
 n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , 
 n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , 
 n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , 
 n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , 
 n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , 
 n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , 
 n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , 
 n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , 
 n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , 
 n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , 
 n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , 
 n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , 
 n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , 
 n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , 
 n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , 
 n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , 
 n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , 
 n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , 
 n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , 
 n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , 
 n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , 
 n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , 
 n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , 
 n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , 
 n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , 
 n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , 
 n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , 
 n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , 
 n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , 
 n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , 
 n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , 
 n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , 
 n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , 
 n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , 
 n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , 
 n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , 
 n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , 
 n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , 
 n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , 
 n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , 
 n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , 
 n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , 
 n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , 
 n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , 
 n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , 
 n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , 
 n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , 
 n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , 
 n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , 
 n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , 
 n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , 
 n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , 
 n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , 
 n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , 
 n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , 
 n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , 
 n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , 
 n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , 
 n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , 
 n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , 
 n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , 
 n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , 
 n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , 
 n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , 
 n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , 
 n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , 
 n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , 
 n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , 
 n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , 
 n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , 
 n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , 
 n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , 
 n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , 
 n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , 
 n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , 
 n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , 
 n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , 
 n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , 
 n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , 
 n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , 
 n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , 
 n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , 
 n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , 
 n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , 
 n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , 
 n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , 
 n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , 
 n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , 
 n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , 
 n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , 
 n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , 
 n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , 
 n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , 
 n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , 
 n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , 
 n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , 
 n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , 
 n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , 
 n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , 
 n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , 
 n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , 
 n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , 
 n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , 
 n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , 
 n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , 
 n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , 
 n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , 
 n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , 
 n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , 
 n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , 
 n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , 
 n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , 
 n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , 
 n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , 
 n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , 
 n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , 
 n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , 
 n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , 
 n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , 
 n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , 
 n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , 
 n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , 
 n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , 
 n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , 
 n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , 
 n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , 
 n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , 
 n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , 
 n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , 
 n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , 
 n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , 
 n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , 
 n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , 
 n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , 
 n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , 
 n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , 
 n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , 
 n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , 
 n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , 
 n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , 
 n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , 
 n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , 
 n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , 
 n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , 
 n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , 
 n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , 
 n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , 
 n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , 
 n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , 
 n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , 
 n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , 
 n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , 
 n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , 
 n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , 
 n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , 
 n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , 
 n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , 
 n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , 
 n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , 
 n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , 
 n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , 
 n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , 
 n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , 
 n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , 
 n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , 
 n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , 
 n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , 
 n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , 
 n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , 
 n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , 
 n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , 
 n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , 
 n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , 
 n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , 
 n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , 
 n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , 
 n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , 
 n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , 
 n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , 
 n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , 
 n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , 
 n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , 
 n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 ;
buf ( n768 , n0 );
buf ( n769 , n1 );
buf ( n770 , n2 );
buf ( n771 , n3 );
buf ( n772 , n4 );
buf ( n773 , n5 );
buf ( n774 , n6 );
buf ( n775 , n7 );
buf ( n776 , n8 );
buf ( n777 , n9 );
buf ( n778 , n10 );
buf ( n779 , n11 );
buf ( n780 , n12 );
buf ( n781 , n13 );
buf ( n782 , n14 );
buf ( n783 , n15 );
buf ( n784 , n16 );
buf ( n785 , n17 );
buf ( n786 , n18 );
buf ( n787 , n19 );
buf ( n788 , n20 );
buf ( n789 , n21 );
buf ( n790 , n22 );
buf ( n791 , n23 );
buf ( n792 , n24 );
buf ( n793 , n25 );
buf ( n794 , n26 );
buf ( n795 , n27 );
buf ( n796 , n28 );
buf ( n797 , n29 );
buf ( n798 , n30 );
buf ( n799 , n31 );
buf ( n800 , n32 );
buf ( n801 , n33 );
buf ( n802 , n34 );
buf ( n803 , n35 );
buf ( n804 , n36 );
buf ( n805 , n37 );
buf ( n806 , n38 );
buf ( n807 , n39 );
buf ( n808 , n40 );
buf ( n809 , n41 );
buf ( n810 , n42 );
buf ( n811 , n43 );
buf ( n812 , n44 );
buf ( n813 , n45 );
buf ( n814 , n46 );
buf ( n815 , n47 );
buf ( n816 , n48 );
buf ( n817 , n49 );
buf ( n818 , n50 );
buf ( n819 , n51 );
buf ( n820 , n52 );
buf ( n821 , n53 );
buf ( n822 , n54 );
buf ( n823 , n55 );
buf ( n824 , n56 );
buf ( n825 , n57 );
buf ( n826 , n58 );
buf ( n827 , n59 );
buf ( n828 , n60 );
buf ( n829 , n61 );
buf ( n830 , n62 );
buf ( n831 , n63 );
buf ( n832 , n64 );
buf ( n833 , n65 );
buf ( n834 , n66 );
buf ( n835 , n67 );
buf ( n836 , n68 );
buf ( n837 , n69 );
buf ( n838 , n70 );
buf ( n839 , n71 );
buf ( n840 , n72 );
buf ( n841 , n73 );
buf ( n842 , n74 );
buf ( n843 , n75 );
buf ( n844 , n76 );
buf ( n845 , n77 );
buf ( n846 , n78 );
buf ( n847 , n79 );
buf ( n848 , n80 );
buf ( n849 , n81 );
buf ( n850 , n82 );
buf ( n851 , n83 );
buf ( n852 , n84 );
buf ( n853 , n85 );
buf ( n854 , n86 );
buf ( n855 , n87 );
buf ( n856 , n88 );
buf ( n857 , n89 );
buf ( n858 , n90 );
buf ( n859 , n91 );
buf ( n860 , n92 );
buf ( n861 , n93 );
buf ( n862 , n94 );
buf ( n863 , n95 );
buf ( n864 , n96 );
buf ( n865 , n97 );
buf ( n866 , n98 );
buf ( n867 , n99 );
buf ( n868 , n100 );
buf ( n869 , n101 );
buf ( n870 , n102 );
buf ( n871 , n103 );
buf ( n872 , n104 );
buf ( n873 , n105 );
buf ( n874 , n106 );
buf ( n875 , n107 );
buf ( n876 , n108 );
buf ( n877 , n109 );
buf ( n878 , n110 );
buf ( n879 , n111 );
buf ( n880 , n112 );
buf ( n881 , n113 );
buf ( n882 , n114 );
buf ( n883 , n115 );
buf ( n884 , n116 );
buf ( n885 , n117 );
buf ( n886 , n118 );
buf ( n887 , n119 );
buf ( n888 , n120 );
buf ( n889 , n121 );
buf ( n890 , n122 );
buf ( n891 , n123 );
buf ( n892 , n124 );
buf ( n893 , n125 );
buf ( n894 , n126 );
buf ( n895 , n127 );
buf ( n128 , n896 );
buf ( n129 , n897 );
buf ( n130 , n898 );
buf ( n131 , n899 );
buf ( n132 , n900 );
buf ( n133 , n901 );
buf ( n134 , n902 );
buf ( n135 , n903 );
buf ( n136 , n904 );
buf ( n137 , n905 );
buf ( n138 , n906 );
buf ( n139 , n907 );
buf ( n140 , n908 );
buf ( n141 , n909 );
buf ( n142 , n910 );
buf ( n143 , n911 );
buf ( n144 , n912 );
buf ( n145 , n913 );
buf ( n146 , n914 );
buf ( n147 , n915 );
buf ( n148 , n916 );
buf ( n149 , n917 );
buf ( n150 , n918 );
buf ( n151 , n919 );
buf ( n152 , n920 );
buf ( n153 , n921 );
buf ( n154 , n922 );
buf ( n155 , n923 );
buf ( n156 , n924 );
buf ( n157 , n925 );
buf ( n158 , n926 );
buf ( n159 , n927 );
buf ( n160 , n928 );
buf ( n161 , n929 );
buf ( n162 , n930 );
buf ( n163 , n931 );
buf ( n164 , n932 );
buf ( n165 , n933 );
buf ( n166 , n934 );
buf ( n167 , n935 );
buf ( n168 , n936 );
buf ( n169 , n937 );
buf ( n170 , n938 );
buf ( n171 , n939 );
buf ( n172 , n940 );
buf ( n173 , n941 );
buf ( n174 , n942 );
buf ( n175 , n943 );
buf ( n176 , n944 );
buf ( n177 , n945 );
buf ( n178 , n946 );
buf ( n179 , n947 );
buf ( n180 , n948 );
buf ( n181 , n949 );
buf ( n182 , n950 );
buf ( n183 , n951 );
buf ( n184 , n952 );
buf ( n185 , n953 );
buf ( n186 , n954 );
buf ( n187 , n955 );
buf ( n188 , n956 );
buf ( n189 , n957 );
buf ( n190 , n958 );
buf ( n191 , n959 );
buf ( n192 , n960 );
buf ( n193 , n961 );
buf ( n194 , n962 );
buf ( n195 , n963 );
buf ( n196 , n964 );
buf ( n197 , n965 );
buf ( n198 , n966 );
buf ( n199 , n967 );
buf ( n200 , n968 );
buf ( n201 , n969 );
buf ( n202 , n970 );
buf ( n203 , n971 );
buf ( n204 , n972 );
buf ( n205 , n973 );
buf ( n206 , n974 );
buf ( n207 , n975 );
buf ( n208 , n976 );
buf ( n209 , n977 );
buf ( n210 , n978 );
buf ( n211 , n979 );
buf ( n212 , n980 );
buf ( n213 , n981 );
buf ( n214 , n982 );
buf ( n215 , n983 );
buf ( n216 , n984 );
buf ( n217 , n985 );
buf ( n218 , n986 );
buf ( n219 , n987 );
buf ( n220 , n988 );
buf ( n221 , n989 );
buf ( n222 , n990 );
buf ( n223 , n991 );
buf ( n224 , n992 );
buf ( n225 , n993 );
buf ( n226 , n994 );
buf ( n227 , n995 );
buf ( n228 , n996 );
buf ( n229 , n997 );
buf ( n230 , n998 );
buf ( n231 , n999 );
buf ( n232 , n1000 );
buf ( n233 , n1001 );
buf ( n234 , n1002 );
buf ( n235 , n1003 );
buf ( n236 , n1004 );
buf ( n237 , n1005 );
buf ( n238 , n1006 );
buf ( n239 , n1007 );
buf ( n240 , n1008 );
buf ( n241 , n1009 );
buf ( n242 , n1010 );
buf ( n243 , n1011 );
buf ( n244 , n1012 );
buf ( n245 , n1013 );
buf ( n246 , n1014 );
buf ( n247 , n1015 );
buf ( n248 , n1016 );
buf ( n249 , n1017 );
buf ( n250 , n1018 );
buf ( n251 , n1019 );
buf ( n252 , n1020 );
buf ( n253 , n1021 );
buf ( n254 , n1022 );
buf ( n255 , n1023 );
buf ( n256 , n1024 );
buf ( n257 , n1025 );
buf ( n258 , n1026 );
buf ( n259 , n1027 );
buf ( n260 , n1028 );
buf ( n261 , n1029 );
buf ( n262 , n1030 );
buf ( n263 , n1031 );
buf ( n264 , n1032 );
buf ( n265 , n1033 );
buf ( n266 , n1034 );
buf ( n267 , n1035 );
buf ( n268 , n1036 );
buf ( n269 , n1037 );
buf ( n270 , n1038 );
buf ( n271 , n1039 );
buf ( n272 , n1040 );
buf ( n273 , n1041 );
buf ( n274 , n1042 );
buf ( n275 , n1043 );
buf ( n276 , n1044 );
buf ( n277 , n1045 );
buf ( n278 , n1046 );
buf ( n279 , n1047 );
buf ( n280 , n1048 );
buf ( n281 , n1049 );
buf ( n282 , n1050 );
buf ( n283 , n1051 );
buf ( n284 , n1052 );
buf ( n285 , n1053 );
buf ( n286 , n1054 );
buf ( n287 , n1055 );
buf ( n288 , n1056 );
buf ( n289 , n1057 );
buf ( n290 , n1058 );
buf ( n291 , n1059 );
buf ( n292 , n1060 );
buf ( n293 , n1061 );
buf ( n294 , n1062 );
buf ( n295 , n1063 );
buf ( n296 , n1064 );
buf ( n297 , n1065 );
buf ( n298 , n1066 );
buf ( n299 , n1067 );
buf ( n300 , n1068 );
buf ( n301 , n1069 );
buf ( n302 , n1070 );
buf ( n303 , n1071 );
buf ( n304 , n1072 );
buf ( n305 , n1073 );
buf ( n306 , n1074 );
buf ( n307 , n1075 );
buf ( n308 , n1076 );
buf ( n309 , n1077 );
buf ( n310 , n1078 );
buf ( n311 , n1079 );
buf ( n312 , n1080 );
buf ( n313 , n1081 );
buf ( n314 , n1082 );
buf ( n315 , n1083 );
buf ( n316 , n1084 );
buf ( n317 , n1085 );
buf ( n318 , n1086 );
buf ( n319 , n1087 );
buf ( n320 , n1088 );
buf ( n321 , n1089 );
buf ( n322 , n1090 );
buf ( n323 , n1091 );
buf ( n324 , n1092 );
buf ( n325 , n1093 );
buf ( n326 , n1094 );
buf ( n327 , n1095 );
buf ( n328 , n1096 );
buf ( n329 , n1097 );
buf ( n330 , n1098 );
buf ( n331 , n1099 );
buf ( n332 , n1100 );
buf ( n333 , n1101 );
buf ( n334 , n1102 );
buf ( n335 , n1103 );
buf ( n336 , n1104 );
buf ( n337 , n1105 );
buf ( n338 , n1106 );
buf ( n339 , n1107 );
buf ( n340 , n1108 );
buf ( n341 , n1109 );
buf ( n342 , n1110 );
buf ( n343 , n1111 );
buf ( n344 , n1112 );
buf ( n345 , n1113 );
buf ( n346 , n1114 );
buf ( n347 , n1115 );
buf ( n348 , n1116 );
buf ( n349 , n1117 );
buf ( n350 , n1118 );
buf ( n351 , n1119 );
buf ( n352 , n1120 );
buf ( n353 , n1121 );
buf ( n354 , n1122 );
buf ( n355 , n1123 );
buf ( n356 , n1124 );
buf ( n357 , n1125 );
buf ( n358 , n1126 );
buf ( n359 , n1127 );
buf ( n360 , n1128 );
buf ( n361 , n1129 );
buf ( n362 , n1130 );
buf ( n363 , n1131 );
buf ( n364 , n1132 );
buf ( n365 , n1133 );
buf ( n366 , n1134 );
buf ( n367 , n1135 );
buf ( n368 , n1136 );
buf ( n369 , n1137 );
buf ( n370 , n1138 );
buf ( n371 , n1139 );
buf ( n372 , n1140 );
buf ( n373 , n1141 );
buf ( n374 , n1142 );
buf ( n375 , n1143 );
buf ( n376 , n1144 );
buf ( n377 , n1145 );
buf ( n378 , n1146 );
buf ( n379 , n1147 );
buf ( n380 , n1148 );
buf ( n381 , n1149 );
buf ( n382 , n1150 );
buf ( n383 , n1151 );
buf ( n896 , n41801 );
buf ( n897 , n41803 );
buf ( n898 , n41805 );
buf ( n899 , n41807 );
buf ( n900 , n41809 );
buf ( n901 , n41812 );
buf ( n902 , n41815 );
buf ( n903 , n41818 );
buf ( n904 , n41821 );
buf ( n905 , n41824 );
buf ( n906 , n41827 );
buf ( n907 , n41830 );
buf ( n908 , n41833 );
buf ( n909 , n41836 );
buf ( n910 , n41839 );
buf ( n911 , n41842 );
buf ( n912 , n41845 );
buf ( n913 , n41848 );
buf ( n914 , n41851 );
buf ( n915 , n41854 );
buf ( n916 , n41857 );
buf ( n917 , n41860 );
buf ( n918 , n41863 );
buf ( n919 , n41866 );
buf ( n920 , n41869 );
buf ( n921 , n41872 );
buf ( n922 , n41875 );
buf ( n923 , n41878 );
buf ( n924 , n41881 );
buf ( n925 , n41884 );
buf ( n926 , n41887 );
buf ( n927 , n41890 );
buf ( n928 , n41893 );
buf ( n929 , n41896 );
buf ( n930 , n41899 );
buf ( n931 , n41902 );
buf ( n932 , n41905 );
buf ( n933 , n41908 );
buf ( n934 , n41911 );
buf ( n935 , n41914 );
buf ( n936 , n41917 );
buf ( n937 , n41920 );
buf ( n938 , n41923 );
buf ( n939 , n41926 );
buf ( n940 , n41929 );
buf ( n941 , n41932 );
buf ( n942 , n41935 );
buf ( n943 , n41938 );
buf ( n944 , n41941 );
buf ( n945 , n41944 );
buf ( n946 , n41947 );
buf ( n947 , n41950 );
buf ( n948 , n41953 );
buf ( n949 , n41956 );
buf ( n950 , n41959 );
buf ( n951 , n41962 );
buf ( n952 , n41965 );
buf ( n953 , n41968 );
buf ( n954 , n41971 );
buf ( n955 , n41974 );
buf ( n956 , n41977 );
buf ( n957 , n41980 );
buf ( n958 , n41983 );
buf ( n959 , n41985 );
buf ( n960 , n41255 );
buf ( n961 , n41257 );
buf ( n962 , n41259 );
buf ( n963 , n41261 );
buf ( n964 , n41263 );
buf ( n965 , n41266 );
buf ( n966 , n41269 );
buf ( n967 , n41272 );
buf ( n968 , n41275 );
buf ( n969 , n41278 );
buf ( n970 , n41281 );
buf ( n971 , n41284 );
buf ( n972 , n41287 );
buf ( n973 , n41290 );
buf ( n974 , n41293 );
buf ( n975 , n41296 );
buf ( n976 , n41299 );
buf ( n977 , n41302 );
buf ( n978 , n41305 );
buf ( n979 , n41308 );
buf ( n980 , n41311 );
buf ( n981 , n41314 );
buf ( n982 , n41317 );
buf ( n983 , n41320 );
buf ( n984 , n41323 );
buf ( n985 , n41326 );
buf ( n986 , n41329 );
buf ( n987 , n41332 );
buf ( n988 , n41335 );
buf ( n989 , n41338 );
buf ( n990 , n41341 );
buf ( n991 , n41344 );
buf ( n992 , n41347 );
buf ( n993 , n41350 );
buf ( n994 , n41353 );
buf ( n995 , n41356 );
buf ( n996 , n41359 );
buf ( n997 , n41362 );
buf ( n998 , n41365 );
buf ( n999 , n41368 );
buf ( n1000 , n41371 );
buf ( n1001 , n41374 );
buf ( n1002 , n41377 );
buf ( n1003 , n41380 );
buf ( n1004 , n41383 );
buf ( n1005 , n41386 );
buf ( n1006 , n41389 );
buf ( n1007 , n41392 );
buf ( n1008 , n41395 );
buf ( n1009 , n41398 );
buf ( n1010 , n41401 );
buf ( n1011 , n41404 );
buf ( n1012 , n41407 );
buf ( n1013 , n41410 );
buf ( n1014 , n41413 );
buf ( n1015 , n41416 );
buf ( n1016 , n41419 );
buf ( n1017 , n41422 );
buf ( n1018 , n41425 );
buf ( n1019 , n41428 );
buf ( n1020 , n41431 );
buf ( n1021 , n41434 );
buf ( n1022 , n41437 );
buf ( n1023 , n41439 );
buf ( n1024 , n40639 );
buf ( n1025 , n40641 );
buf ( n1026 , n40643 );
buf ( n1027 , n40645 );
buf ( n1028 , n40647 );
buf ( n1029 , n40649 );
buf ( n1030 , n40651 );
buf ( n1031 , n40653 );
buf ( n1032 , n40655 );
buf ( n1033 , n40657 );
buf ( n1034 , n40659 );
buf ( n1035 , n40661 );
buf ( n1036 , n40663 );
buf ( n1037 , n40665 );
buf ( n1038 , n40667 );
buf ( n1039 , n40669 );
buf ( n1040 , n40671 );
buf ( n1041 , n40673 );
buf ( n1042 , n40675 );
buf ( n1043 , n40677 );
buf ( n1044 , n40679 );
buf ( n1045 , n40681 );
buf ( n1046 , n40683 );
buf ( n1047 , n40685 );
buf ( n1048 , n40687 );
buf ( n1049 , n40689 );
buf ( n1050 , n40691 );
buf ( n1051 , n40693 );
buf ( n1052 , n40695 );
buf ( n1053 , n40697 );
buf ( n1054 , n40699 );
buf ( n1055 , n40701 );
buf ( n1056 , n40703 );
buf ( n1057 , n40705 );
buf ( n1058 , n40707 );
buf ( n1059 , n40709 );
buf ( n1060 , n40711 );
buf ( n1061 , n40713 );
buf ( n1062 , n40715 );
buf ( n1063 , n40717 );
buf ( n1064 , n40719 );
buf ( n1065 , n40721 );
buf ( n1066 , n40723 );
buf ( n1067 , n40725 );
buf ( n1068 , n40727 );
buf ( n1069 , n40729 );
buf ( n1070 , n40731 );
buf ( n1071 , n40733 );
buf ( n1072 , n40735 );
buf ( n1073 , n40737 );
buf ( n1074 , n40739 );
buf ( n1075 , n40741 );
buf ( n1076 , n40743 );
buf ( n1077 , n40745 );
buf ( n1078 , n40747 );
buf ( n1079 , n40749 );
buf ( n1080 , n40751 );
buf ( n1081 , n40753 );
buf ( n1082 , n40755 );
buf ( n1083 , n40757 );
buf ( n1084 , n40759 );
buf ( n1085 , n40761 );
buf ( n1086 , n40763 );
buf ( n1087 , n40765 );
buf ( n1088 , n40767 );
buf ( n1089 , n40769 );
buf ( n1090 , n40771 );
buf ( n1091 , n40773 );
buf ( n1092 , n40775 );
buf ( n1093 , n40777 );
buf ( n1094 , n40779 );
buf ( n1095 , n40781 );
buf ( n1096 , n40783 );
buf ( n1097 , n40785 );
buf ( n1098 , n40787 );
buf ( n1099 , n40789 );
buf ( n1100 , n40791 );
buf ( n1101 , n40793 );
buf ( n1102 , n40795 );
buf ( n1103 , n40797 );
buf ( n1104 , n40799 );
buf ( n1105 , n40801 );
buf ( n1106 , n40803 );
buf ( n1107 , n40805 );
buf ( n1108 , n40807 );
buf ( n1109 , n40809 );
buf ( n1110 , n40811 );
buf ( n1111 , n40813 );
buf ( n1112 , n40815 );
buf ( n1113 , n40817 );
buf ( n1114 , n40819 );
buf ( n1115 , n40821 );
buf ( n1116 , n40823 );
buf ( n1117 , n40825 );
buf ( n1118 , n40827 );
buf ( n1119 , n40829 );
buf ( n1120 , n40831 );
buf ( n1121 , n40833 );
buf ( n1122 , n40835 );
buf ( n1123 , n40837 );
buf ( n1124 , n40839 );
buf ( n1125 , n40841 );
buf ( n1126 , n40843 );
buf ( n1127 , n40845 );
buf ( n1128 , n40847 );
buf ( n1129 , n40849 );
buf ( n1130 , n40851 );
buf ( n1131 , n40853 );
buf ( n1132 , n40855 );
buf ( n1133 , n40857 );
buf ( n1134 , n40859 );
buf ( n1135 , n40861 );
buf ( n1136 , n40863 );
buf ( n1137 , n40865 );
buf ( n1138 , n40867 );
buf ( n1139 , n40869 );
buf ( n1140 , n40871 );
buf ( n1141 , n40873 );
buf ( n1142 , n40875 );
buf ( n1143 , n40877 );
buf ( n1144 , n40879 );
buf ( n1145 , n40881 );
buf ( n1146 , n40883 );
buf ( n1147 , n40885 );
buf ( n1148 , n40887 );
buf ( n1149 , n40889 );
buf ( n1150 , n40891 );
buf ( n1151 , n40893 );
buf ( n1152 , n832 );
buf ( n1153 , n833 );
buf ( n1154 , n834 );
buf ( n1155 , n835 );
buf ( n1156 , n836 );
buf ( n1157 , n837 );
buf ( n1158 , n838 );
buf ( n1159 , n839 );
buf ( n1160 , n840 );
buf ( n1161 , n841 );
buf ( n1162 , n842 );
buf ( n1163 , n843 );
buf ( n1164 , n844 );
buf ( n1165 , n845 );
buf ( n1166 , n846 );
buf ( n1167 , n847 );
buf ( n1168 , n848 );
buf ( n1169 , n849 );
buf ( n1170 , n850 );
buf ( n1171 , n851 );
buf ( n1172 , n852 );
buf ( n1173 , n853 );
buf ( n1174 , n854 );
buf ( n1175 , n855 );
buf ( n1176 , n856 );
buf ( n1177 , n857 );
buf ( n1178 , n858 );
buf ( n1179 , n859 );
buf ( n1180 , n860 );
buf ( n1181 , n861 );
buf ( n1182 , n862 );
buf ( n1183 , n863 );
buf ( n1184 , n864 );
buf ( n1185 , n865 );
buf ( n1186 , n866 );
buf ( n1187 , n867 );
buf ( n1188 , n868 );
buf ( n1189 , n869 );
buf ( n1190 , n870 );
buf ( n1191 , n871 );
buf ( n1192 , n872 );
buf ( n1193 , n873 );
buf ( n1194 , n874 );
buf ( n1195 , n875 );
buf ( n1196 , n876 );
buf ( n1197 , n877 );
buf ( n1198 , n878 );
buf ( n1199 , n879 );
buf ( n1200 , n880 );
buf ( n1201 , n881 );
buf ( n1202 , n882 );
buf ( n1203 , n883 );
buf ( n1204 , n884 );
buf ( n1205 , n885 );
buf ( n1206 , n886 );
buf ( n1207 , n887 );
buf ( n1208 , n888 );
buf ( n1209 , n889 );
buf ( n1210 , n890 );
buf ( n1211 , n891 );
buf ( n1212 , n892 );
buf ( n1213 , n893 );
buf ( n1214 , n894 );
buf ( n1215 , n895 );
buf ( n1216 , n1186 );
buf ( n1217 , n1187 );
buf ( n1218 , n1188 );
and ( n1219 , n1217 , n1218 );
not ( n1220 , n1219 );
and ( n1221 , n1216 , n1220 );
not ( n1222 , n1221 );
buf ( n1223 , n1153 );
buf ( n1224 , n1184 );
buf ( n1225 , n1185 );
xor ( n1226 , n1224 , n1225 );
xor ( n1227 , n1225 , n1216 );
not ( n1228 , n1227 );
and ( n1229 , n1226 , n1228 );
and ( n1230 , n1223 , n1229 );
buf ( n1231 , n1152 );
and ( n1232 , n1231 , n1227 );
nor ( n1233 , n1230 , n1232 );
and ( n1234 , n1225 , n1216 );
not ( n1235 , n1234 );
and ( n1236 , n1224 , n1235 );
xnor ( n1237 , n1233 , n1236 );
and ( n1238 , n1222 , n1237 );
buf ( n1239 , n1154 );
and ( n1240 , n1239 , n1224 );
and ( n1241 , n1237 , n1240 );
and ( n1242 , n1222 , n1240 );
or ( n1243 , n1238 , n1241 , n1242 );
and ( n1244 , n1231 , n1229 );
not ( n1245 , n1244 );
xnor ( n1246 , n1245 , n1236 );
and ( n1247 , n1243 , n1246 );
and ( n1248 , n1223 , n1224 );
not ( n1249 , n1248 );
and ( n1250 , n1246 , n1249 );
and ( n1251 , n1243 , n1249 );
or ( n1252 , n1247 , n1250 , n1251 );
buf ( n1253 , n1248 );
not ( n1254 , n1236 );
xor ( n1255 , n1253 , n1254 );
and ( n1256 , n1231 , n1224 );
xor ( n1257 , n1255 , n1256 );
xor ( n1258 , n1252 , n1257 );
xor ( n1259 , n1243 , n1246 );
xor ( n1260 , n1259 , n1249 );
xor ( n1261 , n1216 , n1217 );
xor ( n1262 , n1217 , n1218 );
not ( n1263 , n1262 );
and ( n1264 , n1261 , n1263 );
and ( n1265 , n1231 , n1264 );
not ( n1266 , n1265 );
xnor ( n1267 , n1266 , n1221 );
not ( n1268 , n1267 );
and ( n1269 , n1239 , n1229 );
and ( n1270 , n1223 , n1227 );
nor ( n1271 , n1269 , n1270 );
xnor ( n1272 , n1271 , n1236 );
and ( n1273 , n1268 , n1272 );
buf ( n1274 , n1155 );
and ( n1275 , n1274 , n1224 );
and ( n1276 , n1272 , n1275 );
and ( n1277 , n1268 , n1275 );
or ( n1278 , n1273 , n1276 , n1277 );
buf ( n1279 , n1267 );
and ( n1280 , n1278 , n1279 );
xor ( n1281 , n1222 , n1237 );
xor ( n1282 , n1281 , n1240 );
and ( n1283 , n1279 , n1282 );
and ( n1284 , n1278 , n1282 );
or ( n1285 , n1280 , n1283 , n1284 );
and ( n1286 , n1260 , n1285 );
xor ( n1287 , n1278 , n1279 );
xor ( n1288 , n1287 , n1282 );
buf ( n1289 , n1189 );
buf ( n1290 , n1190 );
and ( n1291 , n1289 , n1290 );
not ( n1292 , n1291 );
and ( n1293 , n1218 , n1292 );
not ( n1294 , n1293 );
and ( n1295 , n1223 , n1264 );
and ( n1296 , n1231 , n1262 );
nor ( n1297 , n1295 , n1296 );
xnor ( n1298 , n1297 , n1221 );
and ( n1299 , n1294 , n1298 );
buf ( n1300 , n1156 );
and ( n1301 , n1300 , n1224 );
and ( n1302 , n1298 , n1301 );
and ( n1303 , n1294 , n1301 );
or ( n1304 , n1299 , n1302 , n1303 );
and ( n1305 , n1239 , n1264 );
and ( n1306 , n1223 , n1262 );
nor ( n1307 , n1305 , n1306 );
xnor ( n1308 , n1307 , n1221 );
and ( n1309 , n1300 , n1229 );
and ( n1310 , n1274 , n1227 );
nor ( n1311 , n1309 , n1310 );
xnor ( n1312 , n1311 , n1236 );
and ( n1313 , n1308 , n1312 );
buf ( n1314 , n1157 );
and ( n1315 , n1314 , n1224 );
and ( n1316 , n1312 , n1315 );
and ( n1317 , n1308 , n1315 );
or ( n1318 , n1313 , n1316 , n1317 );
xor ( n1319 , n1218 , n1289 );
xor ( n1320 , n1289 , n1290 );
not ( n1321 , n1320 );
and ( n1322 , n1319 , n1321 );
and ( n1323 , n1231 , n1322 );
not ( n1324 , n1323 );
xnor ( n1325 , n1324 , n1293 );
buf ( n1326 , n1325 );
and ( n1327 , n1318 , n1326 );
and ( n1328 , n1274 , n1229 );
and ( n1329 , n1239 , n1227 );
nor ( n1330 , n1328 , n1329 );
xnor ( n1331 , n1330 , n1236 );
and ( n1332 , n1326 , n1331 );
and ( n1333 , n1318 , n1331 );
or ( n1334 , n1327 , n1332 , n1333 );
and ( n1335 , n1304 , n1334 );
xor ( n1336 , n1268 , n1272 );
xor ( n1337 , n1336 , n1275 );
and ( n1338 , n1334 , n1337 );
and ( n1339 , n1304 , n1337 );
or ( n1340 , n1335 , n1338 , n1339 );
and ( n1341 , n1288 , n1340 );
xor ( n1342 , n1304 , n1334 );
xor ( n1343 , n1342 , n1337 );
buf ( n1344 , n1191 );
buf ( n1345 , n1192 );
and ( n1346 , n1344 , n1345 );
not ( n1347 , n1346 );
and ( n1348 , n1290 , n1347 );
not ( n1349 , n1348 );
and ( n1350 , n1223 , n1322 );
and ( n1351 , n1231 , n1320 );
nor ( n1352 , n1350 , n1351 );
xnor ( n1353 , n1352 , n1293 );
and ( n1354 , n1349 , n1353 );
and ( n1355 , n1314 , n1229 );
and ( n1356 , n1300 , n1227 );
nor ( n1357 , n1355 , n1356 );
xnor ( n1358 , n1357 , n1236 );
and ( n1359 , n1353 , n1358 );
and ( n1360 , n1349 , n1358 );
or ( n1361 , n1354 , n1359 , n1360 );
not ( n1362 , n1325 );
and ( n1363 , n1361 , n1362 );
xor ( n1364 , n1308 , n1312 );
xor ( n1365 , n1364 , n1315 );
and ( n1366 , n1362 , n1365 );
and ( n1367 , n1361 , n1365 );
or ( n1368 , n1363 , n1366 , n1367 );
xor ( n1369 , n1294 , n1298 );
xor ( n1370 , n1369 , n1301 );
and ( n1371 , n1368 , n1370 );
xor ( n1372 , n1318 , n1326 );
xor ( n1373 , n1372 , n1331 );
and ( n1374 , n1370 , n1373 );
and ( n1375 , n1368 , n1373 );
or ( n1376 , n1371 , n1374 , n1375 );
and ( n1377 , n1343 , n1376 );
xor ( n1378 , n1368 , n1370 );
xor ( n1379 , n1378 , n1373 );
and ( n1380 , n1239 , n1322 );
and ( n1381 , n1223 , n1320 );
nor ( n1382 , n1380 , n1381 );
xnor ( n1383 , n1382 , n1293 );
buf ( n1384 , n1383 );
and ( n1385 , n1274 , n1264 );
and ( n1386 , n1239 , n1262 );
nor ( n1387 , n1385 , n1386 );
xnor ( n1388 , n1387 , n1221 );
and ( n1389 , n1384 , n1388 );
buf ( n1390 , n1158 );
and ( n1391 , n1390 , n1224 );
and ( n1392 , n1388 , n1391 );
and ( n1393 , n1384 , n1391 );
or ( n1394 , n1389 , n1392 , n1393 );
xor ( n1395 , n1290 , n1344 );
xor ( n1396 , n1344 , n1345 );
not ( n1397 , n1396 );
and ( n1398 , n1395 , n1397 );
and ( n1399 , n1231 , n1398 );
not ( n1400 , n1399 );
xnor ( n1401 , n1400 , n1348 );
and ( n1402 , n1390 , n1229 );
and ( n1403 , n1314 , n1227 );
nor ( n1404 , n1402 , n1403 );
xnor ( n1405 , n1404 , n1236 );
and ( n1406 , n1401 , n1405 );
buf ( n1407 , n1159 );
and ( n1408 , n1407 , n1224 );
and ( n1409 , n1405 , n1408 );
and ( n1410 , n1401 , n1408 );
or ( n1411 , n1406 , n1409 , n1410 );
xor ( n1412 , n1349 , n1353 );
xor ( n1413 , n1412 , n1358 );
and ( n1414 , n1411 , n1413 );
xor ( n1415 , n1384 , n1388 );
xor ( n1416 , n1415 , n1391 );
and ( n1417 , n1413 , n1416 );
and ( n1418 , n1411 , n1416 );
or ( n1419 , n1414 , n1417 , n1418 );
and ( n1420 , n1394 , n1419 );
xor ( n1421 , n1361 , n1362 );
xor ( n1422 , n1421 , n1365 );
and ( n1423 , n1419 , n1422 );
and ( n1424 , n1394 , n1422 );
or ( n1425 , n1420 , n1423 , n1424 );
and ( n1426 , n1379 , n1425 );
xor ( n1427 , n1394 , n1419 );
xor ( n1428 , n1427 , n1422 );
and ( n1429 , n1274 , n1322 );
and ( n1430 , n1239 , n1320 );
nor ( n1431 , n1429 , n1430 );
xnor ( n1432 , n1431 , n1293 );
and ( n1433 , n1407 , n1229 );
and ( n1434 , n1390 , n1227 );
nor ( n1435 , n1433 , n1434 );
xnor ( n1436 , n1435 , n1236 );
and ( n1437 , n1432 , n1436 );
buf ( n1438 , n1160 );
and ( n1439 , n1438 , n1224 );
and ( n1440 , n1436 , n1439 );
and ( n1441 , n1432 , n1439 );
or ( n1442 , n1437 , n1440 , n1441 );
not ( n1443 , n1383 );
and ( n1444 , n1442 , n1443 );
and ( n1445 , n1300 , n1264 );
and ( n1446 , n1274 , n1262 );
nor ( n1447 , n1445 , n1446 );
xnor ( n1448 , n1447 , n1221 );
and ( n1449 , n1443 , n1448 );
and ( n1450 , n1442 , n1448 );
or ( n1451 , n1444 , n1449 , n1450 );
buf ( n1452 , n1193 );
buf ( n1453 , n1194 );
and ( n1454 , n1452 , n1453 );
not ( n1455 , n1454 );
and ( n1456 , n1345 , n1455 );
not ( n1457 , n1456 );
and ( n1458 , n1223 , n1398 );
and ( n1459 , n1231 , n1396 );
nor ( n1460 , n1458 , n1459 );
xnor ( n1461 , n1460 , n1348 );
and ( n1462 , n1457 , n1461 );
and ( n1463 , n1314 , n1264 );
and ( n1464 , n1300 , n1262 );
nor ( n1465 , n1463 , n1464 );
xnor ( n1466 , n1465 , n1221 );
and ( n1467 , n1461 , n1466 );
and ( n1468 , n1457 , n1466 );
or ( n1469 , n1462 , n1467 , n1468 );
xor ( n1470 , n1401 , n1405 );
xor ( n1471 , n1470 , n1408 );
and ( n1472 , n1469 , n1471 );
xor ( n1473 , n1442 , n1443 );
xor ( n1474 , n1473 , n1448 );
and ( n1475 , n1471 , n1474 );
and ( n1476 , n1469 , n1474 );
or ( n1477 , n1472 , n1475 , n1476 );
and ( n1478 , n1451 , n1477 );
xor ( n1479 , n1411 , n1413 );
xor ( n1480 , n1479 , n1416 );
and ( n1481 , n1477 , n1480 );
and ( n1482 , n1451 , n1480 );
or ( n1483 , n1478 , n1481 , n1482 );
and ( n1484 , n1428 , n1483 );
xor ( n1485 , n1345 , n1452 );
xor ( n1486 , n1452 , n1453 );
not ( n1487 , n1486 );
and ( n1488 , n1485 , n1487 );
and ( n1489 , n1231 , n1488 );
not ( n1490 , n1489 );
xnor ( n1491 , n1490 , n1456 );
and ( n1492 , n1390 , n1264 );
and ( n1493 , n1314 , n1262 );
nor ( n1494 , n1492 , n1493 );
xnor ( n1495 , n1494 , n1221 );
and ( n1496 , n1491 , n1495 );
and ( n1497 , n1438 , n1229 );
and ( n1498 , n1407 , n1227 );
nor ( n1499 , n1497 , n1498 );
xnor ( n1500 , n1499 , n1236 );
and ( n1501 , n1495 , n1500 );
and ( n1502 , n1491 , n1500 );
or ( n1503 , n1496 , n1501 , n1502 );
and ( n1504 , n1239 , n1398 );
and ( n1505 , n1223 , n1396 );
nor ( n1506 , n1504 , n1505 );
xnor ( n1507 , n1506 , n1348 );
buf ( n1508 , n1507 );
and ( n1509 , n1503 , n1508 );
xor ( n1510 , n1432 , n1436 );
xor ( n1511 , n1510 , n1439 );
and ( n1512 , n1508 , n1511 );
and ( n1513 , n1503 , n1511 );
or ( n1514 , n1509 , n1512 , n1513 );
not ( n1515 , n1507 );
and ( n1516 , n1300 , n1322 );
and ( n1517 , n1274 , n1320 );
nor ( n1518 , n1516 , n1517 );
xnor ( n1519 , n1518 , n1293 );
and ( n1520 , n1515 , n1519 );
buf ( n1521 , n1161 );
and ( n1522 , n1521 , n1224 );
and ( n1523 , n1519 , n1522 );
and ( n1524 , n1515 , n1522 );
or ( n1525 , n1520 , n1523 , n1524 );
xor ( n1526 , n1457 , n1461 );
xor ( n1527 , n1526 , n1466 );
and ( n1528 , n1525 , n1527 );
xor ( n1529 , n1503 , n1508 );
xor ( n1530 , n1529 , n1511 );
and ( n1531 , n1527 , n1530 );
and ( n1532 , n1525 , n1530 );
or ( n1533 , n1528 , n1531 , n1532 );
and ( n1534 , n1514 , n1533 );
xor ( n1535 , n1469 , n1471 );
xor ( n1536 , n1535 , n1474 );
and ( n1537 , n1533 , n1536 );
and ( n1538 , n1514 , n1536 );
or ( n1539 , n1534 , n1537 , n1538 );
xor ( n1540 , n1451 , n1477 );
xor ( n1541 , n1540 , n1480 );
and ( n1542 , n1539 , n1541 );
xor ( n1543 , n1514 , n1533 );
xor ( n1544 , n1543 , n1536 );
buf ( n1545 , n1195 );
buf ( n1546 , n1196 );
and ( n1547 , n1545 , n1546 );
not ( n1548 , n1547 );
and ( n1549 , n1453 , n1548 );
not ( n1550 , n1549 );
and ( n1551 , n1223 , n1488 );
and ( n1552 , n1231 , n1486 );
nor ( n1553 , n1551 , n1552 );
xnor ( n1554 , n1553 , n1456 );
and ( n1555 , n1550 , n1554 );
and ( n1556 , n1314 , n1322 );
and ( n1557 , n1300 , n1320 );
nor ( n1558 , n1556 , n1557 );
xnor ( n1559 , n1558 , n1293 );
and ( n1560 , n1554 , n1559 );
and ( n1561 , n1550 , n1559 );
or ( n1562 , n1555 , n1560 , n1561 );
and ( n1563 , n1274 , n1398 );
and ( n1564 , n1239 , n1396 );
nor ( n1565 , n1563 , n1564 );
xnor ( n1566 , n1565 , n1348 );
and ( n1567 , n1407 , n1264 );
and ( n1568 , n1390 , n1262 );
nor ( n1569 , n1567 , n1568 );
xnor ( n1570 , n1569 , n1221 );
and ( n1571 , n1566 , n1570 );
and ( n1572 , n1521 , n1229 );
and ( n1573 , n1438 , n1227 );
nor ( n1574 , n1572 , n1573 );
xnor ( n1575 , n1574 , n1236 );
and ( n1576 , n1570 , n1575 );
and ( n1577 , n1566 , n1575 );
or ( n1578 , n1571 , n1576 , n1577 );
and ( n1579 , n1562 , n1578 );
xor ( n1580 , n1491 , n1495 );
xor ( n1581 , n1580 , n1500 );
and ( n1582 , n1578 , n1581 );
and ( n1583 , n1562 , n1581 );
or ( n1584 , n1579 , n1582 , n1583 );
and ( n1585 , n1239 , n1488 );
and ( n1586 , n1223 , n1486 );
nor ( n1587 , n1585 , n1586 );
xnor ( n1588 , n1587 , n1456 );
and ( n1589 , n1390 , n1322 );
and ( n1590 , n1314 , n1320 );
nor ( n1591 , n1589 , n1590 );
xnor ( n1592 , n1591 , n1293 );
and ( n1593 , n1588 , n1592 );
and ( n1594 , n1438 , n1264 );
and ( n1595 , n1407 , n1262 );
nor ( n1596 , n1594 , n1595 );
xnor ( n1597 , n1596 , n1221 );
and ( n1598 , n1592 , n1597 );
and ( n1599 , n1588 , n1597 );
or ( n1600 , n1593 , n1598 , n1599 );
xor ( n1601 , n1453 , n1545 );
xor ( n1602 , n1545 , n1546 );
not ( n1603 , n1602 );
and ( n1604 , n1601 , n1603 );
and ( n1605 , n1231 , n1604 );
not ( n1606 , n1605 );
xnor ( n1607 , n1606 , n1549 );
buf ( n1608 , n1607 );
and ( n1609 , n1600 , n1608 );
buf ( n1610 , n1162 );
and ( n1611 , n1610 , n1224 );
and ( n1612 , n1608 , n1611 );
and ( n1613 , n1600 , n1611 );
or ( n1614 , n1609 , n1612 , n1613 );
and ( n1615 , n1300 , n1398 );
and ( n1616 , n1274 , n1396 );
nor ( n1617 , n1615 , n1616 );
xnor ( n1618 , n1617 , n1348 );
and ( n1619 , n1610 , n1229 );
and ( n1620 , n1521 , n1227 );
nor ( n1621 , n1619 , n1620 );
xnor ( n1622 , n1621 , n1236 );
and ( n1623 , n1618 , n1622 );
buf ( n1624 , n1163 );
and ( n1625 , n1624 , n1224 );
and ( n1626 , n1622 , n1625 );
and ( n1627 , n1618 , n1625 );
or ( n1628 , n1623 , n1626 , n1627 );
xor ( n1629 , n1550 , n1554 );
xor ( n1630 , n1629 , n1559 );
and ( n1631 , n1628 , n1630 );
xor ( n1632 , n1566 , n1570 );
xor ( n1633 , n1632 , n1575 );
and ( n1634 , n1630 , n1633 );
and ( n1635 , n1628 , n1633 );
or ( n1636 , n1631 , n1634 , n1635 );
and ( n1637 , n1614 , n1636 );
xor ( n1638 , n1515 , n1519 );
xor ( n1639 , n1638 , n1522 );
and ( n1640 , n1636 , n1639 );
and ( n1641 , n1614 , n1639 );
or ( n1642 , n1637 , n1640 , n1641 );
and ( n1643 , n1584 , n1642 );
xor ( n1644 , n1525 , n1527 );
xor ( n1645 , n1644 , n1530 );
and ( n1646 , n1642 , n1645 );
and ( n1647 , n1584 , n1645 );
or ( n1648 , n1643 , n1646 , n1647 );
and ( n1649 , n1544 , n1648 );
xor ( n1650 , n1584 , n1642 );
xor ( n1651 , n1650 , n1645 );
and ( n1652 , n1274 , n1488 );
and ( n1653 , n1239 , n1486 );
nor ( n1654 , n1652 , n1653 );
xnor ( n1655 , n1654 , n1456 );
and ( n1656 , n1407 , n1322 );
and ( n1657 , n1390 , n1320 );
nor ( n1658 , n1656 , n1657 );
xnor ( n1659 , n1658 , n1293 );
and ( n1660 , n1655 , n1659 );
buf ( n1661 , n1164 );
and ( n1662 , n1661 , n1224 );
and ( n1663 , n1659 , n1662 );
and ( n1664 , n1655 , n1662 );
or ( n1665 , n1660 , n1663 , n1664 );
buf ( n1666 , n1197 );
buf ( n1667 , n1198 );
and ( n1668 , n1666 , n1667 );
not ( n1669 , n1668 );
and ( n1670 , n1546 , n1669 );
not ( n1671 , n1670 );
and ( n1672 , n1223 , n1604 );
and ( n1673 , n1231 , n1602 );
nor ( n1674 , n1672 , n1673 );
xnor ( n1675 , n1674 , n1549 );
and ( n1676 , n1671 , n1675 );
and ( n1677 , n1314 , n1398 );
and ( n1678 , n1300 , n1396 );
nor ( n1679 , n1677 , n1678 );
xnor ( n1680 , n1679 , n1348 );
and ( n1681 , n1675 , n1680 );
and ( n1682 , n1671 , n1680 );
or ( n1683 , n1676 , n1681 , n1682 );
and ( n1684 , n1665 , n1683 );
not ( n1685 , n1607 );
and ( n1686 , n1683 , n1685 );
and ( n1687 , n1665 , n1685 );
or ( n1688 , n1684 , n1686 , n1687 );
xor ( n1689 , n1546 , n1666 );
xor ( n1690 , n1666 , n1667 );
not ( n1691 , n1690 );
and ( n1692 , n1689 , n1691 );
and ( n1693 , n1231 , n1692 );
not ( n1694 , n1693 );
xnor ( n1695 , n1694 , n1670 );
buf ( n1696 , n1695 );
and ( n1697 , n1521 , n1264 );
and ( n1698 , n1438 , n1262 );
nor ( n1699 , n1697 , n1698 );
xnor ( n1700 , n1699 , n1221 );
and ( n1701 , n1696 , n1700 );
and ( n1702 , n1624 , n1229 );
and ( n1703 , n1610 , n1227 );
nor ( n1704 , n1702 , n1703 );
xnor ( n1705 , n1704 , n1236 );
and ( n1706 , n1700 , n1705 );
and ( n1707 , n1696 , n1705 );
or ( n1708 , n1701 , n1706 , n1707 );
xor ( n1709 , n1618 , n1622 );
xor ( n1710 , n1709 , n1625 );
and ( n1711 , n1708 , n1710 );
xor ( n1712 , n1588 , n1592 );
xor ( n1713 , n1712 , n1597 );
and ( n1714 , n1710 , n1713 );
and ( n1715 , n1708 , n1713 );
or ( n1716 , n1711 , n1714 , n1715 );
and ( n1717 , n1688 , n1716 );
xor ( n1718 , n1600 , n1608 );
xor ( n1719 , n1718 , n1611 );
and ( n1720 , n1716 , n1719 );
and ( n1721 , n1688 , n1719 );
or ( n1722 , n1717 , n1720 , n1721 );
xor ( n1723 , n1562 , n1578 );
xor ( n1724 , n1723 , n1581 );
and ( n1725 , n1722 , n1724 );
xor ( n1726 , n1614 , n1636 );
xor ( n1727 , n1726 , n1639 );
and ( n1728 , n1724 , n1727 );
and ( n1729 , n1722 , n1727 );
or ( n1730 , n1725 , n1728 , n1729 );
and ( n1731 , n1651 , n1730 );
xor ( n1732 , n1722 , n1724 );
xor ( n1733 , n1732 , n1727 );
and ( n1734 , n1300 , n1488 );
and ( n1735 , n1274 , n1486 );
nor ( n1736 , n1734 , n1735 );
xnor ( n1737 , n1736 , n1456 );
and ( n1738 , n1438 , n1322 );
and ( n1739 , n1407 , n1320 );
nor ( n1740 , n1738 , n1739 );
xnor ( n1741 , n1740 , n1293 );
and ( n1742 , n1737 , n1741 );
and ( n1743 , n1610 , n1264 );
and ( n1744 , n1521 , n1262 );
nor ( n1745 , n1743 , n1744 );
xnor ( n1746 , n1745 , n1221 );
and ( n1747 , n1741 , n1746 );
and ( n1748 , n1737 , n1746 );
or ( n1749 , n1742 , n1747 , n1748 );
and ( n1750 , n1239 , n1604 );
and ( n1751 , n1223 , n1602 );
nor ( n1752 , n1750 , n1751 );
xnor ( n1753 , n1752 , n1549 );
and ( n1754 , n1390 , n1398 );
and ( n1755 , n1314 , n1396 );
nor ( n1756 , n1754 , n1755 );
xnor ( n1757 , n1756 , n1348 );
and ( n1758 , n1753 , n1757 );
buf ( n1759 , n1165 );
and ( n1760 , n1759 , n1224 );
and ( n1761 , n1757 , n1760 );
and ( n1762 , n1753 , n1760 );
or ( n1763 , n1758 , n1761 , n1762 );
and ( n1764 , n1749 , n1763 );
xor ( n1765 , n1671 , n1675 );
xor ( n1766 , n1765 , n1680 );
and ( n1767 , n1763 , n1766 );
and ( n1768 , n1749 , n1766 );
or ( n1769 , n1764 , n1767 , n1768 );
xor ( n1770 , n1665 , n1683 );
xor ( n1771 , n1770 , n1685 );
and ( n1772 , n1769 , n1771 );
xor ( n1773 , n1708 , n1710 );
xor ( n1774 , n1773 , n1713 );
and ( n1775 , n1771 , n1774 );
and ( n1776 , n1769 , n1774 );
or ( n1777 , n1772 , n1775 , n1776 );
xor ( n1778 , n1628 , n1630 );
xor ( n1779 , n1778 , n1633 );
and ( n1780 , n1777 , n1779 );
xor ( n1781 , n1688 , n1716 );
xor ( n1782 , n1781 , n1719 );
and ( n1783 , n1779 , n1782 );
and ( n1784 , n1777 , n1782 );
or ( n1785 , n1780 , n1783 , n1784 );
and ( n1786 , n1733 , n1785 );
xor ( n1787 , n1777 , n1779 );
xor ( n1788 , n1787 , n1782 );
buf ( n1789 , n1199 );
buf ( n1790 , n1200 );
and ( n1791 , n1789 , n1790 );
not ( n1792 , n1791 );
and ( n1793 , n1667 , n1792 );
not ( n1794 , n1793 );
and ( n1795 , n1223 , n1692 );
and ( n1796 , n1231 , n1690 );
nor ( n1797 , n1795 , n1796 );
xnor ( n1798 , n1797 , n1670 );
and ( n1799 , n1794 , n1798 );
and ( n1800 , n1314 , n1488 );
and ( n1801 , n1300 , n1486 );
nor ( n1802 , n1800 , n1801 );
xnor ( n1803 , n1802 , n1456 );
and ( n1804 , n1798 , n1803 );
and ( n1805 , n1794 , n1803 );
or ( n1806 , n1799 , n1804 , n1805 );
not ( n1807 , n1695 );
and ( n1808 , n1806 , n1807 );
and ( n1809 , n1661 , n1229 );
and ( n1810 , n1624 , n1227 );
nor ( n1811 , n1809 , n1810 );
xnor ( n1812 , n1811 , n1236 );
and ( n1813 , n1807 , n1812 );
and ( n1814 , n1806 , n1812 );
or ( n1815 , n1808 , n1813 , n1814 );
xor ( n1816 , n1655 , n1659 );
xor ( n1817 , n1816 , n1662 );
and ( n1818 , n1815 , n1817 );
xor ( n1819 , n1696 , n1700 );
xor ( n1820 , n1819 , n1705 );
and ( n1821 , n1817 , n1820 );
and ( n1822 , n1815 , n1820 );
or ( n1823 , n1818 , n1821 , n1822 );
and ( n1824 , n1407 , n1398 );
and ( n1825 , n1390 , n1396 );
nor ( n1826 , n1824 , n1825 );
xnor ( n1827 , n1826 , n1348 );
and ( n1828 , n1759 , n1229 );
and ( n1829 , n1661 , n1227 );
nor ( n1830 , n1828 , n1829 );
xnor ( n1831 , n1830 , n1236 );
and ( n1832 , n1827 , n1831 );
buf ( n1833 , n1166 );
and ( n1834 , n1833 , n1224 );
and ( n1835 , n1831 , n1834 );
and ( n1836 , n1827 , n1834 );
or ( n1837 , n1832 , n1835 , n1836 );
and ( n1838 , n1274 , n1604 );
and ( n1839 , n1239 , n1602 );
nor ( n1840 , n1838 , n1839 );
xnor ( n1841 , n1840 , n1549 );
and ( n1842 , n1521 , n1322 );
and ( n1843 , n1438 , n1320 );
nor ( n1844 , n1842 , n1843 );
xnor ( n1845 , n1844 , n1293 );
and ( n1846 , n1841 , n1845 );
and ( n1847 , n1624 , n1264 );
and ( n1848 , n1610 , n1262 );
nor ( n1849 , n1847 , n1848 );
xnor ( n1850 , n1849 , n1221 );
and ( n1851 , n1845 , n1850 );
and ( n1852 , n1841 , n1850 );
or ( n1853 , n1846 , n1851 , n1852 );
and ( n1854 , n1837 , n1853 );
xor ( n1855 , n1737 , n1741 );
xor ( n1856 , n1855 , n1746 );
and ( n1857 , n1853 , n1856 );
and ( n1858 , n1837 , n1856 );
or ( n1859 , n1854 , n1857 , n1858 );
and ( n1860 , n1390 , n1488 );
and ( n1861 , n1314 , n1486 );
nor ( n1862 , n1860 , n1861 );
xnor ( n1863 , n1862 , n1456 );
and ( n1864 , n1833 , n1229 );
and ( n1865 , n1759 , n1227 );
nor ( n1866 , n1864 , n1865 );
xnor ( n1867 , n1866 , n1236 );
and ( n1868 , n1863 , n1867 );
buf ( n1869 , n1167 );
and ( n1870 , n1869 , n1224 );
and ( n1871 , n1867 , n1870 );
and ( n1872 , n1863 , n1870 );
or ( n1873 , n1868 , n1871 , n1872 );
and ( n1874 , n1239 , n1692 );
and ( n1875 , n1223 , n1690 );
nor ( n1876 , n1874 , n1875 );
xnor ( n1877 , n1876 , n1670 );
and ( n1878 , n1300 , n1604 );
and ( n1879 , n1274 , n1602 );
nor ( n1880 , n1878 , n1879 );
xnor ( n1881 , n1880 , n1549 );
and ( n1882 , n1877 , n1881 );
and ( n1883 , n1438 , n1398 );
and ( n1884 , n1407 , n1396 );
nor ( n1885 , n1883 , n1884 );
xnor ( n1886 , n1885 , n1348 );
and ( n1887 , n1881 , n1886 );
and ( n1888 , n1877 , n1886 );
or ( n1889 , n1882 , n1887 , n1888 );
and ( n1890 , n1873 , n1889 );
xor ( n1891 , n1667 , n1789 );
xor ( n1892 , n1789 , n1790 );
not ( n1893 , n1892 );
and ( n1894 , n1891 , n1893 );
and ( n1895 , n1231 , n1894 );
not ( n1896 , n1895 );
xnor ( n1897 , n1896 , n1793 );
buf ( n1898 , n1897 );
and ( n1899 , n1889 , n1898 );
and ( n1900 , n1873 , n1898 );
or ( n1901 , n1890 , n1899 , n1900 );
xor ( n1902 , n1753 , n1757 );
xor ( n1903 , n1902 , n1760 );
and ( n1904 , n1901 , n1903 );
xor ( n1905 , n1806 , n1807 );
xor ( n1906 , n1905 , n1812 );
and ( n1907 , n1903 , n1906 );
and ( n1908 , n1901 , n1906 );
or ( n1909 , n1904 , n1907 , n1908 );
and ( n1910 , n1859 , n1909 );
xor ( n1911 , n1749 , n1763 );
xor ( n1912 , n1911 , n1766 );
and ( n1913 , n1909 , n1912 );
and ( n1914 , n1859 , n1912 );
or ( n1915 , n1910 , n1913 , n1914 );
and ( n1916 , n1823 , n1915 );
xor ( n1917 , n1769 , n1771 );
xor ( n1918 , n1917 , n1774 );
and ( n1919 , n1915 , n1918 );
and ( n1920 , n1823 , n1918 );
or ( n1921 , n1916 , n1919 , n1920 );
and ( n1922 , n1788 , n1921 );
xor ( n1923 , n1827 , n1831 );
xor ( n1924 , n1923 , n1834 );
xor ( n1925 , n1841 , n1845 );
xor ( n1926 , n1925 , n1850 );
and ( n1927 , n1924 , n1926 );
xor ( n1928 , n1794 , n1798 );
xor ( n1929 , n1928 , n1803 );
and ( n1930 , n1926 , n1929 );
and ( n1931 , n1924 , n1929 );
or ( n1932 , n1927 , n1930 , n1931 );
xor ( n1933 , n1837 , n1853 );
xor ( n1934 , n1933 , n1856 );
and ( n1935 , n1932 , n1934 );
xor ( n1936 , n1901 , n1903 );
xor ( n1937 , n1936 , n1906 );
and ( n1938 , n1934 , n1937 );
and ( n1939 , n1932 , n1937 );
or ( n1940 , n1935 , n1938 , n1939 );
xor ( n1941 , n1815 , n1817 );
xor ( n1942 , n1941 , n1820 );
and ( n1943 , n1940 , n1942 );
xor ( n1944 , n1859 , n1909 );
xor ( n1945 , n1944 , n1912 );
and ( n1946 , n1942 , n1945 );
and ( n1947 , n1940 , n1945 );
or ( n1948 , n1943 , n1946 , n1947 );
xor ( n1949 , n1823 , n1915 );
xor ( n1950 , n1949 , n1918 );
and ( n1951 , n1948 , n1950 );
xor ( n1952 , n1940 , n1942 );
xor ( n1953 , n1952 , n1945 );
and ( n1954 , n1274 , n1692 );
and ( n1955 , n1239 , n1690 );
nor ( n1956 , n1954 , n1955 );
xnor ( n1957 , n1956 , n1670 );
and ( n1958 , n1521 , n1398 );
and ( n1959 , n1438 , n1396 );
nor ( n1960 , n1958 , n1959 );
xnor ( n1961 , n1960 , n1348 );
and ( n1962 , n1957 , n1961 );
buf ( n1963 , n1168 );
and ( n1964 , n1963 , n1224 );
and ( n1965 , n1961 , n1964 );
and ( n1966 , n1957 , n1964 );
or ( n1967 , n1962 , n1965 , n1966 );
and ( n1968 , n1407 , n1488 );
and ( n1969 , n1390 , n1486 );
nor ( n1970 , n1968 , n1969 );
xnor ( n1971 , n1970 , n1456 );
and ( n1972 , n1759 , n1264 );
and ( n1973 , n1661 , n1262 );
nor ( n1974 , n1972 , n1973 );
xnor ( n1975 , n1974 , n1221 );
and ( n1976 , n1971 , n1975 );
and ( n1977 , n1869 , n1229 );
and ( n1978 , n1833 , n1227 );
nor ( n1979 , n1977 , n1978 );
xnor ( n1980 , n1979 , n1236 );
and ( n1981 , n1975 , n1980 );
and ( n1982 , n1971 , n1980 );
or ( n1983 , n1976 , n1981 , n1982 );
and ( n1984 , n1967 , n1983 );
buf ( n1985 , n1201 );
buf ( n1986 , n1202 );
and ( n1987 , n1985 , n1986 );
not ( n1988 , n1987 );
and ( n1989 , n1790 , n1988 );
not ( n1990 , n1989 );
and ( n1991 , n1223 , n1894 );
and ( n1992 , n1231 , n1892 );
nor ( n1993 , n1991 , n1992 );
xnor ( n1994 , n1993 , n1793 );
and ( n1995 , n1990 , n1994 );
and ( n1996 , n1314 , n1604 );
and ( n1997 , n1300 , n1602 );
nor ( n1998 , n1996 , n1997 );
xnor ( n1999 , n1998 , n1549 );
and ( n2000 , n1994 , n1999 );
and ( n2001 , n1990 , n1999 );
or ( n2002 , n1995 , n2000 , n2001 );
and ( n2003 , n1983 , n2002 );
and ( n2004 , n1967 , n2002 );
or ( n2005 , n1984 , n2003 , n2004 );
not ( n2006 , n1897 );
and ( n2007 , n1610 , n1322 );
and ( n2008 , n1521 , n1320 );
nor ( n2009 , n2007 , n2008 );
xnor ( n2010 , n2009 , n1293 );
and ( n2011 , n2006 , n2010 );
and ( n2012 , n1661 , n1264 );
and ( n2013 , n1624 , n1262 );
nor ( n2014 , n2012 , n2013 );
xnor ( n2015 , n2014 , n1221 );
and ( n2016 , n2010 , n2015 );
and ( n2017 , n2006 , n2015 );
or ( n2018 , n2011 , n2016 , n2017 );
and ( n2019 , n2005 , n2018 );
xor ( n2020 , n1873 , n1889 );
xor ( n2021 , n2020 , n1898 );
and ( n2022 , n2018 , n2021 );
and ( n2023 , n2005 , n2021 );
or ( n2024 , n2019 , n2022 , n2023 );
xor ( n2025 , n1863 , n1867 );
xor ( n2026 , n2025 , n1870 );
xor ( n2027 , n1877 , n1881 );
xor ( n2028 , n2027 , n1886 );
and ( n2029 , n2026 , n2028 );
xor ( n2030 , n2006 , n2010 );
xor ( n2031 , n2030 , n2015 );
and ( n2032 , n2028 , n2031 );
and ( n2033 , n2026 , n2031 );
or ( n2034 , n2029 , n2032 , n2033 );
and ( n2035 , n1390 , n1604 );
and ( n2036 , n1314 , n1602 );
nor ( n2037 , n2035 , n2036 );
xnor ( n2038 , n2037 , n1549 );
and ( n2039 , n1833 , n1264 );
and ( n2040 , n1759 , n1262 );
nor ( n2041 , n2039 , n2040 );
xnor ( n2042 , n2041 , n1221 );
and ( n2043 , n2038 , n2042 );
and ( n2044 , n1963 , n1229 );
and ( n2045 , n1869 , n1227 );
nor ( n2046 , n2044 , n2045 );
xnor ( n2047 , n2046 , n1236 );
and ( n2048 , n2042 , n2047 );
and ( n2049 , n2038 , n2047 );
or ( n2050 , n2043 , n2048 , n2049 );
xor ( n2051 , n1790 , n1985 );
xor ( n2052 , n1985 , n1986 );
not ( n2053 , n2052 );
and ( n2054 , n2051 , n2053 );
and ( n2055 , n1231 , n2054 );
not ( n2056 , n2055 );
xnor ( n2057 , n2056 , n1989 );
buf ( n2058 , n2057 );
and ( n2059 , n2050 , n2058 );
and ( n2060 , n1624 , n1322 );
and ( n2061 , n1610 , n1320 );
nor ( n2062 , n2060 , n2061 );
xnor ( n2063 , n2062 , n1293 );
and ( n2064 , n2058 , n2063 );
and ( n2065 , n2050 , n2063 );
or ( n2066 , n2059 , n2064 , n2065 );
and ( n2067 , n1239 , n1894 );
and ( n2068 , n1223 , n1892 );
nor ( n2069 , n2067 , n2068 );
xnor ( n2070 , n2069 , n1793 );
and ( n2071 , n1438 , n1488 );
and ( n2072 , n1407 , n1486 );
nor ( n2073 , n2071 , n2072 );
xnor ( n2074 , n2073 , n1456 );
and ( n2075 , n2070 , n2074 );
buf ( n2076 , n1169 );
and ( n2077 , n2076 , n1224 );
and ( n2078 , n2074 , n2077 );
and ( n2079 , n2070 , n2077 );
or ( n2080 , n2075 , n2078 , n2079 );
and ( n2081 , n1300 , n1692 );
and ( n2082 , n1274 , n1690 );
nor ( n2083 , n2081 , n2082 );
xnor ( n2084 , n2083 , n1670 );
and ( n2085 , n1610 , n1398 );
and ( n2086 , n1521 , n1396 );
nor ( n2087 , n2085 , n2086 );
xnor ( n2088 , n2087 , n1348 );
and ( n2089 , n2084 , n2088 );
and ( n2090 , n1661 , n1322 );
and ( n2091 , n1624 , n1320 );
nor ( n2092 , n2090 , n2091 );
xnor ( n2093 , n2092 , n1293 );
and ( n2094 , n2088 , n2093 );
and ( n2095 , n2084 , n2093 );
or ( n2096 , n2089 , n2094 , n2095 );
and ( n2097 , n2080 , n2096 );
xor ( n2098 , n1957 , n1961 );
xor ( n2099 , n2098 , n1964 );
and ( n2100 , n2096 , n2099 );
and ( n2101 , n2080 , n2099 );
or ( n2102 , n2097 , n2100 , n2101 );
and ( n2103 , n2066 , n2102 );
xor ( n2104 , n1967 , n1983 );
xor ( n2105 , n2104 , n2002 );
and ( n2106 , n2102 , n2105 );
and ( n2107 , n2066 , n2105 );
or ( n2108 , n2103 , n2106 , n2107 );
and ( n2109 , n2034 , n2108 );
xor ( n2110 , n1924 , n1926 );
xor ( n2111 , n2110 , n1929 );
and ( n2112 , n2108 , n2111 );
and ( n2113 , n2034 , n2111 );
or ( n2114 , n2109 , n2112 , n2113 );
and ( n2115 , n2024 , n2114 );
xor ( n2116 , n1932 , n1934 );
xor ( n2117 , n2116 , n1937 );
and ( n2118 , n2114 , n2117 );
and ( n2119 , n2024 , n2117 );
or ( n2120 , n2115 , n2118 , n2119 );
and ( n2121 , n1953 , n2120 );
xor ( n2122 , n2024 , n2114 );
xor ( n2123 , n2122 , n2117 );
xor ( n2124 , n1971 , n1975 );
xor ( n2125 , n2124 , n1980 );
xor ( n2126 , n1990 , n1994 );
xor ( n2127 , n2126 , n1999 );
and ( n2128 , n2125 , n2127 );
xor ( n2129 , n2050 , n2058 );
xor ( n2130 , n2129 , n2063 );
and ( n2131 , n2127 , n2130 );
and ( n2132 , n2125 , n2130 );
or ( n2133 , n2128 , n2131 , n2132 );
buf ( n2134 , n1203 );
buf ( n2135 , n1204 );
and ( n2136 , n2134 , n2135 );
not ( n2137 , n2136 );
and ( n2138 , n1986 , n2137 );
not ( n2139 , n2138 );
and ( n2140 , n1223 , n2054 );
and ( n2141 , n1231 , n2052 );
nor ( n2142 , n2140 , n2141 );
xnor ( n2143 , n2142 , n1989 );
and ( n2144 , n2139 , n2143 );
and ( n2145 , n1314 , n1692 );
and ( n2146 , n1300 , n1690 );
nor ( n2147 , n2145 , n2146 );
xnor ( n2148 , n2147 , n1670 );
and ( n2149 , n2143 , n2148 );
and ( n2150 , n2139 , n2148 );
or ( n2151 , n2144 , n2149 , n2150 );
and ( n2152 , n1407 , n1604 );
and ( n2153 , n1390 , n1602 );
nor ( n2154 , n2152 , n2153 );
xnor ( n2155 , n2154 , n1549 );
and ( n2156 , n1759 , n1322 );
and ( n2157 , n1661 , n1320 );
nor ( n2158 , n2156 , n2157 );
xnor ( n2159 , n2158 , n1293 );
and ( n2160 , n2155 , n2159 );
and ( n2161 , n1869 , n1264 );
and ( n2162 , n1833 , n1262 );
nor ( n2163 , n2161 , n2162 );
xnor ( n2164 , n2163 , n1221 );
and ( n2165 , n2159 , n2164 );
and ( n2166 , n2155 , n2164 );
or ( n2167 , n2160 , n2165 , n2166 );
and ( n2168 , n2151 , n2167 );
not ( n2169 , n2057 );
and ( n2170 , n2167 , n2169 );
and ( n2171 , n2151 , n2169 );
or ( n2172 , n2168 , n2170 , n2171 );
and ( n2173 , n1274 , n1894 );
and ( n2174 , n1239 , n1892 );
nor ( n2175 , n2173 , n2174 );
xnor ( n2176 , n2175 , n1793 );
and ( n2177 , n2076 , n1229 );
and ( n2178 , n1963 , n1227 );
nor ( n2179 , n2177 , n2178 );
xnor ( n2180 , n2179 , n1236 );
and ( n2181 , n2176 , n2180 );
buf ( n2182 , n1170 );
and ( n2183 , n2182 , n1224 );
and ( n2184 , n2180 , n2183 );
and ( n2185 , n2176 , n2183 );
or ( n2186 , n2181 , n2184 , n2185 );
xor ( n2187 , n2070 , n2074 );
xor ( n2188 , n2187 , n2077 );
and ( n2189 , n2186 , n2188 );
xor ( n2190 , n2038 , n2042 );
xor ( n2191 , n2190 , n2047 );
and ( n2192 , n2188 , n2191 );
and ( n2193 , n2186 , n2191 );
or ( n2194 , n2189 , n2192 , n2193 );
and ( n2195 , n2172 , n2194 );
xor ( n2196 , n2080 , n2096 );
xor ( n2197 , n2196 , n2099 );
and ( n2198 , n2194 , n2197 );
and ( n2199 , n2172 , n2197 );
or ( n2200 , n2195 , n2198 , n2199 );
and ( n2201 , n2133 , n2200 );
xor ( n2202 , n2026 , n2028 );
xor ( n2203 , n2202 , n2031 );
and ( n2204 , n2200 , n2203 );
and ( n2205 , n2133 , n2203 );
or ( n2206 , n2201 , n2204 , n2205 );
xor ( n2207 , n2005 , n2018 );
xor ( n2208 , n2207 , n2021 );
and ( n2209 , n2206 , n2208 );
xor ( n2210 , n2034 , n2108 );
xor ( n2211 , n2210 , n2111 );
and ( n2212 , n2208 , n2211 );
and ( n2213 , n2206 , n2211 );
or ( n2214 , n2209 , n2212 , n2213 );
and ( n2215 , n2123 , n2214 );
xor ( n2216 , n2206 , n2208 );
xor ( n2217 , n2216 , n2211 );
xor ( n2218 , n1986 , n2134 );
xor ( n2219 , n2134 , n2135 );
not ( n2220 , n2219 );
and ( n2221 , n2218 , n2220 );
and ( n2222 , n1231 , n2221 );
not ( n2223 , n2222 );
xnor ( n2224 , n2223 , n2138 );
and ( n2225 , n1300 , n1894 );
and ( n2226 , n1274 , n1892 );
nor ( n2227 , n2225 , n2226 );
xnor ( n2228 , n2227 , n1793 );
and ( n2229 , n2224 , n2228 );
and ( n2230 , n1610 , n1488 );
and ( n2231 , n1521 , n1486 );
nor ( n2232 , n2230 , n2231 );
xnor ( n2233 , n2232 , n1456 );
and ( n2234 , n2228 , n2233 );
and ( n2235 , n2224 , n2233 );
or ( n2236 , n2229 , n2234 , n2235 );
and ( n2237 , n1390 , n1692 );
and ( n2238 , n1314 , n1690 );
nor ( n2239 , n2237 , n2238 );
xnor ( n2240 , n2239 , n1670 );
and ( n2241 , n1833 , n1322 );
and ( n2242 , n1759 , n1320 );
nor ( n2243 , n2241 , n2242 );
xnor ( n2244 , n2243 , n1293 );
and ( n2245 , n2240 , n2244 );
and ( n2246 , n1963 , n1264 );
and ( n2247 , n1869 , n1262 );
nor ( n2248 , n2246 , n2247 );
xnor ( n2249 , n2248 , n1221 );
and ( n2250 , n2244 , n2249 );
and ( n2251 , n2240 , n2249 );
or ( n2252 , n2245 , n2250 , n2251 );
and ( n2253 , n2236 , n2252 );
and ( n2254 , n1438 , n1604 );
and ( n2255 , n1407 , n1602 );
nor ( n2256 , n2254 , n2255 );
xnor ( n2257 , n2256 , n1549 );
and ( n2258 , n2182 , n1229 );
and ( n2259 , n2076 , n1227 );
nor ( n2260 , n2258 , n2259 );
xnor ( n2261 , n2260 , n1236 );
and ( n2262 , n2257 , n2261 );
buf ( n2263 , n1171 );
and ( n2264 , n2263 , n1224 );
and ( n2265 , n2261 , n2264 );
and ( n2266 , n2257 , n2264 );
or ( n2267 , n2262 , n2265 , n2266 );
and ( n2268 , n2252 , n2267 );
and ( n2269 , n2236 , n2267 );
or ( n2270 , n2253 , n2268 , n2269 );
and ( n2271 , n1239 , n2054 );
and ( n2272 , n1223 , n2052 );
nor ( n2273 , n2271 , n2272 );
xnor ( n2274 , n2273 , n1989 );
buf ( n2275 , n2274 );
and ( n2276 , n1521 , n1488 );
and ( n2277 , n1438 , n1486 );
nor ( n2278 , n2276 , n2277 );
xnor ( n2279 , n2278 , n1456 );
and ( n2280 , n2275 , n2279 );
and ( n2281 , n1624 , n1398 );
and ( n2282 , n1610 , n1396 );
nor ( n2283 , n2281 , n2282 );
xnor ( n2284 , n2283 , n1348 );
and ( n2285 , n2279 , n2284 );
and ( n2286 , n2275 , n2284 );
or ( n2287 , n2280 , n2285 , n2286 );
and ( n2288 , n2270 , n2287 );
xor ( n2289 , n2084 , n2088 );
xor ( n2290 , n2289 , n2093 );
and ( n2291 , n2287 , n2290 );
and ( n2292 , n2270 , n2290 );
or ( n2293 , n2288 , n2291 , n2292 );
xor ( n2294 , n2176 , n2180 );
xor ( n2295 , n2294 , n2183 );
xor ( n2296 , n2139 , n2143 );
xor ( n2297 , n2296 , n2148 );
and ( n2298 , n2295 , n2297 );
xor ( n2299 , n2155 , n2159 );
xor ( n2300 , n2299 , n2164 );
and ( n2301 , n2297 , n2300 );
and ( n2302 , n2295 , n2300 );
or ( n2303 , n2298 , n2301 , n2302 );
xor ( n2304 , n2151 , n2167 );
xor ( n2305 , n2304 , n2169 );
and ( n2306 , n2303 , n2305 );
xor ( n2307 , n2186 , n2188 );
xor ( n2308 , n2307 , n2191 );
and ( n2309 , n2305 , n2308 );
and ( n2310 , n2303 , n2308 );
or ( n2311 , n2306 , n2309 , n2310 );
and ( n2312 , n2293 , n2311 );
xor ( n2313 , n2125 , n2127 );
xor ( n2314 , n2313 , n2130 );
and ( n2315 , n2311 , n2314 );
and ( n2316 , n2293 , n2314 );
or ( n2317 , n2312 , n2315 , n2316 );
xor ( n2318 , n2066 , n2102 );
xor ( n2319 , n2318 , n2105 );
and ( n2320 , n2317 , n2319 );
xor ( n2321 , n2133 , n2200 );
xor ( n2322 , n2321 , n2203 );
and ( n2323 , n2319 , n2322 );
and ( n2324 , n2317 , n2322 );
or ( n2325 , n2320 , n2323 , n2324 );
and ( n2326 , n2217 , n2325 );
xor ( n2327 , n2317 , n2319 );
xor ( n2328 , n2327 , n2322 );
and ( n2329 , n1521 , n1604 );
and ( n2330 , n1438 , n1602 );
nor ( n2331 , n2329 , n2330 );
xnor ( n2332 , n2331 , n1549 );
and ( n2333 , n1624 , n1488 );
and ( n2334 , n1610 , n1486 );
nor ( n2335 , n2333 , n2334 );
xnor ( n2336 , n2335 , n1456 );
and ( n2337 , n2332 , n2336 );
buf ( n2338 , n1172 );
and ( n2339 , n2338 , n1224 );
and ( n2340 , n2336 , n2339 );
and ( n2341 , n2332 , n2339 );
or ( n2342 , n2337 , n2340 , n2341 );
and ( n2343 , n1407 , n1692 );
and ( n2344 , n1390 , n1690 );
nor ( n2345 , n2343 , n2344 );
xnor ( n2346 , n2345 , n1670 );
and ( n2347 , n1759 , n1398 );
and ( n2348 , n1661 , n1396 );
nor ( n2349 , n2347 , n2348 );
xnor ( n2350 , n2349 , n1348 );
and ( n2351 , n2346 , n2350 );
and ( n2352 , n1869 , n1322 );
and ( n2353 , n1833 , n1320 );
nor ( n2354 , n2352 , n2353 );
xnor ( n2355 , n2354 , n1293 );
and ( n2356 , n2350 , n2355 );
and ( n2357 , n2346 , n2355 );
or ( n2358 , n2351 , n2356 , n2357 );
and ( n2359 , n2342 , n2358 );
buf ( n2360 , n1205 );
buf ( n2361 , n1206 );
and ( n2362 , n2360 , n2361 );
not ( n2363 , n2362 );
and ( n2364 , n2135 , n2363 );
not ( n2365 , n2364 );
and ( n2366 , n1223 , n2221 );
and ( n2367 , n1231 , n2219 );
nor ( n2368 , n2366 , n2367 );
xnor ( n2369 , n2368 , n2138 );
and ( n2370 , n2365 , n2369 );
and ( n2371 , n1314 , n1894 );
and ( n2372 , n1300 , n1892 );
nor ( n2373 , n2371 , n2372 );
xnor ( n2374 , n2373 , n1793 );
and ( n2375 , n2369 , n2374 );
and ( n2376 , n2365 , n2374 );
or ( n2377 , n2370 , n2375 , n2376 );
and ( n2378 , n2358 , n2377 );
and ( n2379 , n2342 , n2377 );
or ( n2380 , n2359 , n2378 , n2379 );
and ( n2381 , n1274 , n2054 );
and ( n2382 , n1239 , n2052 );
nor ( n2383 , n2381 , n2382 );
xnor ( n2384 , n2383 , n1989 );
and ( n2385 , n2076 , n1264 );
and ( n2386 , n1963 , n1262 );
nor ( n2387 , n2385 , n2386 );
xnor ( n2388 , n2387 , n1221 );
and ( n2389 , n2384 , n2388 );
and ( n2390 , n2263 , n1229 );
and ( n2391 , n2182 , n1227 );
nor ( n2392 , n2390 , n2391 );
xnor ( n2393 , n2392 , n1236 );
and ( n2394 , n2388 , n2393 );
and ( n2395 , n2384 , n2393 );
or ( n2396 , n2389 , n2394 , n2395 );
not ( n2397 , n2274 );
and ( n2398 , n2396 , n2397 );
and ( n2399 , n1661 , n1398 );
and ( n2400 , n1624 , n1396 );
nor ( n2401 , n2399 , n2400 );
xnor ( n2402 , n2401 , n1348 );
and ( n2403 , n2397 , n2402 );
and ( n2404 , n2396 , n2402 );
or ( n2405 , n2398 , n2403 , n2404 );
and ( n2406 , n2380 , n2405 );
xor ( n2407 , n2275 , n2279 );
xor ( n2408 , n2407 , n2284 );
and ( n2409 , n2405 , n2408 );
and ( n2410 , n2380 , n2408 );
or ( n2411 , n2406 , n2409 , n2410 );
xor ( n2412 , n2224 , n2228 );
xor ( n2413 , n2412 , n2233 );
xor ( n2414 , n2240 , n2244 );
xor ( n2415 , n2414 , n2249 );
and ( n2416 , n2413 , n2415 );
xor ( n2417 , n2257 , n2261 );
xor ( n2418 , n2417 , n2264 );
and ( n2419 , n2415 , n2418 );
and ( n2420 , n2413 , n2418 );
or ( n2421 , n2416 , n2419 , n2420 );
xor ( n2422 , n2236 , n2252 );
xor ( n2423 , n2422 , n2267 );
and ( n2424 , n2421 , n2423 );
xor ( n2425 , n2295 , n2297 );
xor ( n2426 , n2425 , n2300 );
and ( n2427 , n2423 , n2426 );
and ( n2428 , n2421 , n2426 );
or ( n2429 , n2424 , n2427 , n2428 );
and ( n2430 , n2411 , n2429 );
xor ( n2431 , n2270 , n2287 );
xor ( n2432 , n2431 , n2290 );
and ( n2433 , n2429 , n2432 );
and ( n2434 , n2411 , n2432 );
or ( n2435 , n2430 , n2433 , n2434 );
xor ( n2436 , n2172 , n2194 );
xor ( n2437 , n2436 , n2197 );
and ( n2438 , n2435 , n2437 );
xor ( n2439 , n2293 , n2311 );
xor ( n2440 , n2439 , n2314 );
and ( n2441 , n2437 , n2440 );
and ( n2442 , n2435 , n2440 );
or ( n2443 , n2438 , n2441 , n2442 );
and ( n2444 , n2328 , n2443 );
xor ( n2445 , n2435 , n2437 );
xor ( n2446 , n2445 , n2440 );
xor ( n2447 , n2135 , n2360 );
xor ( n2448 , n2360 , n2361 );
not ( n2449 , n2448 );
and ( n2450 , n2447 , n2449 );
and ( n2451 , n1231 , n2450 );
not ( n2452 , n2451 );
xnor ( n2453 , n2452 , n2364 );
and ( n2454 , n1300 , n2054 );
and ( n2455 , n1274 , n2052 );
nor ( n2456 , n2454 , n2455 );
xnor ( n2457 , n2456 , n1989 );
and ( n2458 , n2453 , n2457 );
buf ( n2459 , n1173 );
and ( n2460 , n2459 , n1224 );
and ( n2461 , n2457 , n2460 );
and ( n2462 , n2453 , n2460 );
or ( n2463 , n2458 , n2461 , n2462 );
and ( n2464 , n1390 , n1894 );
and ( n2465 , n1314 , n1892 );
nor ( n2466 , n2464 , n2465 );
xnor ( n2467 , n2466 , n1793 );
and ( n2468 , n1833 , n1398 );
and ( n2469 , n1759 , n1396 );
nor ( n2470 , n2468 , n2469 );
xnor ( n2471 , n2470 , n1348 );
and ( n2472 , n2467 , n2471 );
and ( n2473 , n1963 , n1322 );
and ( n2474 , n1869 , n1320 );
nor ( n2475 , n2473 , n2474 );
xnor ( n2476 , n2475 , n1293 );
and ( n2477 , n2471 , n2476 );
and ( n2478 , n2467 , n2476 );
or ( n2479 , n2472 , n2477 , n2478 );
and ( n2480 , n2463 , n2479 );
and ( n2481 , n1239 , n2221 );
and ( n2482 , n1223 , n2219 );
nor ( n2483 , n2481 , n2482 );
xnor ( n2484 , n2483 , n2138 );
buf ( n2485 , n2484 );
and ( n2486 , n2479 , n2485 );
and ( n2487 , n2463 , n2485 );
or ( n2488 , n2480 , n2486 , n2487 );
xor ( n2489 , n2342 , n2358 );
xor ( n2490 , n2489 , n2377 );
and ( n2491 , n2488 , n2490 );
xor ( n2492 , n2396 , n2397 );
xor ( n2493 , n2492 , n2402 );
and ( n2494 , n2490 , n2493 );
and ( n2495 , n2488 , n2493 );
or ( n2496 , n2491 , n2494 , n2495 );
xor ( n2497 , n2380 , n2405 );
xor ( n2498 , n2497 , n2408 );
and ( n2499 , n2496 , n2498 );
xor ( n2500 , n2421 , n2423 );
xor ( n2501 , n2500 , n2426 );
and ( n2502 , n2498 , n2501 );
and ( n2503 , n2496 , n2501 );
or ( n2504 , n2499 , n2502 , n2503 );
xor ( n2505 , n2303 , n2305 );
xor ( n2506 , n2505 , n2308 );
and ( n2507 , n2504 , n2506 );
xor ( n2508 , n2411 , n2429 );
xor ( n2509 , n2508 , n2432 );
and ( n2510 , n2506 , n2509 );
and ( n2511 , n2504 , n2509 );
or ( n2512 , n2507 , n2510 , n2511 );
and ( n2513 , n2446 , n2512 );
xor ( n2514 , n2504 , n2506 );
xor ( n2515 , n2514 , n2509 );
not ( n2516 , n2484 );
and ( n2517 , n1610 , n1604 );
and ( n2518 , n1521 , n1602 );
nor ( n2519 , n2517 , n2518 );
xnor ( n2520 , n2519 , n1549 );
and ( n2521 , n2516 , n2520 );
and ( n2522 , n1661 , n1488 );
and ( n2523 , n1624 , n1486 );
nor ( n2524 , n2522 , n2523 );
xnor ( n2525 , n2524 , n1456 );
and ( n2526 , n2520 , n2525 );
and ( n2527 , n2516 , n2525 );
or ( n2528 , n2521 , n2526 , n2527 );
xor ( n2529 , n2346 , n2350 );
xor ( n2530 , n2529 , n2355 );
and ( n2531 , n2528 , n2530 );
xor ( n2532 , n2365 , n2369 );
xor ( n2533 , n2532 , n2374 );
and ( n2534 , n2530 , n2533 );
and ( n2535 , n2528 , n2533 );
or ( n2536 , n2531 , n2534 , n2535 );
and ( n2537 , n1438 , n1692 );
and ( n2538 , n1407 , n1690 );
nor ( n2539 , n2537 , n2538 );
xnor ( n2540 , n2539 , n1670 );
and ( n2541 , n2182 , n1264 );
and ( n2542 , n2076 , n1262 );
nor ( n2543 , n2541 , n2542 );
xnor ( n2544 , n2543 , n1221 );
and ( n2545 , n2540 , n2544 );
and ( n2546 , n2338 , n1229 );
and ( n2547 , n2263 , n1227 );
nor ( n2548 , n2546 , n2547 );
xnor ( n2549 , n2548 , n1236 );
and ( n2550 , n2544 , n2549 );
and ( n2551 , n2540 , n2549 );
or ( n2552 , n2545 , n2550 , n2551 );
xor ( n2553 , n2332 , n2336 );
xor ( n2554 , n2553 , n2339 );
and ( n2555 , n2552 , n2554 );
xor ( n2556 , n2384 , n2388 );
xor ( n2557 , n2556 , n2393 );
and ( n2558 , n2554 , n2557 );
and ( n2559 , n2552 , n2557 );
or ( n2560 , n2555 , n2558 , n2559 );
and ( n2561 , n2536 , n2560 );
xor ( n2562 , n2413 , n2415 );
xor ( n2563 , n2562 , n2418 );
and ( n2564 , n2560 , n2563 );
and ( n2565 , n2536 , n2563 );
or ( n2566 , n2561 , n2564 , n2565 );
and ( n2567 , n1274 , n2221 );
and ( n2568 , n1239 , n2219 );
nor ( n2569 , n2567 , n2568 );
xnor ( n2570 , n2569 , n2138 );
and ( n2571 , n2076 , n1322 );
and ( n2572 , n1963 , n1320 );
nor ( n2573 , n2571 , n2572 );
xnor ( n2574 , n2573 , n1293 );
and ( n2575 , n2570 , n2574 );
and ( n2576 , n2263 , n1264 );
and ( n2577 , n2182 , n1262 );
nor ( n2578 , n2576 , n2577 );
xnor ( n2579 , n2578 , n1221 );
and ( n2580 , n2574 , n2579 );
and ( n2581 , n2570 , n2579 );
or ( n2582 , n2575 , n2580 , n2581 );
buf ( n2583 , n1207 );
buf ( n2584 , n1208 );
and ( n2585 , n2583 , n2584 );
not ( n2586 , n2585 );
and ( n2587 , n2361 , n2586 );
not ( n2588 , n2587 );
and ( n2589 , n1223 , n2450 );
and ( n2590 , n1231 , n2448 );
nor ( n2591 , n2589 , n2590 );
xnor ( n2592 , n2591 , n2364 );
and ( n2593 , n2588 , n2592 );
and ( n2594 , n1314 , n2054 );
and ( n2595 , n1300 , n2052 );
nor ( n2596 , n2594 , n2595 );
xnor ( n2597 , n2596 , n1989 );
and ( n2598 , n2592 , n2597 );
and ( n2599 , n2588 , n2597 );
or ( n2600 , n2593 , n2598 , n2599 );
and ( n2601 , n2582 , n2600 );
and ( n2602 , n1521 , n1692 );
and ( n2603 , n1438 , n1690 );
nor ( n2604 , n2602 , n2603 );
xnor ( n2605 , n2604 , n1670 );
and ( n2606 , n2459 , n1229 );
and ( n2607 , n2338 , n1227 );
nor ( n2608 , n2606 , n2607 );
xnor ( n2609 , n2608 , n1236 );
and ( n2610 , n2605 , n2609 );
buf ( n2611 , n1174 );
and ( n2612 , n2611 , n1224 );
and ( n2613 , n2609 , n2612 );
and ( n2614 , n2605 , n2612 );
or ( n2615 , n2610 , n2613 , n2614 );
and ( n2616 , n2600 , n2615 );
and ( n2617 , n2582 , n2615 );
or ( n2618 , n2601 , n2616 , n2617 );
and ( n2619 , n1407 , n1894 );
and ( n2620 , n1390 , n1892 );
nor ( n2621 , n2619 , n2620 );
xnor ( n2622 , n2621 , n1793 );
and ( n2623 , n1759 , n1488 );
and ( n2624 , n1661 , n1486 );
nor ( n2625 , n2623 , n2624 );
xnor ( n2626 , n2625 , n1456 );
and ( n2627 , n2622 , n2626 );
and ( n2628 , n1869 , n1398 );
and ( n2629 , n1833 , n1396 );
nor ( n2630 , n2628 , n2629 );
xnor ( n2631 , n2630 , n1348 );
and ( n2632 , n2626 , n2631 );
and ( n2633 , n2622 , n2631 );
or ( n2634 , n2627 , n2632 , n2633 );
xor ( n2635 , n2453 , n2457 );
xor ( n2636 , n2635 , n2460 );
and ( n2637 , n2634 , n2636 );
xor ( n2638 , n2467 , n2471 );
xor ( n2639 , n2638 , n2476 );
and ( n2640 , n2636 , n2639 );
and ( n2641 , n2634 , n2639 );
or ( n2642 , n2637 , n2640 , n2641 );
and ( n2643 , n2618 , n2642 );
xor ( n2644 , n2463 , n2479 );
xor ( n2645 , n2644 , n2485 );
and ( n2646 , n2642 , n2645 );
and ( n2647 , n2618 , n2645 );
or ( n2648 , n2643 , n2646 , n2647 );
and ( n2649 , n1300 , n2221 );
and ( n2650 , n1274 , n2219 );
nor ( n2651 , n2649 , n2650 );
xnor ( n2652 , n2651 , n2138 );
and ( n2653 , n1661 , n1604 );
and ( n2654 , n1624 , n1602 );
nor ( n2655 , n2653 , n2654 );
xnor ( n2656 , n2655 , n1549 );
and ( n2657 , n2652 , n2656 );
buf ( n2658 , n1175 );
and ( n2659 , n2658 , n1224 );
and ( n2660 , n2656 , n2659 );
and ( n2661 , n2652 , n2659 );
or ( n2662 , n2657 , n2660 , n2661 );
xor ( n2663 , n2361 , n2583 );
xor ( n2664 , n2583 , n2584 );
not ( n2665 , n2664 );
and ( n2666 , n2663 , n2665 );
and ( n2667 , n1231 , n2666 );
not ( n2668 , n2667 );
xnor ( n2669 , n2668 , n2587 );
and ( n2670 , n1610 , n1692 );
and ( n2671 , n1521 , n1690 );
nor ( n2672 , n2670 , n2671 );
xnor ( n2673 , n2672 , n1670 );
and ( n2674 , n2669 , n2673 );
and ( n2675 , n2611 , n1229 );
and ( n2676 , n2459 , n1227 );
nor ( n2677 , n2675 , n2676 );
xnor ( n2678 , n2677 , n1236 );
and ( n2679 , n2673 , n2678 );
and ( n2680 , n2669 , n2678 );
or ( n2681 , n2674 , n2679 , n2680 );
and ( n2682 , n2662 , n2681 );
and ( n2683 , n1390 , n2054 );
and ( n2684 , n1314 , n2052 );
nor ( n2685 , n2683 , n2684 );
xnor ( n2686 , n2685 , n1989 );
and ( n2687 , n1833 , n1488 );
and ( n2688 , n1759 , n1486 );
nor ( n2689 , n2687 , n2688 );
xnor ( n2690 , n2689 , n1456 );
and ( n2691 , n2686 , n2690 );
and ( n2692 , n1963 , n1398 );
and ( n2693 , n1869 , n1396 );
nor ( n2694 , n2692 , n2693 );
xnor ( n2695 , n2694 , n1348 );
and ( n2696 , n2690 , n2695 );
and ( n2697 , n2686 , n2695 );
or ( n2698 , n2691 , n2696 , n2697 );
and ( n2699 , n2681 , n2698 );
and ( n2700 , n2662 , n2698 );
or ( n2701 , n2682 , n2699 , n2700 );
xor ( n2702 , n2540 , n2544 );
xor ( n2703 , n2702 , n2549 );
and ( n2704 , n2701 , n2703 );
xor ( n2705 , n2516 , n2520 );
xor ( n2706 , n2705 , n2525 );
and ( n2707 , n2703 , n2706 );
and ( n2708 , n2701 , n2706 );
or ( n2709 , n2704 , n2707 , n2708 );
xor ( n2710 , n2528 , n2530 );
xor ( n2711 , n2710 , n2533 );
and ( n2712 , n2709 , n2711 );
xor ( n2713 , n2552 , n2554 );
xor ( n2714 , n2713 , n2557 );
and ( n2715 , n2711 , n2714 );
and ( n2716 , n2709 , n2714 );
or ( n2717 , n2712 , n2715 , n2716 );
and ( n2718 , n2648 , n2717 );
xor ( n2719 , n2488 , n2490 );
xor ( n2720 , n2719 , n2493 );
and ( n2721 , n2717 , n2720 );
and ( n2722 , n2648 , n2720 );
or ( n2723 , n2718 , n2721 , n2722 );
and ( n2724 , n2566 , n2723 );
xor ( n2725 , n2496 , n2498 );
xor ( n2726 , n2725 , n2501 );
and ( n2727 , n2723 , n2726 );
and ( n2728 , n2566 , n2726 );
or ( n2729 , n2724 , n2727 , n2728 );
and ( n2730 , n2515 , n2729 );
xor ( n2731 , n2566 , n2723 );
xor ( n2732 , n2731 , n2726 );
and ( n2733 , n1438 , n1894 );
and ( n2734 , n1407 , n1892 );
nor ( n2735 , n2733 , n2734 );
xnor ( n2736 , n2735 , n1793 );
and ( n2737 , n2182 , n1322 );
and ( n2738 , n2076 , n1320 );
nor ( n2739 , n2737 , n2738 );
xnor ( n2740 , n2739 , n1293 );
and ( n2741 , n2736 , n2740 );
and ( n2742 , n2338 , n1264 );
and ( n2743 , n2263 , n1262 );
nor ( n2744 , n2742 , n2743 );
xnor ( n2745 , n2744 , n1221 );
and ( n2746 , n2740 , n2745 );
and ( n2747 , n2736 , n2745 );
or ( n2748 , n2741 , n2746 , n2747 );
and ( n2749 , n1239 , n2450 );
and ( n2750 , n1223 , n2448 );
nor ( n2751 , n2749 , n2750 );
xnor ( n2752 , n2751 , n2364 );
buf ( n2753 , n2752 );
and ( n2754 , n2748 , n2753 );
and ( n2755 , n1624 , n1604 );
and ( n2756 , n1610 , n1602 );
nor ( n2757 , n2755 , n2756 );
xnor ( n2758 , n2757 , n1549 );
and ( n2759 , n2753 , n2758 );
and ( n2760 , n2748 , n2758 );
or ( n2761 , n2754 , n2759 , n2760 );
xor ( n2762 , n2570 , n2574 );
xor ( n2763 , n2762 , n2579 );
xor ( n2764 , n2622 , n2626 );
xor ( n2765 , n2764 , n2631 );
and ( n2766 , n2763 , n2765 );
xor ( n2767 , n2588 , n2592 );
xor ( n2768 , n2767 , n2597 );
and ( n2769 , n2765 , n2768 );
and ( n2770 , n2763 , n2768 );
or ( n2771 , n2766 , n2769 , n2770 );
and ( n2772 , n2761 , n2771 );
xor ( n2773 , n2582 , n2600 );
xor ( n2774 , n2773 , n2615 );
and ( n2775 , n2771 , n2774 );
and ( n2776 , n2761 , n2774 );
or ( n2777 , n2772 , n2775 , n2776 );
and ( n2778 , n1274 , n2450 );
and ( n2779 , n1239 , n2448 );
nor ( n2780 , n2778 , n2779 );
xnor ( n2781 , n2780 , n2364 );
and ( n2782 , n2076 , n1398 );
and ( n2783 , n1963 , n1396 );
nor ( n2784 , n2782 , n2783 );
xnor ( n2785 , n2784 , n1348 );
and ( n2786 , n2781 , n2785 );
and ( n2787 , n2263 , n1322 );
and ( n2788 , n2182 , n1320 );
nor ( n2789 , n2787 , n2788 );
xnor ( n2790 , n2789 , n1293 );
and ( n2791 , n2785 , n2790 );
and ( n2792 , n2781 , n2790 );
or ( n2793 , n2786 , n2791 , n2792 );
and ( n2794 , n1407 , n2054 );
and ( n2795 , n1390 , n2052 );
nor ( n2796 , n2794 , n2795 );
xnor ( n2797 , n2796 , n1989 );
and ( n2798 , n1759 , n1604 );
and ( n2799 , n1661 , n1602 );
nor ( n2800 , n2798 , n2799 );
xnor ( n2801 , n2800 , n1549 );
and ( n2802 , n2797 , n2801 );
and ( n2803 , n1869 , n1488 );
and ( n2804 , n1833 , n1486 );
nor ( n2805 , n2803 , n2804 );
xnor ( n2806 , n2805 , n1456 );
and ( n2807 , n2801 , n2806 );
and ( n2808 , n2797 , n2806 );
or ( n2809 , n2802 , n2807 , n2808 );
and ( n2810 , n2793 , n2809 );
not ( n2811 , n2752 );
and ( n2812 , n2809 , n2811 );
and ( n2813 , n2793 , n2811 );
or ( n2814 , n2810 , n2812 , n2813 );
xor ( n2815 , n2605 , n2609 );
xor ( n2816 , n2815 , n2612 );
and ( n2817 , n2814 , n2816 );
xor ( n2818 , n2748 , n2753 );
xor ( n2819 , n2818 , n2758 );
and ( n2820 , n2816 , n2819 );
and ( n2821 , n2814 , n2819 );
or ( n2822 , n2817 , n2820 , n2821 );
xor ( n2823 , n2634 , n2636 );
xor ( n2824 , n2823 , n2639 );
and ( n2825 , n2822 , n2824 );
xor ( n2826 , n2701 , n2703 );
xor ( n2827 , n2826 , n2706 );
and ( n2828 , n2824 , n2827 );
and ( n2829 , n2822 , n2827 );
or ( n2830 , n2825 , n2828 , n2829 );
and ( n2831 , n2777 , n2830 );
xor ( n2832 , n2618 , n2642 );
xor ( n2833 , n2832 , n2645 );
and ( n2834 , n2830 , n2833 );
and ( n2835 , n2777 , n2833 );
or ( n2836 , n2831 , n2834 , n2835 );
xor ( n2837 , n2536 , n2560 );
xor ( n2838 , n2837 , n2563 );
and ( n2839 , n2836 , n2838 );
xor ( n2840 , n2648 , n2717 );
xor ( n2841 , n2840 , n2720 );
and ( n2842 , n2838 , n2841 );
and ( n2843 , n2836 , n2841 );
or ( n2844 , n2839 , n2842 , n2843 );
and ( n2845 , n2732 , n2844 );
xor ( n2846 , n2836 , n2838 );
xor ( n2847 , n2846 , n2841 );
and ( n2848 , n1521 , n1894 );
and ( n2849 , n1438 , n1892 );
nor ( n2850 , n2848 , n2849 );
xnor ( n2851 , n2850 , n1793 );
and ( n2852 , n2459 , n1264 );
and ( n2853 , n2338 , n1262 );
nor ( n2854 , n2852 , n2853 );
xnor ( n2855 , n2854 , n1221 );
and ( n2856 , n2851 , n2855 );
and ( n2857 , n2658 , n1229 );
and ( n2858 , n2611 , n1227 );
nor ( n2859 , n2857 , n2858 );
xnor ( n2860 , n2859 , n1236 );
and ( n2861 , n2855 , n2860 );
and ( n2862 , n2851 , n2860 );
or ( n2863 , n2856 , n2861 , n2862 );
buf ( n2864 , n1209 );
buf ( n2865 , n1210 );
and ( n2866 , n2864 , n2865 );
not ( n2867 , n2866 );
and ( n2868 , n2584 , n2867 );
not ( n2869 , n2868 );
and ( n2870 , n1223 , n2666 );
and ( n2871 , n1231 , n2664 );
nor ( n2872 , n2870 , n2871 );
xnor ( n2873 , n2872 , n2587 );
and ( n2874 , n2869 , n2873 );
and ( n2875 , n1314 , n2221 );
and ( n2876 , n1300 , n2219 );
nor ( n2877 , n2875 , n2876 );
xnor ( n2878 , n2877 , n2138 );
and ( n2879 , n2873 , n2878 );
and ( n2880 , n2869 , n2878 );
or ( n2881 , n2874 , n2879 , n2880 );
and ( n2882 , n2863 , n2881 );
xor ( n2883 , n2652 , n2656 );
xor ( n2884 , n2883 , n2659 );
and ( n2885 , n2881 , n2884 );
and ( n2886 , n2863 , n2884 );
or ( n2887 , n2882 , n2885 , n2886 );
xor ( n2888 , n2669 , n2673 );
xor ( n2889 , n2888 , n2678 );
xor ( n2890 , n2736 , n2740 );
xor ( n2891 , n2890 , n2745 );
and ( n2892 , n2889 , n2891 );
xor ( n2893 , n2686 , n2690 );
xor ( n2894 , n2893 , n2695 );
and ( n2895 , n2891 , n2894 );
and ( n2896 , n2889 , n2894 );
or ( n2897 , n2892 , n2895 , n2896 );
and ( n2898 , n2887 , n2897 );
xor ( n2899 , n2662 , n2681 );
xor ( n2900 , n2899 , n2698 );
and ( n2901 , n2897 , n2900 );
and ( n2902 , n2887 , n2900 );
or ( n2903 , n2898 , n2901 , n2902 );
and ( n2904 , n1390 , n2221 );
and ( n2905 , n1314 , n2219 );
nor ( n2906 , n2904 , n2905 );
xnor ( n2907 , n2906 , n2138 );
and ( n2908 , n1833 , n1604 );
and ( n2909 , n1759 , n1602 );
nor ( n2910 , n2908 , n2909 );
xnor ( n2911 , n2910 , n1549 );
and ( n2912 , n2907 , n2911 );
and ( n2913 , n1963 , n1488 );
and ( n2914 , n1869 , n1486 );
nor ( n2915 , n2913 , n2914 );
xnor ( n2916 , n2915 , n1456 );
and ( n2917 , n2911 , n2916 );
and ( n2918 , n2907 , n2916 );
or ( n2919 , n2912 , n2917 , n2918 );
and ( n2920 , n1438 , n2054 );
and ( n2921 , n1407 , n2052 );
nor ( n2922 , n2920 , n2921 );
xnor ( n2923 , n2922 , n1989 );
and ( n2924 , n2182 , n1398 );
and ( n2925 , n2076 , n1396 );
nor ( n2926 , n2924 , n2925 );
xnor ( n2927 , n2926 , n1348 );
and ( n2928 , n2923 , n2927 );
and ( n2929 , n2338 , n1322 );
and ( n2930 , n2263 , n1320 );
nor ( n2931 , n2929 , n2930 );
xnor ( n2932 , n2931 , n1293 );
and ( n2933 , n2927 , n2932 );
and ( n2934 , n2923 , n2932 );
or ( n2935 , n2928 , n2933 , n2934 );
and ( n2936 , n2919 , n2935 );
xor ( n2937 , n2584 , n2864 );
xor ( n2938 , n2864 , n2865 );
not ( n2939 , n2938 );
and ( n2940 , n2937 , n2939 );
and ( n2941 , n1231 , n2940 );
not ( n2942 , n2941 );
xnor ( n2943 , n2942 , n2868 );
and ( n2944 , n1610 , n1894 );
and ( n2945 , n1521 , n1892 );
nor ( n2946 , n2944 , n2945 );
xnor ( n2947 , n2946 , n1793 );
and ( n2948 , n2943 , n2947 );
and ( n2949 , n2611 , n1264 );
and ( n2950 , n2459 , n1262 );
nor ( n2951 , n2949 , n2950 );
xnor ( n2952 , n2951 , n1221 );
and ( n2953 , n2947 , n2952 );
and ( n2954 , n2943 , n2952 );
or ( n2955 , n2948 , n2953 , n2954 );
and ( n2956 , n2935 , n2955 );
and ( n2957 , n2919 , n2955 );
or ( n2958 , n2936 , n2956 , n2957 );
and ( n2959 , n1239 , n2666 );
and ( n2960 , n1223 , n2664 );
nor ( n2961 , n2959 , n2960 );
xnor ( n2962 , n2961 , n2587 );
buf ( n2963 , n2962 );
and ( n2964 , n1624 , n1692 );
and ( n2965 , n1610 , n1690 );
nor ( n2966 , n2964 , n2965 );
xnor ( n2967 , n2966 , n1670 );
and ( n2968 , n2963 , n2967 );
buf ( n2969 , n1176 );
and ( n2970 , n2969 , n1224 );
and ( n2971 , n2967 , n2970 );
and ( n2972 , n2963 , n2970 );
or ( n2973 , n2968 , n2971 , n2972 );
and ( n2974 , n2958 , n2973 );
xor ( n2975 , n2793 , n2809 );
xor ( n2976 , n2975 , n2811 );
and ( n2977 , n2973 , n2976 );
and ( n2978 , n2958 , n2976 );
or ( n2979 , n2974 , n2977 , n2978 );
xor ( n2980 , n2763 , n2765 );
xor ( n2981 , n2980 , n2768 );
and ( n2982 , n2979 , n2981 );
xor ( n2983 , n2814 , n2816 );
xor ( n2984 , n2983 , n2819 );
and ( n2985 , n2981 , n2984 );
and ( n2986 , n2979 , n2984 );
or ( n2987 , n2982 , n2985 , n2986 );
and ( n2988 , n2903 , n2987 );
xor ( n2989 , n2761 , n2771 );
xor ( n2990 , n2989 , n2774 );
and ( n2991 , n2987 , n2990 );
and ( n2992 , n2903 , n2990 );
or ( n2993 , n2988 , n2991 , n2992 );
xor ( n2994 , n2709 , n2711 );
xor ( n2995 , n2994 , n2714 );
and ( n2996 , n2993 , n2995 );
xor ( n2997 , n2777 , n2830 );
xor ( n2998 , n2997 , n2833 );
and ( n2999 , n2995 , n2998 );
and ( n3000 , n2993 , n2998 );
or ( n3001 , n2996 , n2999 , n3000 );
and ( n3002 , n2847 , n3001 );
xor ( n3003 , n2993 , n2995 );
xor ( n3004 , n3003 , n2998 );
xor ( n3005 , n2822 , n2824 );
xor ( n3006 , n3005 , n2827 );
xor ( n3007 , n2903 , n2987 );
xor ( n3008 , n3007 , n2990 );
and ( n3009 , n3006 , n3008 );
and ( n3010 , n1300 , n2450 );
and ( n3011 , n1274 , n2448 );
nor ( n3012 , n3010 , n3011 );
xnor ( n3013 , n3012 , n2364 );
and ( n3014 , n2969 , n1229 );
and ( n3015 , n2658 , n1227 );
nor ( n3016 , n3014 , n3015 );
xnor ( n3017 , n3016 , n1236 );
and ( n3018 , n3013 , n3017 );
buf ( n3019 , n1177 );
and ( n3020 , n3019 , n1224 );
and ( n3021 , n3017 , n3020 );
and ( n3022 , n3013 , n3020 );
or ( n3023 , n3018 , n3021 , n3022 );
xor ( n3024 , n2797 , n2801 );
xor ( n3025 , n3024 , n2806 );
and ( n3026 , n3023 , n3025 );
xor ( n3027 , n2869 , n2873 );
xor ( n3028 , n3027 , n2878 );
and ( n3029 , n3025 , n3028 );
and ( n3030 , n3023 , n3028 );
or ( n3031 , n3026 , n3029 , n3030 );
xor ( n3032 , n2851 , n2855 );
xor ( n3033 , n3032 , n2860 );
xor ( n3034 , n2781 , n2785 );
xor ( n3035 , n3034 , n2790 );
and ( n3036 , n3033 , n3035 );
xor ( n3037 , n2963 , n2967 );
xor ( n3038 , n3037 , n2970 );
and ( n3039 , n3035 , n3038 );
and ( n3040 , n3033 , n3038 );
or ( n3041 , n3036 , n3039 , n3040 );
and ( n3042 , n3031 , n3041 );
xor ( n3043 , n2863 , n2881 );
xor ( n3044 , n3043 , n2884 );
and ( n3045 , n3041 , n3044 );
and ( n3046 , n3031 , n3044 );
or ( n3047 , n3042 , n3045 , n3046 );
xor ( n3048 , n2887 , n2897 );
xor ( n3049 , n3048 , n2900 );
and ( n3050 , n3047 , n3049 );
and ( n3051 , n3008 , n3050 );
and ( n3052 , n3006 , n3050 );
or ( n3053 , n3009 , n3051 , n3052 );
and ( n3054 , n3004 , n3053 );
xor ( n3055 , n2979 , n2981 );
xor ( n3056 , n3055 , n2984 );
xor ( n3057 , n2889 , n2891 );
xor ( n3058 , n3057 , n2894 );
xor ( n3059 , n2958 , n2973 );
xor ( n3060 , n3059 , n2976 );
and ( n3061 , n3058 , n3060 );
and ( n3062 , n3056 , n3061 );
xor ( n3063 , n3047 , n3049 );
and ( n3064 , n3061 , n3063 );
and ( n3065 , n3056 , n3063 );
or ( n3066 , n3062 , n3064 , n3065 );
xor ( n3067 , n3006 , n3008 );
xor ( n3068 , n3067 , n3050 );
and ( n3069 , n3066 , n3068 );
and ( n3070 , n1624 , n1894 );
and ( n3071 , n1610 , n1892 );
nor ( n3072 , n3070 , n3071 );
xnor ( n3073 , n3072 , n1793 );
and ( n3074 , n3019 , n1229 );
and ( n3075 , n2969 , n1227 );
nor ( n3076 , n3074 , n3075 );
xnor ( n3077 , n3076 , n1236 );
and ( n3078 , n3073 , n3077 );
buf ( n3079 , n1178 );
and ( n3080 , n3079 , n1224 );
and ( n3081 , n3077 , n3080 );
and ( n3082 , n3073 , n3080 );
or ( n3083 , n3078 , n3081 , n3082 );
xor ( n3084 , n3013 , n3017 );
xor ( n3085 , n3084 , n3020 );
and ( n3086 , n3083 , n3085 );
xor ( n3087 , n2907 , n2911 );
xor ( n3088 , n3087 , n2916 );
and ( n3089 , n3085 , n3088 );
and ( n3090 , n3083 , n3088 );
or ( n3091 , n3086 , n3089 , n3090 );
xor ( n3092 , n3023 , n3025 );
xor ( n3093 , n3092 , n3028 );
and ( n3094 , n3091 , n3093 );
xor ( n3095 , n3033 , n3035 );
xor ( n3096 , n3095 , n3038 );
and ( n3097 , n3093 , n3096 );
and ( n3098 , n3091 , n3096 );
or ( n3099 , n3094 , n3097 , n3098 );
xor ( n3100 , n3031 , n3041 );
xor ( n3101 , n3100 , n3044 );
and ( n3102 , n3099 , n3101 );
xor ( n3103 , n2919 , n2935 );
xor ( n3104 , n3103 , n2955 );
and ( n3105 , n1521 , n2054 );
and ( n3106 , n1438 , n2052 );
nor ( n3107 , n3105 , n3106 );
xnor ( n3108 , n3107 , n1989 );
and ( n3109 , n2459 , n1322 );
and ( n3110 , n2338 , n1320 );
nor ( n3111 , n3109 , n3110 );
xnor ( n3112 , n3111 , n1293 );
and ( n3113 , n3108 , n3112 );
and ( n3114 , n2658 , n1264 );
and ( n3115 , n2611 , n1262 );
nor ( n3116 , n3114 , n3115 );
xnor ( n3117 , n3116 , n1221 );
and ( n3118 , n3112 , n3117 );
and ( n3119 , n3108 , n3117 );
or ( n3120 , n3113 , n3118 , n3119 );
not ( n3121 , n2962 );
and ( n3122 , n3120 , n3121 );
and ( n3123 , n1661 , n1692 );
and ( n3124 , n1624 , n1690 );
nor ( n3125 , n3123 , n3124 );
xnor ( n3126 , n3125 , n1670 );
and ( n3127 , n3121 , n3126 );
and ( n3128 , n3120 , n3126 );
or ( n3129 , n3122 , n3127 , n3128 );
and ( n3130 , n3104 , n3129 );
and ( n3131 , n1407 , n2221 );
and ( n3132 , n1390 , n2219 );
nor ( n3133 , n3131 , n3132 );
xnor ( n3134 , n3133 , n2138 );
and ( n3135 , n1759 , n1692 );
and ( n3136 , n1661 , n1690 );
nor ( n3137 , n3135 , n3136 );
xnor ( n3138 , n3137 , n1670 );
and ( n3139 , n3134 , n3138 );
and ( n3140 , n1869 , n1604 );
and ( n3141 , n1833 , n1602 );
nor ( n3142 , n3140 , n3141 );
xnor ( n3143 , n3142 , n1549 );
and ( n3144 , n3138 , n3143 );
and ( n3145 , n3134 , n3143 );
or ( n3146 , n3139 , n3144 , n3145 );
and ( n3147 , n1274 , n2666 );
and ( n3148 , n1239 , n2664 );
nor ( n3149 , n3147 , n3148 );
xnor ( n3150 , n3149 , n2587 );
and ( n3151 , n2076 , n1488 );
and ( n3152 , n1963 , n1486 );
nor ( n3153 , n3151 , n3152 );
xnor ( n3154 , n3153 , n1456 );
and ( n3155 , n3150 , n3154 );
and ( n3156 , n2263 , n1398 );
and ( n3157 , n2182 , n1396 );
nor ( n3158 , n3156 , n3157 );
xnor ( n3159 , n3158 , n1348 );
and ( n3160 , n3154 , n3159 );
and ( n3161 , n3150 , n3159 );
or ( n3162 , n3155 , n3160 , n3161 );
and ( n3163 , n3146 , n3162 );
buf ( n3164 , n1211 );
buf ( n3165 , n1212 );
and ( n3166 , n3164 , n3165 );
not ( n3167 , n3166 );
and ( n3168 , n2865 , n3167 );
not ( n3169 , n3168 );
and ( n3170 , n1223 , n2940 );
and ( n3171 , n1231 , n2938 );
nor ( n3172 , n3170 , n3171 );
xnor ( n3173 , n3172 , n2868 );
and ( n3174 , n3169 , n3173 );
and ( n3175 , n3162 , n3174 );
and ( n3176 , n3146 , n3174 );
or ( n3177 , n3163 , n3175 , n3176 );
and ( n3178 , n3129 , n3177 );
and ( n3179 , n3104 , n3177 );
or ( n3180 , n3130 , n3178 , n3179 );
xor ( n3181 , n2923 , n2927 );
xor ( n3182 , n3181 , n2932 );
xor ( n3183 , n2943 , n2947 );
xor ( n3184 , n3183 , n2952 );
and ( n3185 , n3182 , n3184 );
xor ( n3186 , n3120 , n3121 );
xor ( n3187 , n3186 , n3126 );
and ( n3188 , n3184 , n3187 );
and ( n3189 , n3182 , n3187 );
or ( n3190 , n3185 , n3188 , n3189 );
and ( n3191 , n1239 , n2940 );
and ( n3192 , n1223 , n2938 );
nor ( n3193 , n3191 , n3192 );
xnor ( n3194 , n3193 , n2868 );
and ( n3195 , n1390 , n2450 );
and ( n3196 , n1314 , n2448 );
nor ( n3197 , n3195 , n3196 );
xnor ( n3198 , n3197 , n2364 );
and ( n3199 , n3194 , n3198 );
and ( n3200 , n1833 , n1692 );
and ( n3201 , n1759 , n1690 );
nor ( n3202 , n3200 , n3201 );
xnor ( n3203 , n3202 , n1670 );
and ( n3204 , n3198 , n3203 );
and ( n3205 , n3194 , n3203 );
or ( n3206 , n3199 , n3204 , n3205 );
and ( n3207 , n1438 , n2221 );
and ( n3208 , n1407 , n2219 );
nor ( n3209 , n3207 , n3208 );
xnor ( n3210 , n3209 , n2138 );
and ( n3211 , n1963 , n1604 );
and ( n3212 , n1869 , n1602 );
nor ( n3213 , n3211 , n3212 );
xnor ( n3214 , n3213 , n1549 );
and ( n3215 , n3210 , n3214 );
and ( n3216 , n2182 , n1488 );
and ( n3217 , n2076 , n1486 );
nor ( n3218 , n3216 , n3217 );
xnor ( n3219 , n3218 , n1456 );
and ( n3220 , n3214 , n3219 );
and ( n3221 , n3210 , n3219 );
or ( n3222 , n3215 , n3220 , n3221 );
and ( n3223 , n3206 , n3222 );
xor ( n3224 , n2865 , n3164 );
xor ( n3225 , n3164 , n3165 );
not ( n3226 , n3225 );
and ( n3227 , n3224 , n3226 );
and ( n3228 , n1231 , n3227 );
not ( n3229 , n3228 );
xnor ( n3230 , n3229 , n3168 );
buf ( n3231 , n3230 );
and ( n3232 , n3222 , n3231 );
and ( n3233 , n3206 , n3231 );
or ( n3234 , n3223 , n3232 , n3233 );
and ( n3235 , n1661 , n1894 );
and ( n3236 , n1624 , n1892 );
nor ( n3237 , n3235 , n3236 );
xnor ( n3238 , n3237 , n1793 );
and ( n3239 , n2611 , n1322 );
and ( n3240 , n2459 , n1320 );
nor ( n3241 , n3239 , n3240 );
xnor ( n3242 , n3241 , n1293 );
and ( n3243 , n3238 , n3242 );
and ( n3244 , n2969 , n1264 );
and ( n3245 , n2658 , n1262 );
nor ( n3246 , n3244 , n3245 );
xnor ( n3247 , n3246 , n1221 );
and ( n3248 , n3242 , n3247 );
and ( n3249 , n3238 , n3247 );
or ( n3250 , n3243 , n3248 , n3249 );
and ( n3251 , n1300 , n2666 );
and ( n3252 , n1274 , n2664 );
nor ( n3253 , n3251 , n3252 );
xnor ( n3254 , n3253 , n2587 );
and ( n3255 , n1610 , n2054 );
and ( n3256 , n1521 , n2052 );
nor ( n3257 , n3255 , n3256 );
xnor ( n3258 , n3257 , n1989 );
and ( n3259 , n3254 , n3258 );
and ( n3260 , n2338 , n1398 );
and ( n3261 , n2263 , n1396 );
nor ( n3262 , n3260 , n3261 );
xnor ( n3263 , n3262 , n1348 );
and ( n3264 , n3258 , n3263 );
and ( n3265 , n3254 , n3263 );
or ( n3266 , n3259 , n3264 , n3265 );
and ( n3267 , n3250 , n3266 );
xor ( n3268 , n3134 , n3138 );
xor ( n3269 , n3268 , n3143 );
and ( n3270 , n3266 , n3269 );
and ( n3271 , n3250 , n3269 );
or ( n3272 , n3267 , n3270 , n3271 );
and ( n3273 , n3234 , n3272 );
and ( n3274 , n3190 , n3273 );
xor ( n3275 , n3083 , n3085 );
xor ( n3276 , n3275 , n3088 );
and ( n3277 , n1314 , n2450 );
and ( n3278 , n1300 , n2448 );
nor ( n3279 , n3277 , n3278 );
xnor ( n3280 , n3279 , n2364 );
xor ( n3281 , n3073 , n3077 );
xor ( n3282 , n3281 , n3080 );
and ( n3283 , n3280 , n3282 );
xor ( n3284 , n3108 , n3112 );
xor ( n3285 , n3284 , n3117 );
and ( n3286 , n3282 , n3285 );
and ( n3287 , n3280 , n3285 );
or ( n3288 , n3283 , n3286 , n3287 );
and ( n3289 , n3276 , n3288 );
xor ( n3290 , n3146 , n3162 );
xor ( n3291 , n3290 , n3174 );
and ( n3292 , n3288 , n3291 );
and ( n3293 , n3276 , n3291 );
or ( n3294 , n3289 , n3292 , n3293 );
and ( n3295 , n3273 , n3294 );
and ( n3296 , n3190 , n3294 );
or ( n3297 , n3274 , n3295 , n3296 );
and ( n3298 , n3180 , n3297 );
xor ( n3299 , n3058 , n3060 );
and ( n3300 , n3297 , n3299 );
and ( n3301 , n3180 , n3299 );
or ( n3302 , n3298 , n3300 , n3301 );
and ( n3303 , n3102 , n3302 );
xor ( n3304 , n3104 , n3129 );
xor ( n3305 , n3304 , n3177 );
and ( n3306 , n1624 , n2054 );
and ( n3307 , n1610 , n2052 );
nor ( n3308 , n3306 , n3307 );
xnor ( n3309 , n3308 , n1989 );
and ( n3310 , n2658 , n1322 );
and ( n3311 , n2611 , n1320 );
nor ( n3312 , n3310 , n3311 );
xnor ( n3313 , n3312 , n1293 );
and ( n3314 , n3309 , n3313 );
and ( n3315 , n3019 , n1264 );
and ( n3316 , n2969 , n1262 );
nor ( n3317 , n3315 , n3316 );
xnor ( n3318 , n3317 , n1221 );
and ( n3319 , n3313 , n3318 );
and ( n3320 , n3309 , n3318 );
or ( n3321 , n3314 , n3319 , n3320 );
and ( n3322 , n1274 , n2940 );
and ( n3323 , n1239 , n2938 );
nor ( n3324 , n3322 , n3323 );
xnor ( n3325 , n3324 , n2868 );
and ( n3326 , n1521 , n2221 );
and ( n3327 , n1438 , n2219 );
nor ( n3328 , n3326 , n3327 );
xnor ( n3329 , n3328 , n2138 );
and ( n3330 , n3325 , n3329 );
and ( n3331 , n2459 , n1398 );
and ( n3332 , n2338 , n1396 );
nor ( n3333 , n3331 , n3332 );
xnor ( n3334 , n3333 , n1348 );
and ( n3335 , n3329 , n3334 );
and ( n3336 , n3325 , n3334 );
or ( n3337 , n3330 , n3335 , n3336 );
and ( n3338 , n3321 , n3337 );
xor ( n3339 , n3194 , n3198 );
xor ( n3340 , n3339 , n3203 );
and ( n3341 , n3337 , n3340 );
and ( n3342 , n3321 , n3340 );
or ( n3343 , n3338 , n3341 , n3342 );
xor ( n3344 , n3206 , n3222 );
xor ( n3345 , n3344 , n3231 );
and ( n3346 , n3343 , n3345 );
xor ( n3347 , n3250 , n3266 );
xor ( n3348 , n3347 , n3269 );
and ( n3349 , n3345 , n3348 );
and ( n3350 , n3343 , n3348 );
or ( n3351 , n3346 , n3349 , n3350 );
xor ( n3352 , n3182 , n3184 );
xor ( n3353 , n3352 , n3187 );
and ( n3354 , n3351 , n3353 );
and ( n3355 , n3305 , n3354 );
xor ( n3356 , n3234 , n3272 );
and ( n3357 , n1759 , n1894 );
and ( n3358 , n1661 , n1892 );
nor ( n3359 , n3357 , n3358 );
xnor ( n3360 , n3359 , n1793 );
and ( n3361 , n1869 , n1692 );
and ( n3362 , n1833 , n1690 );
nor ( n3363 , n3361 , n3362 );
xnor ( n3364 , n3363 , n1670 );
and ( n3365 , n3360 , n3364 );
buf ( n3366 , n1180 );
and ( n3367 , n3366 , n1224 );
and ( n3368 , n3364 , n3367 );
and ( n3369 , n3360 , n3367 );
or ( n3370 , n3365 , n3368 , n3369 );
buf ( n3371 , n1213 );
buf ( n3372 , n1214 );
and ( n3373 , n3371 , n3372 );
not ( n3374 , n3373 );
and ( n3375 , n3165 , n3374 );
not ( n3376 , n3375 );
and ( n3377 , n1223 , n3227 );
and ( n3378 , n1231 , n3225 );
nor ( n3379 , n3377 , n3378 );
xnor ( n3380 , n3379 , n3168 );
and ( n3381 , n3376 , n3380 );
and ( n3382 , n1314 , n2666 );
and ( n3383 , n1300 , n2664 );
nor ( n3384 , n3382 , n3383 );
xnor ( n3385 , n3384 , n2587 );
and ( n3386 , n3380 , n3385 );
and ( n3387 , n3376 , n3385 );
or ( n3388 , n3381 , n3386 , n3387 );
and ( n3389 , n3370 , n3388 );
and ( n3390 , n1407 , n2450 );
and ( n3391 , n1390 , n2448 );
nor ( n3392 , n3390 , n3391 );
xnor ( n3393 , n3392 , n2364 );
and ( n3394 , n2076 , n1604 );
and ( n3395 , n1963 , n1602 );
nor ( n3396 , n3394 , n3395 );
xnor ( n3397 , n3396 , n1549 );
and ( n3398 , n3393 , n3397 );
and ( n3399 , n2263 , n1488 );
and ( n3400 , n2182 , n1486 );
nor ( n3401 , n3399 , n3400 );
xnor ( n3402 , n3401 , n1456 );
and ( n3403 , n3397 , n3402 );
and ( n3404 , n3393 , n3402 );
or ( n3405 , n3398 , n3403 , n3404 );
and ( n3406 , n3388 , n3405 );
and ( n3407 , n3370 , n3405 );
or ( n3408 , n3389 , n3406 , n3407 );
not ( n3409 , n3230 );
and ( n3410 , n3079 , n1229 );
and ( n3411 , n3019 , n1227 );
nor ( n3412 , n3410 , n3411 );
xnor ( n3413 , n3412 , n1236 );
and ( n3414 , n3409 , n3413 );
buf ( n3415 , n1179 );
and ( n3416 , n3415 , n1224 );
and ( n3417 , n3413 , n3416 );
and ( n3418 , n3409 , n3416 );
or ( n3419 , n3414 , n3417 , n3418 );
and ( n3420 , n3408 , n3419 );
xor ( n3421 , n3150 , n3154 );
xor ( n3422 , n3421 , n3159 );
and ( n3423 , n3419 , n3422 );
and ( n3424 , n3408 , n3422 );
or ( n3425 , n3420 , n3423 , n3424 );
and ( n3426 , n3356 , n3425 );
xor ( n3427 , n3169 , n3173 );
xor ( n3428 , n3238 , n3242 );
xor ( n3429 , n3428 , n3247 );
xor ( n3430 , n3210 , n3214 );
xor ( n3431 , n3430 , n3219 );
and ( n3432 , n3429 , n3431 );
xor ( n3433 , n3254 , n3258 );
xor ( n3434 , n3433 , n3263 );
and ( n3435 , n3431 , n3434 );
and ( n3436 , n3429 , n3434 );
or ( n3437 , n3432 , n3435 , n3436 );
and ( n3438 , n3427 , n3437 );
xor ( n3439 , n3280 , n3282 );
xor ( n3440 , n3439 , n3285 );
and ( n3441 , n3437 , n3440 );
and ( n3442 , n3427 , n3440 );
or ( n3443 , n3438 , n3441 , n3442 );
and ( n3444 , n3425 , n3443 );
and ( n3445 , n3356 , n3443 );
or ( n3446 , n3426 , n3444 , n3445 );
and ( n3447 , n3354 , n3446 );
and ( n3448 , n3305 , n3446 );
or ( n3449 , n3355 , n3447 , n3448 );
xor ( n3450 , n3099 , n3101 );
and ( n3451 , n3449 , n3450 );
xor ( n3452 , n3190 , n3273 );
xor ( n3453 , n3452 , n3294 );
xor ( n3454 , n3091 , n3093 );
xor ( n3455 , n3454 , n3096 );
and ( n3456 , n3453 , n3455 );
xor ( n3457 , n3276 , n3288 );
xor ( n3458 , n3457 , n3291 );
xor ( n3459 , n3351 , n3353 );
and ( n3460 , n3458 , n3459 );
xor ( n3461 , n3408 , n3419 );
xor ( n3462 , n3461 , n3422 );
xor ( n3463 , n3343 , n3345 );
xor ( n3464 , n3463 , n3348 );
and ( n3465 , n3462 , n3464 );
and ( n3466 , n1661 , n2054 );
and ( n3467 , n1624 , n2052 );
nor ( n3468 , n3466 , n3467 );
xnor ( n3469 , n3468 , n1989 );
and ( n3470 , n3079 , n1264 );
and ( n3471 , n3019 , n1262 );
nor ( n3472 , n3470 , n3471 );
xnor ( n3473 , n3472 , n1221 );
and ( n3474 , n3469 , n3473 );
and ( n3475 , n3366 , n1229 );
and ( n3476 , n3415 , n1227 );
nor ( n3477 , n3475 , n3476 );
xnor ( n3478 , n3477 , n1236 );
and ( n3479 , n3473 , n3478 );
and ( n3480 , n3469 , n3478 );
or ( n3481 , n3474 , n3479 , n3480 );
xor ( n3482 , n3360 , n3364 );
xor ( n3483 , n3482 , n3367 );
and ( n3484 , n3481 , n3483 );
xor ( n3485 , n3376 , n3380 );
xor ( n3486 , n3485 , n3385 );
and ( n3487 , n3483 , n3486 );
and ( n3488 , n3481 , n3486 );
or ( n3489 , n3484 , n3487 , n3488 );
xor ( n3490 , n3370 , n3388 );
xor ( n3491 , n3490 , n3405 );
and ( n3492 , n3489 , n3491 );
xor ( n3493 , n3321 , n3337 );
xor ( n3494 , n3493 , n3340 );
and ( n3495 , n3491 , n3494 );
and ( n3496 , n3489 , n3494 );
or ( n3497 , n3492 , n3495 , n3496 );
and ( n3498 , n3464 , n3497 );
and ( n3499 , n3462 , n3497 );
or ( n3500 , n3465 , n3498 , n3499 );
and ( n3501 , n3459 , n3500 );
and ( n3502 , n3458 , n3500 );
or ( n3503 , n3460 , n3501 , n3502 );
and ( n3504 , n3455 , n3503 );
and ( n3505 , n3453 , n3503 );
or ( n3506 , n3456 , n3504 , n3505 );
and ( n3507 , n3450 , n3506 );
and ( n3508 , n3449 , n3506 );
or ( n3509 , n3451 , n3507 , n3508 );
and ( n3510 , n3302 , n3509 );
and ( n3511 , n3102 , n3509 );
or ( n3512 , n3303 , n3510 , n3511 );
and ( n3513 , n3068 , n3512 );
and ( n3514 , n3066 , n3512 );
or ( n3515 , n3069 , n3513 , n3514 );
and ( n3516 , n3053 , n3515 );
and ( n3517 , n3004 , n3515 );
or ( n3518 , n3054 , n3516 , n3517 );
and ( n3519 , n3001 , n3518 );
and ( n3520 , n2847 , n3518 );
or ( n3521 , n3002 , n3519 , n3520 );
and ( n3522 , n2844 , n3521 );
and ( n3523 , n2732 , n3521 );
or ( n3524 , n2845 , n3522 , n3523 );
and ( n3525 , n2729 , n3524 );
and ( n3526 , n2515 , n3524 );
or ( n3527 , n2730 , n3525 , n3526 );
and ( n3528 , n2512 , n3527 );
and ( n3529 , n2446 , n3527 );
or ( n3530 , n2513 , n3528 , n3529 );
and ( n3531 , n2443 , n3530 );
and ( n3532 , n2328 , n3530 );
or ( n3533 , n2444 , n3531 , n3532 );
and ( n3534 , n2325 , n3533 );
and ( n3535 , n2217 , n3533 );
or ( n3536 , n2326 , n3534 , n3535 );
and ( n3537 , n2214 , n3536 );
and ( n3538 , n2123 , n3536 );
or ( n3539 , n2215 , n3537 , n3538 );
and ( n3540 , n2120 , n3539 );
and ( n3541 , n1953 , n3539 );
or ( n3542 , n2121 , n3540 , n3541 );
and ( n3543 , n1950 , n3542 );
and ( n3544 , n1948 , n3542 );
or ( n3545 , n1951 , n3543 , n3544 );
and ( n3546 , n1921 , n3545 );
and ( n3547 , n1788 , n3545 );
or ( n3548 , n1922 , n3546 , n3547 );
and ( n3549 , n1785 , n3548 );
and ( n3550 , n1733 , n3548 );
or ( n3551 , n1786 , n3549 , n3550 );
and ( n3552 , n1730 , n3551 );
and ( n3553 , n1651 , n3551 );
or ( n3554 , n1731 , n3552 , n3553 );
and ( n3555 , n1648 , n3554 );
and ( n3556 , n1544 , n3554 );
or ( n3557 , n1649 , n3555 , n3556 );
and ( n3558 , n1541 , n3557 );
and ( n3559 , n1539 , n3557 );
or ( n3560 , n1542 , n3558 , n3559 );
and ( n3561 , n1483 , n3560 );
and ( n3562 , n1428 , n3560 );
or ( n3563 , n1484 , n3561 , n3562 );
and ( n3564 , n1425 , n3563 );
and ( n3565 , n1379 , n3563 );
or ( n3566 , n1426 , n3564 , n3565 );
and ( n3567 , n1376 , n3566 );
and ( n3568 , n1343 , n3566 );
or ( n3569 , n1377 , n3567 , n3568 );
and ( n3570 , n1340 , n3569 );
and ( n3571 , n1288 , n3569 );
or ( n3572 , n1341 , n3570 , n3571 );
and ( n3573 , n1285 , n3572 );
and ( n3574 , n1260 , n3572 );
or ( n3575 , n1286 , n3573 , n3574 );
xor ( n3576 , n1258 , n3575 );
xor ( n3577 , n1260 , n1285 );
xor ( n3578 , n3577 , n3572 );
xor ( n3579 , n1288 , n1340 );
xor ( n3580 , n3579 , n3569 );
xor ( n3581 , n1343 , n1376 );
xor ( n3582 , n3581 , n3566 );
xor ( n3583 , n1379 , n1425 );
xor ( n3584 , n3583 , n3563 );
xor ( n3585 , n1428 , n1483 );
xor ( n3586 , n3585 , n3560 );
xor ( n3587 , n1539 , n1541 );
xor ( n3588 , n3587 , n3557 );
xor ( n3589 , n1544 , n1648 );
xor ( n3590 , n3589 , n3554 );
xor ( n3591 , n1651 , n1730 );
xor ( n3592 , n3591 , n3551 );
xor ( n3593 , n1733 , n1785 );
xor ( n3594 , n3593 , n3548 );
xor ( n3595 , n1788 , n1921 );
xor ( n3596 , n3595 , n3545 );
xor ( n3597 , n1948 , n1950 );
xor ( n3598 , n3597 , n3542 );
xor ( n3599 , n1953 , n2120 );
xor ( n3600 , n3599 , n3539 );
xor ( n3601 , n2123 , n2214 );
xor ( n3602 , n3601 , n3536 );
xor ( n3603 , n2217 , n2325 );
xor ( n3604 , n3603 , n3533 );
xor ( n3605 , n2328 , n2443 );
xor ( n3606 , n3605 , n3530 );
xor ( n3607 , n2446 , n2512 );
xor ( n3608 , n3607 , n3527 );
xor ( n3609 , n2515 , n2729 );
xor ( n3610 , n3609 , n3524 );
xor ( n3611 , n2732 , n2844 );
xor ( n3612 , n3611 , n3521 );
xor ( n3613 , n2847 , n3001 );
xor ( n3614 , n3613 , n3518 );
xor ( n3615 , n3004 , n3053 );
xor ( n3616 , n3615 , n3515 );
xor ( n3617 , n3056 , n3061 );
xor ( n3618 , n3617 , n3063 );
xor ( n3619 , n3180 , n3297 );
xor ( n3620 , n3619 , n3299 );
xor ( n3621 , n3305 , n3354 );
xor ( n3622 , n3621 , n3446 );
xor ( n3623 , n3356 , n3425 );
xor ( n3624 , n3623 , n3443 );
xor ( n3625 , n3309 , n3313 );
xor ( n3626 , n3625 , n3318 );
xor ( n3627 , n3325 , n3329 );
xor ( n3628 , n3627 , n3334 );
and ( n3629 , n3626 , n3628 );
xor ( n3630 , n3393 , n3397 );
xor ( n3631 , n3630 , n3402 );
and ( n3632 , n3628 , n3631 );
and ( n3633 , n3626 , n3631 );
or ( n3634 , n3629 , n3632 , n3633 );
xor ( n3635 , n3429 , n3431 );
xor ( n3636 , n3635 , n3434 );
and ( n3637 , n3634 , n3636 );
xor ( n3638 , n3427 , n3437 );
xor ( n3639 , n3638 , n3440 );
and ( n3640 , n3637 , n3639 );
xor ( n3641 , n3409 , n3413 );
xor ( n3642 , n3641 , n3416 );
and ( n3643 , n1300 , n2940 );
and ( n3644 , n1274 , n2938 );
nor ( n3645 , n3643 , n3644 );
xnor ( n3646 , n3645 , n2868 );
and ( n3647 , n2182 , n1604 );
and ( n3648 , n2076 , n1602 );
nor ( n3649 , n3647 , n3648 );
xnor ( n3650 , n3649 , n1549 );
and ( n3651 , n3646 , n3650 );
and ( n3652 , n2338 , n1488 );
and ( n3653 , n2263 , n1486 );
nor ( n3654 , n3652 , n3653 );
xnor ( n3655 , n3654 , n1456 );
and ( n3656 , n3650 , n3655 );
and ( n3657 , n3646 , n3655 );
or ( n3658 , n3651 , n3656 , n3657 );
and ( n3659 , n1610 , n2221 );
and ( n3660 , n1521 , n2219 );
nor ( n3661 , n3659 , n3660 );
xnor ( n3662 , n3661 , n2138 );
and ( n3663 , n2611 , n1398 );
and ( n3664 , n2459 , n1396 );
nor ( n3665 , n3663 , n3664 );
xnor ( n3666 , n3665 , n1348 );
and ( n3667 , n3662 , n3666 );
and ( n3668 , n2969 , n1322 );
and ( n3669 , n2658 , n1320 );
nor ( n3670 , n3668 , n3669 );
xnor ( n3671 , n3670 , n1293 );
and ( n3672 , n3666 , n3671 );
and ( n3673 , n3662 , n3671 );
or ( n3674 , n3667 , n3672 , n3673 );
and ( n3675 , n3658 , n3674 );
and ( n3676 , n1438 , n2450 );
and ( n3677 , n1407 , n2448 );
nor ( n3678 , n3676 , n3677 );
xnor ( n3679 , n3678 , n2364 );
and ( n3680 , n1833 , n1894 );
and ( n3681 , n1759 , n1892 );
nor ( n3682 , n3680 , n3681 );
xnor ( n3683 , n3682 , n1793 );
and ( n3684 , n3679 , n3683 );
and ( n3685 , n1963 , n1692 );
and ( n3686 , n1869 , n1690 );
nor ( n3687 , n3685 , n3686 );
xnor ( n3688 , n3687 , n1670 );
and ( n3689 , n3683 , n3688 );
and ( n3690 , n3679 , n3688 );
or ( n3691 , n3684 , n3689 , n3690 );
and ( n3692 , n3674 , n3691 );
and ( n3693 , n3658 , n3691 );
or ( n3694 , n3675 , n3692 , n3693 );
and ( n3695 , n3642 , n3694 );
xor ( n3696 , n3489 , n3491 );
xor ( n3697 , n3696 , n3494 );
and ( n3698 , n3694 , n3697 );
and ( n3699 , n3642 , n3697 );
or ( n3700 , n3695 , n3698 , n3699 );
and ( n3701 , n3639 , n3700 );
and ( n3702 , n3637 , n3700 );
or ( n3703 , n3640 , n3701 , n3702 );
and ( n3704 , n3624 , n3703 );
xor ( n3705 , n3458 , n3459 );
xor ( n3706 , n3705 , n3500 );
and ( n3707 , n3703 , n3706 );
and ( n3708 , n3624 , n3706 );
or ( n3709 , n3704 , n3707 , n3708 );
and ( n3710 , n3622 , n3709 );
xor ( n3711 , n3453 , n3455 );
xor ( n3712 , n3711 , n3503 );
and ( n3713 , n3709 , n3712 );
and ( n3714 , n3622 , n3712 );
or ( n3715 , n3710 , n3713 , n3714 );
and ( n3716 , n3620 , n3715 );
xor ( n3717 , n3449 , n3450 );
xor ( n3718 , n3717 , n3506 );
and ( n3719 , n3715 , n3718 );
and ( n3720 , n3620 , n3718 );
or ( n3721 , n3716 , n3719 , n3720 );
and ( n3722 , n3618 , n3721 );
xor ( n3723 , n3102 , n3302 );
xor ( n3724 , n3723 , n3509 );
and ( n3725 , n3721 , n3724 );
and ( n3726 , n3618 , n3724 );
or ( n3727 , n3722 , n3725 , n3726 );
xor ( n3728 , n3066 , n3068 );
xor ( n3729 , n3728 , n3512 );
and ( n3730 , n3727 , n3729 );
xor ( n3731 , n3727 , n3729 );
xor ( n3732 , n3618 , n3721 );
xor ( n3733 , n3732 , n3724 );
xor ( n3734 , n3620 , n3715 );
xor ( n3735 , n3734 , n3718 );
xor ( n3736 , n3622 , n3709 );
xor ( n3737 , n3736 , n3712 );
xor ( n3738 , n3634 , n3636 );
and ( n3739 , n1239 , n3227 );
and ( n3740 , n1223 , n3225 );
nor ( n3741 , n3739 , n3740 );
xnor ( n3742 , n3741 , n3168 );
and ( n3743 , n1390 , n2666 );
and ( n3744 , n1314 , n2664 );
nor ( n3745 , n3743 , n3744 );
xnor ( n3746 , n3745 , n2587 );
xor ( n3747 , n3742 , n3746 );
buf ( n3748 , n1181 );
and ( n3749 , n3748 , n1224 );
xor ( n3750 , n3747 , n3749 );
xor ( n3751 , n3646 , n3650 );
xor ( n3752 , n3751 , n3655 );
and ( n3753 , n3750 , n3752 );
xor ( n3754 , n3662 , n3666 );
xor ( n3755 , n3754 , n3671 );
and ( n3756 , n3752 , n3755 );
and ( n3757 , n3750 , n3755 );
or ( n3758 , n3753 , n3756 , n3757 );
and ( n3759 , n1624 , n2221 );
and ( n3760 , n1610 , n2219 );
nor ( n3761 , n3759 , n3760 );
xnor ( n3762 , n3761 , n2138 );
and ( n3763 , n2658 , n1398 );
and ( n3764 , n2611 , n1396 );
nor ( n3765 , n3763 , n3764 );
xnor ( n3766 , n3765 , n1348 );
and ( n3767 , n3762 , n3766 );
and ( n3768 , n3019 , n1322 );
and ( n3769 , n2969 , n1320 );
nor ( n3770 , n3768 , n3769 );
xnor ( n3771 , n3770 , n1293 );
and ( n3772 , n3766 , n3771 );
and ( n3773 , n3762 , n3771 );
or ( n3774 , n3767 , n3772 , n3773 );
xor ( n3775 , n3679 , n3683 );
xor ( n3776 , n3775 , n3688 );
and ( n3777 , n3774 , n3776 );
xor ( n3778 , n3469 , n3473 );
xor ( n3779 , n3778 , n3478 );
and ( n3780 , n3776 , n3779 );
and ( n3781 , n3774 , n3779 );
or ( n3782 , n3777 , n3780 , n3781 );
and ( n3783 , n3758 , n3782 );
xor ( n3784 , n3658 , n3674 );
xor ( n3785 , n3784 , n3691 );
and ( n3786 , n3782 , n3785 );
and ( n3787 , n3758 , n3785 );
or ( n3788 , n3783 , n3786 , n3787 );
and ( n3789 , n3738 , n3788 );
xor ( n3790 , n3481 , n3483 );
xor ( n3791 , n3790 , n3486 );
xor ( n3792 , n3626 , n3628 );
xor ( n3793 , n3792 , n3631 );
and ( n3794 , n3791 , n3793 );
and ( n3795 , n3788 , n3794 );
and ( n3796 , n3738 , n3794 );
or ( n3797 , n3789 , n3795 , n3796 );
xor ( n3798 , n3462 , n3464 );
xor ( n3799 , n3798 , n3497 );
and ( n3800 , n3797 , n3799 );
and ( n3801 , n3415 , n1229 );
and ( n3802 , n3079 , n1227 );
nor ( n3803 , n3801 , n3802 );
xnor ( n3804 , n3803 , n1236 );
and ( n3805 , n3742 , n3746 );
and ( n3806 , n3746 , n3749 );
and ( n3807 , n3742 , n3749 );
or ( n3808 , n3805 , n3806 , n3807 );
and ( n3809 , n3804 , n3808 );
xor ( n3810 , n3165 , n3371 );
xor ( n3811 , n3371 , n3372 );
not ( n3812 , n3811 );
and ( n3813 , n3810 , n3812 );
and ( n3814 , n1223 , n3813 );
and ( n3815 , n1231 , n3811 );
nor ( n3816 , n3814 , n3815 );
xnor ( n3817 , n3816 , n3375 );
and ( n3818 , n1314 , n2940 );
and ( n3819 , n1300 , n2938 );
nor ( n3820 , n3818 , n3819 );
xnor ( n3821 , n3820 , n2868 );
and ( n3822 , n3817 , n3821 );
and ( n3823 , n1869 , n1894 );
and ( n3824 , n1833 , n1892 );
nor ( n3825 , n3823 , n3824 );
xnor ( n3826 , n3825 , n1793 );
and ( n3827 , n3821 , n3826 );
and ( n3828 , n3817 , n3826 );
or ( n3829 , n3822 , n3827 , n3828 );
and ( n3830 , n1274 , n3227 );
and ( n3831 , n1239 , n3225 );
nor ( n3832 , n3830 , n3831 );
xnor ( n3833 , n3832 , n3168 );
and ( n3834 , n1521 , n2450 );
and ( n3835 , n1438 , n2448 );
nor ( n3836 , n3834 , n3835 );
xnor ( n3837 , n3836 , n2364 );
and ( n3838 , n3833 , n3837 );
and ( n3839 , n2459 , n1488 );
and ( n3840 , n2338 , n1486 );
nor ( n3841 , n3839 , n3840 );
xnor ( n3842 , n3841 , n1456 );
and ( n3843 , n3837 , n3842 );
and ( n3844 , n3833 , n3842 );
or ( n3845 , n3838 , n3843 , n3844 );
and ( n3846 , n3829 , n3845 );
and ( n3847 , n1407 , n2666 );
and ( n3848 , n1390 , n2664 );
nor ( n3849 , n3847 , n3848 );
xnor ( n3850 , n3849 , n2587 );
and ( n3851 , n2076 , n1692 );
and ( n3852 , n1963 , n1690 );
nor ( n3853 , n3851 , n3852 );
xnor ( n3854 , n3853 , n1670 );
and ( n3855 , n3850 , n3854 );
and ( n3856 , n2263 , n1604 );
and ( n3857 , n2182 , n1602 );
nor ( n3858 , n3856 , n3857 );
xnor ( n3859 , n3858 , n1549 );
and ( n3860 , n3854 , n3859 );
and ( n3861 , n3850 , n3859 );
or ( n3862 , n3855 , n3860 , n3861 );
and ( n3863 , n3845 , n3862 );
and ( n3864 , n3829 , n3862 );
or ( n3865 , n3846 , n3863 , n3864 );
and ( n3866 , n3808 , n3865 );
and ( n3867 , n3804 , n3865 );
or ( n3868 , n3809 , n3866 , n3867 );
xor ( n3869 , n3758 , n3782 );
xor ( n3870 , n3869 , n3785 );
xor ( n3871 , n3791 , n3793 );
and ( n3872 , n3870 , n3871 );
and ( n3873 , n1390 , n2940 );
and ( n3874 , n1314 , n2938 );
nor ( n3875 , n3873 , n3874 );
xnor ( n3876 , n3875 , n2868 );
and ( n3877 , n1833 , n2054 );
and ( n3878 , n1759 , n2052 );
nor ( n3879 , n3877 , n3878 );
xnor ( n3880 , n3879 , n1989 );
and ( n3881 , n3876 , n3880 );
buf ( n3882 , n1182 );
and ( n3883 , n3882 , n1229 );
and ( n3884 , n3748 , n1227 );
nor ( n3885 , n3883 , n3884 );
xnor ( n3886 , n3885 , n1236 );
and ( n3887 , n3880 , n3886 );
and ( n3888 , n3876 , n3886 );
or ( n3889 , n3881 , n3887 , n3888 );
and ( n3890 , n1661 , n2221 );
and ( n3891 , n1624 , n2219 );
nor ( n3892 , n3890 , n3891 );
xnor ( n3893 , n3892 , n2138 );
and ( n3894 , n2611 , n1488 );
and ( n3895 , n2459 , n1486 );
nor ( n3896 , n3894 , n3895 );
xnor ( n3897 , n3896 , n1456 );
and ( n3898 , n3893 , n3897 );
and ( n3899 , n2969 , n1398 );
and ( n3900 , n2658 , n1396 );
nor ( n3901 , n3899 , n3900 );
xnor ( n3902 , n3901 , n1348 );
and ( n3903 , n3897 , n3902 );
and ( n3904 , n3893 , n3902 );
or ( n3905 , n3898 , n3903 , n3904 );
and ( n3906 , n3889 , n3905 );
and ( n3907 , n1438 , n2666 );
and ( n3908 , n1407 , n2664 );
nor ( n3909 , n3907 , n3908 );
xnor ( n3910 , n3909 , n2587 );
and ( n3911 , n1963 , n1894 );
and ( n3912 , n1869 , n1892 );
nor ( n3913 , n3911 , n3912 );
xnor ( n3914 , n3913 , n1793 );
and ( n3915 , n3910 , n3914 );
and ( n3916 , n2182 , n1692 );
and ( n3917 , n2076 , n1690 );
nor ( n3918 , n3916 , n3917 );
xnor ( n3919 , n3918 , n1670 );
and ( n3920 , n3914 , n3919 );
and ( n3921 , n3910 , n3919 );
or ( n3922 , n3915 , n3920 , n3921 );
and ( n3923 , n3905 , n3922 );
and ( n3924 , n3889 , n3922 );
or ( n3925 , n3906 , n3923 , n3924 );
buf ( n3926 , n1215 );
xor ( n3927 , n3372 , n3926 );
not ( n3928 , n3926 );
and ( n3929 , n3927 , n3928 );
and ( n3930 , n1231 , n3929 );
not ( n3931 , n3930 );
xnor ( n3932 , n3931 , n3372 );
and ( n3933 , n1239 , n3813 );
and ( n3934 , n1223 , n3811 );
nor ( n3935 , n3933 , n3934 );
xnor ( n3936 , n3935 , n3375 );
and ( n3937 , n3932 , n3936 );
buf ( n3938 , n1183 );
and ( n3939 , n3938 , n1224 );
and ( n3940 , n3936 , n3939 );
and ( n3941 , n3932 , n3939 );
or ( n3942 , n3937 , n3940 , n3941 );
and ( n3943 , n3942 , n3372 );
and ( n3944 , n3415 , n1264 );
and ( n3945 , n3079 , n1262 );
nor ( n3946 , n3944 , n3945 );
xnor ( n3947 , n3946 , n1221 );
and ( n3948 , n3372 , n3947 );
and ( n3949 , n3942 , n3947 );
or ( n3950 , n3943 , n3948 , n3949 );
and ( n3951 , n3925 , n3950 );
xor ( n3952 , n3829 , n3845 );
xor ( n3953 , n3952 , n3862 );
and ( n3954 , n3950 , n3953 );
and ( n3955 , n3925 , n3953 );
or ( n3956 , n3951 , n3954 , n3955 );
and ( n3957 , n3871 , n3956 );
and ( n3958 , n3870 , n3956 );
or ( n3959 , n3872 , n3957 , n3958 );
and ( n3960 , n3868 , n3959 );
xor ( n3961 , n3642 , n3694 );
xor ( n3962 , n3961 , n3697 );
and ( n3963 , n3959 , n3962 );
and ( n3964 , n3868 , n3962 );
or ( n3965 , n3960 , n3963 , n3964 );
and ( n3966 , n3799 , n3965 );
and ( n3967 , n3797 , n3965 );
or ( n3968 , n3800 , n3966 , n3967 );
xor ( n3969 , n3624 , n3703 );
xor ( n3970 , n3969 , n3706 );
and ( n3971 , n3968 , n3970 );
xor ( n3972 , n3637 , n3639 );
xor ( n3973 , n3972 , n3700 );
xor ( n3974 , n3738 , n3788 );
xor ( n3975 , n3974 , n3794 );
and ( n3976 , n1231 , n3813 );
not ( n3977 , n3976 );
xnor ( n3978 , n3977 , n3375 );
and ( n3979 , n1759 , n2054 );
and ( n3980 , n1661 , n2052 );
nor ( n3981 , n3979 , n3980 );
xnor ( n3982 , n3981 , n1989 );
and ( n3983 , n3748 , n1229 );
and ( n3984 , n3366 , n1227 );
nor ( n3985 , n3983 , n3984 );
xnor ( n3986 , n3985 , n1236 );
and ( n3987 , n3982 , n3986 );
and ( n3988 , n3882 , n1224 );
and ( n3989 , n3986 , n3988 );
and ( n3990 , n3982 , n3988 );
or ( n3991 , n3987 , n3989 , n3990 );
and ( n3992 , n3978 , n3991 );
not ( n3993 , n3372 );
buf ( n3994 , n3993 );
and ( n3995 , n3991 , n3994 );
and ( n3996 , n3978 , n3994 );
or ( n3997 , n3992 , n3995 , n3996 );
xor ( n3998 , n3804 , n3808 );
xor ( n3999 , n3998 , n3865 );
and ( n4000 , n3997 , n3999 );
and ( n4001 , n1300 , n3227 );
and ( n4002 , n1274 , n3225 );
nor ( n4003 , n4001 , n4002 );
xnor ( n4004 , n4003 , n3168 );
and ( n4005 , n1610 , n2450 );
and ( n4006 , n1521 , n2448 );
nor ( n4007 , n4005 , n4006 );
xnor ( n4008 , n4007 , n2364 );
xor ( n4009 , n4004 , n4008 );
and ( n4010 , n2338 , n1604 );
and ( n4011 , n2263 , n1602 );
nor ( n4012 , n4010 , n4011 );
xnor ( n4013 , n4012 , n1549 );
xor ( n4014 , n4009 , n4013 );
xor ( n4015 , n3893 , n3897 );
xor ( n4016 , n4015 , n3902 );
and ( n4017 , n4014 , n4016 );
xor ( n4018 , n3910 , n3914 );
xor ( n4019 , n4018 , n3919 );
and ( n4020 , n4016 , n4019 );
and ( n4021 , n4014 , n4019 );
or ( n4022 , n4017 , n4020 , n4021 );
xor ( n4023 , n3889 , n3905 );
xor ( n4024 , n4023 , n3922 );
and ( n4025 , n4022 , n4024 );
xor ( n4026 , n3942 , n3372 );
xor ( n4027 , n4026 , n3947 );
and ( n4028 , n4024 , n4027 );
and ( n4029 , n4022 , n4027 );
or ( n4030 , n4025 , n4028 , n4029 );
xor ( n4031 , n3750 , n3752 );
xor ( n4032 , n4031 , n3755 );
and ( n4033 , n4030 , n4032 );
xor ( n4034 , n3774 , n3776 );
xor ( n4035 , n4034 , n3779 );
and ( n4036 , n4032 , n4035 );
and ( n4037 , n4030 , n4035 );
or ( n4038 , n4033 , n4036 , n4037 );
and ( n4039 , n3999 , n4038 );
and ( n4040 , n3997 , n4038 );
or ( n4041 , n4000 , n4039 , n4040 );
and ( n4042 , n3975 , n4041 );
and ( n4043 , n1223 , n3929 );
and ( n4044 , n1231 , n3926 );
nor ( n4045 , n4043 , n4044 );
xnor ( n4046 , n4045 , n3372 );
and ( n4047 , n3938 , n1227 );
not ( n4048 , n4047 );
and ( n4049 , n4048 , n1236 );
and ( n4050 , n4046 , n4049 );
and ( n4051 , n3079 , n1322 );
and ( n4052 , n3019 , n1320 );
nor ( n4053 , n4051 , n4052 );
xnor ( n4054 , n4053 , n1293 );
and ( n4055 , n4050 , n4054 );
and ( n4056 , n3366 , n1264 );
and ( n4057 , n3415 , n1262 );
nor ( n4058 , n4056 , n4057 );
xnor ( n4059 , n4058 , n1221 );
and ( n4060 , n4054 , n4059 );
and ( n4061 , n4050 , n4059 );
or ( n4062 , n4055 , n4060 , n4061 );
and ( n4063 , n1274 , n3813 );
and ( n4064 , n1239 , n3811 );
nor ( n4065 , n4063 , n4064 );
xnor ( n4066 , n4065 , n3375 );
and ( n4067 , n1407 , n2940 );
and ( n4068 , n1390 , n2938 );
nor ( n4069 , n4067 , n4068 );
xnor ( n4070 , n4069 , n2868 );
and ( n4071 , n4066 , n4070 );
and ( n4072 , n3938 , n1229 );
and ( n4073 , n3882 , n1227 );
nor ( n4074 , n4072 , n4073 );
xnor ( n4075 , n4074 , n1236 );
and ( n4076 , n4070 , n4075 );
and ( n4077 , n4066 , n4075 );
or ( n4078 , n4071 , n4076 , n4077 );
and ( n4079 , n1521 , n2666 );
and ( n4080 , n1438 , n2664 );
nor ( n4081 , n4079 , n4080 );
xnor ( n4082 , n4081 , n2587 );
and ( n4083 , n1869 , n2054 );
and ( n4084 , n1833 , n2052 );
nor ( n4085 , n4083 , n4084 );
xnor ( n4086 , n4085 , n1989 );
and ( n4087 , n4082 , n4086 );
and ( n4088 , n2076 , n1894 );
and ( n4089 , n1963 , n1892 );
nor ( n4090 , n4088 , n4089 );
xnor ( n4091 , n4090 , n1793 );
and ( n4092 , n4086 , n4091 );
and ( n4093 , n4082 , n4091 );
or ( n4094 , n4087 , n4092 , n4093 );
and ( n4095 , n4078 , n4094 );
and ( n4096 , n1314 , n3227 );
and ( n4097 , n1300 , n3225 );
nor ( n4098 , n4096 , n4097 );
xnor ( n4099 , n4098 , n3168 );
and ( n4100 , n2263 , n1692 );
and ( n4101 , n2182 , n1690 );
nor ( n4102 , n4100 , n4101 );
xnor ( n4103 , n4102 , n1670 );
and ( n4104 , n4099 , n4103 );
and ( n4105 , n2459 , n1604 );
and ( n4106 , n2338 , n1602 );
nor ( n4107 , n4105 , n4106 );
xnor ( n4108 , n4107 , n1549 );
and ( n4109 , n4103 , n4108 );
and ( n4110 , n4099 , n4108 );
or ( n4111 , n4104 , n4109 , n4110 );
and ( n4112 , n4094 , n4111 );
and ( n4113 , n4078 , n4111 );
or ( n4114 , n4095 , n4112 , n4113 );
and ( n4115 , n4062 , n4114 );
and ( n4116 , n1759 , n2221 );
and ( n4117 , n1661 , n2219 );
nor ( n4118 , n4116 , n4117 );
xnor ( n4119 , n4118 , n2138 );
and ( n4120 , n3415 , n1322 );
and ( n4121 , n3079 , n1320 );
nor ( n4122 , n4120 , n4121 );
xnor ( n4123 , n4122 , n1293 );
and ( n4124 , n4119 , n4123 );
and ( n4125 , n3748 , n1264 );
and ( n4126 , n3366 , n1262 );
nor ( n4127 , n4125 , n4126 );
xnor ( n4128 , n4127 , n1221 );
and ( n4129 , n4123 , n4128 );
and ( n4130 , n4119 , n4128 );
or ( n4131 , n4124 , n4129 , n4130 );
and ( n4132 , n1624 , n2450 );
and ( n4133 , n1610 , n2448 );
nor ( n4134 , n4132 , n4133 );
xnor ( n4135 , n4134 , n2364 );
and ( n4136 , n2658 , n1488 );
and ( n4137 , n2611 , n1486 );
nor ( n4138 , n4136 , n4137 );
xnor ( n4139 , n4138 , n1456 );
and ( n4140 , n4135 , n4139 );
and ( n4141 , n3019 , n1398 );
and ( n4142 , n2969 , n1396 );
nor ( n4143 , n4141 , n4142 );
xnor ( n4144 , n4143 , n1348 );
and ( n4145 , n4139 , n4144 );
and ( n4146 , n4135 , n4144 );
or ( n4147 , n4140 , n4145 , n4146 );
and ( n4148 , n4131 , n4147 );
xor ( n4149 , n3932 , n3936 );
xor ( n4150 , n4149 , n3939 );
and ( n4151 , n4147 , n4150 );
and ( n4152 , n4131 , n4150 );
or ( n4153 , n4148 , n4151 , n4152 );
and ( n4154 , n4114 , n4153 );
and ( n4155 , n4062 , n4153 );
or ( n4156 , n4115 , n4154 , n4155 );
not ( n4157 , n4156 );
xor ( n4158 , n3925 , n3950 );
xor ( n4159 , n4158 , n3953 );
and ( n4160 , n4157 , n4159 );
buf ( n4161 , n4156 );
and ( n4162 , n4160 , n4161 );
xor ( n4163 , n3817 , n3821 );
xor ( n4164 , n4163 , n3826 );
xor ( n4165 , n3833 , n3837 );
xor ( n4166 , n4165 , n3842 );
and ( n4167 , n4164 , n4166 );
xor ( n4168 , n3850 , n3854 );
xor ( n4169 , n4168 , n3859 );
and ( n4170 , n4166 , n4169 );
and ( n4171 , n4164 , n4169 );
or ( n4172 , n4167 , n4170 , n4171 );
xor ( n4173 , n3762 , n3766 );
xor ( n4174 , n4173 , n3771 );
and ( n4175 , n4004 , n4008 );
and ( n4176 , n4008 , n4013 );
and ( n4177 , n4004 , n4013 );
or ( n4178 , n4175 , n4176 , n4177 );
and ( n4179 , n4174 , n4178 );
xor ( n4180 , n3982 , n3986 );
xor ( n4181 , n4180 , n3988 );
and ( n4182 , n4178 , n4181 );
and ( n4183 , n4174 , n4181 );
or ( n4184 , n4179 , n4182 , n4183 );
and ( n4185 , n4172 , n4184 );
xor ( n4186 , n3978 , n3991 );
xor ( n4187 , n4186 , n3994 );
and ( n4188 , n4184 , n4187 );
and ( n4189 , n4172 , n4187 );
or ( n4190 , n4185 , n4188 , n4189 );
and ( n4191 , n4161 , n4190 );
and ( n4192 , n4160 , n4190 );
or ( n4193 , n4162 , n4191 , n4192 );
and ( n4194 , n4041 , n4193 );
and ( n4195 , n3975 , n4193 );
or ( n4196 , n4042 , n4194 , n4195 );
and ( n4197 , n3973 , n4196 );
xor ( n4198 , n3797 , n3799 );
xor ( n4199 , n4198 , n3965 );
and ( n4200 , n4196 , n4199 );
and ( n4201 , n3973 , n4199 );
or ( n4202 , n4197 , n4200 , n4201 );
and ( n4203 , n3970 , n4202 );
and ( n4204 , n3968 , n4202 );
or ( n4205 , n3971 , n4203 , n4204 );
and ( n4206 , n3737 , n4205 );
xor ( n4207 , n3737 , n4205 );
xor ( n4208 , n3968 , n3970 );
xor ( n4209 , n4208 , n4202 );
xor ( n4210 , n3868 , n3959 );
xor ( n4211 , n4210 , n3962 );
xor ( n4212 , n3870 , n3871 );
xor ( n4213 , n4212 , n3956 );
xor ( n4214 , n4030 , n4032 );
xor ( n4215 , n4214 , n4035 );
xor ( n4216 , n4157 , n4159 );
and ( n4217 , n4215 , n4216 );
xor ( n4218 , n4046 , n4049 );
and ( n4219 , n1239 , n3929 );
and ( n4220 , n1223 , n3926 );
nor ( n4221 , n4219 , n4220 );
xnor ( n4222 , n4221 , n3372 );
and ( n4223 , n1300 , n3813 );
and ( n4224 , n1274 , n3811 );
nor ( n4225 , n4223 , n4224 );
xnor ( n4226 , n4225 , n3375 );
and ( n4227 , n4222 , n4226 );
and ( n4228 , n4226 , n4047 );
and ( n4229 , n4222 , n4047 );
or ( n4230 , n4227 , n4228 , n4229 );
and ( n4231 , n4218 , n4230 );
and ( n4232 , n1438 , n2940 );
and ( n4233 , n1407 , n2938 );
nor ( n4234 , n4232 , n4233 );
xnor ( n4235 , n4234 , n2868 );
and ( n4236 , n1963 , n2054 );
and ( n4237 , n1869 , n2052 );
nor ( n4238 , n4236 , n4237 );
xnor ( n4239 , n4238 , n1989 );
and ( n4240 , n4235 , n4239 );
and ( n4241 , n2182 , n1894 );
and ( n4242 , n2076 , n1892 );
nor ( n4243 , n4241 , n4242 );
xnor ( n4244 , n4243 , n1793 );
and ( n4245 , n4239 , n4244 );
and ( n4246 , n4235 , n4244 );
or ( n4247 , n4240 , n4245 , n4246 );
and ( n4248 , n4230 , n4247 );
and ( n4249 , n4218 , n4247 );
or ( n4250 , n4231 , n4248 , n4249 );
xor ( n4251 , n4066 , n4070 );
xor ( n4252 , n4251 , n4075 );
xor ( n4253 , n4119 , n4123 );
xor ( n4254 , n4253 , n4128 );
and ( n4255 , n4252 , n4254 );
xor ( n4256 , n4082 , n4086 );
xor ( n4257 , n4256 , n4091 );
and ( n4258 , n4254 , n4257 );
and ( n4259 , n4252 , n4257 );
or ( n4260 , n4255 , n4258 , n4259 );
and ( n4261 , n4250 , n4260 );
xor ( n4262 , n4131 , n4147 );
xor ( n4263 , n4262 , n4150 );
and ( n4264 , n4260 , n4263 );
and ( n4265 , n4250 , n4263 );
or ( n4266 , n4261 , n4264 , n4265 );
xor ( n4267 , n4062 , n4114 );
xor ( n4268 , n4267 , n4153 );
and ( n4269 , n4266 , n4268 );
xor ( n4270 , n4022 , n4024 );
xor ( n4271 , n4270 , n4027 );
and ( n4272 , n4268 , n4271 );
and ( n4273 , n4266 , n4271 );
or ( n4274 , n4269 , n4272 , n4273 );
and ( n4275 , n4216 , n4274 );
and ( n4276 , n4215 , n4274 );
or ( n4277 , n4217 , n4275 , n4276 );
and ( n4278 , n4213 , n4277 );
xor ( n4279 , n3997 , n3999 );
xor ( n4280 , n4279 , n4038 );
and ( n4281 , n4277 , n4280 );
and ( n4282 , n4213 , n4280 );
or ( n4283 , n4278 , n4281 , n4282 );
and ( n4284 , n4211 , n4283 );
xor ( n4285 , n3975 , n4041 );
xor ( n4286 , n4285 , n4193 );
and ( n4287 , n4283 , n4286 );
and ( n4288 , n4211 , n4286 );
or ( n4289 , n4284 , n4287 , n4288 );
xor ( n4290 , n3973 , n4196 );
xor ( n4291 , n4290 , n4199 );
and ( n4292 , n4289 , n4291 );
xor ( n4293 , n4289 , n4291 );
xor ( n4294 , n4160 , n4161 );
xor ( n4295 , n4294 , n4190 );
xor ( n4296 , n4164 , n4166 );
xor ( n4297 , n4296 , n4169 );
xor ( n4298 , n4174 , n4178 );
xor ( n4299 , n4298 , n4181 );
and ( n4300 , n4297 , n4299 );
and ( n4301 , n1390 , n3227 );
and ( n4302 , n1314 , n3225 );
nor ( n4303 , n4301 , n4302 );
xnor ( n4304 , n4303 , n3168 );
and ( n4305 , n1661 , n2450 );
and ( n4306 , n1624 , n2448 );
nor ( n4307 , n4305 , n4306 );
xnor ( n4308 , n4307 , n2364 );
and ( n4309 , n4304 , n4308 );
and ( n4310 , n2969 , n1488 );
and ( n4311 , n2658 , n1486 );
nor ( n4312 , n4310 , n4311 );
xnor ( n4313 , n4312 , n1456 );
and ( n4314 , n4308 , n4313 );
and ( n4315 , n4304 , n4313 );
or ( n4316 , n4309 , n4314 , n4315 );
and ( n4317 , n1833 , n2221 );
and ( n4318 , n1759 , n2219 );
nor ( n4319 , n4317 , n4318 );
xnor ( n4320 , n4319 , n2138 );
and ( n4321 , n3079 , n1398 );
and ( n4322 , n3019 , n1396 );
nor ( n4323 , n4321 , n4322 );
xnor ( n4324 , n4323 , n1348 );
and ( n4325 , n4320 , n4324 );
and ( n4326 , n3366 , n1322 );
and ( n4327 , n3415 , n1320 );
nor ( n4328 , n4326 , n4327 );
xnor ( n4329 , n4328 , n1293 );
and ( n4330 , n4324 , n4329 );
and ( n4331 , n4320 , n4329 );
or ( n4332 , n4325 , n4330 , n4331 );
and ( n4333 , n4316 , n4332 );
and ( n4334 , n1610 , n2666 );
and ( n4335 , n1521 , n2664 );
nor ( n4336 , n4334 , n4335 );
xnor ( n4337 , n4336 , n2587 );
and ( n4338 , n2338 , n1692 );
and ( n4339 , n2263 , n1690 );
nor ( n4340 , n4338 , n4339 );
xnor ( n4341 , n4340 , n1670 );
and ( n4342 , n4337 , n4341 );
and ( n4343 , n2611 , n1604 );
and ( n4344 , n2459 , n1602 );
nor ( n4345 , n4343 , n4344 );
xnor ( n4346 , n4345 , n1549 );
and ( n4347 , n4341 , n4346 );
and ( n4348 , n4337 , n4346 );
or ( n4349 , n4342 , n4347 , n4348 );
and ( n4350 , n4332 , n4349 );
and ( n4351 , n4316 , n4349 );
or ( n4352 , n4333 , n4350 , n4351 );
xor ( n4353 , n3876 , n3880 );
xor ( n4354 , n4353 , n3886 );
and ( n4355 , n4352 , n4354 );
xor ( n4356 , n4050 , n4054 );
xor ( n4357 , n4356 , n4059 );
and ( n4358 , n4354 , n4357 );
and ( n4359 , n4352 , n4357 );
or ( n4360 , n4355 , n4358 , n4359 );
and ( n4361 , n4299 , n4360 );
and ( n4362 , n4297 , n4360 );
or ( n4363 , n4300 , n4361 , n4362 );
xor ( n4364 , n4172 , n4184 );
xor ( n4365 , n4364 , n4187 );
and ( n4366 , n4363 , n4365 );
xor ( n4367 , n4078 , n4094 );
xor ( n4368 , n4367 , n4111 );
xor ( n4369 , n4014 , n4016 );
xor ( n4370 , n4369 , n4019 );
and ( n4371 , n4368 , n4370 );
xor ( n4372 , n4099 , n4103 );
xor ( n4373 , n4372 , n4108 );
xor ( n4374 , n4135 , n4139 );
xor ( n4375 , n4374 , n4144 );
and ( n4376 , n4373 , n4375 );
and ( n4377 , n4370 , n4376 );
and ( n4378 , n4368 , n4376 );
or ( n4379 , n4371 , n4377 , n4378 );
xor ( n4380 , n4266 , n4268 );
xor ( n4381 , n4380 , n4271 );
and ( n4382 , n4379 , n4381 );
xor ( n4383 , n4297 , n4299 );
xor ( n4384 , n4383 , n4360 );
and ( n4385 , n4381 , n4384 );
and ( n4386 , n4379 , n4384 );
or ( n4387 , n4382 , n4385 , n4386 );
and ( n4388 , n4365 , n4387 );
and ( n4389 , n4363 , n4387 );
or ( n4390 , n4366 , n4388 , n4389 );
and ( n4391 , n4295 , n4390 );
xor ( n4392 , n4213 , n4277 );
xor ( n4393 , n4392 , n4280 );
and ( n4394 , n4390 , n4393 );
and ( n4395 , n4295 , n4393 );
or ( n4396 , n4391 , n4394 , n4395 );
xor ( n4397 , n4211 , n4283 );
xor ( n4398 , n4397 , n4286 );
and ( n4399 , n4396 , n4398 );
xor ( n4400 , n4396 , n4398 );
xor ( n4401 , n4215 , n4216 );
xor ( n4402 , n4401 , n4274 );
and ( n4403 , n1314 , n3813 );
and ( n4404 , n1300 , n3811 );
nor ( n4405 , n4403 , n4404 );
xnor ( n4406 , n4405 , n3375 );
and ( n4407 , n1521 , n2940 );
and ( n4408 , n1438 , n2938 );
nor ( n4409 , n4407 , n4408 );
xnor ( n4410 , n4409 , n2868 );
and ( n4411 , n4406 , n4410 );
and ( n4412 , n2076 , n2054 );
and ( n4413 , n1963 , n2052 );
nor ( n4414 , n4412 , n4413 );
xnor ( n4415 , n4414 , n1989 );
and ( n4416 , n4410 , n4415 );
and ( n4417 , n4406 , n4415 );
or ( n4418 , n4411 , n4416 , n4417 );
and ( n4419 , n1274 , n3929 );
and ( n4420 , n1239 , n3926 );
nor ( n4421 , n4419 , n4420 );
xnor ( n4422 , n4421 , n3372 );
and ( n4423 , n3938 , n1262 );
not ( n4424 , n4423 );
and ( n4425 , n4424 , n1221 );
and ( n4426 , n4422 , n4425 );
and ( n4427 , n4418 , n4426 );
and ( n4428 , n3882 , n1264 );
and ( n4429 , n3748 , n1262 );
nor ( n4430 , n4428 , n4429 );
xnor ( n4431 , n4430 , n1221 );
and ( n4432 , n4426 , n4431 );
and ( n4433 , n4418 , n4431 );
or ( n4434 , n4427 , n4432 , n4433 );
xor ( n4435 , n4316 , n4332 );
xor ( n4436 , n4435 , n4349 );
and ( n4437 , n4434 , n4436 );
xor ( n4438 , n4218 , n4230 );
xor ( n4439 , n4438 , n4247 );
and ( n4440 , n4436 , n4439 );
and ( n4441 , n4434 , n4439 );
or ( n4442 , n4437 , n4440 , n4441 );
xor ( n4443 , n4304 , n4308 );
xor ( n4444 , n4443 , n4313 );
xor ( n4445 , n4222 , n4226 );
xor ( n4446 , n4445 , n4047 );
and ( n4447 , n4444 , n4446 );
xor ( n4448 , n4320 , n4324 );
xor ( n4449 , n4448 , n4329 );
and ( n4450 , n4446 , n4449 );
and ( n4451 , n4444 , n4449 );
or ( n4452 , n4447 , n4450 , n4451 );
xor ( n4453 , n4422 , n4425 );
and ( n4454 , n3748 , n1322 );
and ( n4455 , n3366 , n1320 );
nor ( n4456 , n4454 , n4455 );
xnor ( n4457 , n4456 , n1293 );
and ( n4458 , n4453 , n4457 );
and ( n4459 , n3938 , n1264 );
and ( n4460 , n3882 , n1262 );
nor ( n4461 , n4459 , n4460 );
xnor ( n4462 , n4461 , n1221 );
and ( n4463 , n4457 , n4462 );
and ( n4464 , n4453 , n4462 );
or ( n4465 , n4458 , n4463 , n4464 );
xor ( n4466 , n4337 , n4341 );
xor ( n4467 , n4466 , n4346 );
and ( n4468 , n4465 , n4467 );
xor ( n4469 , n4235 , n4239 );
xor ( n4470 , n4469 , n4244 );
and ( n4471 , n4467 , n4470 );
and ( n4472 , n4465 , n4470 );
or ( n4473 , n4468 , n4471 , n4472 );
and ( n4474 , n4452 , n4473 );
xor ( n4475 , n4252 , n4254 );
xor ( n4476 , n4475 , n4257 );
and ( n4477 , n4473 , n4476 );
and ( n4478 , n4452 , n4476 );
or ( n4479 , n4474 , n4477 , n4478 );
and ( n4480 , n4442 , n4479 );
xor ( n4481 , n4352 , n4354 );
xor ( n4482 , n4481 , n4357 );
and ( n4483 , n4479 , n4482 );
and ( n4484 , n4442 , n4482 );
or ( n4485 , n4480 , n4483 , n4484 );
xor ( n4486 , n4250 , n4260 );
xor ( n4487 , n4486 , n4263 );
xor ( n4488 , n4368 , n4370 );
xor ( n4489 , n4488 , n4376 );
and ( n4490 , n4487 , n4489 );
xor ( n4491 , n4373 , n4375 );
and ( n4492 , n1869 , n2221 );
and ( n4493 , n1833 , n2219 );
nor ( n4494 , n4492 , n4493 );
xnor ( n4495 , n4494 , n2138 );
and ( n4496 , n3019 , n1488 );
and ( n4497 , n2969 , n1486 );
nor ( n4498 , n4496 , n4497 );
xnor ( n4499 , n4498 , n1456 );
and ( n4500 , n4495 , n4499 );
and ( n4501 , n3415 , n1398 );
and ( n4502 , n3079 , n1396 );
nor ( n4503 , n4501 , n4502 );
xnor ( n4504 , n4503 , n1348 );
and ( n4505 , n4499 , n4504 );
and ( n4506 , n4495 , n4504 );
or ( n4507 , n4500 , n4505 , n4506 );
and ( n4508 , n1407 , n3227 );
and ( n4509 , n1390 , n3225 );
nor ( n4510 , n4508 , n4509 );
xnor ( n4511 , n4510 , n3168 );
and ( n4512 , n1759 , n2450 );
and ( n4513 , n1661 , n2448 );
nor ( n4514 , n4512 , n4513 );
xnor ( n4515 , n4514 , n2364 );
and ( n4516 , n4511 , n4515 );
and ( n4517 , n2658 , n1604 );
and ( n4518 , n2611 , n1602 );
nor ( n4519 , n4517 , n4518 );
xnor ( n4520 , n4519 , n1549 );
and ( n4521 , n4515 , n4520 );
and ( n4522 , n4511 , n4520 );
or ( n4523 , n4516 , n4521 , n4522 );
and ( n4524 , n4507 , n4523 );
and ( n4525 , n1624 , n2666 );
and ( n4526 , n1610 , n2664 );
nor ( n4527 , n4525 , n4526 );
xnor ( n4528 , n4527 , n2587 );
and ( n4529 , n2459 , n1692 );
and ( n4530 , n2338 , n1690 );
nor ( n4531 , n4529 , n4530 );
xnor ( n4532 , n4531 , n1670 );
and ( n4533 , n4528 , n4532 );
and ( n4534 , n4523 , n4533 );
and ( n4535 , n4507 , n4533 );
or ( n4536 , n4524 , n4534 , n4535 );
and ( n4537 , n4491 , n4536 );
and ( n4538 , n1390 , n3813 );
and ( n4539 , n1314 , n3811 );
nor ( n4540 , n4538 , n4539 );
xnor ( n4541 , n4540 , n3375 );
and ( n4542 , n1610 , n2940 );
and ( n4543 , n1521 , n2938 );
nor ( n4544 , n4542 , n4543 );
xnor ( n4545 , n4544 , n2868 );
and ( n4546 , n4541 , n4545 );
and ( n4547 , n4545 , n4423 );
and ( n4548 , n4541 , n4423 );
or ( n4549 , n4546 , n4547 , n4548 );
and ( n4550 , n1300 , n3929 );
and ( n4551 , n1274 , n3926 );
nor ( n4552 , n4550 , n4551 );
xnor ( n4553 , n4552 , n3372 );
and ( n4554 , n2611 , n1692 );
and ( n4555 , n2459 , n1690 );
nor ( n4556 , n4554 , n4555 );
xnor ( n4557 , n4556 , n1670 );
and ( n4558 , n4553 , n4557 );
and ( n4559 , n2969 , n1604 );
and ( n4560 , n2658 , n1602 );
nor ( n4561 , n4559 , n4560 );
xnor ( n4562 , n4561 , n1549 );
and ( n4563 , n4557 , n4562 );
and ( n4564 , n4553 , n4562 );
or ( n4565 , n4558 , n4563 , n4564 );
and ( n4566 , n4549 , n4565 );
and ( n4567 , n1661 , n2666 );
and ( n4568 , n1624 , n2664 );
nor ( n4569 , n4567 , n4568 );
xnor ( n4570 , n4569 , n2587 );
and ( n4571 , n2182 , n2054 );
and ( n4572 , n2076 , n2052 );
nor ( n4573 , n4571 , n4572 );
xnor ( n4574 , n4573 , n1989 );
and ( n4575 , n4570 , n4574 );
and ( n4576 , n2338 , n1894 );
and ( n4577 , n2263 , n1892 );
nor ( n4578 , n4576 , n4577 );
xnor ( n4579 , n4578 , n1793 );
and ( n4580 , n4574 , n4579 );
and ( n4581 , n4570 , n4579 );
or ( n4582 , n4575 , n4580 , n4581 );
and ( n4583 , n4565 , n4582 );
and ( n4584 , n4549 , n4582 );
or ( n4585 , n4566 , n4583 , n4584 );
xor ( n4586 , n4418 , n4426 );
xor ( n4587 , n4586 , n4431 );
and ( n4588 , n4585 , n4587 );
and ( n4589 , n4536 , n4588 );
and ( n4590 , n4491 , n4588 );
or ( n4591 , n4537 , n4589 , n4590 );
and ( n4592 , n4489 , n4591 );
and ( n4593 , n4487 , n4591 );
or ( n4594 , n4490 , n4592 , n4593 );
and ( n4595 , n4485 , n4594 );
xor ( n4596 , n4379 , n4381 );
xor ( n4597 , n4596 , n4384 );
and ( n4598 , n4594 , n4597 );
and ( n4599 , n4485 , n4597 );
or ( n4600 , n4595 , n4598 , n4599 );
and ( n4601 , n4402 , n4600 );
xor ( n4602 , n4363 , n4365 );
xor ( n4603 , n4602 , n4387 );
and ( n4604 , n4600 , n4603 );
and ( n4605 , n4402 , n4603 );
or ( n4606 , n4601 , n4604 , n4605 );
xor ( n4607 , n4295 , n4390 );
xor ( n4608 , n4607 , n4393 );
and ( n4609 , n4606 , n4608 );
xor ( n4610 , n4606 , n4608 );
xor ( n4611 , n4402 , n4600 );
xor ( n4612 , n4611 , n4603 );
xor ( n4613 , n4442 , n4479 );
xor ( n4614 , n4613 , n4482 );
and ( n4615 , n1624 , n2940 );
and ( n4616 , n1610 , n2938 );
nor ( n4617 , n4615 , n4616 );
xnor ( n4618 , n4617 , n2868 );
and ( n4619 , n2263 , n2054 );
and ( n4620 , n2182 , n2052 );
nor ( n4621 , n4619 , n4620 );
xnor ( n4622 , n4621 , n1989 );
and ( n4623 , n4618 , n4622 );
and ( n4624 , n2459 , n1894 );
and ( n4625 , n2338 , n1892 );
nor ( n4626 , n4624 , n4625 );
xnor ( n4627 , n4626 , n1793 );
and ( n4628 , n4622 , n4627 );
and ( n4629 , n4618 , n4627 );
or ( n4630 , n4623 , n4628 , n4629 );
and ( n4631 , n1759 , n2666 );
and ( n4632 , n1661 , n2664 );
nor ( n4633 , n4631 , n4632 );
xnor ( n4634 , n4633 , n2587 );
and ( n4635 , n2658 , n1692 );
and ( n4636 , n2611 , n1690 );
nor ( n4637 , n4635 , n4636 );
xnor ( n4638 , n4637 , n1670 );
and ( n4639 , n4634 , n4638 );
and ( n4640 , n3019 , n1604 );
and ( n4641 , n2969 , n1602 );
nor ( n4642 , n4640 , n4641 );
xnor ( n4643 , n4642 , n1549 );
and ( n4644 , n4638 , n4643 );
and ( n4645 , n4634 , n4643 );
or ( n4646 , n4639 , n4644 , n4645 );
and ( n4647 , n4630 , n4646 );
and ( n4648 , n1407 , n3813 );
and ( n4649 , n1390 , n3811 );
nor ( n4650 , n4648 , n4649 );
xnor ( n4651 , n4650 , n3375 );
and ( n4652 , n3938 , n1320 );
not ( n4653 , n4652 );
and ( n4654 , n4653 , n1293 );
and ( n4655 , n4651 , n4654 );
and ( n4656 , n4646 , n4655 );
and ( n4657 , n4630 , n4655 );
or ( n4658 , n4647 , n4656 , n4657 );
xor ( n4659 , n4541 , n4545 );
xor ( n4660 , n4659 , n4423 );
and ( n4661 , n1438 , n3227 );
and ( n4662 , n1407 , n3225 );
nor ( n4663 , n4661 , n4662 );
xnor ( n4664 , n4663 , n3168 );
and ( n4665 , n1963 , n2221 );
and ( n4666 , n1869 , n2219 );
nor ( n4667 , n4665 , n4666 );
xnor ( n4668 , n4667 , n2138 );
xor ( n4669 , n4664 , n4668 );
and ( n4670 , n3882 , n1322 );
and ( n4671 , n3748 , n1320 );
nor ( n4672 , n4670 , n4671 );
xnor ( n4673 , n4672 , n1293 );
xor ( n4674 , n4669 , n4673 );
and ( n4675 , n4660 , n4674 );
xor ( n4676 , n4553 , n4557 );
xor ( n4677 , n4676 , n4562 );
and ( n4678 , n4674 , n4677 );
and ( n4679 , n4660 , n4677 );
or ( n4680 , n4675 , n4678 , n4679 );
and ( n4681 , n4658 , n4680 );
xor ( n4682 , n4453 , n4457 );
xor ( n4683 , n4682 , n4462 );
and ( n4684 , n4680 , n4683 );
and ( n4685 , n4658 , n4683 );
or ( n4686 , n4681 , n4684 , n4685 );
and ( n4687 , n1314 , n3929 );
and ( n4688 , n1300 , n3926 );
nor ( n4689 , n4687 , n4688 );
xnor ( n4690 , n4689 , n3372 );
and ( n4691 , n1869 , n2450 );
and ( n4692 , n1833 , n2448 );
nor ( n4693 , n4691 , n4692 );
xnor ( n4694 , n4693 , n2364 );
and ( n4695 , n4690 , n4694 );
and ( n4696 , n3415 , n1488 );
and ( n4697 , n3079 , n1486 );
nor ( n4698 , n4696 , n4697 );
xnor ( n4699 , n4698 , n1456 );
and ( n4700 , n4694 , n4699 );
and ( n4701 , n4690 , n4699 );
or ( n4702 , n4695 , n4700 , n4701 );
and ( n4703 , n1521 , n3227 );
and ( n4704 , n1438 , n3225 );
nor ( n4705 , n4703 , n4704 );
xnor ( n4706 , n4705 , n3168 );
and ( n4707 , n3748 , n1398 );
and ( n4708 , n3366 , n1396 );
nor ( n4709 , n4707 , n4708 );
xnor ( n4710 , n4709 , n1348 );
and ( n4711 , n4706 , n4710 );
and ( n4712 , n3938 , n1322 );
and ( n4713 , n3882 , n1320 );
nor ( n4714 , n4712 , n4713 );
xnor ( n4715 , n4714 , n1293 );
and ( n4716 , n4710 , n4715 );
and ( n4717 , n4706 , n4715 );
or ( n4718 , n4711 , n4716 , n4717 );
and ( n4719 , n4702 , n4718 );
xor ( n4720 , n4570 , n4574 );
xor ( n4721 , n4720 , n4579 );
and ( n4722 , n4718 , n4721 );
and ( n4723 , n4702 , n4721 );
or ( n4724 , n4719 , n4722 , n4723 );
xor ( n4725 , n4549 , n4565 );
xor ( n4726 , n4725 , n4582 );
and ( n4727 , n4724 , n4726 );
and ( n4728 , n4664 , n4668 );
and ( n4729 , n4668 , n4673 );
and ( n4730 , n4664 , n4673 );
or ( n4731 , n4728 , n4729 , n4730 );
and ( n4732 , n1833 , n2450 );
and ( n4733 , n1759 , n2448 );
nor ( n4734 , n4732 , n4733 );
xnor ( n4735 , n4734 , n2364 );
and ( n4736 , n3079 , n1488 );
and ( n4737 , n3019 , n1486 );
nor ( n4738 , n4736 , n4737 );
xnor ( n4739 , n4738 , n1456 );
and ( n4740 , n4735 , n4739 );
and ( n4741 , n3366 , n1398 );
and ( n4742 , n3415 , n1396 );
nor ( n4743 , n4741 , n4742 );
xnor ( n4744 , n4743 , n1348 );
and ( n4745 , n4739 , n4744 );
and ( n4746 , n4735 , n4744 );
or ( n4747 , n4740 , n4745 , n4746 );
xor ( n4748 , n4731 , n4747 );
xor ( n4749 , n4406 , n4410 );
xor ( n4750 , n4749 , n4415 );
xor ( n4751 , n4748 , n4750 );
and ( n4752 , n4726 , n4751 );
and ( n4753 , n4724 , n4751 );
or ( n4754 , n4727 , n4752 , n4753 );
and ( n4755 , n4686 , n4754 );
xor ( n4756 , n4444 , n4446 );
xor ( n4757 , n4756 , n4449 );
and ( n4758 , n4754 , n4757 );
and ( n4759 , n4686 , n4757 );
or ( n4760 , n4755 , n4758 , n4759 );
xor ( n4761 , n4434 , n4436 );
xor ( n4762 , n4761 , n4439 );
and ( n4763 , n4760 , n4762 );
xor ( n4764 , n4452 , n4473 );
xor ( n4765 , n4764 , n4476 );
and ( n4766 , n4762 , n4765 );
and ( n4767 , n4760 , n4765 );
or ( n4768 , n4763 , n4766 , n4767 );
and ( n4769 , n4614 , n4768 );
and ( n4770 , n4731 , n4747 );
and ( n4771 , n4747 , n4750 );
and ( n4772 , n4731 , n4750 );
or ( n4773 , n4770 , n4771 , n4772 );
and ( n4774 , n2263 , n1894 );
and ( n4775 , n2182 , n1892 );
nor ( n4776 , n4774 , n4775 );
xnor ( n4777 , n4776 , n1793 );
xor ( n4778 , n4495 , n4499 );
xor ( n4779 , n4778 , n4504 );
and ( n4780 , n4777 , n4779 );
xor ( n4781 , n4511 , n4515 );
xor ( n4782 , n4781 , n4520 );
and ( n4783 , n4779 , n4782 );
and ( n4784 , n4777 , n4782 );
or ( n4785 , n4780 , n4783 , n4784 );
and ( n4786 , n4773 , n4785 );
xor ( n4787 , n4507 , n4523 );
xor ( n4788 , n4787 , n4533 );
and ( n4789 , n4785 , n4788 );
and ( n4790 , n4773 , n4788 );
or ( n4791 , n4786 , n4789 , n4790 );
xor ( n4792 , n4465 , n4467 );
xor ( n4793 , n4792 , n4470 );
xor ( n4794 , n4585 , n4587 );
and ( n4795 , n4793 , n4794 );
xor ( n4796 , n4773 , n4785 );
xor ( n4797 , n4796 , n4788 );
and ( n4798 , n4794 , n4797 );
and ( n4799 , n4793 , n4797 );
or ( n4800 , n4795 , n4798 , n4799 );
and ( n4801 , n4791 , n4800 );
xor ( n4802 , n4491 , n4536 );
xor ( n4803 , n4802 , n4588 );
and ( n4804 , n4800 , n4803 );
and ( n4805 , n4791 , n4803 );
or ( n4806 , n4801 , n4804 , n4805 );
and ( n4807 , n4768 , n4806 );
and ( n4808 , n4614 , n4806 );
or ( n4809 , n4769 , n4807 , n4808 );
xor ( n4810 , n4485 , n4594 );
xor ( n4811 , n4810 , n4597 );
and ( n4812 , n4809 , n4811 );
xor ( n4813 , n4487 , n4489 );
xor ( n4814 , n4813 , n4591 );
xor ( n4815 , n4760 , n4762 );
xor ( n4816 , n4815 , n4765 );
xor ( n4817 , n4686 , n4754 );
xor ( n4818 , n4817 , n4757 );
xor ( n4819 , n4658 , n4680 );
xor ( n4820 , n4819 , n4683 );
xor ( n4821 , n4724 , n4726 );
xor ( n4822 , n4821 , n4751 );
and ( n4823 , n4820 , n4822 );
and ( n4824 , n4818 , n4823 );
xor ( n4825 , n4528 , n4532 );
xor ( n4826 , n4777 , n4779 );
xor ( n4827 , n4826 , n4782 );
and ( n4828 , n4825 , n4827 );
and ( n4829 , n1963 , n2450 );
and ( n4830 , n1869 , n2448 );
nor ( n4831 , n4829 , n4830 );
xnor ( n4832 , n4831 , n2364 );
and ( n4833 , n3366 , n1488 );
and ( n4834 , n3415 , n1486 );
nor ( n4835 , n4833 , n4834 );
xnor ( n4836 , n4835 , n1456 );
and ( n4837 , n4832 , n4836 );
and ( n4838 , n3882 , n1398 );
and ( n4839 , n3748 , n1396 );
nor ( n4840 , n4838 , n4839 );
xnor ( n4841 , n4840 , n1348 );
and ( n4842 , n4836 , n4841 );
and ( n4843 , n4832 , n4841 );
or ( n4844 , n4837 , n4842 , n4843 );
and ( n4845 , n1833 , n2666 );
and ( n4846 , n1759 , n2664 );
nor ( n4847 , n4845 , n4846 );
xnor ( n4848 , n4847 , n2587 );
and ( n4849 , n2338 , n2054 );
and ( n4850 , n2263 , n2052 );
nor ( n4851 , n4849 , n4850 );
xnor ( n4852 , n4851 , n1989 );
and ( n4853 , n4848 , n4852 );
and ( n4854 , n2611 , n1894 );
and ( n4855 , n2459 , n1892 );
nor ( n4856 , n4854 , n4855 );
xnor ( n4857 , n4856 , n1793 );
and ( n4858 , n4852 , n4857 );
and ( n4859 , n4848 , n4857 );
or ( n4860 , n4853 , n4858 , n4859 );
and ( n4861 , n4844 , n4860 );
and ( n4862 , n1390 , n3929 );
and ( n4863 , n1314 , n3926 );
nor ( n4864 , n4862 , n4863 );
xnor ( n4865 , n4864 , n3372 );
and ( n4866 , n2969 , n1692 );
and ( n4867 , n2658 , n1690 );
nor ( n4868 , n4866 , n4867 );
xnor ( n4869 , n4868 , n1670 );
and ( n4870 , n4865 , n4869 );
and ( n4871 , n3079 , n1604 );
and ( n4872 , n3019 , n1602 );
nor ( n4873 , n4871 , n4872 );
xnor ( n4874 , n4873 , n1549 );
and ( n4875 , n4869 , n4874 );
and ( n4876 , n4865 , n4874 );
or ( n4877 , n4870 , n4875 , n4876 );
and ( n4878 , n4860 , n4877 );
and ( n4879 , n4844 , n4877 );
or ( n4880 , n4861 , n4878 , n4879 );
xor ( n4881 , n4651 , n4654 );
and ( n4882 , n1438 , n3813 );
and ( n4883 , n1407 , n3811 );
nor ( n4884 , n4882 , n4883 );
xnor ( n4885 , n4884 , n3375 );
and ( n4886 , n1661 , n2940 );
and ( n4887 , n1624 , n2938 );
nor ( n4888 , n4886 , n4887 );
xnor ( n4889 , n4888 , n2868 );
and ( n4890 , n4885 , n4889 );
and ( n4891 , n4889 , n4652 );
and ( n4892 , n4885 , n4652 );
or ( n4893 , n4890 , n4891 , n4892 );
and ( n4894 , n4881 , n4893 );
and ( n4895 , n2076 , n2221 );
and ( n4896 , n1963 , n2219 );
nor ( n4897 , n4895 , n4896 );
xnor ( n4898 , n4897 , n2138 );
and ( n4899 , n4893 , n4898 );
and ( n4900 , n4881 , n4898 );
or ( n4901 , n4894 , n4899 , n4900 );
and ( n4902 , n4880 , n4901 );
xor ( n4903 , n4735 , n4739 );
xor ( n4904 , n4903 , n4744 );
and ( n4905 , n4901 , n4904 );
and ( n4906 , n4880 , n4904 );
or ( n4907 , n4902 , n4905 , n4906 );
and ( n4908 , n4827 , n4907 );
and ( n4909 , n4825 , n4907 );
or ( n4910 , n4828 , n4908 , n4909 );
and ( n4911 , n4823 , n4910 );
and ( n4912 , n4818 , n4910 );
or ( n4913 , n4824 , n4911 , n4912 );
and ( n4914 , n4816 , n4913 );
xor ( n4915 , n4791 , n4800 );
xor ( n4916 , n4915 , n4803 );
and ( n4917 , n4913 , n4916 );
and ( n4918 , n4816 , n4916 );
or ( n4919 , n4914 , n4917 , n4918 );
and ( n4920 , n4814 , n4919 );
xor ( n4921 , n4614 , n4768 );
xor ( n4922 , n4921 , n4806 );
and ( n4923 , n4919 , n4922 );
and ( n4924 , n4814 , n4922 );
or ( n4925 , n4920 , n4923 , n4924 );
and ( n4926 , n4811 , n4925 );
and ( n4927 , n4809 , n4925 );
or ( n4928 , n4812 , n4926 , n4927 );
and ( n4929 , n4612 , n4928 );
xor ( n4930 , n4612 , n4928 );
xor ( n4931 , n4809 , n4811 );
xor ( n4932 , n4931 , n4925 );
xor ( n4933 , n4814 , n4919 );
xor ( n4934 , n4933 , n4922 );
xor ( n4935 , n4793 , n4794 );
xor ( n4936 , n4935 , n4797 );
xor ( n4937 , n4618 , n4622 );
xor ( n4938 , n4937 , n4627 );
xor ( n4939 , n4690 , n4694 );
xor ( n4940 , n4939 , n4699 );
and ( n4941 , n4938 , n4940 );
xor ( n4942 , n4706 , n4710 );
xor ( n4943 , n4942 , n4715 );
and ( n4944 , n4940 , n4943 );
and ( n4945 , n4938 , n4943 );
or ( n4946 , n4941 , n4944 , n4945 );
xor ( n4947 , n4630 , n4646 );
xor ( n4948 , n4947 , n4655 );
and ( n4949 , n4946 , n4948 );
xor ( n4950 , n4702 , n4718 );
xor ( n4951 , n4950 , n4721 );
and ( n4952 , n4948 , n4951 );
and ( n4953 , n4946 , n4951 );
or ( n4954 , n4949 , n4952 , n4953 );
xor ( n4955 , n4820 , n4822 );
and ( n4956 , n4954 , n4955 );
xor ( n4957 , n4825 , n4827 );
xor ( n4958 , n4957 , n4907 );
and ( n4959 , n4955 , n4958 );
and ( n4960 , n4954 , n4958 );
or ( n4961 , n4956 , n4959 , n4960 );
and ( n4962 , n4936 , n4961 );
xor ( n4963 , n4818 , n4823 );
xor ( n4964 , n4963 , n4910 );
and ( n4965 , n4961 , n4964 );
and ( n4966 , n4936 , n4964 );
or ( n4967 , n4962 , n4965 , n4966 );
xor ( n4968 , n4816 , n4913 );
xor ( n4969 , n4968 , n4916 );
and ( n4970 , n4967 , n4969 );
and ( n4971 , n1521 , n3813 );
and ( n4972 , n1438 , n3811 );
nor ( n4973 , n4971 , n4972 );
xnor ( n4974 , n4973 , n3375 );
and ( n4975 , n3938 , n1396 );
not ( n4976 , n4975 );
and ( n4977 , n4976 , n1348 );
and ( n4978 , n4974 , n4977 );
and ( n4979 , n1610 , n3227 );
and ( n4980 , n1521 , n3225 );
nor ( n4981 , n4979 , n4980 );
xnor ( n4982 , n4981 , n3168 );
and ( n4983 , n4978 , n4982 );
and ( n4984 , n2182 , n2221 );
and ( n4985 , n2076 , n2219 );
nor ( n4986 , n4984 , n4985 );
xnor ( n4987 , n4986 , n2138 );
and ( n4988 , n4982 , n4987 );
and ( n4989 , n4978 , n4987 );
or ( n4990 , n4983 , n4988 , n4989 );
xor ( n4991 , n4634 , n4638 );
xor ( n4992 , n4991 , n4643 );
and ( n4993 , n4990 , n4992 );
xor ( n4994 , n4881 , n4893 );
xor ( n4995 , n4994 , n4898 );
and ( n4996 , n4992 , n4995 );
and ( n4997 , n4990 , n4995 );
or ( n4998 , n4993 , n4996 , n4997 );
and ( n4999 , n1407 , n3929 );
and ( n5000 , n1390 , n3926 );
nor ( n5001 , n4999 , n5000 );
xnor ( n5002 , n5001 , n3372 );
and ( n5003 , n2076 , n2450 );
and ( n5004 , n1963 , n2448 );
nor ( n5005 , n5003 , n5004 );
xnor ( n5006 , n5005 , n2364 );
and ( n5007 , n5002 , n5006 );
and ( n5008 , n3748 , n1488 );
and ( n5009 , n3366 , n1486 );
nor ( n5010 , n5008 , n5009 );
xnor ( n5011 , n5010 , n1456 );
and ( n5012 , n5006 , n5011 );
and ( n5013 , n5002 , n5011 );
or ( n5014 , n5007 , n5012 , n5013 );
and ( n5015 , n1759 , n2940 );
and ( n5016 , n1661 , n2938 );
nor ( n5017 , n5015 , n5016 );
xnor ( n5018 , n5017 , n2868 );
and ( n5019 , n2459 , n2054 );
and ( n5020 , n2338 , n2052 );
nor ( n5021 , n5019 , n5020 );
xnor ( n5022 , n5021 , n1989 );
and ( n5023 , n5018 , n5022 );
and ( n5024 , n2658 , n1894 );
and ( n5025 , n2611 , n1892 );
nor ( n5026 , n5024 , n5025 );
xnor ( n5027 , n5026 , n1793 );
and ( n5028 , n5022 , n5027 );
and ( n5029 , n5018 , n5027 );
or ( n5030 , n5023 , n5028 , n5029 );
and ( n5031 , n5014 , n5030 );
and ( n5032 , n1869 , n2666 );
and ( n5033 , n1833 , n2664 );
nor ( n5034 , n5032 , n5033 );
xnor ( n5035 , n5034 , n2587 );
and ( n5036 , n3019 , n1692 );
and ( n5037 , n2969 , n1690 );
nor ( n5038 , n5036 , n5037 );
xnor ( n5039 , n5038 , n1670 );
and ( n5040 , n5035 , n5039 );
and ( n5041 , n3415 , n1604 );
and ( n5042 , n3079 , n1602 );
nor ( n5043 , n5041 , n5042 );
xnor ( n5044 , n5043 , n1549 );
and ( n5045 , n5039 , n5044 );
and ( n5046 , n5035 , n5044 );
or ( n5047 , n5040 , n5045 , n5046 );
and ( n5048 , n5030 , n5047 );
and ( n5049 , n5014 , n5047 );
or ( n5050 , n5031 , n5048 , n5049 );
and ( n5051 , n1624 , n3227 );
and ( n5052 , n1610 , n3225 );
nor ( n5053 , n5051 , n5052 );
xnor ( n5054 , n5053 , n3168 );
and ( n5055 , n2263 , n2221 );
and ( n5056 , n2182 , n2219 );
nor ( n5057 , n5055 , n5056 );
xnor ( n5058 , n5057 , n2138 );
and ( n5059 , n5054 , n5058 );
and ( n5060 , n3938 , n1398 );
and ( n5061 , n3882 , n1396 );
nor ( n5062 , n5060 , n5061 );
xnor ( n5063 , n5062 , n1348 );
and ( n5064 , n5058 , n5063 );
and ( n5065 , n5054 , n5063 );
or ( n5066 , n5059 , n5064 , n5065 );
xor ( n5067 , n4885 , n4889 );
xor ( n5068 , n5067 , n4652 );
and ( n5069 , n5066 , n5068 );
xor ( n5070 , n4865 , n4869 );
xor ( n5071 , n5070 , n4874 );
and ( n5072 , n5068 , n5071 );
and ( n5073 , n5066 , n5071 );
or ( n5074 , n5069 , n5072 , n5073 );
and ( n5075 , n5050 , n5074 );
xor ( n5076 , n4844 , n4860 );
xor ( n5077 , n5076 , n4877 );
and ( n5078 , n5074 , n5077 );
and ( n5079 , n5050 , n5077 );
or ( n5080 , n5075 , n5078 , n5079 );
and ( n5081 , n4998 , n5080 );
xor ( n5082 , n4660 , n4674 );
xor ( n5083 , n5082 , n4677 );
and ( n5084 , n5080 , n5083 );
and ( n5085 , n4998 , n5083 );
or ( n5086 , n5081 , n5084 , n5085 );
xor ( n5087 , n4832 , n4836 );
xor ( n5088 , n5087 , n4841 );
xor ( n5089 , n4848 , n4852 );
xor ( n5090 , n5089 , n4857 );
and ( n5091 , n5088 , n5090 );
xor ( n5092 , n4978 , n4982 );
xor ( n5093 , n5092 , n4987 );
and ( n5094 , n5090 , n5093 );
and ( n5095 , n5088 , n5093 );
or ( n5096 , n5091 , n5094 , n5095 );
xor ( n5097 , n4938 , n4940 );
xor ( n5098 , n5097 , n4943 );
and ( n5099 , n5096 , n5098 );
xor ( n5100 , n4990 , n4992 );
xor ( n5101 , n5100 , n4995 );
and ( n5102 , n5098 , n5101 );
and ( n5103 , n5096 , n5101 );
or ( n5104 , n5099 , n5102 , n5103 );
xor ( n5105 , n4880 , n4901 );
xor ( n5106 , n5105 , n4904 );
and ( n5107 , n5104 , n5106 );
xor ( n5108 , n4946 , n4948 );
xor ( n5109 , n5108 , n4951 );
and ( n5110 , n5106 , n5109 );
and ( n5111 , n5104 , n5109 );
or ( n5112 , n5107 , n5110 , n5111 );
and ( n5113 , n5086 , n5112 );
xor ( n5114 , n4936 , n4961 );
xor ( n5115 , n5114 , n4964 );
and ( n5116 , n5113 , n5115 );
xor ( n5117 , n4954 , n4955 );
xor ( n5118 , n5117 , n4958 );
xor ( n5119 , n5086 , n5112 );
and ( n5120 , n5118 , n5119 );
xor ( n5121 , n4974 , n4977 );
and ( n5122 , n1963 , n2666 );
and ( n5123 , n1869 , n2664 );
nor ( n5124 , n5122 , n5123 );
xnor ( n5125 , n5124 , n2587 );
and ( n5126 , n2611 , n2054 );
and ( n5127 , n2459 , n2052 );
nor ( n5128 , n5126 , n5127 );
xnor ( n5129 , n5128 , n1989 );
and ( n5130 , n5125 , n5129 );
and ( n5131 , n2969 , n1894 );
and ( n5132 , n2658 , n1892 );
nor ( n5133 , n5131 , n5132 );
xnor ( n5134 , n5133 , n1793 );
and ( n5135 , n5129 , n5134 );
and ( n5136 , n5125 , n5134 );
or ( n5137 , n5130 , n5135 , n5136 );
and ( n5138 , n5121 , n5137 );
and ( n5139 , n1438 , n3929 );
and ( n5140 , n1407 , n3926 );
nor ( n5141 , n5139 , n5140 );
xnor ( n5142 , n5141 , n3372 );
and ( n5143 , n3079 , n1692 );
and ( n5144 , n3019 , n1690 );
nor ( n5145 , n5143 , n5144 );
xnor ( n5146 , n5145 , n1670 );
and ( n5147 , n5142 , n5146 );
and ( n5148 , n3366 , n1604 );
and ( n5149 , n3415 , n1602 );
nor ( n5150 , n5148 , n5149 );
xnor ( n5151 , n5150 , n1549 );
and ( n5152 , n5146 , n5151 );
and ( n5153 , n5142 , n5151 );
or ( n5154 , n5147 , n5152 , n5153 );
and ( n5155 , n5137 , n5154 );
and ( n5156 , n5121 , n5154 );
or ( n5157 , n5138 , n5155 , n5156 );
and ( n5158 , n1610 , n3813 );
and ( n5159 , n1521 , n3811 );
nor ( n5160 , n5158 , n5159 );
xnor ( n5161 , n5160 , n3375 );
and ( n5162 , n1833 , n2940 );
and ( n5163 , n1759 , n2938 );
nor ( n5164 , n5162 , n5163 );
xnor ( n5165 , n5164 , n2868 );
and ( n5166 , n5161 , n5165 );
and ( n5167 , n5165 , n4975 );
and ( n5168 , n5161 , n4975 );
or ( n5169 , n5166 , n5167 , n5168 );
and ( n5170 , n1661 , n3227 );
and ( n5171 , n1624 , n3225 );
nor ( n5172 , n5170 , n5171 );
xnor ( n5173 , n5172 , n3168 );
and ( n5174 , n2182 , n2450 );
and ( n5175 , n2076 , n2448 );
nor ( n5176 , n5174 , n5175 );
xnor ( n5177 , n5176 , n2364 );
and ( n5178 , n5173 , n5177 );
and ( n5179 , n3882 , n1488 );
and ( n5180 , n3748 , n1486 );
nor ( n5181 , n5179 , n5180 );
xnor ( n5182 , n5181 , n1456 );
and ( n5183 , n5177 , n5182 );
and ( n5184 , n5173 , n5182 );
or ( n5185 , n5178 , n5183 , n5184 );
and ( n5186 , n5169 , n5185 );
xor ( n5187 , n5054 , n5058 );
xor ( n5188 , n5187 , n5063 );
and ( n5189 , n5185 , n5188 );
and ( n5190 , n5169 , n5188 );
or ( n5191 , n5186 , n5189 , n5190 );
and ( n5192 , n5157 , n5191 );
xor ( n5193 , n5002 , n5006 );
xor ( n5194 , n5193 , n5011 );
xor ( n5195 , n5018 , n5022 );
xor ( n5196 , n5195 , n5027 );
and ( n5197 , n5194 , n5196 );
xor ( n5198 , n5035 , n5039 );
xor ( n5199 , n5198 , n5044 );
and ( n5200 , n5196 , n5199 );
and ( n5201 , n5194 , n5199 );
or ( n5202 , n5197 , n5200 , n5201 );
and ( n5203 , n5191 , n5202 );
and ( n5204 , n5157 , n5202 );
or ( n5205 , n5192 , n5203 , n5204 );
xor ( n5206 , n5014 , n5030 );
xor ( n5207 , n5206 , n5047 );
xor ( n5208 , n5066 , n5068 );
xor ( n5209 , n5208 , n5071 );
and ( n5210 , n5207 , n5209 );
xor ( n5211 , n5088 , n5090 );
xor ( n5212 , n5211 , n5093 );
and ( n5213 , n5209 , n5212 );
and ( n5214 , n5207 , n5212 );
or ( n5215 , n5210 , n5213 , n5214 );
and ( n5216 , n5205 , n5215 );
xor ( n5217 , n5050 , n5074 );
xor ( n5218 , n5217 , n5077 );
and ( n5219 , n5215 , n5218 );
and ( n5220 , n5205 , n5218 );
or ( n5221 , n5216 , n5219 , n5220 );
xor ( n5222 , n4998 , n5080 );
xor ( n5223 , n5222 , n5083 );
and ( n5224 , n5221 , n5223 );
xor ( n5225 , n5104 , n5106 );
xor ( n5226 , n5225 , n5109 );
and ( n5227 , n5223 , n5226 );
and ( n5228 , n5221 , n5226 );
or ( n5229 , n5224 , n5227 , n5228 );
and ( n5230 , n5119 , n5229 );
and ( n5231 , n5118 , n5229 );
or ( n5232 , n5120 , n5230 , n5231 );
and ( n5233 , n5115 , n5232 );
and ( n5234 , n5113 , n5232 );
or ( n5235 , n5116 , n5233 , n5234 );
and ( n5236 , n4969 , n5235 );
and ( n5237 , n4967 , n5235 );
or ( n5238 , n4970 , n5236 , n5237 );
and ( n5239 , n4934 , n5238 );
xor ( n5240 , n4934 , n5238 );
xor ( n5241 , n4967 , n4969 );
xor ( n5242 , n5241 , n5235 );
xor ( n5243 , n5113 , n5115 );
xor ( n5244 , n5243 , n5232 );
xor ( n5245 , n5118 , n5119 );
xor ( n5246 , n5245 , n5229 );
xor ( n5247 , n5221 , n5223 );
xor ( n5248 , n5247 , n5226 );
and ( n5249 , n2076 , n2666 );
and ( n5250 , n1963 , n2664 );
nor ( n5251 , n5249 , n5250 );
xnor ( n5252 , n5251 , n2587 );
and ( n5253 , n3415 , n1692 );
and ( n5254 , n3079 , n1690 );
nor ( n5255 , n5253 , n5254 );
xnor ( n5256 , n5255 , n1670 );
and ( n5257 , n5252 , n5256 );
and ( n5258 , n3748 , n1604 );
and ( n5259 , n3366 , n1602 );
nor ( n5260 , n5258 , n5259 );
xnor ( n5261 , n5260 , n1549 );
and ( n5262 , n5256 , n5261 );
and ( n5263 , n5252 , n5261 );
or ( n5264 , n5257 , n5262 , n5263 );
and ( n5265 , n1624 , n3813 );
and ( n5266 , n1610 , n3811 );
nor ( n5267 , n5265 , n5266 );
xnor ( n5268 , n5267 , n3375 );
and ( n5269 , n3938 , n1486 );
not ( n5270 , n5269 );
and ( n5271 , n5270 , n1456 );
and ( n5272 , n5268 , n5271 );
and ( n5273 , n5264 , n5272 );
and ( n5274 , n2338 , n2221 );
and ( n5275 , n2263 , n2219 );
nor ( n5276 , n5274 , n5275 );
xnor ( n5277 , n5276 , n2138 );
and ( n5278 , n5272 , n5277 );
and ( n5279 , n5264 , n5277 );
or ( n5280 , n5273 , n5278 , n5279 );
xor ( n5281 , n5161 , n5165 );
xor ( n5282 , n5281 , n4975 );
xor ( n5283 , n5125 , n5129 );
xor ( n5284 , n5283 , n5134 );
and ( n5285 , n5282 , n5284 );
xor ( n5286 , n5142 , n5146 );
xor ( n5287 , n5286 , n5151 );
and ( n5288 , n5284 , n5287 );
and ( n5289 , n5282 , n5287 );
or ( n5290 , n5285 , n5288 , n5289 );
and ( n5291 , n5280 , n5290 );
xor ( n5292 , n5169 , n5185 );
xor ( n5293 , n5292 , n5188 );
and ( n5294 , n5290 , n5293 );
and ( n5295 , n5280 , n5293 );
or ( n5296 , n5291 , n5294 , n5295 );
and ( n5297 , n1521 , n3929 );
and ( n5298 , n1438 , n3926 );
nor ( n5299 , n5297 , n5298 );
xnor ( n5300 , n5299 , n3372 );
and ( n5301 , n1759 , n3227 );
and ( n5302 , n1661 , n3225 );
nor ( n5303 , n5301 , n5302 );
xnor ( n5304 , n5303 , n3168 );
and ( n5305 , n5300 , n5304 );
and ( n5306 , n3938 , n1488 );
and ( n5307 , n3882 , n1486 );
nor ( n5308 , n5306 , n5307 );
xnor ( n5309 , n5308 , n1456 );
and ( n5310 , n5304 , n5309 );
and ( n5311 , n5300 , n5309 );
or ( n5312 , n5305 , n5310 , n5311 );
and ( n5313 , n1869 , n2940 );
and ( n5314 , n1833 , n2938 );
nor ( n5315 , n5313 , n5314 );
xnor ( n5316 , n5315 , n2868 );
and ( n5317 , n2658 , n2054 );
and ( n5318 , n2611 , n2052 );
nor ( n5319 , n5317 , n5318 );
xnor ( n5320 , n5319 , n1989 );
and ( n5321 , n5316 , n5320 );
and ( n5322 , n3019 , n1894 );
and ( n5323 , n2969 , n1892 );
nor ( n5324 , n5322 , n5323 );
xnor ( n5325 , n5324 , n1793 );
and ( n5326 , n5320 , n5325 );
and ( n5327 , n5316 , n5325 );
or ( n5328 , n5321 , n5326 , n5327 );
and ( n5329 , n5312 , n5328 );
xor ( n5330 , n5173 , n5177 );
xor ( n5331 , n5330 , n5182 );
and ( n5332 , n5328 , n5331 );
and ( n5333 , n5312 , n5331 );
or ( n5334 , n5329 , n5332 , n5333 );
xor ( n5335 , n5121 , n5137 );
xor ( n5336 , n5335 , n5154 );
and ( n5337 , n5334 , n5336 );
xor ( n5338 , n5194 , n5196 );
xor ( n5339 , n5338 , n5199 );
and ( n5340 , n5336 , n5339 );
and ( n5341 , n5334 , n5339 );
or ( n5342 , n5337 , n5340 , n5341 );
and ( n5343 , n5296 , n5342 );
xor ( n5344 , n5157 , n5191 );
xor ( n5345 , n5344 , n5202 );
and ( n5346 , n5342 , n5345 );
and ( n5347 , n5296 , n5345 );
or ( n5348 , n5343 , n5346 , n5347 );
xor ( n5349 , n5096 , n5098 );
xor ( n5350 , n5349 , n5101 );
and ( n5351 , n5348 , n5350 );
xor ( n5352 , n5205 , n5215 );
xor ( n5353 , n5352 , n5218 );
and ( n5354 , n5350 , n5353 );
and ( n5355 , n5348 , n5353 );
or ( n5356 , n5351 , n5354 , n5355 );
and ( n5357 , n5248 , n5356 );
xor ( n5358 , n5248 , n5356 );
and ( n5359 , n1833 , n3227 );
and ( n5360 , n1759 , n3225 );
nor ( n5361 , n5359 , n5360 );
xnor ( n5362 , n5361 , n3168 );
and ( n5363 , n2338 , n2450 );
and ( n5364 , n2263 , n2448 );
nor ( n5365 , n5363 , n5364 );
xnor ( n5366 , n5365 , n2364 );
and ( n5367 , n5362 , n5366 );
and ( n5368 , n2611 , n2221 );
and ( n5369 , n2459 , n2219 );
nor ( n5370 , n5368 , n5369 );
xnor ( n5371 , n5370 , n2138 );
and ( n5372 , n5366 , n5371 );
and ( n5373 , n5362 , n5371 );
or ( n5374 , n5367 , n5372 , n5373 );
and ( n5375 , n1661 , n3813 );
and ( n5376 , n1624 , n3811 );
nor ( n5377 , n5375 , n5376 );
xnor ( n5378 , n5377 , n3375 );
and ( n5379 , n1963 , n2940 );
and ( n5380 , n1869 , n2938 );
nor ( n5381 , n5379 , n5380 );
xnor ( n5382 , n5381 , n2868 );
and ( n5383 , n5378 , n5382 );
and ( n5384 , n5382 , n5269 );
and ( n5385 , n5378 , n5269 );
or ( n5386 , n5383 , n5384 , n5385 );
and ( n5387 , n5374 , n5386 );
and ( n5388 , n1610 , n3929 );
and ( n5389 , n1521 , n3926 );
nor ( n5390 , n5388 , n5389 );
xnor ( n5391 , n5390 , n3372 );
and ( n5392 , n3366 , n1692 );
and ( n5393 , n3415 , n1690 );
nor ( n5394 , n5392 , n5393 );
xnor ( n5395 , n5394 , n1670 );
and ( n5396 , n5391 , n5395 );
and ( n5397 , n3882 , n1604 );
and ( n5398 , n3748 , n1602 );
nor ( n5399 , n5397 , n5398 );
xnor ( n5400 , n5399 , n1549 );
and ( n5401 , n5395 , n5400 );
and ( n5402 , n5391 , n5400 );
or ( n5403 , n5396 , n5401 , n5402 );
and ( n5404 , n5386 , n5403 );
and ( n5405 , n5374 , n5403 );
or ( n5406 , n5387 , n5404 , n5405 );
xor ( n5407 , n5268 , n5271 );
and ( n5408 , n2263 , n2450 );
and ( n5409 , n2182 , n2448 );
nor ( n5410 , n5408 , n5409 );
xnor ( n5411 , n5410 , n2364 );
and ( n5412 , n5407 , n5411 );
and ( n5413 , n2459 , n2221 );
and ( n5414 , n2338 , n2219 );
nor ( n5415 , n5413 , n5414 );
xnor ( n5416 , n5415 , n2138 );
and ( n5417 , n5411 , n5416 );
and ( n5418 , n5407 , n5416 );
or ( n5419 , n5412 , n5417 , n5418 );
and ( n5420 , n5406 , n5419 );
xor ( n5421 , n5264 , n5272 );
xor ( n5422 , n5421 , n5277 );
and ( n5423 , n5419 , n5422 );
and ( n5424 , n5406 , n5422 );
or ( n5425 , n5420 , n5423 , n5424 );
and ( n5426 , n2182 , n2666 );
and ( n5427 , n2076 , n2664 );
nor ( n5428 , n5426 , n5427 );
xnor ( n5429 , n5428 , n2587 );
and ( n5430 , n2969 , n2054 );
and ( n5431 , n2658 , n2052 );
nor ( n5432 , n5430 , n5431 );
xnor ( n5433 , n5432 , n1989 );
and ( n5434 , n5429 , n5433 );
and ( n5435 , n3079 , n1894 );
and ( n5436 , n3019 , n1892 );
nor ( n5437 , n5435 , n5436 );
xnor ( n5438 , n5437 , n1793 );
and ( n5439 , n5433 , n5438 );
and ( n5440 , n5429 , n5438 );
or ( n5441 , n5434 , n5439 , n5440 );
xor ( n5442 , n5300 , n5304 );
xor ( n5443 , n5442 , n5309 );
and ( n5444 , n5441 , n5443 );
xor ( n5445 , n5252 , n5256 );
xor ( n5446 , n5445 , n5261 );
and ( n5447 , n5443 , n5446 );
and ( n5448 , n5441 , n5446 );
or ( n5449 , n5444 , n5447 , n5448 );
xor ( n5450 , n5312 , n5328 );
xor ( n5451 , n5450 , n5331 );
and ( n5452 , n5449 , n5451 );
xor ( n5453 , n5282 , n5284 );
xor ( n5454 , n5453 , n5287 );
and ( n5455 , n5451 , n5454 );
and ( n5456 , n5449 , n5454 );
or ( n5457 , n5452 , n5455 , n5456 );
and ( n5458 , n5425 , n5457 );
xor ( n5459 , n5280 , n5290 );
xor ( n5460 , n5459 , n5293 );
and ( n5461 , n5457 , n5460 );
and ( n5462 , n5425 , n5460 );
or ( n5463 , n5458 , n5461 , n5462 );
xor ( n5464 , n5296 , n5342 );
xor ( n5465 , n5464 , n5345 );
and ( n5466 , n5463 , n5465 );
xor ( n5467 , n5207 , n5209 );
xor ( n5468 , n5467 , n5212 );
and ( n5469 , n5465 , n5468 );
and ( n5470 , n5463 , n5468 );
or ( n5471 , n5466 , n5469 , n5470 );
xor ( n5472 , n5348 , n5350 );
xor ( n5473 , n5472 , n5353 );
and ( n5474 , n5471 , n5473 );
xor ( n5475 , n5471 , n5473 );
xor ( n5476 , n5463 , n5465 );
xor ( n5477 , n5476 , n5468 );
and ( n5478 , n2263 , n2666 );
and ( n5479 , n2182 , n2664 );
nor ( n5480 , n5478 , n5479 );
xnor ( n5481 , n5480 , n2587 );
and ( n5482 , n3748 , n1692 );
and ( n5483 , n3366 , n1690 );
nor ( n5484 , n5482 , n5483 );
xnor ( n5485 , n5484 , n1670 );
and ( n5486 , n5481 , n5485 );
and ( n5487 , n3938 , n1604 );
and ( n5488 , n3882 , n1602 );
nor ( n5489 , n5487 , n5488 );
xnor ( n5490 , n5489 , n1549 );
and ( n5491 , n5485 , n5490 );
and ( n5492 , n5481 , n5490 );
or ( n5493 , n5486 , n5491 , n5492 );
and ( n5494 , n1624 , n3929 );
and ( n5495 , n1610 , n3926 );
nor ( n5496 , n5494 , n5495 );
xnor ( n5497 , n5496 , n3372 );
and ( n5498 , n1869 , n3227 );
and ( n5499 , n1833 , n3225 );
nor ( n5500 , n5498 , n5499 );
xnor ( n5501 , n5500 , n3168 );
and ( n5502 , n5497 , n5501 );
and ( n5503 , n2459 , n2450 );
and ( n5504 , n2338 , n2448 );
nor ( n5505 , n5503 , n5504 );
xnor ( n5506 , n5505 , n2364 );
and ( n5507 , n5501 , n5506 );
and ( n5508 , n5497 , n5506 );
or ( n5509 , n5502 , n5507 , n5508 );
and ( n5510 , n5493 , n5509 );
and ( n5511 , n1759 , n3813 );
and ( n5512 , n1661 , n3811 );
nor ( n5513 , n5511 , n5512 );
xnor ( n5514 , n5513 , n3375 );
and ( n5515 , n3938 , n1602 );
not ( n5516 , n5515 );
and ( n5517 , n5516 , n1549 );
and ( n5518 , n5514 , n5517 );
and ( n5519 , n5509 , n5518 );
and ( n5520 , n5493 , n5518 );
or ( n5521 , n5510 , n5519 , n5520 );
xor ( n5522 , n5316 , n5320 );
xor ( n5523 , n5522 , n5325 );
and ( n5524 , n5521 , n5523 );
xor ( n5525 , n5407 , n5411 );
xor ( n5526 , n5525 , n5416 );
and ( n5527 , n5523 , n5526 );
and ( n5528 , n5521 , n5526 );
or ( n5529 , n5524 , n5527 , n5528 );
and ( n5530 , n2076 , n2940 );
and ( n5531 , n1963 , n2938 );
nor ( n5532 , n5530 , n5531 );
xnor ( n5533 , n5532 , n2868 );
and ( n5534 , n3019 , n2054 );
and ( n5535 , n2969 , n2052 );
nor ( n5536 , n5534 , n5535 );
xnor ( n5537 , n5536 , n1989 );
and ( n5538 , n5533 , n5537 );
and ( n5539 , n3415 , n1894 );
and ( n5540 , n3079 , n1892 );
nor ( n5541 , n5539 , n5540 );
xnor ( n5542 , n5541 , n1793 );
and ( n5543 , n5537 , n5542 );
and ( n5544 , n5533 , n5542 );
or ( n5545 , n5538 , n5543 , n5544 );
xor ( n5546 , n5362 , n5366 );
xor ( n5547 , n5546 , n5371 );
and ( n5548 , n5545 , n5547 );
xor ( n5549 , n5429 , n5433 );
xor ( n5550 , n5549 , n5438 );
and ( n5551 , n5547 , n5550 );
and ( n5552 , n5545 , n5550 );
or ( n5553 , n5548 , n5551 , n5552 );
xor ( n5554 , n5374 , n5386 );
xor ( n5555 , n5554 , n5403 );
and ( n5556 , n5553 , n5555 );
xor ( n5557 , n5441 , n5443 );
xor ( n5558 , n5557 , n5446 );
and ( n5559 , n5555 , n5558 );
and ( n5560 , n5553 , n5558 );
or ( n5561 , n5556 , n5559 , n5560 );
and ( n5562 , n5529 , n5561 );
xor ( n5563 , n5406 , n5419 );
xor ( n5564 , n5563 , n5422 );
and ( n5565 , n5561 , n5564 );
and ( n5566 , n5529 , n5564 );
or ( n5567 , n5562 , n5565 , n5566 );
xor ( n5568 , n5334 , n5336 );
xor ( n5569 , n5568 , n5339 );
and ( n5570 , n5567 , n5569 );
xor ( n5571 , n5425 , n5457 );
xor ( n5572 , n5571 , n5460 );
and ( n5573 , n5569 , n5572 );
and ( n5574 , n5567 , n5572 );
or ( n5575 , n5570 , n5573 , n5574 );
and ( n5576 , n5477 , n5575 );
xor ( n5577 , n5477 , n5575 );
xor ( n5578 , n5567 , n5569 );
xor ( n5579 , n5578 , n5572 );
xor ( n5580 , n5514 , n5517 );
and ( n5581 , n1833 , n3813 );
and ( n5582 , n1759 , n3811 );
nor ( n5583 , n5581 , n5582 );
xnor ( n5584 , n5583 , n3375 );
and ( n5585 , n3079 , n2054 );
and ( n5586 , n3019 , n2052 );
nor ( n5587 , n5585 , n5586 );
xnor ( n5588 , n5587 , n1989 );
and ( n5589 , n5584 , n5588 );
and ( n5590 , n3366 , n1894 );
and ( n5591 , n3415 , n1892 );
nor ( n5592 , n5590 , n5591 );
xnor ( n5593 , n5592 , n1793 );
and ( n5594 , n5588 , n5593 );
and ( n5595 , n5584 , n5593 );
or ( n5596 , n5589 , n5594 , n5595 );
and ( n5597 , n5580 , n5596 );
and ( n5598 , n2658 , n2221 );
and ( n5599 , n2611 , n2219 );
nor ( n5600 , n5598 , n5599 );
xnor ( n5601 , n5600 , n2138 );
and ( n5602 , n5596 , n5601 );
and ( n5603 , n5580 , n5601 );
or ( n5604 , n5597 , n5602 , n5603 );
xor ( n5605 , n5378 , n5382 );
xor ( n5606 , n5605 , n5269 );
and ( n5607 , n5604 , n5606 );
xor ( n5608 , n5391 , n5395 );
xor ( n5609 , n5608 , n5400 );
and ( n5610 , n5606 , n5609 );
and ( n5611 , n5604 , n5609 );
or ( n5612 , n5607 , n5610 , n5611 );
xor ( n5613 , n5521 , n5523 );
xor ( n5614 , n5613 , n5526 );
and ( n5615 , n5612 , n5614 );
xor ( n5616 , n5553 , n5555 );
xor ( n5617 , n5616 , n5558 );
and ( n5618 , n5614 , n5617 );
and ( n5619 , n5612 , n5617 );
or ( n5620 , n5615 , n5618 , n5619 );
xor ( n5621 , n5449 , n5451 );
xor ( n5622 , n5621 , n5454 );
and ( n5623 , n5620 , n5622 );
xor ( n5624 , n5529 , n5561 );
xor ( n5625 , n5624 , n5564 );
and ( n5626 , n5622 , n5625 );
and ( n5627 , n5620 , n5625 );
or ( n5628 , n5623 , n5626 , n5627 );
and ( n5629 , n5579 , n5628 );
xor ( n5630 , n5579 , n5628 );
xor ( n5631 , n5620 , n5622 );
xor ( n5632 , n5631 , n5625 );
and ( n5633 , n1661 , n3929 );
and ( n5634 , n1624 , n3926 );
nor ( n5635 , n5633 , n5634 );
xnor ( n5636 , n5635 , n3372 );
and ( n5637 , n2182 , n2940 );
and ( n5638 , n2076 , n2938 );
nor ( n5639 , n5637 , n5638 );
xnor ( n5640 , n5639 , n2868 );
and ( n5641 , n5636 , n5640 );
and ( n5642 , n5640 , n5515 );
and ( n5643 , n5636 , n5515 );
or ( n5644 , n5641 , n5642 , n5643 );
and ( n5645 , n1963 , n3227 );
and ( n5646 , n1869 , n3225 );
nor ( n5647 , n5645 , n5646 );
xnor ( n5648 , n5647 , n3168 );
and ( n5649 , n2338 , n2666 );
and ( n5650 , n2263 , n2664 );
nor ( n5651 , n5649 , n5650 );
xnor ( n5652 , n5651 , n2587 );
and ( n5653 , n5648 , n5652 );
and ( n5654 , n3882 , n1692 );
and ( n5655 , n3748 , n1690 );
nor ( n5656 , n5654 , n5655 );
xnor ( n5657 , n5656 , n1670 );
and ( n5658 , n5652 , n5657 );
and ( n5659 , n5648 , n5657 );
or ( n5660 , n5653 , n5658 , n5659 );
and ( n5661 , n5644 , n5660 );
xor ( n5662 , n5497 , n5501 );
xor ( n5663 , n5662 , n5506 );
and ( n5664 , n5660 , n5663 );
and ( n5665 , n5644 , n5663 );
or ( n5666 , n5661 , n5664 , n5665 );
and ( n5667 , n1759 , n3929 );
and ( n5668 , n1661 , n3926 );
nor ( n5669 , n5667 , n5668 );
xnor ( n5670 , n5669 , n3372 );
and ( n5671 , n3938 , n1690 );
not ( n5672 , n5671 );
and ( n5673 , n5672 , n1670 );
and ( n5674 , n5670 , n5673 );
and ( n5675 , n2611 , n2450 );
and ( n5676 , n2459 , n2448 );
nor ( n5677 , n5675 , n5676 );
xnor ( n5678 , n5677 , n2364 );
and ( n5679 , n5674 , n5678 );
and ( n5680 , n2969 , n2221 );
and ( n5681 , n2658 , n2219 );
nor ( n5682 , n5680 , n5681 );
xnor ( n5683 , n5682 , n2138 );
and ( n5684 , n5678 , n5683 );
and ( n5685 , n5674 , n5683 );
or ( n5686 , n5679 , n5684 , n5685 );
xor ( n5687 , n5481 , n5485 );
xor ( n5688 , n5687 , n5490 );
and ( n5689 , n5686 , n5688 );
xor ( n5690 , n5533 , n5537 );
xor ( n5691 , n5690 , n5542 );
and ( n5692 , n5688 , n5691 );
and ( n5693 , n5686 , n5691 );
or ( n5694 , n5689 , n5692 , n5693 );
and ( n5695 , n5666 , n5694 );
xor ( n5696 , n5493 , n5509 );
xor ( n5697 , n5696 , n5518 );
and ( n5698 , n5694 , n5697 );
and ( n5699 , n5666 , n5697 );
or ( n5700 , n5695 , n5698 , n5699 );
and ( n5701 , n2263 , n2940 );
and ( n5702 , n2182 , n2938 );
nor ( n5703 , n5701 , n5702 );
xnor ( n5704 , n5703 , n2868 );
and ( n5705 , n3415 , n2054 );
and ( n5706 , n3079 , n2052 );
nor ( n5707 , n5705 , n5706 );
xnor ( n5708 , n5707 , n1989 );
and ( n5709 , n5704 , n5708 );
and ( n5710 , n3748 , n1894 );
and ( n5711 , n3366 , n1892 );
nor ( n5712 , n5710 , n5711 );
xnor ( n5713 , n5712 , n1793 );
and ( n5714 , n5708 , n5713 );
and ( n5715 , n5704 , n5713 );
or ( n5716 , n5709 , n5714 , n5715 );
and ( n5717 , n2076 , n3227 );
and ( n5718 , n1963 , n3225 );
nor ( n5719 , n5717 , n5718 );
xnor ( n5720 , n5719 , n3168 );
and ( n5721 , n2658 , n2450 );
and ( n5722 , n2611 , n2448 );
nor ( n5723 , n5721 , n5722 );
xnor ( n5724 , n5723 , n2364 );
and ( n5725 , n5720 , n5724 );
and ( n5726 , n3019 , n2221 );
and ( n5727 , n2969 , n2219 );
nor ( n5728 , n5726 , n5727 );
xnor ( n5729 , n5728 , n2138 );
and ( n5730 , n5724 , n5729 );
and ( n5731 , n5720 , n5729 );
or ( n5732 , n5725 , n5730 , n5731 );
and ( n5733 , n5716 , n5732 );
and ( n5734 , n1869 , n3813 );
and ( n5735 , n1833 , n3811 );
nor ( n5736 , n5734 , n5735 );
xnor ( n5737 , n5736 , n3375 );
and ( n5738 , n2459 , n2666 );
and ( n5739 , n2338 , n2664 );
nor ( n5740 , n5738 , n5739 );
xnor ( n5741 , n5740 , n2587 );
and ( n5742 , n5737 , n5741 );
and ( n5743 , n3938 , n1692 );
and ( n5744 , n3882 , n1690 );
nor ( n5745 , n5743 , n5744 );
xnor ( n5746 , n5745 , n1670 );
and ( n5747 , n5741 , n5746 );
and ( n5748 , n5737 , n5746 );
or ( n5749 , n5742 , n5747 , n5748 );
and ( n5750 , n5732 , n5749 );
and ( n5751 , n5716 , n5749 );
or ( n5752 , n5733 , n5750 , n5751 );
xor ( n5753 , n5580 , n5596 );
xor ( n5754 , n5753 , n5601 );
and ( n5755 , n5752 , n5754 );
xor ( n5756 , n5644 , n5660 );
xor ( n5757 , n5756 , n5663 );
and ( n5758 , n5754 , n5757 );
and ( n5759 , n5752 , n5757 );
or ( n5760 , n5755 , n5758 , n5759 );
xor ( n5761 , n5545 , n5547 );
xor ( n5762 , n5761 , n5550 );
and ( n5763 , n5760 , n5762 );
xor ( n5764 , n5604 , n5606 );
xor ( n5765 , n5764 , n5609 );
and ( n5766 , n5762 , n5765 );
and ( n5767 , n5760 , n5765 );
or ( n5768 , n5763 , n5766 , n5767 );
and ( n5769 , n5700 , n5768 );
xor ( n5770 , n5612 , n5614 );
xor ( n5771 , n5770 , n5617 );
and ( n5772 , n5768 , n5771 );
and ( n5773 , n5700 , n5771 );
or ( n5774 , n5769 , n5772 , n5773 );
and ( n5775 , n5632 , n5774 );
xor ( n5776 , n5632 , n5774 );
xor ( n5777 , n5700 , n5768 );
xor ( n5778 , n5777 , n5771 );
xor ( n5779 , n5636 , n5640 );
xor ( n5780 , n5779 , n5515 );
xor ( n5781 , n5648 , n5652 );
xor ( n5782 , n5781 , n5657 );
and ( n5783 , n5780 , n5782 );
xor ( n5784 , n5584 , n5588 );
xor ( n5785 , n5784 , n5593 );
and ( n5786 , n5782 , n5785 );
and ( n5787 , n5780 , n5785 );
or ( n5788 , n5783 , n5786 , n5787 );
xor ( n5789 , n5686 , n5688 );
xor ( n5790 , n5789 , n5691 );
and ( n5791 , n5788 , n5790 );
xor ( n5792 , n5752 , n5754 );
xor ( n5793 , n5792 , n5757 );
and ( n5794 , n5790 , n5793 );
and ( n5795 , n5788 , n5793 );
or ( n5796 , n5791 , n5794 , n5795 );
xor ( n5797 , n5666 , n5694 );
xor ( n5798 , n5797 , n5697 );
and ( n5799 , n5796 , n5798 );
xor ( n5800 , n5760 , n5762 );
xor ( n5801 , n5800 , n5765 );
and ( n5802 , n5798 , n5801 );
and ( n5803 , n5796 , n5801 );
or ( n5804 , n5799 , n5802 , n5803 );
and ( n5805 , n5778 , n5804 );
xor ( n5806 , n5778 , n5804 );
xor ( n5807 , n5796 , n5798 );
xor ( n5808 , n5807 , n5801 );
xor ( n5809 , n5670 , n5673 );
and ( n5810 , n1963 , n3813 );
and ( n5811 , n1869 , n3811 );
nor ( n5812 , n5810 , n5811 );
xnor ( n5813 , n5812 , n3375 );
and ( n5814 , n3366 , n2054 );
and ( n5815 , n3415 , n2052 );
nor ( n5816 , n5814 , n5815 );
xnor ( n5817 , n5816 , n1989 );
and ( n5818 , n5813 , n5817 );
and ( n5819 , n3882 , n1894 );
and ( n5820 , n3748 , n1892 );
nor ( n5821 , n5819 , n5820 );
xnor ( n5822 , n5821 , n1793 );
and ( n5823 , n5817 , n5822 );
and ( n5824 , n5813 , n5822 );
or ( n5825 , n5818 , n5823 , n5824 );
and ( n5826 , n5809 , n5825 );
and ( n5827 , n1833 , n3929 );
and ( n5828 , n1759 , n3926 );
nor ( n5829 , n5827 , n5828 );
xnor ( n5830 , n5829 , n3372 );
and ( n5831 , n2338 , n2940 );
and ( n5832 , n2263 , n2938 );
nor ( n5833 , n5831 , n5832 );
xnor ( n5834 , n5833 , n2868 );
and ( n5835 , n5830 , n5834 );
and ( n5836 , n5834 , n5671 );
and ( n5837 , n5830 , n5671 );
or ( n5838 , n5835 , n5836 , n5837 );
and ( n5839 , n5825 , n5838 );
and ( n5840 , n5809 , n5838 );
or ( n5841 , n5826 , n5839 , n5840 );
and ( n5842 , n2182 , n3227 );
and ( n5843 , n2076 , n3225 );
nor ( n5844 , n5842 , n5843 );
xnor ( n5845 , n5844 , n3168 );
and ( n5846 , n2611 , n2666 );
and ( n5847 , n2459 , n2664 );
nor ( n5848 , n5846 , n5847 );
xnor ( n5849 , n5848 , n2587 );
and ( n5850 , n5845 , n5849 );
and ( n5851 , n2969 , n2450 );
and ( n5852 , n2658 , n2448 );
nor ( n5853 , n5851 , n5852 );
xnor ( n5854 , n5853 , n2364 );
and ( n5855 , n5849 , n5854 );
and ( n5856 , n5845 , n5854 );
or ( n5857 , n5850 , n5855 , n5856 );
xor ( n5858 , n5704 , n5708 );
xor ( n5859 , n5858 , n5713 );
and ( n5860 , n5857 , n5859 );
xor ( n5861 , n5720 , n5724 );
xor ( n5862 , n5861 , n5729 );
and ( n5863 , n5859 , n5862 );
and ( n5864 , n5857 , n5862 );
or ( n5865 , n5860 , n5863 , n5864 );
and ( n5866 , n5841 , n5865 );
xor ( n5867 , n5674 , n5678 );
xor ( n5868 , n5867 , n5683 );
and ( n5869 , n5865 , n5868 );
and ( n5870 , n5841 , n5868 );
or ( n5871 , n5866 , n5869 , n5870 );
xor ( n5872 , n5716 , n5732 );
xor ( n5873 , n5872 , n5749 );
xor ( n5874 , n5780 , n5782 );
xor ( n5875 , n5874 , n5785 );
and ( n5876 , n5873 , n5875 );
xor ( n5877 , n5841 , n5865 );
xor ( n5878 , n5877 , n5868 );
and ( n5879 , n5875 , n5878 );
and ( n5880 , n5873 , n5878 );
or ( n5881 , n5876 , n5879 , n5880 );
and ( n5882 , n5871 , n5881 );
xor ( n5883 , n5788 , n5790 );
xor ( n5884 , n5883 , n5793 );
and ( n5885 , n5881 , n5884 );
and ( n5886 , n5871 , n5884 );
or ( n5887 , n5882 , n5885 , n5886 );
and ( n5888 , n5808 , n5887 );
xor ( n5889 , n5808 , n5887 );
xor ( n5890 , n5871 , n5881 );
xor ( n5891 , n5890 , n5884 );
and ( n5892 , n2459 , n2940 );
and ( n5893 , n2338 , n2938 );
nor ( n5894 , n5892 , n5893 );
xnor ( n5895 , n5894 , n2868 );
and ( n5896 , n3748 , n2054 );
and ( n5897 , n3366 , n2052 );
nor ( n5898 , n5896 , n5897 );
xnor ( n5899 , n5898 , n1989 );
and ( n5900 , n5895 , n5899 );
and ( n5901 , n3938 , n1894 );
and ( n5902 , n3882 , n1892 );
nor ( n5903 , n5901 , n5902 );
xnor ( n5904 , n5903 , n1793 );
and ( n5905 , n5899 , n5904 );
and ( n5906 , n5895 , n5904 );
or ( n5907 , n5900 , n5905 , n5906 );
and ( n5908 , n1869 , n3929 );
and ( n5909 , n1833 , n3926 );
nor ( n5910 , n5908 , n5909 );
xnor ( n5911 , n5910 , n3372 );
and ( n5912 , n3938 , n1892 );
not ( n5913 , n5912 );
and ( n5914 , n5913 , n1793 );
and ( n5915 , n5911 , n5914 );
and ( n5916 , n5907 , n5915 );
and ( n5917 , n3079 , n2221 );
and ( n5918 , n3019 , n2219 );
nor ( n5919 , n5917 , n5918 );
xnor ( n5920 , n5919 , n2138 );
and ( n5921 , n5915 , n5920 );
and ( n5922 , n5907 , n5920 );
or ( n5923 , n5916 , n5921 , n5922 );
xor ( n5924 , n5737 , n5741 );
xor ( n5925 , n5924 , n5746 );
and ( n5926 , n5923 , n5925 );
xor ( n5927 , n5809 , n5825 );
xor ( n5928 , n5927 , n5838 );
and ( n5929 , n5925 , n5928 );
and ( n5930 , n5923 , n5928 );
or ( n5931 , n5926 , n5929 , n5930 );
and ( n5932 , n2076 , n3813 );
and ( n5933 , n1963 , n3811 );
nor ( n5934 , n5932 , n5933 );
xnor ( n5935 , n5934 , n3375 );
and ( n5936 , n2263 , n3227 );
and ( n5937 , n2182 , n3225 );
nor ( n5938 , n5936 , n5937 );
xnor ( n5939 , n5938 , n3168 );
and ( n5940 , n5935 , n5939 );
and ( n5941 , n2658 , n2666 );
and ( n5942 , n2611 , n2664 );
nor ( n5943 , n5941 , n5942 );
xnor ( n5944 , n5943 , n2587 );
and ( n5945 , n5939 , n5944 );
and ( n5946 , n5935 , n5944 );
or ( n5947 , n5940 , n5945 , n5946 );
xor ( n5948 , n5830 , n5834 );
xor ( n5949 , n5948 , n5671 );
and ( n5950 , n5947 , n5949 );
xor ( n5951 , n5845 , n5849 );
xor ( n5952 , n5951 , n5854 );
and ( n5953 , n5949 , n5952 );
and ( n5954 , n5947 , n5952 );
or ( n5955 , n5950 , n5953 , n5954 );
xor ( n5956 , n5911 , n5914 );
and ( n5957 , n3019 , n2450 );
and ( n5958 , n2969 , n2448 );
nor ( n5959 , n5957 , n5958 );
xnor ( n5960 , n5959 , n2364 );
and ( n5961 , n5956 , n5960 );
and ( n5962 , n3415 , n2221 );
and ( n5963 , n3079 , n2219 );
nor ( n5964 , n5962 , n5963 );
xnor ( n5965 , n5964 , n2138 );
and ( n5966 , n5960 , n5965 );
and ( n5967 , n5956 , n5965 );
or ( n5968 , n5961 , n5966 , n5967 );
xor ( n5969 , n5813 , n5817 );
xor ( n5970 , n5969 , n5822 );
and ( n5971 , n5968 , n5970 );
xor ( n5972 , n5907 , n5915 );
xor ( n5973 , n5972 , n5920 );
and ( n5974 , n5970 , n5973 );
and ( n5975 , n5968 , n5973 );
or ( n5976 , n5971 , n5974 , n5975 );
and ( n5977 , n5955 , n5976 );
xor ( n5978 , n5857 , n5859 );
xor ( n5979 , n5978 , n5862 );
and ( n5980 , n5976 , n5979 );
and ( n5981 , n5955 , n5979 );
or ( n5982 , n5977 , n5980 , n5981 );
and ( n5983 , n5931 , n5982 );
xor ( n5984 , n5873 , n5875 );
xor ( n5985 , n5984 , n5878 );
and ( n5986 , n5982 , n5985 );
and ( n5987 , n5931 , n5985 );
or ( n5988 , n5983 , n5986 , n5987 );
and ( n5989 , n5891 , n5988 );
xor ( n5990 , n5891 , n5988 );
xor ( n5991 , n5931 , n5982 );
xor ( n5992 , n5991 , n5985 );
and ( n5993 , n2611 , n2940 );
and ( n5994 , n2459 , n2938 );
nor ( n5995 , n5993 , n5994 );
xnor ( n5996 , n5995 , n2868 );
and ( n5997 , n2969 , n2666 );
and ( n5998 , n2658 , n2664 );
nor ( n5999 , n5997 , n5998 );
xnor ( n6000 , n5999 , n2587 );
and ( n6001 , n5996 , n6000 );
and ( n6002 , n3882 , n2054 );
and ( n6003 , n3748 , n2052 );
nor ( n6004 , n6002 , n6003 );
xnor ( n6005 , n6004 , n1989 );
and ( n6006 , n6000 , n6005 );
and ( n6007 , n5996 , n6005 );
or ( n6008 , n6001 , n6006 , n6007 );
and ( n6009 , n1963 , n3929 );
and ( n6010 , n1869 , n3926 );
nor ( n6011 , n6009 , n6010 );
xnor ( n6012 , n6011 , n3372 );
and ( n6013 , n2182 , n3813 );
and ( n6014 , n2076 , n3811 );
nor ( n6015 , n6013 , n6014 );
xnor ( n6016 , n6015 , n3375 );
and ( n6017 , n6012 , n6016 );
and ( n6018 , n6016 , n5912 );
and ( n6019 , n6012 , n5912 );
or ( n6020 , n6017 , n6018 , n6019 );
and ( n6021 , n6008 , n6020 );
and ( n6022 , n2338 , n3227 );
and ( n6023 , n2263 , n3225 );
nor ( n6024 , n6022 , n6023 );
xnor ( n6025 , n6024 , n3168 );
and ( n6026 , n3079 , n2450 );
and ( n6027 , n3019 , n2448 );
nor ( n6028 , n6026 , n6027 );
xnor ( n6029 , n6028 , n2364 );
and ( n6030 , n6025 , n6029 );
and ( n6031 , n3366 , n2221 );
and ( n6032 , n3415 , n2219 );
nor ( n6033 , n6031 , n6032 );
xnor ( n6034 , n6033 , n2138 );
and ( n6035 , n6029 , n6034 );
and ( n6036 , n6025 , n6034 );
or ( n6037 , n6030 , n6035 , n6036 );
and ( n6038 , n6020 , n6037 );
and ( n6039 , n6008 , n6037 );
or ( n6040 , n6021 , n6038 , n6039 );
xor ( n6041 , n5895 , n5899 );
xor ( n6042 , n6041 , n5904 );
xor ( n6043 , n5935 , n5939 );
xor ( n6044 , n6043 , n5944 );
and ( n6045 , n6042 , n6044 );
xor ( n6046 , n5956 , n5960 );
xor ( n6047 , n6046 , n5965 );
and ( n6048 , n6044 , n6047 );
and ( n6049 , n6042 , n6047 );
or ( n6050 , n6045 , n6048 , n6049 );
and ( n6051 , n6040 , n6050 );
xor ( n6052 , n5947 , n5949 );
xor ( n6053 , n6052 , n5952 );
and ( n6054 , n6050 , n6053 );
and ( n6055 , n6040 , n6053 );
or ( n6056 , n6051 , n6054 , n6055 );
xor ( n6057 , n5923 , n5925 );
xor ( n6058 , n6057 , n5928 );
and ( n6059 , n6056 , n6058 );
xor ( n6060 , n5955 , n5976 );
xor ( n6061 , n6060 , n5979 );
and ( n6062 , n6058 , n6061 );
and ( n6063 , n6056 , n6061 );
or ( n6064 , n6059 , n6062 , n6063 );
and ( n6065 , n5992 , n6064 );
xor ( n6066 , n5992 , n6064 );
xor ( n6067 , n6056 , n6058 );
xor ( n6068 , n6067 , n6061 );
and ( n6069 , n2263 , n3813 );
and ( n6070 , n2182 , n3811 );
nor ( n6071 , n6069 , n6070 );
xnor ( n6072 , n6071 , n3375 );
and ( n6073 , n2658 , n2940 );
and ( n6074 , n2611 , n2938 );
nor ( n6075 , n6073 , n6074 );
xnor ( n6076 , n6075 , n2868 );
and ( n6077 , n6072 , n6076 );
and ( n6078 , n3938 , n2054 );
and ( n6079 , n3882 , n2052 );
nor ( n6080 , n6078 , n6079 );
xnor ( n6081 , n6080 , n1989 );
and ( n6082 , n6076 , n6081 );
and ( n6083 , n6072 , n6081 );
or ( n6084 , n6077 , n6082 , n6083 );
and ( n6085 , n2459 , n3227 );
and ( n6086 , n2338 , n3225 );
nor ( n6087 , n6085 , n6086 );
xnor ( n6088 , n6087 , n3168 );
and ( n6089 , n3019 , n2666 );
and ( n6090 , n2969 , n2664 );
nor ( n6091 , n6089 , n6090 );
xnor ( n6092 , n6091 , n2587 );
and ( n6093 , n6088 , n6092 );
and ( n6094 , n3415 , n2450 );
and ( n6095 , n3079 , n2448 );
nor ( n6096 , n6094 , n6095 );
xnor ( n6097 , n6096 , n2364 );
and ( n6098 , n6092 , n6097 );
and ( n6099 , n6088 , n6097 );
or ( n6100 , n6093 , n6098 , n6099 );
and ( n6101 , n6084 , n6100 );
and ( n6102 , n2076 , n3929 );
and ( n6103 , n1963 , n3926 );
nor ( n6104 , n6102 , n6103 );
xnor ( n6105 , n6104 , n3372 );
and ( n6106 , n3938 , n2052 );
not ( n6107 , n6106 );
and ( n6108 , n6107 , n1989 );
and ( n6109 , n6105 , n6108 );
and ( n6110 , n6100 , n6109 );
and ( n6111 , n6084 , n6109 );
or ( n6112 , n6101 , n6110 , n6111 );
xor ( n6113 , n5996 , n6000 );
xor ( n6114 , n6113 , n6005 );
xor ( n6115 , n6012 , n6016 );
xor ( n6116 , n6115 , n5912 );
and ( n6117 , n6114 , n6116 );
xor ( n6118 , n6025 , n6029 );
xor ( n6119 , n6118 , n6034 );
and ( n6120 , n6116 , n6119 );
and ( n6121 , n6114 , n6119 );
or ( n6122 , n6117 , n6120 , n6121 );
and ( n6123 , n6112 , n6122 );
xor ( n6124 , n6008 , n6020 );
xor ( n6125 , n6124 , n6037 );
and ( n6126 , n6122 , n6125 );
and ( n6127 , n6112 , n6125 );
or ( n6128 , n6123 , n6126 , n6127 );
xor ( n6129 , n5968 , n5970 );
xor ( n6130 , n6129 , n5973 );
and ( n6131 , n6128 , n6130 );
xor ( n6132 , n6040 , n6050 );
xor ( n6133 , n6132 , n6053 );
and ( n6134 , n6130 , n6133 );
and ( n6135 , n6128 , n6133 );
or ( n6136 , n6131 , n6134 , n6135 );
and ( n6137 , n6068 , n6136 );
xor ( n6138 , n6068 , n6136 );
xor ( n6139 , n6105 , n6108 );
and ( n6140 , n2182 , n3929 );
and ( n6141 , n2076 , n3926 );
nor ( n6142 , n6140 , n6141 );
xnor ( n6143 , n6142 , n3372 );
and ( n6144 , n2338 , n3813 );
and ( n6145 , n2263 , n3811 );
nor ( n6146 , n6144 , n6145 );
xnor ( n6147 , n6146 , n3375 );
and ( n6148 , n6143 , n6147 );
and ( n6149 , n6147 , n6106 );
and ( n6150 , n6143 , n6106 );
or ( n6151 , n6148 , n6149 , n6150 );
and ( n6152 , n6139 , n6151 );
and ( n6153 , n3748 , n2221 );
and ( n6154 , n3366 , n2219 );
nor ( n6155 , n6153 , n6154 );
xnor ( n6156 , n6155 , n2138 );
and ( n6157 , n6151 , n6156 );
and ( n6158 , n6139 , n6156 );
or ( n6159 , n6152 , n6157 , n6158 );
and ( n6160 , n2611 , n3227 );
and ( n6161 , n2459 , n3225 );
nor ( n6162 , n6160 , n6161 );
xnor ( n6163 , n6162 , n3168 );
and ( n6164 , n2969 , n2940 );
and ( n6165 , n2658 , n2938 );
nor ( n6166 , n6164 , n6165 );
xnor ( n6167 , n6166 , n2868 );
and ( n6168 , n6163 , n6167 );
and ( n6169 , n3079 , n2666 );
and ( n6170 , n3019 , n2664 );
nor ( n6171 , n6169 , n6170 );
xnor ( n6172 , n6171 , n2587 );
and ( n6173 , n6167 , n6172 );
and ( n6174 , n6163 , n6172 );
or ( n6175 , n6168 , n6173 , n6174 );
xor ( n6176 , n6072 , n6076 );
xor ( n6177 , n6176 , n6081 );
and ( n6178 , n6175 , n6177 );
xor ( n6179 , n6088 , n6092 );
xor ( n6180 , n6179 , n6097 );
and ( n6181 , n6177 , n6180 );
and ( n6182 , n6175 , n6180 );
or ( n6183 , n6178 , n6181 , n6182 );
and ( n6184 , n6159 , n6183 );
xor ( n6185 , n6084 , n6100 );
xor ( n6186 , n6185 , n6109 );
and ( n6187 , n6183 , n6186 );
and ( n6188 , n6159 , n6186 );
or ( n6189 , n6184 , n6187 , n6188 );
xor ( n6190 , n6042 , n6044 );
xor ( n6191 , n6190 , n6047 );
and ( n6192 , n6189 , n6191 );
xor ( n6193 , n6112 , n6122 );
xor ( n6194 , n6193 , n6125 );
and ( n6195 , n6191 , n6194 );
and ( n6196 , n6189 , n6194 );
or ( n6197 , n6192 , n6195 , n6196 );
xor ( n6198 , n6128 , n6130 );
xor ( n6199 , n6198 , n6133 );
and ( n6200 , n6197 , n6199 );
xor ( n6201 , n6197 , n6199 );
xor ( n6202 , n6189 , n6191 );
xor ( n6203 , n6202 , n6194 );
and ( n6204 , n2263 , n3929 );
and ( n6205 , n2182 , n3926 );
nor ( n6206 , n6204 , n6205 );
xnor ( n6207 , n6206 , n3372 );
and ( n6208 , n3938 , n2219 );
not ( n6209 , n6208 );
and ( n6210 , n6209 , n2138 );
and ( n6211 , n6207 , n6210 );
and ( n6212 , n3366 , n2450 );
and ( n6213 , n3415 , n2448 );
nor ( n6214 , n6212 , n6213 );
xnor ( n6215 , n6214 , n2364 );
and ( n6216 , n6211 , n6215 );
and ( n6217 , n3882 , n2221 );
and ( n6218 , n3748 , n2219 );
nor ( n6219 , n6217 , n6218 );
xnor ( n6220 , n6219 , n2138 );
and ( n6221 , n6215 , n6220 );
and ( n6222 , n6211 , n6220 );
or ( n6223 , n6216 , n6221 , n6222 );
and ( n6224 , n2459 , n3813 );
and ( n6225 , n2338 , n3811 );
nor ( n6226 , n6224 , n6225 );
xnor ( n6227 , n6226 , n3375 );
and ( n6228 , n3019 , n2940 );
and ( n6229 , n2969 , n2938 );
nor ( n6230 , n6228 , n6229 );
xnor ( n6231 , n6230 , n2868 );
and ( n6232 , n6227 , n6231 );
and ( n6233 , n3415 , n2666 );
and ( n6234 , n3079 , n2664 );
nor ( n6235 , n6233 , n6234 );
xnor ( n6236 , n6235 , n2587 );
and ( n6237 , n6231 , n6236 );
and ( n6238 , n6227 , n6236 );
or ( n6239 , n6232 , n6237 , n6238 );
and ( n6240 , n2658 , n3227 );
and ( n6241 , n2611 , n3225 );
nor ( n6242 , n6240 , n6241 );
xnor ( n6243 , n6242 , n3168 );
and ( n6244 , n3748 , n2450 );
and ( n6245 , n3366 , n2448 );
nor ( n6246 , n6244 , n6245 );
xnor ( n6247 , n6246 , n2364 );
and ( n6248 , n6243 , n6247 );
and ( n6249 , n3938 , n2221 );
and ( n6250 , n3882 , n2219 );
nor ( n6251 , n6249 , n6250 );
xnor ( n6252 , n6251 , n2138 );
and ( n6253 , n6247 , n6252 );
and ( n6254 , n6243 , n6252 );
or ( n6255 , n6248 , n6253 , n6254 );
and ( n6256 , n6239 , n6255 );
xor ( n6257 , n6143 , n6147 );
xor ( n6258 , n6257 , n6106 );
and ( n6259 , n6255 , n6258 );
and ( n6260 , n6239 , n6258 );
or ( n6261 , n6256 , n6259 , n6260 );
and ( n6262 , n6223 , n6261 );
xor ( n6263 , n6139 , n6151 );
xor ( n6264 , n6263 , n6156 );
and ( n6265 , n6261 , n6264 );
and ( n6266 , n6223 , n6264 );
or ( n6267 , n6262 , n6265 , n6266 );
xor ( n6268 , n6114 , n6116 );
xor ( n6269 , n6268 , n6119 );
and ( n6270 , n6267 , n6269 );
xor ( n6271 , n6159 , n6183 );
xor ( n6272 , n6271 , n6186 );
and ( n6273 , n6269 , n6272 );
and ( n6274 , n6267 , n6272 );
or ( n6275 , n6270 , n6273 , n6274 );
and ( n6276 , n6203 , n6275 );
xor ( n6277 , n6203 , n6275 );
xor ( n6278 , n6267 , n6269 );
xor ( n6279 , n6278 , n6272 );
xor ( n6280 , n6207 , n6210 );
and ( n6281 , n2611 , n3813 );
and ( n6282 , n2459 , n3811 );
nor ( n6283 , n6281 , n6282 );
xnor ( n6284 , n6283 , n3375 );
and ( n6285 , n3079 , n2940 );
and ( n6286 , n3019 , n2938 );
nor ( n6287 , n6285 , n6286 );
xnor ( n6288 , n6287 , n2868 );
and ( n6289 , n6284 , n6288 );
and ( n6290 , n6288 , n6208 );
and ( n6291 , n6284 , n6208 );
or ( n6292 , n6289 , n6290 , n6291 );
and ( n6293 , n6280 , n6292 );
and ( n6294 , n2338 , n3929 );
and ( n6295 , n2263 , n3926 );
nor ( n6296 , n6294 , n6295 );
xnor ( n6297 , n6296 , n3372 );
and ( n6298 , n3366 , n2666 );
and ( n6299 , n3415 , n2664 );
nor ( n6300 , n6298 , n6299 );
xnor ( n6301 , n6300 , n2587 );
and ( n6302 , n6297 , n6301 );
and ( n6303 , n3882 , n2450 );
and ( n6304 , n3748 , n2448 );
nor ( n6305 , n6303 , n6304 );
xnor ( n6306 , n6305 , n2364 );
and ( n6307 , n6301 , n6306 );
and ( n6308 , n6297 , n6306 );
or ( n6309 , n6302 , n6307 , n6308 );
and ( n6310 , n6292 , n6309 );
and ( n6311 , n6280 , n6309 );
or ( n6312 , n6293 , n6310 , n6311 );
xor ( n6313 , n6163 , n6167 );
xor ( n6314 , n6313 , n6172 );
and ( n6315 , n6312 , n6314 );
xor ( n6316 , n6211 , n6215 );
xor ( n6317 , n6316 , n6220 );
and ( n6318 , n6314 , n6317 );
and ( n6319 , n6312 , n6317 );
or ( n6320 , n6315 , n6318 , n6319 );
xor ( n6321 , n6175 , n6177 );
xor ( n6322 , n6321 , n6180 );
and ( n6323 , n6320 , n6322 );
xor ( n6324 , n6223 , n6261 );
xor ( n6325 , n6324 , n6264 );
and ( n6326 , n6322 , n6325 );
and ( n6327 , n6320 , n6325 );
or ( n6328 , n6323 , n6326 , n6327 );
and ( n6329 , n6279 , n6328 );
xor ( n6330 , n6279 , n6328 );
xor ( n6331 , n6320 , n6322 );
xor ( n6332 , n6331 , n6325 );
and ( n6333 , n2459 , n3929 );
and ( n6334 , n2338 , n3926 );
nor ( n6335 , n6333 , n6334 );
xnor ( n6336 , n6335 , n3372 );
and ( n6337 , n3415 , n2940 );
and ( n6338 , n3079 , n2938 );
nor ( n6339 , n6337 , n6338 );
xnor ( n6340 , n6339 , n2868 );
and ( n6341 , n6336 , n6340 );
and ( n6342 , n3748 , n2666 );
and ( n6343 , n3366 , n2664 );
nor ( n6344 , n6342 , n6343 );
xnor ( n6345 , n6344 , n2587 );
and ( n6346 , n6340 , n6345 );
and ( n6347 , n6336 , n6345 );
or ( n6348 , n6341 , n6346 , n6347 );
and ( n6349 , n2658 , n3813 );
and ( n6350 , n2611 , n3811 );
nor ( n6351 , n6349 , n6350 );
xnor ( n6352 , n6351 , n3375 );
and ( n6353 , n3938 , n2448 );
not ( n6354 , n6353 );
and ( n6355 , n6354 , n2364 );
and ( n6356 , n6352 , n6355 );
and ( n6357 , n6348 , n6356 );
and ( n6358 , n2969 , n3227 );
and ( n6359 , n2658 , n3225 );
nor ( n6360 , n6358 , n6359 );
xnor ( n6361 , n6360 , n3168 );
and ( n6362 , n6356 , n6361 );
and ( n6363 , n6348 , n6361 );
or ( n6364 , n6357 , n6362 , n6363 );
xor ( n6365 , n6227 , n6231 );
xor ( n6366 , n6365 , n6236 );
and ( n6367 , n6364 , n6366 );
xor ( n6368 , n6243 , n6247 );
xor ( n6369 , n6368 , n6252 );
and ( n6370 , n6366 , n6369 );
and ( n6371 , n6364 , n6369 );
or ( n6372 , n6367 , n6370 , n6371 );
xor ( n6373 , n6239 , n6255 );
xor ( n6374 , n6373 , n6258 );
and ( n6375 , n6372 , n6374 );
xor ( n6376 , n6312 , n6314 );
xor ( n6377 , n6376 , n6317 );
and ( n6378 , n6374 , n6377 );
and ( n6379 , n6372 , n6377 );
or ( n6380 , n6375 , n6378 , n6379 );
and ( n6381 , n6332 , n6380 );
xor ( n6382 , n6332 , n6380 );
xor ( n6383 , n6372 , n6374 );
xor ( n6384 , n6383 , n6377 );
xor ( n6385 , n6352 , n6355 );
and ( n6386 , n3019 , n3227 );
and ( n6387 , n2969 , n3225 );
nor ( n6388 , n6386 , n6387 );
xnor ( n6389 , n6388 , n3168 );
and ( n6390 , n6385 , n6389 );
and ( n6391 , n3938 , n2450 );
and ( n6392 , n3882 , n2448 );
nor ( n6393 , n6391 , n6392 );
xnor ( n6394 , n6393 , n2364 );
and ( n6395 , n6389 , n6394 );
and ( n6396 , n6385 , n6394 );
or ( n6397 , n6390 , n6395 , n6396 );
xor ( n6398 , n6284 , n6288 );
xor ( n6399 , n6398 , n6208 );
and ( n6400 , n6397 , n6399 );
xor ( n6401 , n6297 , n6301 );
xor ( n6402 , n6401 , n6306 );
and ( n6403 , n6399 , n6402 );
and ( n6404 , n6397 , n6402 );
or ( n6405 , n6400 , n6403 , n6404 );
xor ( n6406 , n6280 , n6292 );
xor ( n6407 , n6406 , n6309 );
and ( n6408 , n6405 , n6407 );
xor ( n6409 , n6364 , n6366 );
xor ( n6410 , n6409 , n6369 );
and ( n6411 , n6407 , n6410 );
and ( n6412 , n6405 , n6410 );
or ( n6413 , n6408 , n6411 , n6412 );
and ( n6414 , n6384 , n6413 );
xor ( n6415 , n6384 , n6413 );
xor ( n6416 , n6405 , n6407 );
xor ( n6417 , n6416 , n6410 );
and ( n6418 , n2611 , n3929 );
and ( n6419 , n2459 , n3926 );
nor ( n6420 , n6418 , n6419 );
xnor ( n6421 , n6420 , n3372 );
and ( n6422 , n3079 , n3227 );
and ( n6423 , n3019 , n3225 );
nor ( n6424 , n6422 , n6423 );
xnor ( n6425 , n6424 , n3168 );
and ( n6426 , n6421 , n6425 );
and ( n6427 , n3882 , n2666 );
and ( n6428 , n3748 , n2664 );
nor ( n6429 , n6427 , n6428 );
xnor ( n6430 , n6429 , n2587 );
and ( n6431 , n6425 , n6430 );
and ( n6432 , n6421 , n6430 );
or ( n6433 , n6426 , n6431 , n6432 );
and ( n6434 , n2969 , n3813 );
and ( n6435 , n2658 , n3811 );
nor ( n6436 , n6434 , n6435 );
xnor ( n6437 , n6436 , n3375 );
and ( n6438 , n3366 , n2940 );
and ( n6439 , n3415 , n2938 );
nor ( n6440 , n6438 , n6439 );
xnor ( n6441 , n6440 , n2868 );
and ( n6442 , n6437 , n6441 );
and ( n6443 , n6441 , n6353 );
and ( n6444 , n6437 , n6353 );
or ( n6445 , n6442 , n6443 , n6444 );
and ( n6446 , n6433 , n6445 );
xor ( n6447 , n6336 , n6340 );
xor ( n6448 , n6447 , n6345 );
and ( n6449 , n6445 , n6448 );
and ( n6450 , n6433 , n6448 );
or ( n6451 , n6446 , n6449 , n6450 );
xor ( n6452 , n6348 , n6356 );
xor ( n6453 , n6452 , n6361 );
and ( n6454 , n6451 , n6453 );
xor ( n6455 , n6397 , n6399 );
xor ( n6456 , n6455 , n6402 );
and ( n6457 , n6453 , n6456 );
and ( n6458 , n6451 , n6456 );
or ( n6459 , n6454 , n6457 , n6458 );
and ( n6460 , n6417 , n6459 );
xor ( n6461 , n6417 , n6459 );
and ( n6462 , n2658 , n3929 );
and ( n6463 , n2611 , n3926 );
nor ( n6464 , n6462 , n6463 );
xnor ( n6465 , n6464 , n3372 );
and ( n6466 , n3748 , n2940 );
and ( n6467 , n3366 , n2938 );
nor ( n6468 , n6466 , n6467 );
xnor ( n6469 , n6468 , n2868 );
and ( n6470 , n6465 , n6469 );
and ( n6471 , n3938 , n2666 );
and ( n6472 , n3882 , n2664 );
nor ( n6473 , n6471 , n6472 );
xnor ( n6474 , n6473 , n2587 );
and ( n6475 , n6469 , n6474 );
and ( n6476 , n6465 , n6474 );
or ( n6477 , n6470 , n6475 , n6476 );
and ( n6478 , n3019 , n3813 );
and ( n6479 , n2969 , n3811 );
nor ( n6480 , n6478 , n6479 );
xnor ( n6481 , n6480 , n3375 );
and ( n6482 , n3938 , n2664 );
not ( n6483 , n6482 );
and ( n6484 , n6483 , n2587 );
and ( n6485 , n6481 , n6484 );
and ( n6486 , n6477 , n6485 );
xor ( n6487 , n6437 , n6441 );
xor ( n6488 , n6487 , n6353 );
and ( n6489 , n6485 , n6488 );
and ( n6490 , n6477 , n6488 );
or ( n6491 , n6486 , n6489 , n6490 );
xor ( n6492 , n6385 , n6389 );
xor ( n6493 , n6492 , n6394 );
and ( n6494 , n6491 , n6493 );
xor ( n6495 , n6433 , n6445 );
xor ( n6496 , n6495 , n6448 );
and ( n6497 , n6493 , n6496 );
and ( n6498 , n6491 , n6496 );
or ( n6499 , n6494 , n6497 , n6498 );
xor ( n6500 , n6451 , n6453 );
xor ( n6501 , n6500 , n6456 );
and ( n6502 , n6499 , n6501 );
xor ( n6503 , n6499 , n6501 );
xor ( n6504 , n6491 , n6493 );
xor ( n6505 , n6504 , n6496 );
xor ( n6506 , n6481 , n6484 );
and ( n6507 , n2969 , n3929 );
and ( n6508 , n2658 , n3926 );
nor ( n6509 , n6507 , n6508 );
xnor ( n6510 , n6509 , n3372 );
and ( n6511 , n3882 , n2940 );
and ( n6512 , n3748 , n2938 );
nor ( n6513 , n6511 , n6512 );
xnor ( n6514 , n6513 , n2868 );
and ( n6515 , n6510 , n6514 );
and ( n6516 , n6514 , n6482 );
and ( n6517 , n6510 , n6482 );
or ( n6518 , n6515 , n6516 , n6517 );
and ( n6519 , n6506 , n6518 );
and ( n6520 , n3415 , n3227 );
and ( n6521 , n3079 , n3225 );
nor ( n6522 , n6520 , n6521 );
xnor ( n6523 , n6522 , n3168 );
and ( n6524 , n6518 , n6523 );
and ( n6525 , n6506 , n6523 );
or ( n6526 , n6519 , n6524 , n6525 );
xor ( n6527 , n6421 , n6425 );
xor ( n6528 , n6527 , n6430 );
and ( n6529 , n6526 , n6528 );
xor ( n6530 , n6477 , n6485 );
xor ( n6531 , n6530 , n6488 );
and ( n6532 , n6528 , n6531 );
and ( n6533 , n6526 , n6531 );
or ( n6534 , n6529 , n6532 , n6533 );
and ( n6535 , n6505 , n6534 );
xor ( n6536 , n6505 , n6534 );
xor ( n6537 , n6526 , n6528 );
xor ( n6538 , n6537 , n6531 );
and ( n6539 , n3019 , n3929 );
and ( n6540 , n2969 , n3926 );
nor ( n6541 , n6539 , n6540 );
xnor ( n6542 , n6541 , n3372 );
and ( n6543 , n3938 , n2938 );
not ( n6544 , n6543 );
and ( n6545 , n6544 , n2868 );
and ( n6546 , n6542 , n6545 );
and ( n6547 , n3079 , n3813 );
and ( n6548 , n3019 , n3811 );
nor ( n6549 , n6547 , n6548 );
xnor ( n6550 , n6549 , n3375 );
and ( n6551 , n6546 , n6550 );
and ( n6552 , n3366 , n3227 );
and ( n6553 , n3415 , n3225 );
nor ( n6554 , n6552 , n6553 );
xnor ( n6555 , n6554 , n3168 );
and ( n6556 , n6550 , n6555 );
and ( n6557 , n6546 , n6555 );
or ( n6558 , n6551 , n6556 , n6557 );
xor ( n6559 , n6465 , n6469 );
xor ( n6560 , n6559 , n6474 );
and ( n6561 , n6558 , n6560 );
xor ( n6562 , n6506 , n6518 );
xor ( n6563 , n6562 , n6523 );
and ( n6564 , n6560 , n6563 );
and ( n6565 , n6558 , n6563 );
or ( n6566 , n6561 , n6564 , n6565 );
and ( n6567 , n6538 , n6566 );
xor ( n6568 , n6538 , n6566 );
xor ( n6569 , n6558 , n6560 );
xor ( n6570 , n6569 , n6563 );
and ( n6571 , n3415 , n3813 );
and ( n6572 , n3079 , n3811 );
nor ( n6573 , n6571 , n6572 );
xnor ( n6574 , n6573 , n3375 );
and ( n6575 , n3748 , n3227 );
and ( n6576 , n3366 , n3225 );
nor ( n6577 , n6575 , n6576 );
xnor ( n6578 , n6577 , n3168 );
and ( n6579 , n6574 , n6578 );
and ( n6580 , n3938 , n2940 );
and ( n6581 , n3882 , n2938 );
nor ( n6582 , n6580 , n6581 );
xnor ( n6583 , n6582 , n2868 );
and ( n6584 , n6578 , n6583 );
and ( n6585 , n6574 , n6583 );
or ( n6586 , n6579 , n6584 , n6585 );
xor ( n6587 , n6510 , n6514 );
xor ( n6588 , n6587 , n6482 );
and ( n6589 , n6586 , n6588 );
xor ( n6590 , n6546 , n6550 );
xor ( n6591 , n6590 , n6555 );
and ( n6592 , n6588 , n6591 );
and ( n6593 , n6586 , n6591 );
or ( n6594 , n6589 , n6592 , n6593 );
and ( n6595 , n6570 , n6594 );
xor ( n6596 , n6570 , n6594 );
xor ( n6597 , n6542 , n6545 );
and ( n6598 , n3079 , n3929 );
and ( n6599 , n3019 , n3926 );
nor ( n6600 , n6598 , n6599 );
xnor ( n6601 , n6600 , n3372 );
and ( n6602 , n3366 , n3813 );
and ( n6603 , n3415 , n3811 );
nor ( n6604 , n6602 , n6603 );
xnor ( n6605 , n6604 , n3375 );
and ( n6606 , n6601 , n6605 );
and ( n6607 , n6605 , n6543 );
and ( n6608 , n6601 , n6543 );
or ( n6609 , n6606 , n6607 , n6608 );
and ( n6610 , n6597 , n6609 );
xor ( n6611 , n6574 , n6578 );
xor ( n6612 , n6611 , n6583 );
and ( n6613 , n6609 , n6612 );
and ( n6614 , n6597 , n6612 );
or ( n6615 , n6610 , n6613 , n6614 );
xor ( n6616 , n6586 , n6588 );
xor ( n6617 , n6616 , n6591 );
and ( n6618 , n6615 , n6617 );
xor ( n6619 , n6615 , n6617 );
xor ( n6620 , n6597 , n6609 );
xor ( n6621 , n6620 , n6612 );
and ( n6622 , n3415 , n3929 );
and ( n6623 , n3079 , n3926 );
nor ( n6624 , n6622 , n6623 );
xnor ( n6625 , n6624 , n3372 );
and ( n6626 , n3938 , n3225 );
not ( n6627 , n6626 );
and ( n6628 , n6627 , n3168 );
and ( n6629 , n6625 , n6628 );
and ( n6630 , n3882 , n3227 );
and ( n6631 , n3748 , n3225 );
nor ( n6632 , n6630 , n6631 );
xnor ( n6633 , n6632 , n3168 );
and ( n6634 , n6629 , n6633 );
xor ( n6635 , n6601 , n6605 );
xor ( n6636 , n6635 , n6543 );
and ( n6637 , n6633 , n6636 );
and ( n6638 , n6629 , n6636 );
or ( n6639 , n6634 , n6637 , n6638 );
and ( n6640 , n6621 , n6639 );
xor ( n6641 , n6621 , n6639 );
xor ( n6642 , n6629 , n6633 );
xor ( n6643 , n6642 , n6636 );
xor ( n6644 , n6625 , n6628 );
and ( n6645 , n3748 , n3813 );
and ( n6646 , n3366 , n3811 );
nor ( n6647 , n6645 , n6646 );
xnor ( n6648 , n6647 , n3375 );
and ( n6649 , n6644 , n6648 );
and ( n6650 , n3938 , n3227 );
and ( n6651 , n3882 , n3225 );
nor ( n6652 , n6650 , n6651 );
xnor ( n6653 , n6652 , n3168 );
and ( n6654 , n6648 , n6653 );
and ( n6655 , n6644 , n6653 );
or ( n6656 , n6649 , n6654 , n6655 );
and ( n6657 , n6643 , n6656 );
xor ( n6658 , n6643 , n6656 );
and ( n6659 , n3366 , n3929 );
and ( n6660 , n3415 , n3926 );
nor ( n6661 , n6659 , n6660 );
xnor ( n6662 , n6661 , n3372 );
and ( n6663 , n3882 , n3813 );
and ( n6664 , n3748 , n3811 );
nor ( n6665 , n6663 , n6664 );
xnor ( n6666 , n6665 , n3375 );
and ( n6667 , n6662 , n6666 );
and ( n6668 , n6666 , n6626 );
and ( n6669 , n6662 , n6626 );
or ( n6670 , n6667 , n6668 , n6669 );
xor ( n6671 , n6644 , n6648 );
xor ( n6672 , n6671 , n6653 );
and ( n6673 , n6670 , n6672 );
xor ( n6674 , n6670 , n6672 );
xor ( n6675 , n6662 , n6666 );
xor ( n6676 , n6675 , n6626 );
and ( n6677 , n3748 , n3929 );
and ( n6678 , n3366 , n3926 );
nor ( n6679 , n6677 , n6678 );
xnor ( n6680 , n6679 , n3372 );
and ( n6681 , n3938 , n3811 );
not ( n6682 , n6681 );
and ( n6683 , n6682 , n3375 );
and ( n6684 , n6680 , n6683 );
and ( n6685 , n6676 , n6684 );
xor ( n6686 , n6676 , n6684 );
and ( n6687 , n3938 , n3813 );
and ( n6688 , n3882 , n3811 );
nor ( n6689 , n6687 , n6688 );
xnor ( n6690 , n6689 , n3375 );
xor ( n6691 , n6680 , n6683 );
and ( n6692 , n6690 , n6691 );
xor ( n6693 , n6690 , n6691 );
and ( n6694 , n3882 , n3929 );
and ( n6695 , n3748 , n3926 );
nor ( n6696 , n6694 , n6695 );
xnor ( n6697 , n6696 , n3372 );
and ( n6698 , n6697 , n6681 );
xor ( n6699 , n6697 , n6681 );
and ( n6700 , n3938 , n3929 );
and ( n6701 , n3882 , n3926 );
nor ( n6702 , n6700 , n6701 );
xnor ( n6703 , n6702 , n3372 );
and ( n6704 , n3938 , n3926 );
not ( n6705 , n6704 );
and ( n6706 , n6705 , n3372 );
and ( n6707 , n6703 , n6706 );
and ( n6708 , n6699 , n6707 );
or ( n6709 , n6698 , n6708 );
and ( n6710 , n6693 , n6709 );
or ( n6711 , n6692 , n6710 );
and ( n6712 , n6686 , n6711 );
or ( n6713 , n6685 , n6712 );
and ( n6714 , n6674 , n6713 );
or ( n6715 , n6673 , n6714 );
and ( n6716 , n6658 , n6715 );
or ( n6717 , n6657 , n6716 );
and ( n6718 , n6641 , n6717 );
or ( n6719 , n6640 , n6718 );
and ( n6720 , n6619 , n6719 );
or ( n6721 , n6618 , n6720 );
and ( n6722 , n6596 , n6721 );
or ( n6723 , n6595 , n6722 );
and ( n6724 , n6568 , n6723 );
or ( n6725 , n6567 , n6724 );
and ( n6726 , n6536 , n6725 );
or ( n6727 , n6535 , n6726 );
and ( n6728 , n6503 , n6727 );
or ( n6729 , n6502 , n6728 );
and ( n6730 , n6461 , n6729 );
or ( n6731 , n6460 , n6730 );
and ( n6732 , n6415 , n6731 );
or ( n6733 , n6414 , n6732 );
and ( n6734 , n6382 , n6733 );
or ( n6735 , n6381 , n6734 );
and ( n6736 , n6330 , n6735 );
or ( n6737 , n6329 , n6736 );
and ( n6738 , n6277 , n6737 );
or ( n6739 , n6276 , n6738 );
and ( n6740 , n6201 , n6739 );
or ( n6741 , n6200 , n6740 );
and ( n6742 , n6138 , n6741 );
or ( n6743 , n6137 , n6742 );
and ( n6744 , n6066 , n6743 );
or ( n6745 , n6065 , n6744 );
and ( n6746 , n5990 , n6745 );
or ( n6747 , n5989 , n6746 );
and ( n6748 , n5889 , n6747 );
or ( n6749 , n5888 , n6748 );
and ( n6750 , n5806 , n6749 );
or ( n6751 , n5805 , n6750 );
and ( n6752 , n5776 , n6751 );
or ( n6753 , n5775 , n6752 );
and ( n6754 , n5630 , n6753 );
or ( n6755 , n5629 , n6754 );
and ( n6756 , n5577 , n6755 );
or ( n6757 , n5576 , n6756 );
and ( n6758 , n5475 , n6757 );
or ( n6759 , n5474 , n6758 );
and ( n6760 , n5358 , n6759 );
or ( n6761 , n5357 , n6760 );
and ( n6762 , n5246 , n6761 );
and ( n6763 , n5244 , n6762 );
and ( n6764 , n5242 , n6763 );
and ( n6765 , n5240 , n6764 );
or ( n6766 , n5239 , n6765 );
and ( n6767 , n4932 , n6766 );
and ( n6768 , n4930 , n6767 );
or ( n6769 , n4929 , n6768 );
and ( n6770 , n4610 , n6769 );
or ( n6771 , n4609 , n6770 );
and ( n6772 , n4400 , n6771 );
or ( n6773 , n4399 , n6772 );
and ( n6774 , n4293 , n6773 );
or ( n6775 , n4292 , n6774 );
and ( n6776 , n4209 , n6775 );
and ( n6777 , n4207 , n6776 );
or ( n6778 , n4206 , n6777 );
and ( n6779 , n3735 , n6778 );
and ( n6780 , n3733 , n6779 );
and ( n6781 , n3731 , n6780 );
or ( n6782 , n3730 , n6781 );
and ( n6783 , n3616 , n6782 );
and ( n6784 , n3614 , n6783 );
and ( n6785 , n3612 , n6784 );
and ( n6786 , n3610 , n6785 );
and ( n6787 , n3608 , n6786 );
and ( n6788 , n3606 , n6787 );
and ( n6789 , n3604 , n6788 );
and ( n6790 , n3602 , n6789 );
and ( n6791 , n3600 , n6790 );
and ( n6792 , n3598 , n6791 );
and ( n6793 , n3596 , n6792 );
and ( n6794 , n3594 , n6793 );
and ( n6795 , n3592 , n6794 );
and ( n6796 , n3590 , n6795 );
and ( n6797 , n3588 , n6796 );
and ( n6798 , n3586 , n6797 );
and ( n6799 , n3584 , n6798 );
and ( n6800 , n3582 , n6799 );
and ( n6801 , n3580 , n6800 );
and ( n6802 , n3578 , n6801 );
xor ( n6803 , n3576 , n6802 );
buf ( n6804 , n6803 );
xor ( n6805 , n3578 , n6801 );
buf ( n6806 , n6805 );
xor ( n6807 , n3580 , n6800 );
buf ( n6808 , n6807 );
xor ( n6809 , n3582 , n6799 );
buf ( n6810 , n6809 );
xor ( n6811 , n3584 , n6798 );
buf ( n6812 , n6811 );
xor ( n6813 , n3586 , n6797 );
buf ( n6814 , n6813 );
xor ( n6815 , n3588 , n6796 );
buf ( n6816 , n6815 );
xor ( n6817 , n3590 , n6795 );
buf ( n6818 , n6817 );
xor ( n6819 , n3592 , n6794 );
buf ( n6820 , n6819 );
xor ( n6821 , n3594 , n6793 );
buf ( n6822 , n6821 );
xor ( n6823 , n3596 , n6792 );
buf ( n6824 , n6823 );
xor ( n6825 , n3598 , n6791 );
buf ( n6826 , n6825 );
xor ( n6827 , n3600 , n6790 );
buf ( n6828 , n6827 );
xor ( n6829 , n3602 , n6789 );
buf ( n6830 , n6829 );
xor ( n6831 , n3604 , n6788 );
buf ( n6832 , n6831 );
xor ( n6833 , n3606 , n6787 );
buf ( n6834 , n6833 );
xor ( n6835 , n3608 , n6786 );
buf ( n6836 , n6835 );
xor ( n6837 , n3610 , n6785 );
buf ( n6838 , n6837 );
xor ( n6839 , n3612 , n6784 );
buf ( n6840 , n6839 );
xor ( n6841 , n3614 , n6783 );
buf ( n6842 , n6841 );
xor ( n6843 , n3616 , n6782 );
buf ( n6844 , n6843 );
xor ( n6845 , n3731 , n6780 );
buf ( n6846 , n6845 );
xor ( n6847 , n3733 , n6779 );
buf ( n6848 , n6847 );
xor ( n6849 , n3735 , n6778 );
buf ( n6850 , n6849 );
xor ( n6851 , n4207 , n6776 );
buf ( n6852 , n6851 );
xor ( n6853 , n4209 , n6775 );
buf ( n6854 , n6853 );
xor ( n6855 , n4293 , n6773 );
buf ( n6856 , n6855 );
xor ( n6857 , n4400 , n6771 );
buf ( n6858 , n6857 );
xor ( n6859 , n4610 , n6769 );
buf ( n6860 , n6859 );
xor ( n6861 , n4930 , n6767 );
buf ( n6862 , n6861 );
xor ( n6863 , n4932 , n6766 );
buf ( n6864 , n6863 );
xor ( n6865 , n5240 , n6764 );
buf ( n6866 , n6865 );
xor ( n6867 , n5242 , n6763 );
buf ( n6868 , n6867 );
xor ( n6869 , n5244 , n6762 );
buf ( n6870 , n6869 );
xor ( n6871 , n5246 , n6761 );
buf ( n6872 , n6871 );
xor ( n6873 , n5358 , n6759 );
buf ( n6874 , n6873 );
xor ( n6875 , n5475 , n6757 );
buf ( n6876 , n6875 );
xor ( n6877 , n5577 , n6755 );
buf ( n6878 , n6877 );
xor ( n6879 , n5630 , n6753 );
buf ( n6880 , n6879 );
xor ( n6881 , n5776 , n6751 );
buf ( n6882 , n6881 );
xor ( n6883 , n5806 , n6749 );
buf ( n6884 , n6883 );
xor ( n6885 , n5889 , n6747 );
buf ( n6886 , n6885 );
xor ( n6887 , n5990 , n6745 );
buf ( n6888 , n6887 );
xor ( n6889 , n6066 , n6743 );
buf ( n6890 , n6889 );
xor ( n6891 , n6138 , n6741 );
buf ( n6892 , n6891 );
xor ( n6893 , n6201 , n6739 );
buf ( n6894 , n6893 );
xor ( n6895 , n6277 , n6737 );
buf ( n6896 , n6895 );
xor ( n6897 , n6330 , n6735 );
buf ( n6898 , n6897 );
xor ( n6899 , n6382 , n6733 );
buf ( n6900 , n6899 );
xor ( n6901 , n6415 , n6731 );
buf ( n6902 , n6901 );
xor ( n6903 , n6461 , n6729 );
buf ( n6904 , n6903 );
xor ( n6905 , n6503 , n6727 );
buf ( n6906 , n6905 );
xor ( n6907 , n6536 , n6725 );
buf ( n6908 , n6907 );
xor ( n6909 , n6568 , n6723 );
buf ( n6910 , n6909 );
xor ( n6911 , n6596 , n6721 );
buf ( n6912 , n6911 );
xor ( n6913 , n6619 , n6719 );
buf ( n6914 , n6913 );
xor ( n6915 , n6641 , n6717 );
buf ( n6916 , n6915 );
xor ( n6917 , n6658 , n6715 );
buf ( n6918 , n6917 );
xor ( n6919 , n6674 , n6713 );
buf ( n6920 , n6919 );
xor ( n6921 , n6686 , n6711 );
buf ( n6922 , n6921 );
xor ( n6923 , n6693 , n6709 );
buf ( n6924 , n6923 );
xor ( n6925 , n6699 , n6707 );
buf ( n6926 , n6925 );
xor ( n6927 , n6703 , n6706 );
buf ( n6928 , n6927 );
buf ( n6929 , n6704 );
buf ( n6930 , n6929 );
buf ( n6931 , n799 );
buf ( n6932 , n6931 );
buf ( n6933 , n831 );
buf ( n6934 , n6933 );
and ( n6935 , n6932 , n6934 );
buf ( n6936 , n895 );
buf ( n6937 , n6936 );
xor ( n6938 , n6935 , n6937 );
buf ( n6939 , n6938 );
buf ( n6940 , n799 );
buf ( n6941 , n6940 );
buf ( n6942 , n831 );
buf ( n6943 , n6942 );
and ( n6944 , n6941 , n6943 );
buf ( n6945 , n863 );
buf ( n6946 , n6945 );
xor ( n6947 , n6944 , n6946 );
buf ( n6948 , n6947 );
not ( n6949 , n831 );
and ( n6950 , n6949 , n6939 );
and ( n6951 , n6948 , n831 );
or ( n6952 , n6950 , n6951 );
buf ( n6953 , n830 );
buf ( n6954 , n6953 );
xor ( n6955 , n6954 , n6934 );
not ( n6956 , n6934 );
and ( n6957 , n6955 , n6956 );
and ( n6958 , n6932 , n6957 );
buf ( n6959 , n798 );
buf ( n6960 , n6959 );
and ( n6961 , n6960 , n6934 );
nor ( n6962 , n6958 , n6961 );
xnor ( n6963 , n6962 , n6954 );
not ( n6964 , n6935 );
and ( n6965 , n6964 , n6954 );
buf ( n6966 , n894 );
buf ( n6967 , n6966 );
xor ( n6968 , n6965 , n6967 );
xor ( n6969 , n6963 , n6968 );
and ( n6970 , n6935 , n6937 );
xor ( n6971 , n6969 , n6970 );
buf ( n6972 , n6971 );
buf ( n6973 , n830 );
buf ( n6974 , n6973 );
xor ( n6975 , n6974 , n6943 );
not ( n6976 , n6943 );
and ( n6977 , n6975 , n6976 );
and ( n6978 , n6941 , n6977 );
buf ( n6979 , n798 );
buf ( n6980 , n6979 );
and ( n6981 , n6980 , n6943 );
nor ( n6982 , n6978 , n6981 );
xnor ( n6983 , n6982 , n6974 );
not ( n6984 , n6944 );
and ( n6985 , n6984 , n6974 );
buf ( n6986 , n862 );
buf ( n6987 , n6986 );
xor ( n6988 , n6985 , n6987 );
xor ( n6989 , n6983 , n6988 );
and ( n6990 , n6944 , n6946 );
xor ( n6991 , n6989 , n6990 );
buf ( n6992 , n6991 );
not ( n6993 , n831 );
and ( n6994 , n6993 , n6972 );
and ( n6995 , n6992 , n831 );
or ( n6996 , n6994 , n6995 );
and ( n6997 , n6960 , n6957 );
buf ( n6998 , n797 );
buf ( n6999 , n6998 );
and ( n7000 , n6999 , n6934 );
nor ( n7001 , n6997 , n7000 );
xnor ( n7002 , n7001 , n6954 );
buf ( n7003 , n829 );
buf ( n7004 , n7003 );
xor ( n7005 , n7004 , n6954 );
and ( n7006 , n6932 , n7005 );
xor ( n7007 , n7002 , n7006 );
buf ( n7008 , n893 );
buf ( n7009 , n7008 );
xor ( n7010 , n7007 , n7009 );
and ( n7011 , n6965 , n6967 );
xor ( n7012 , n7010 , n7011 );
and ( n7013 , n6963 , n6968 );
and ( n7014 , n6969 , n6970 );
or ( n7015 , n7013 , n7014 );
xor ( n7016 , n7012 , n7015 );
buf ( n7017 , n7016 );
and ( n7018 , n6980 , n6977 );
buf ( n7019 , n797 );
buf ( n7020 , n7019 );
and ( n7021 , n7020 , n6943 );
nor ( n7022 , n7018 , n7021 );
xnor ( n7023 , n7022 , n6974 );
buf ( n7024 , n829 );
buf ( n7025 , n7024 );
xor ( n7026 , n7025 , n6974 );
and ( n7027 , n6941 , n7026 );
xor ( n7028 , n7023 , n7027 );
buf ( n7029 , n861 );
buf ( n7030 , n7029 );
xor ( n7031 , n7028 , n7030 );
and ( n7032 , n6985 , n6987 );
xor ( n7033 , n7031 , n7032 );
and ( n7034 , n6983 , n6988 );
and ( n7035 , n6989 , n6990 );
or ( n7036 , n7034 , n7035 );
xor ( n7037 , n7033 , n7036 );
buf ( n7038 , n7037 );
not ( n7039 , n831 );
and ( n7040 , n7039 , n7017 );
and ( n7041 , n7038 , n831 );
or ( n7042 , n7040 , n7041 );
and ( n7043 , n7002 , n7006 );
and ( n7044 , n7006 , n7009 );
and ( n7045 , n7002 , n7009 );
or ( n7046 , n7043 , n7044 , n7045 );
and ( n7047 , n6999 , n6957 );
buf ( n7048 , n796 );
buf ( n7049 , n7048 );
and ( n7050 , n7049 , n6934 );
nor ( n7051 , n7047 , n7050 );
xnor ( n7052 , n7051 , n6954 );
not ( n7053 , n7006 );
buf ( n7054 , n828 );
buf ( n7055 , n7054 );
and ( n7056 , n7004 , n6954 );
not ( n7057 , n7056 );
and ( n7058 , n7055 , n7057 );
and ( n7059 , n7053 , n7058 );
xor ( n7060 , n7052 , n7059 );
xor ( n7061 , n7055 , n7004 );
not ( n7062 , n7005 );
and ( n7063 , n7061 , n7062 );
and ( n7064 , n6932 , n7063 );
and ( n7065 , n6960 , n7005 );
nor ( n7066 , n7064 , n7065 );
xnor ( n7067 , n7066 , n7058 );
buf ( n7068 , n892 );
buf ( n7069 , n7068 );
xor ( n7070 , n7067 , n7069 );
xor ( n7071 , n7060 , n7070 );
xor ( n7072 , n7046 , n7071 );
and ( n7073 , n7010 , n7011 );
and ( n7074 , n7012 , n7015 );
or ( n7075 , n7073 , n7074 );
xor ( n7076 , n7072 , n7075 );
buf ( n7077 , n7076 );
and ( n7078 , n7023 , n7027 );
and ( n7079 , n7027 , n7030 );
and ( n7080 , n7023 , n7030 );
or ( n7081 , n7078 , n7079 , n7080 );
and ( n7082 , n7020 , n6977 );
buf ( n7083 , n796 );
buf ( n7084 , n7083 );
and ( n7085 , n7084 , n6943 );
nor ( n7086 , n7082 , n7085 );
xnor ( n7087 , n7086 , n6974 );
not ( n7088 , n7027 );
buf ( n7089 , n828 );
buf ( n7090 , n7089 );
and ( n7091 , n7025 , n6974 );
not ( n7092 , n7091 );
and ( n7093 , n7090 , n7092 );
and ( n7094 , n7088 , n7093 );
xor ( n7095 , n7087 , n7094 );
xor ( n7096 , n7090 , n7025 );
not ( n7097 , n7026 );
and ( n7098 , n7096 , n7097 );
and ( n7099 , n6941 , n7098 );
and ( n7100 , n6980 , n7026 );
nor ( n7101 , n7099 , n7100 );
xnor ( n7102 , n7101 , n7093 );
buf ( n7103 , n860 );
buf ( n7104 , n7103 );
xor ( n7105 , n7102 , n7104 );
xor ( n7106 , n7095 , n7105 );
xor ( n7107 , n7081 , n7106 );
and ( n7108 , n7031 , n7032 );
and ( n7109 , n7033 , n7036 );
or ( n7110 , n7108 , n7109 );
xor ( n7111 , n7107 , n7110 );
buf ( n7112 , n7111 );
not ( n7113 , n831 );
and ( n7114 , n7113 , n7077 );
and ( n7115 , n7112 , n831 );
or ( n7116 , n7114 , n7115 );
and ( n7117 , n7052 , n7059 );
and ( n7118 , n7059 , n7070 );
and ( n7119 , n7052 , n7070 );
or ( n7120 , n7117 , n7118 , n7119 );
buf ( n7121 , n891 );
buf ( n7122 , n7121 );
and ( n7123 , n7049 , n6957 );
buf ( n7124 , n795 );
buf ( n7125 , n7124 );
and ( n7126 , n7125 , n6934 );
nor ( n7127 , n7123 , n7126 );
xnor ( n7128 , n7127 , n6954 );
and ( n7129 , n6960 , n7063 );
and ( n7130 , n6999 , n7005 );
nor ( n7131 , n7129 , n7130 );
xnor ( n7132 , n7131 , n7058 );
xor ( n7133 , n7128 , n7132 );
buf ( n7134 , n827 );
buf ( n7135 , n7134 );
xor ( n7136 , n7135 , n7055 );
and ( n7137 , n6932 , n7136 );
xor ( n7138 , n7133 , n7137 );
xor ( n7139 , n7122 , n7138 );
and ( n7140 , n7067 , n7069 );
xor ( n7141 , n7139 , n7140 );
xor ( n7142 , n7120 , n7141 );
and ( n7143 , n7046 , n7071 );
and ( n7144 , n7072 , n7075 );
or ( n7145 , n7143 , n7144 );
xor ( n7146 , n7142 , n7145 );
buf ( n7147 , n7146 );
and ( n7148 , n7087 , n7094 );
and ( n7149 , n7094 , n7105 );
and ( n7150 , n7087 , n7105 );
or ( n7151 , n7148 , n7149 , n7150 );
buf ( n7152 , n859 );
buf ( n7153 , n7152 );
and ( n7154 , n7084 , n6977 );
buf ( n7155 , n795 );
buf ( n7156 , n7155 );
and ( n7157 , n7156 , n6943 );
nor ( n7158 , n7154 , n7157 );
xnor ( n7159 , n7158 , n6974 );
and ( n7160 , n6980 , n7098 );
and ( n7161 , n7020 , n7026 );
nor ( n7162 , n7160 , n7161 );
xnor ( n7163 , n7162 , n7093 );
xor ( n7164 , n7159 , n7163 );
buf ( n7165 , n827 );
buf ( n7166 , n7165 );
xor ( n7167 , n7166 , n7090 );
and ( n7168 , n6941 , n7167 );
xor ( n7169 , n7164 , n7168 );
xor ( n7170 , n7153 , n7169 );
and ( n7171 , n7102 , n7104 );
xor ( n7172 , n7170 , n7171 );
xor ( n7173 , n7151 , n7172 );
and ( n7174 , n7081 , n7106 );
and ( n7175 , n7107 , n7110 );
or ( n7176 , n7174 , n7175 );
xor ( n7177 , n7173 , n7176 );
buf ( n7178 , n7177 );
not ( n7179 , n831 );
and ( n7180 , n7179 , n7147 );
and ( n7181 , n7178 , n831 );
or ( n7182 , n7180 , n7181 );
and ( n7183 , n7122 , n7138 );
and ( n7184 , n7138 , n7140 );
and ( n7185 , n7122 , n7140 );
or ( n7186 , n7183 , n7184 , n7185 );
and ( n7187 , n7128 , n7132 );
and ( n7188 , n7132 , n7137 );
and ( n7189 , n7128 , n7137 );
or ( n7190 , n7187 , n7188 , n7189 );
buf ( n7191 , n890 );
buf ( n7192 , n7191 );
xor ( n7193 , n7190 , n7192 );
and ( n7194 , n7125 , n6957 );
buf ( n7195 , n794 );
buf ( n7196 , n7195 );
and ( n7197 , n7196 , n6934 );
nor ( n7198 , n7194 , n7197 );
xnor ( n7199 , n7198 , n6954 );
not ( n7200 , n7137 );
buf ( n7201 , n826 );
buf ( n7202 , n7201 );
and ( n7203 , n7135 , n7055 );
not ( n7204 , n7203 );
and ( n7205 , n7202 , n7204 );
and ( n7206 , n7200 , n7205 );
xor ( n7207 , n7199 , n7206 );
and ( n7208 , n6999 , n7063 );
and ( n7209 , n7049 , n7005 );
nor ( n7210 , n7208 , n7209 );
xnor ( n7211 , n7210 , n7058 );
xor ( n7212 , n7207 , n7211 );
xor ( n7213 , n7202 , n7135 );
not ( n7214 , n7136 );
and ( n7215 , n7213 , n7214 );
and ( n7216 , n6932 , n7215 );
and ( n7217 , n6960 , n7136 );
nor ( n7218 , n7216 , n7217 );
xnor ( n7219 , n7218 , n7205 );
xor ( n7220 , n7212 , n7219 );
xor ( n7221 , n7193 , n7220 );
xor ( n7222 , n7186 , n7221 );
and ( n7223 , n7120 , n7141 );
and ( n7224 , n7142 , n7145 );
or ( n7225 , n7223 , n7224 );
xor ( n7226 , n7222 , n7225 );
buf ( n7227 , n7226 );
and ( n7228 , n7153 , n7169 );
and ( n7229 , n7169 , n7171 );
and ( n7230 , n7153 , n7171 );
or ( n7231 , n7228 , n7229 , n7230 );
and ( n7232 , n7159 , n7163 );
and ( n7233 , n7163 , n7168 );
and ( n7234 , n7159 , n7168 );
or ( n7235 , n7232 , n7233 , n7234 );
buf ( n7236 , n858 );
buf ( n7237 , n7236 );
xor ( n7238 , n7235 , n7237 );
and ( n7239 , n7156 , n6977 );
buf ( n7240 , n794 );
buf ( n7241 , n7240 );
and ( n7242 , n7241 , n6943 );
nor ( n7243 , n7239 , n7242 );
xnor ( n7244 , n7243 , n6974 );
not ( n7245 , n7168 );
buf ( n7246 , n826 );
buf ( n7247 , n7246 );
and ( n7248 , n7166 , n7090 );
not ( n7249 , n7248 );
and ( n7250 , n7247 , n7249 );
and ( n7251 , n7245 , n7250 );
xor ( n7252 , n7244 , n7251 );
and ( n7253 , n7020 , n7098 );
and ( n7254 , n7084 , n7026 );
nor ( n7255 , n7253 , n7254 );
xnor ( n7256 , n7255 , n7093 );
xor ( n7257 , n7252 , n7256 );
xor ( n7258 , n7247 , n7166 );
not ( n7259 , n7167 );
and ( n7260 , n7258 , n7259 );
and ( n7261 , n6941 , n7260 );
and ( n7262 , n6980 , n7167 );
nor ( n7263 , n7261 , n7262 );
xnor ( n7264 , n7263 , n7250 );
xor ( n7265 , n7257 , n7264 );
xor ( n7266 , n7238 , n7265 );
xor ( n7267 , n7231 , n7266 );
and ( n7268 , n7151 , n7172 );
and ( n7269 , n7173 , n7176 );
or ( n7270 , n7268 , n7269 );
xor ( n7271 , n7267 , n7270 );
buf ( n7272 , n7271 );
not ( n7273 , n831 );
and ( n7274 , n7273 , n7227 );
and ( n7275 , n7272 , n831 );
or ( n7276 , n7274 , n7275 );
and ( n7277 , n7207 , n7211 );
and ( n7278 , n7211 , n7219 );
and ( n7279 , n7207 , n7219 );
or ( n7280 , n7277 , n7278 , n7279 );
buf ( n7281 , n889 );
buf ( n7282 , n7281 );
xor ( n7283 , n7280 , n7282 );
and ( n7284 , n7199 , n7206 );
and ( n7285 , n6960 , n7215 );
and ( n7286 , n6999 , n7136 );
nor ( n7287 , n7285 , n7286 );
xnor ( n7288 , n7287 , n7205 );
xor ( n7289 , n7284 , n7288 );
and ( n7290 , n7196 , n6957 );
buf ( n7291 , n793 );
buf ( n7292 , n7291 );
and ( n7293 , n7292 , n6934 );
nor ( n7294 , n7290 , n7293 );
xnor ( n7295 , n7294 , n6954 );
and ( n7296 , n7049 , n7063 );
and ( n7297 , n7125 , n7005 );
nor ( n7298 , n7296 , n7297 );
xnor ( n7299 , n7298 , n7058 );
xor ( n7300 , n7295 , n7299 );
buf ( n7301 , n825 );
buf ( n7302 , n7301 );
xor ( n7303 , n7302 , n7202 );
and ( n7304 , n6932 , n7303 );
xor ( n7305 , n7300 , n7304 );
xor ( n7306 , n7289 , n7305 );
xor ( n7307 , n7283 , n7306 );
and ( n7308 , n7190 , n7192 );
and ( n7309 , n7192 , n7220 );
and ( n7310 , n7190 , n7220 );
or ( n7311 , n7308 , n7309 , n7310 );
xor ( n7312 , n7307 , n7311 );
and ( n7313 , n7186 , n7221 );
and ( n7314 , n7222 , n7225 );
or ( n7315 , n7313 , n7314 );
xor ( n7316 , n7312 , n7315 );
buf ( n7317 , n7316 );
and ( n7318 , n7252 , n7256 );
and ( n7319 , n7256 , n7264 );
and ( n7320 , n7252 , n7264 );
or ( n7321 , n7318 , n7319 , n7320 );
buf ( n7322 , n857 );
buf ( n7323 , n7322 );
xor ( n7324 , n7321 , n7323 );
and ( n7325 , n7244 , n7251 );
and ( n7326 , n6980 , n7260 );
and ( n7327 , n7020 , n7167 );
nor ( n7328 , n7326 , n7327 );
xnor ( n7329 , n7328 , n7250 );
xor ( n7330 , n7325 , n7329 );
and ( n7331 , n7241 , n6977 );
buf ( n7332 , n793 );
buf ( n7333 , n7332 );
and ( n7334 , n7333 , n6943 );
nor ( n7335 , n7331 , n7334 );
xnor ( n7336 , n7335 , n6974 );
and ( n7337 , n7084 , n7098 );
and ( n7338 , n7156 , n7026 );
nor ( n7339 , n7337 , n7338 );
xnor ( n7340 , n7339 , n7093 );
xor ( n7341 , n7336 , n7340 );
buf ( n7342 , n825 );
buf ( n7343 , n7342 );
xor ( n7344 , n7343 , n7247 );
and ( n7345 , n6941 , n7344 );
xor ( n7346 , n7341 , n7345 );
xor ( n7347 , n7330 , n7346 );
xor ( n7348 , n7324 , n7347 );
and ( n7349 , n7235 , n7237 );
and ( n7350 , n7237 , n7265 );
and ( n7351 , n7235 , n7265 );
or ( n7352 , n7349 , n7350 , n7351 );
xor ( n7353 , n7348 , n7352 );
and ( n7354 , n7231 , n7266 );
and ( n7355 , n7267 , n7270 );
or ( n7356 , n7354 , n7355 );
xor ( n7357 , n7353 , n7356 );
buf ( n7358 , n7357 );
not ( n7359 , n831 );
and ( n7360 , n7359 , n7317 );
and ( n7361 , n7358 , n831 );
or ( n7362 , n7360 , n7361 );
and ( n7363 , n7284 , n7288 );
and ( n7364 , n7288 , n7305 );
and ( n7365 , n7284 , n7305 );
or ( n7366 , n7363 , n7364 , n7365 );
buf ( n7367 , n888 );
buf ( n7368 , n7367 );
xor ( n7369 , n7366 , n7368 );
and ( n7370 , n7292 , n6957 );
buf ( n7371 , n792 );
buf ( n7372 , n7371 );
and ( n7373 , n7372 , n6934 );
nor ( n7374 , n7370 , n7373 );
xnor ( n7375 , n7374 , n6954 );
not ( n7376 , n7304 );
buf ( n7377 , n824 );
buf ( n7378 , n7377 );
and ( n7379 , n7302 , n7202 );
not ( n7380 , n7379 );
and ( n7381 , n7378 , n7380 );
and ( n7382 , n7376 , n7381 );
xor ( n7383 , n7375 , n7382 );
and ( n7384 , n7295 , n7299 );
and ( n7385 , n7299 , n7304 );
and ( n7386 , n7295 , n7304 );
or ( n7387 , n7384 , n7385 , n7386 );
xor ( n7388 , n7383 , n7387 );
and ( n7389 , n7125 , n7063 );
and ( n7390 , n7196 , n7005 );
nor ( n7391 , n7389 , n7390 );
xnor ( n7392 , n7391 , n7058 );
and ( n7393 , n6999 , n7215 );
and ( n7394 , n7049 , n7136 );
nor ( n7395 , n7393 , n7394 );
xnor ( n7396 , n7395 , n7205 );
xor ( n7397 , n7392 , n7396 );
xor ( n7398 , n7378 , n7302 );
not ( n7399 , n7303 );
and ( n7400 , n7398 , n7399 );
and ( n7401 , n6932 , n7400 );
and ( n7402 , n6960 , n7303 );
nor ( n7403 , n7401 , n7402 );
xnor ( n7404 , n7403 , n7381 );
xor ( n7405 , n7397 , n7404 );
xor ( n7406 , n7388 , n7405 );
xor ( n7407 , n7369 , n7406 );
and ( n7408 , n7280 , n7282 );
and ( n7409 , n7282 , n7306 );
and ( n7410 , n7280 , n7306 );
or ( n7411 , n7408 , n7409 , n7410 );
xor ( n7412 , n7407 , n7411 );
and ( n7413 , n7307 , n7311 );
and ( n7414 , n7312 , n7315 );
or ( n7415 , n7413 , n7414 );
xor ( n7416 , n7412 , n7415 );
buf ( n7417 , n7416 );
and ( n7418 , n7325 , n7329 );
and ( n7419 , n7329 , n7346 );
and ( n7420 , n7325 , n7346 );
or ( n7421 , n7418 , n7419 , n7420 );
buf ( n7422 , n856 );
buf ( n7423 , n7422 );
xor ( n7424 , n7421 , n7423 );
and ( n7425 , n7333 , n6977 );
buf ( n7426 , n792 );
buf ( n7427 , n7426 );
and ( n7428 , n7427 , n6943 );
nor ( n7429 , n7425 , n7428 );
xnor ( n7430 , n7429 , n6974 );
not ( n7431 , n7345 );
buf ( n7432 , n824 );
buf ( n7433 , n7432 );
and ( n7434 , n7343 , n7247 );
not ( n7435 , n7434 );
and ( n7436 , n7433 , n7435 );
and ( n7437 , n7431 , n7436 );
xor ( n7438 , n7430 , n7437 );
and ( n7439 , n7336 , n7340 );
and ( n7440 , n7340 , n7345 );
and ( n7441 , n7336 , n7345 );
or ( n7442 , n7439 , n7440 , n7441 );
xor ( n7443 , n7438 , n7442 );
and ( n7444 , n7156 , n7098 );
and ( n7445 , n7241 , n7026 );
nor ( n7446 , n7444 , n7445 );
xnor ( n7447 , n7446 , n7093 );
and ( n7448 , n7020 , n7260 );
and ( n7449 , n7084 , n7167 );
nor ( n7450 , n7448 , n7449 );
xnor ( n7451 , n7450 , n7250 );
xor ( n7452 , n7447 , n7451 );
xor ( n7453 , n7433 , n7343 );
not ( n7454 , n7344 );
and ( n7455 , n7453 , n7454 );
and ( n7456 , n6941 , n7455 );
and ( n7457 , n6980 , n7344 );
nor ( n7458 , n7456 , n7457 );
xnor ( n7459 , n7458 , n7436 );
xor ( n7460 , n7452 , n7459 );
xor ( n7461 , n7443 , n7460 );
xor ( n7462 , n7424 , n7461 );
and ( n7463 , n7321 , n7323 );
and ( n7464 , n7323 , n7347 );
and ( n7465 , n7321 , n7347 );
or ( n7466 , n7463 , n7464 , n7465 );
xor ( n7467 , n7462 , n7466 );
and ( n7468 , n7348 , n7352 );
and ( n7469 , n7353 , n7356 );
or ( n7470 , n7468 , n7469 );
xor ( n7471 , n7467 , n7470 );
buf ( n7472 , n7471 );
not ( n7473 , n831 );
and ( n7474 , n7473 , n7417 );
and ( n7475 , n7472 , n831 );
or ( n7476 , n7474 , n7475 );
and ( n7477 , n7366 , n7368 );
and ( n7478 , n7368 , n7406 );
and ( n7479 , n7366 , n7406 );
or ( n7480 , n7477 , n7478 , n7479 );
and ( n7481 , n7383 , n7387 );
and ( n7482 , n7387 , n7405 );
and ( n7483 , n7383 , n7405 );
or ( n7484 , n7481 , n7482 , n7483 );
buf ( n7485 , n887 );
buf ( n7486 , n7485 );
xor ( n7487 , n7484 , n7486 );
and ( n7488 , n7392 , n7396 );
and ( n7489 , n7396 , n7404 );
and ( n7490 , n7392 , n7404 );
or ( n7491 , n7488 , n7489 , n7490 );
and ( n7492 , n7372 , n6957 );
buf ( n7493 , n791 );
buf ( n7494 , n7493 );
and ( n7495 , n7494 , n6934 );
nor ( n7496 , n7492 , n7495 );
xnor ( n7497 , n7496 , n6954 );
and ( n7498 , n6960 , n7400 );
and ( n7499 , n6999 , n7303 );
nor ( n7500 , n7498 , n7499 );
xnor ( n7501 , n7500 , n7381 );
xor ( n7502 , n7497 , n7501 );
buf ( n7503 , n823 );
buf ( n7504 , n7503 );
xor ( n7505 , n7504 , n7378 );
and ( n7506 , n6932 , n7505 );
xor ( n7507 , n7502 , n7506 );
xor ( n7508 , n7491 , n7507 );
and ( n7509 , n7375 , n7382 );
and ( n7510 , n7196 , n7063 );
and ( n7511 , n7292 , n7005 );
nor ( n7512 , n7510 , n7511 );
xnor ( n7513 , n7512 , n7058 );
xor ( n7514 , n7509 , n7513 );
and ( n7515 , n7049 , n7215 );
and ( n7516 , n7125 , n7136 );
nor ( n7517 , n7515 , n7516 );
xnor ( n7518 , n7517 , n7205 );
xor ( n7519 , n7514 , n7518 );
xor ( n7520 , n7508 , n7519 );
xor ( n7521 , n7487 , n7520 );
xor ( n7522 , n7480 , n7521 );
and ( n7523 , n7407 , n7411 );
and ( n7524 , n7412 , n7415 );
or ( n7525 , n7523 , n7524 );
xor ( n7526 , n7522 , n7525 );
buf ( n7527 , n7526 );
and ( n7528 , n7421 , n7423 );
and ( n7529 , n7423 , n7461 );
and ( n7530 , n7421 , n7461 );
or ( n7531 , n7528 , n7529 , n7530 );
and ( n7532 , n7438 , n7442 );
and ( n7533 , n7442 , n7460 );
and ( n7534 , n7438 , n7460 );
or ( n7535 , n7532 , n7533 , n7534 );
buf ( n7536 , n855 );
buf ( n7537 , n7536 );
xor ( n7538 , n7535 , n7537 );
and ( n7539 , n7447 , n7451 );
and ( n7540 , n7451 , n7459 );
and ( n7541 , n7447 , n7459 );
or ( n7542 , n7539 , n7540 , n7541 );
and ( n7543 , n7427 , n6977 );
buf ( n7544 , n791 );
buf ( n7545 , n7544 );
and ( n7546 , n7545 , n6943 );
nor ( n7547 , n7543 , n7546 );
xnor ( n7548 , n7547 , n6974 );
and ( n7549 , n6980 , n7455 );
and ( n7550 , n7020 , n7344 );
nor ( n7551 , n7549 , n7550 );
xnor ( n7552 , n7551 , n7436 );
xor ( n7553 , n7548 , n7552 );
buf ( n7554 , n823 );
buf ( n7555 , n7554 );
xor ( n7556 , n7555 , n7433 );
and ( n7557 , n6941 , n7556 );
xor ( n7558 , n7553 , n7557 );
xor ( n7559 , n7542 , n7558 );
and ( n7560 , n7430 , n7437 );
and ( n7561 , n7241 , n7098 );
and ( n7562 , n7333 , n7026 );
nor ( n7563 , n7561 , n7562 );
xnor ( n7564 , n7563 , n7093 );
xor ( n7565 , n7560 , n7564 );
and ( n7566 , n7084 , n7260 );
and ( n7567 , n7156 , n7167 );
nor ( n7568 , n7566 , n7567 );
xnor ( n7569 , n7568 , n7250 );
xor ( n7570 , n7565 , n7569 );
xor ( n7571 , n7559 , n7570 );
xor ( n7572 , n7538 , n7571 );
xor ( n7573 , n7531 , n7572 );
and ( n7574 , n7462 , n7466 );
and ( n7575 , n7467 , n7470 );
or ( n7576 , n7574 , n7575 );
xor ( n7577 , n7573 , n7576 );
buf ( n7578 , n7577 );
not ( n7579 , n831 );
and ( n7580 , n7579 , n7527 );
and ( n7581 , n7578 , n831 );
or ( n7582 , n7580 , n7581 );
and ( n7583 , n7491 , n7507 );
and ( n7584 , n7507 , n7519 );
and ( n7585 , n7491 , n7519 );
or ( n7586 , n7583 , n7584 , n7585 );
buf ( n7587 , n886 );
buf ( n7588 , n7587 );
xor ( n7589 , n7586 , n7588 );
and ( n7590 , n7509 , n7513 );
and ( n7591 , n7513 , n7518 );
and ( n7592 , n7509 , n7518 );
or ( n7593 , n7590 , n7591 , n7592 );
and ( n7594 , n7494 , n6957 );
buf ( n7595 , n790 );
buf ( n7596 , n7595 );
and ( n7597 , n7596 , n6934 );
nor ( n7598 , n7594 , n7597 );
xnor ( n7599 , n7598 , n6954 );
and ( n7600 , n6999 , n7400 );
and ( n7601 , n7049 , n7303 );
nor ( n7602 , n7600 , n7601 );
xnor ( n7603 , n7602 , n7381 );
xor ( n7604 , n7599 , n7603 );
buf ( n7605 , n822 );
buf ( n7606 , n7605 );
xor ( n7607 , n7606 , n7504 );
not ( n7608 , n7505 );
and ( n7609 , n7607 , n7608 );
and ( n7610 , n6932 , n7609 );
and ( n7611 , n6960 , n7505 );
nor ( n7612 , n7610 , n7611 );
and ( n7613 , n7504 , n7378 );
not ( n7614 , n7613 );
and ( n7615 , n7606 , n7614 );
xnor ( n7616 , n7612 , n7615 );
xor ( n7617 , n7604 , n7616 );
xor ( n7618 , n7593 , n7617 );
and ( n7619 , n7292 , n7063 );
and ( n7620 , n7372 , n7005 );
nor ( n7621 , n7619 , n7620 );
xnor ( n7622 , n7621 , n7058 );
not ( n7623 , n7506 );
and ( n7624 , n7623 , n7615 );
xor ( n7625 , n7622 , n7624 );
and ( n7626 , n7497 , n7501 );
and ( n7627 , n7501 , n7506 );
and ( n7628 , n7497 , n7506 );
or ( n7629 , n7626 , n7627 , n7628 );
xor ( n7630 , n7625 , n7629 );
and ( n7631 , n7125 , n7215 );
and ( n7632 , n7196 , n7136 );
nor ( n7633 , n7631 , n7632 );
xnor ( n7634 , n7633 , n7205 );
xor ( n7635 , n7630 , n7634 );
xor ( n7636 , n7618 , n7635 );
xor ( n7637 , n7589 , n7636 );
and ( n7638 , n7484 , n7486 );
and ( n7639 , n7486 , n7520 );
and ( n7640 , n7484 , n7520 );
or ( n7641 , n7638 , n7639 , n7640 );
xor ( n7642 , n7637 , n7641 );
and ( n7643 , n7480 , n7521 );
and ( n7644 , n7522 , n7525 );
or ( n7645 , n7643 , n7644 );
xor ( n7646 , n7642 , n7645 );
buf ( n7647 , n7646 );
and ( n7648 , n7542 , n7558 );
and ( n7649 , n7558 , n7570 );
and ( n7650 , n7542 , n7570 );
or ( n7651 , n7648 , n7649 , n7650 );
buf ( n7652 , n854 );
buf ( n7653 , n7652 );
xor ( n7654 , n7651 , n7653 );
and ( n7655 , n7560 , n7564 );
and ( n7656 , n7564 , n7569 );
and ( n7657 , n7560 , n7569 );
or ( n7658 , n7655 , n7656 , n7657 );
and ( n7659 , n7545 , n6977 );
buf ( n7660 , n790 );
buf ( n7661 , n7660 );
and ( n7662 , n7661 , n6943 );
nor ( n7663 , n7659 , n7662 );
xnor ( n7664 , n7663 , n6974 );
and ( n7665 , n7020 , n7455 );
and ( n7666 , n7084 , n7344 );
nor ( n7667 , n7665 , n7666 );
xnor ( n7668 , n7667 , n7436 );
xor ( n7669 , n7664 , n7668 );
buf ( n7670 , n822 );
buf ( n7671 , n7670 );
xor ( n7672 , n7671 , n7555 );
not ( n7673 , n7556 );
and ( n7674 , n7672 , n7673 );
and ( n7675 , n6941 , n7674 );
and ( n7676 , n6980 , n7556 );
nor ( n7677 , n7675 , n7676 );
and ( n7678 , n7555 , n7433 );
not ( n7679 , n7678 );
and ( n7680 , n7671 , n7679 );
xnor ( n7681 , n7677 , n7680 );
xor ( n7682 , n7669 , n7681 );
xor ( n7683 , n7658 , n7682 );
and ( n7684 , n7333 , n7098 );
and ( n7685 , n7427 , n7026 );
nor ( n7686 , n7684 , n7685 );
xnor ( n7687 , n7686 , n7093 );
not ( n7688 , n7557 );
and ( n7689 , n7688 , n7680 );
xor ( n7690 , n7687 , n7689 );
and ( n7691 , n7548 , n7552 );
and ( n7692 , n7552 , n7557 );
and ( n7693 , n7548 , n7557 );
or ( n7694 , n7691 , n7692 , n7693 );
xor ( n7695 , n7690 , n7694 );
and ( n7696 , n7156 , n7260 );
and ( n7697 , n7241 , n7167 );
nor ( n7698 , n7696 , n7697 );
xnor ( n7699 , n7698 , n7250 );
xor ( n7700 , n7695 , n7699 );
xor ( n7701 , n7683 , n7700 );
xor ( n7702 , n7654 , n7701 );
and ( n7703 , n7535 , n7537 );
and ( n7704 , n7537 , n7571 );
and ( n7705 , n7535 , n7571 );
or ( n7706 , n7703 , n7704 , n7705 );
xor ( n7707 , n7702 , n7706 );
and ( n7708 , n7531 , n7572 );
and ( n7709 , n7573 , n7576 );
or ( n7710 , n7708 , n7709 );
xor ( n7711 , n7707 , n7710 );
buf ( n7712 , n7711 );
not ( n7713 , n831 );
and ( n7714 , n7713 , n7647 );
and ( n7715 , n7712 , n831 );
or ( n7716 , n7714 , n7715 );
and ( n7717 , n7593 , n7617 );
and ( n7718 , n7617 , n7635 );
and ( n7719 , n7593 , n7635 );
or ( n7720 , n7717 , n7718 , n7719 );
buf ( n7721 , n885 );
buf ( n7722 , n7721 );
xor ( n7723 , n7720 , n7722 );
and ( n7724 , n7625 , n7629 );
and ( n7725 , n7629 , n7634 );
and ( n7726 , n7625 , n7634 );
or ( n7727 , n7724 , n7725 , n7726 );
and ( n7728 , n7596 , n6957 );
buf ( n7729 , n789 );
buf ( n7730 , n7729 );
and ( n7731 , n7730 , n6934 );
nor ( n7732 , n7728 , n7731 );
xnor ( n7733 , n7732 , n6954 );
and ( n7734 , n7196 , n7215 );
and ( n7735 , n7292 , n7136 );
nor ( n7736 , n7734 , n7735 );
xnor ( n7737 , n7736 , n7205 );
xor ( n7738 , n7733 , n7737 );
and ( n7739 , n6960 , n7609 );
and ( n7740 , n6999 , n7505 );
nor ( n7741 , n7739 , n7740 );
xnor ( n7742 , n7741 , n7615 );
xor ( n7743 , n7738 , n7742 );
xor ( n7744 , n7727 , n7743 );
and ( n7745 , n7599 , n7603 );
and ( n7746 , n7603 , n7616 );
and ( n7747 , n7599 , n7616 );
or ( n7748 , n7745 , n7746 , n7747 );
and ( n7749 , n7622 , n7624 );
xor ( n7750 , n7748 , n7749 );
and ( n7751 , n7372 , n7063 );
and ( n7752 , n7494 , n7005 );
nor ( n7753 , n7751 , n7752 );
xnor ( n7754 , n7753 , n7058 );
and ( n7755 , n7049 , n7400 );
and ( n7756 , n7125 , n7303 );
nor ( n7757 , n7755 , n7756 );
xnor ( n7758 , n7757 , n7381 );
xor ( n7759 , n7754 , n7758 );
buf ( n7760 , n821 );
buf ( n7761 , n7760 );
xor ( n7762 , n7761 , n7606 );
and ( n7763 , n6932 , n7762 );
xor ( n7764 , n7759 , n7763 );
xor ( n7765 , n7750 , n7764 );
xor ( n7766 , n7744 , n7765 );
xor ( n7767 , n7723 , n7766 );
and ( n7768 , n7586 , n7588 );
and ( n7769 , n7588 , n7636 );
and ( n7770 , n7586 , n7636 );
or ( n7771 , n7768 , n7769 , n7770 );
xor ( n7772 , n7767 , n7771 );
and ( n7773 , n7637 , n7641 );
and ( n7774 , n7642 , n7645 );
or ( n7775 , n7773 , n7774 );
xor ( n7776 , n7772 , n7775 );
buf ( n7777 , n7776 );
and ( n7778 , n7658 , n7682 );
and ( n7779 , n7682 , n7700 );
and ( n7780 , n7658 , n7700 );
or ( n7781 , n7778 , n7779 , n7780 );
buf ( n7782 , n853 );
buf ( n7783 , n7782 );
xor ( n7784 , n7781 , n7783 );
and ( n7785 , n7690 , n7694 );
and ( n7786 , n7694 , n7699 );
and ( n7787 , n7690 , n7699 );
or ( n7788 , n7785 , n7786 , n7787 );
and ( n7789 , n7661 , n6977 );
buf ( n7790 , n789 );
buf ( n7791 , n7790 );
and ( n7792 , n7791 , n6943 );
nor ( n7793 , n7789 , n7792 );
xnor ( n7794 , n7793 , n6974 );
and ( n7795 , n7241 , n7260 );
and ( n7796 , n7333 , n7167 );
nor ( n7797 , n7795 , n7796 );
xnor ( n7798 , n7797 , n7250 );
xor ( n7799 , n7794 , n7798 );
and ( n7800 , n6980 , n7674 );
and ( n7801 , n7020 , n7556 );
nor ( n7802 , n7800 , n7801 );
xnor ( n7803 , n7802 , n7680 );
xor ( n7804 , n7799 , n7803 );
xor ( n7805 , n7788 , n7804 );
and ( n7806 , n7664 , n7668 );
and ( n7807 , n7668 , n7681 );
and ( n7808 , n7664 , n7681 );
or ( n7809 , n7806 , n7807 , n7808 );
and ( n7810 , n7687 , n7689 );
xor ( n7811 , n7809 , n7810 );
and ( n7812 , n7427 , n7098 );
and ( n7813 , n7545 , n7026 );
nor ( n7814 , n7812 , n7813 );
xnor ( n7815 , n7814 , n7093 );
and ( n7816 , n7084 , n7455 );
and ( n7817 , n7156 , n7344 );
nor ( n7818 , n7816 , n7817 );
xnor ( n7819 , n7818 , n7436 );
xor ( n7820 , n7815 , n7819 );
buf ( n7821 , n821 );
buf ( n7822 , n7821 );
xor ( n7823 , n7822 , n7671 );
and ( n7824 , n6941 , n7823 );
xor ( n7825 , n7820 , n7824 );
xor ( n7826 , n7811 , n7825 );
xor ( n7827 , n7805 , n7826 );
xor ( n7828 , n7784 , n7827 );
and ( n7829 , n7651 , n7653 );
and ( n7830 , n7653 , n7701 );
and ( n7831 , n7651 , n7701 );
or ( n7832 , n7829 , n7830 , n7831 );
xor ( n7833 , n7828 , n7832 );
and ( n7834 , n7702 , n7706 );
and ( n7835 , n7707 , n7710 );
or ( n7836 , n7834 , n7835 );
xor ( n7837 , n7833 , n7836 );
buf ( n7838 , n7837 );
not ( n7839 , n831 );
and ( n7840 , n7839 , n7777 );
and ( n7841 , n7838 , n831 );
or ( n7842 , n7840 , n7841 );
and ( n7843 , n7727 , n7743 );
and ( n7844 , n7743 , n7765 );
and ( n7845 , n7727 , n7765 );
or ( n7846 , n7843 , n7844 , n7845 );
buf ( n7847 , n884 );
buf ( n7848 , n7847 );
xor ( n7849 , n7846 , n7848 );
and ( n7850 , n7748 , n7749 );
and ( n7851 , n7749 , n7764 );
and ( n7852 , n7748 , n7764 );
or ( n7853 , n7850 , n7851 , n7852 );
and ( n7854 , n7494 , n7063 );
and ( n7855 , n7596 , n7005 );
nor ( n7856 , n7854 , n7855 );
xnor ( n7857 , n7856 , n7058 );
not ( n7858 , n7763 );
buf ( n7859 , n820 );
buf ( n7860 , n7859 );
and ( n7861 , n7761 , n7606 );
not ( n7862 , n7861 );
and ( n7863 , n7860 , n7862 );
and ( n7864 , n7858 , n7863 );
xor ( n7865 , n7857 , n7864 );
and ( n7866 , n7292 , n7215 );
and ( n7867 , n7372 , n7136 );
nor ( n7868 , n7866 , n7867 );
xnor ( n7869 , n7868 , n7205 );
xor ( n7870 , n7865 , n7869 );
xor ( n7871 , n7860 , n7761 );
not ( n7872 , n7762 );
and ( n7873 , n7871 , n7872 );
and ( n7874 , n6932 , n7873 );
and ( n7875 , n6960 , n7762 );
nor ( n7876 , n7874 , n7875 );
xnor ( n7877 , n7876 , n7863 );
xor ( n7878 , n7870 , n7877 );
xor ( n7879 , n7853 , n7878 );
and ( n7880 , n7754 , n7758 );
and ( n7881 , n7758 , n7763 );
and ( n7882 , n7754 , n7763 );
or ( n7883 , n7880 , n7881 , n7882 );
and ( n7884 , n7733 , n7737 );
and ( n7885 , n7737 , n7742 );
and ( n7886 , n7733 , n7742 );
or ( n7887 , n7884 , n7885 , n7886 );
xor ( n7888 , n7883 , n7887 );
and ( n7889 , n7730 , n6957 );
buf ( n7890 , n788 );
buf ( n7891 , n7890 );
and ( n7892 , n7891 , n6934 );
nor ( n7893 , n7889 , n7892 );
xnor ( n7894 , n7893 , n6954 );
and ( n7895 , n7125 , n7400 );
and ( n7896 , n7196 , n7303 );
nor ( n7897 , n7895 , n7896 );
xnor ( n7898 , n7897 , n7381 );
xor ( n7899 , n7894 , n7898 );
and ( n7900 , n6999 , n7609 );
and ( n7901 , n7049 , n7505 );
nor ( n7902 , n7900 , n7901 );
xnor ( n7903 , n7902 , n7615 );
xor ( n7904 , n7899 , n7903 );
xor ( n7905 , n7888 , n7904 );
xor ( n7906 , n7879 , n7905 );
xor ( n7907 , n7849 , n7906 );
and ( n7908 , n7720 , n7722 );
and ( n7909 , n7722 , n7766 );
and ( n7910 , n7720 , n7766 );
or ( n7911 , n7908 , n7909 , n7910 );
xor ( n7912 , n7907 , n7911 );
and ( n7913 , n7767 , n7771 );
and ( n7914 , n7772 , n7775 );
or ( n7915 , n7913 , n7914 );
xor ( n7916 , n7912 , n7915 );
buf ( n7917 , n7916 );
and ( n7918 , n7788 , n7804 );
and ( n7919 , n7804 , n7826 );
and ( n7920 , n7788 , n7826 );
or ( n7921 , n7918 , n7919 , n7920 );
buf ( n7922 , n852 );
buf ( n7923 , n7922 );
xor ( n7924 , n7921 , n7923 );
and ( n7925 , n7809 , n7810 );
and ( n7926 , n7810 , n7825 );
and ( n7927 , n7809 , n7825 );
or ( n7928 , n7925 , n7926 , n7927 );
and ( n7929 , n7545 , n7098 );
and ( n7930 , n7661 , n7026 );
nor ( n7931 , n7929 , n7930 );
xnor ( n7932 , n7931 , n7093 );
not ( n7933 , n7824 );
buf ( n7934 , n820 );
buf ( n7935 , n7934 );
and ( n7936 , n7822 , n7671 );
not ( n7937 , n7936 );
and ( n7938 , n7935 , n7937 );
and ( n7939 , n7933 , n7938 );
xor ( n7940 , n7932 , n7939 );
and ( n7941 , n7333 , n7260 );
and ( n7942 , n7427 , n7167 );
nor ( n7943 , n7941 , n7942 );
xnor ( n7944 , n7943 , n7250 );
xor ( n7945 , n7940 , n7944 );
xor ( n7946 , n7935 , n7822 );
not ( n7947 , n7823 );
and ( n7948 , n7946 , n7947 );
and ( n7949 , n6941 , n7948 );
and ( n7950 , n6980 , n7823 );
nor ( n7951 , n7949 , n7950 );
xnor ( n7952 , n7951 , n7938 );
xor ( n7953 , n7945 , n7952 );
xor ( n7954 , n7928 , n7953 );
and ( n7955 , n7815 , n7819 );
and ( n7956 , n7819 , n7824 );
and ( n7957 , n7815 , n7824 );
or ( n7958 , n7955 , n7956 , n7957 );
and ( n7959 , n7794 , n7798 );
and ( n7960 , n7798 , n7803 );
and ( n7961 , n7794 , n7803 );
or ( n7962 , n7959 , n7960 , n7961 );
xor ( n7963 , n7958 , n7962 );
and ( n7964 , n7791 , n6977 );
buf ( n7965 , n788 );
buf ( n7966 , n7965 );
and ( n7967 , n7966 , n6943 );
nor ( n7968 , n7964 , n7967 );
xnor ( n7969 , n7968 , n6974 );
and ( n7970 , n7156 , n7455 );
and ( n7971 , n7241 , n7344 );
nor ( n7972 , n7970 , n7971 );
xnor ( n7973 , n7972 , n7436 );
xor ( n7974 , n7969 , n7973 );
and ( n7975 , n7020 , n7674 );
and ( n7976 , n7084 , n7556 );
nor ( n7977 , n7975 , n7976 );
xnor ( n7978 , n7977 , n7680 );
xor ( n7979 , n7974 , n7978 );
xor ( n7980 , n7963 , n7979 );
xor ( n7981 , n7954 , n7980 );
xor ( n7982 , n7924 , n7981 );
and ( n7983 , n7781 , n7783 );
and ( n7984 , n7783 , n7827 );
and ( n7985 , n7781 , n7827 );
or ( n7986 , n7983 , n7984 , n7985 );
xor ( n7987 , n7982 , n7986 );
and ( n7988 , n7828 , n7832 );
and ( n7989 , n7833 , n7836 );
or ( n7990 , n7988 , n7989 );
xor ( n7991 , n7987 , n7990 );
buf ( n7992 , n7991 );
not ( n7993 , n831 );
and ( n7994 , n7993 , n7917 );
and ( n7995 , n7992 , n831 );
or ( n7996 , n7994 , n7995 );
and ( n7997 , n7846 , n7848 );
and ( n7998 , n7848 , n7906 );
and ( n7999 , n7846 , n7906 );
or ( n8000 , n7997 , n7998 , n7999 );
and ( n8001 , n7853 , n7878 );
and ( n8002 , n7878 , n7905 );
and ( n8003 , n7853 , n7905 );
or ( n8004 , n8001 , n8002 , n8003 );
buf ( n8005 , n883 );
buf ( n8006 , n8005 );
xor ( n8007 , n8004 , n8006 );
and ( n8008 , n7883 , n7887 );
and ( n8009 , n7887 , n7904 );
and ( n8010 , n7883 , n7904 );
or ( n8011 , n8008 , n8009 , n8010 );
and ( n8012 , n7894 , n7898 );
and ( n8013 , n7898 , n7903 );
and ( n8014 , n7894 , n7903 );
or ( n8015 , n8012 , n8013 , n8014 );
and ( n8016 , n7857 , n7864 );
xor ( n8017 , n8015 , n8016 );
and ( n8018 , n7372 , n7215 );
and ( n8019 , n7494 , n7136 );
nor ( n8020 , n8018 , n8019 );
xnor ( n8021 , n8020 , n7205 );
xor ( n8022 , n8017 , n8021 );
xor ( n8023 , n8011 , n8022 );
and ( n8024 , n7865 , n7869 );
and ( n8025 , n7869 , n7877 );
and ( n8026 , n7865 , n7877 );
or ( n8027 , n8024 , n8025 , n8026 );
and ( n8028 , n7596 , n7063 );
and ( n8029 , n7730 , n7005 );
nor ( n8030 , n8028 , n8029 );
xnor ( n8031 , n8030 , n7058 );
and ( n8032 , n7196 , n7400 );
and ( n8033 , n7292 , n7303 );
nor ( n8034 , n8032 , n8033 );
xnor ( n8035 , n8034 , n7381 );
xor ( n8036 , n8031 , n8035 );
buf ( n8037 , n819 );
buf ( n8038 , n8037 );
xor ( n8039 , n8038 , n7860 );
and ( n8040 , n6932 , n8039 );
xor ( n8041 , n8036 , n8040 );
xor ( n8042 , n8027 , n8041 );
and ( n8043 , n7891 , n6957 );
buf ( n8044 , n787 );
buf ( n8045 , n8044 );
and ( n8046 , n8045 , n6934 );
nor ( n8047 , n8043 , n8046 );
xnor ( n8048 , n8047 , n6954 );
and ( n8049 , n7049 , n7609 );
and ( n8050 , n7125 , n7505 );
nor ( n8051 , n8049 , n8050 );
xnor ( n8052 , n8051 , n7615 );
xor ( n8053 , n8048 , n8052 );
and ( n8054 , n6960 , n7873 );
and ( n8055 , n6999 , n7762 );
nor ( n8056 , n8054 , n8055 );
xnor ( n8057 , n8056 , n7863 );
xor ( n8058 , n8053 , n8057 );
xor ( n8059 , n8042 , n8058 );
xor ( n8060 , n8023 , n8059 );
xor ( n8061 , n8007 , n8060 );
xor ( n8062 , n8000 , n8061 );
and ( n8063 , n7907 , n7911 );
and ( n8064 , n7912 , n7915 );
or ( n8065 , n8063 , n8064 );
xor ( n8066 , n8062 , n8065 );
buf ( n8067 , n8066 );
and ( n8068 , n7921 , n7923 );
and ( n8069 , n7923 , n7981 );
and ( n8070 , n7921 , n7981 );
or ( n8071 , n8068 , n8069 , n8070 );
and ( n8072 , n7928 , n7953 );
and ( n8073 , n7953 , n7980 );
and ( n8074 , n7928 , n7980 );
or ( n8075 , n8072 , n8073 , n8074 );
buf ( n8076 , n851 );
buf ( n8077 , n8076 );
xor ( n8078 , n8075 , n8077 );
and ( n8079 , n7958 , n7962 );
and ( n8080 , n7962 , n7979 );
and ( n8081 , n7958 , n7979 );
or ( n8082 , n8079 , n8080 , n8081 );
and ( n8083 , n7969 , n7973 );
and ( n8084 , n7973 , n7978 );
and ( n8085 , n7969 , n7978 );
or ( n8086 , n8083 , n8084 , n8085 );
and ( n8087 , n7932 , n7939 );
xor ( n8088 , n8086 , n8087 );
and ( n8089 , n7427 , n7260 );
and ( n8090 , n7545 , n7167 );
nor ( n8091 , n8089 , n8090 );
xnor ( n8092 , n8091 , n7250 );
xor ( n8093 , n8088 , n8092 );
xor ( n8094 , n8082 , n8093 );
and ( n8095 , n7940 , n7944 );
and ( n8096 , n7944 , n7952 );
and ( n8097 , n7940 , n7952 );
or ( n8098 , n8095 , n8096 , n8097 );
and ( n8099 , n7661 , n7098 );
and ( n8100 , n7791 , n7026 );
nor ( n8101 , n8099 , n8100 );
xnor ( n8102 , n8101 , n7093 );
and ( n8103 , n7241 , n7455 );
and ( n8104 , n7333 , n7344 );
nor ( n8105 , n8103 , n8104 );
xnor ( n8106 , n8105 , n7436 );
xor ( n8107 , n8102 , n8106 );
buf ( n8108 , n819 );
buf ( n8109 , n8108 );
xor ( n8110 , n8109 , n7935 );
and ( n8111 , n6941 , n8110 );
xor ( n8112 , n8107 , n8111 );
xor ( n8113 , n8098 , n8112 );
and ( n8114 , n7966 , n6977 );
buf ( n8115 , n787 );
buf ( n8116 , n8115 );
and ( n8117 , n8116 , n6943 );
nor ( n8118 , n8114 , n8117 );
xnor ( n8119 , n8118 , n6974 );
and ( n8120 , n7084 , n7674 );
and ( n8121 , n7156 , n7556 );
nor ( n8122 , n8120 , n8121 );
xnor ( n8123 , n8122 , n7680 );
xor ( n8124 , n8119 , n8123 );
and ( n8125 , n6980 , n7948 );
and ( n8126 , n7020 , n7823 );
nor ( n8127 , n8125 , n8126 );
xnor ( n8128 , n8127 , n7938 );
xor ( n8129 , n8124 , n8128 );
xor ( n8130 , n8113 , n8129 );
xor ( n8131 , n8094 , n8130 );
xor ( n8132 , n8078 , n8131 );
xor ( n8133 , n8071 , n8132 );
and ( n8134 , n7982 , n7986 );
and ( n8135 , n7987 , n7990 );
or ( n8136 , n8134 , n8135 );
xor ( n8137 , n8133 , n8136 );
buf ( n8138 , n8137 );
not ( n8139 , n831 );
and ( n8140 , n8139 , n8067 );
and ( n8141 , n8138 , n831 );
or ( n8142 , n8140 , n8141 );
and ( n8143 , n8011 , n8022 );
and ( n8144 , n8022 , n8059 );
and ( n8145 , n8011 , n8059 );
or ( n8146 , n8143 , n8144 , n8145 );
buf ( n8147 , n882 );
buf ( n8148 , n8147 );
xor ( n8149 , n8146 , n8148 );
and ( n8150 , n8027 , n8041 );
and ( n8151 , n8041 , n8058 );
and ( n8152 , n8027 , n8058 );
or ( n8153 , n8150 , n8151 , n8152 );
and ( n8154 , n8045 , n6957 );
buf ( n8155 , n786 );
buf ( n8156 , n8155 );
and ( n8157 , n8156 , n6934 );
nor ( n8158 , n8154 , n8157 );
xnor ( n8159 , n8158 , n6954 );
not ( n8160 , n8040 );
buf ( n8161 , n818 );
buf ( n8162 , n8161 );
and ( n8163 , n8038 , n7860 );
not ( n8164 , n8163 );
and ( n8165 , n8162 , n8164 );
and ( n8166 , n8160 , n8165 );
xor ( n8167 , n8159 , n8166 );
and ( n8168 , n8031 , n8035 );
and ( n8169 , n8035 , n8040 );
and ( n8170 , n8031 , n8040 );
or ( n8171 , n8168 , n8169 , n8170 );
xor ( n8172 , n8167 , n8171 );
and ( n8173 , n8048 , n8052 );
and ( n8174 , n8052 , n8057 );
and ( n8175 , n8048 , n8057 );
or ( n8176 , n8173 , n8174 , n8175 );
xor ( n8177 , n8172 , n8176 );
xor ( n8178 , n8153 , n8177 );
and ( n8179 , n8015 , n8016 );
and ( n8180 , n8016 , n8021 );
and ( n8181 , n8015 , n8021 );
or ( n8182 , n8179 , n8180 , n8181 );
and ( n8183 , n7730 , n7063 );
and ( n8184 , n7891 , n7005 );
nor ( n8185 , n8183 , n8184 );
xnor ( n8186 , n8185 , n7058 );
and ( n8187 , n7292 , n7400 );
and ( n8188 , n7372 , n7303 );
nor ( n8189 , n8187 , n8188 );
xnor ( n8190 , n8189 , n7381 );
xor ( n8191 , n8186 , n8190 );
and ( n8192 , n7125 , n7609 );
and ( n8193 , n7196 , n7505 );
nor ( n8194 , n8192 , n8193 );
xnor ( n8195 , n8194 , n7615 );
xor ( n8196 , n8191 , n8195 );
xor ( n8197 , n8182 , n8196 );
and ( n8198 , n7494 , n7215 );
and ( n8199 , n7596 , n7136 );
nor ( n8200 , n8198 , n8199 );
xnor ( n8201 , n8200 , n7205 );
and ( n8202 , n6999 , n7873 );
and ( n8203 , n7049 , n7762 );
nor ( n8204 , n8202 , n8203 );
xnor ( n8205 , n8204 , n7863 );
xor ( n8206 , n8201 , n8205 );
xor ( n8207 , n8162 , n8038 );
not ( n8208 , n8039 );
and ( n8209 , n8207 , n8208 );
and ( n8210 , n6932 , n8209 );
and ( n8211 , n6960 , n8039 );
nor ( n8212 , n8210 , n8211 );
xnor ( n8213 , n8212 , n8165 );
xor ( n8214 , n8206 , n8213 );
xor ( n8215 , n8197 , n8214 );
xor ( n8216 , n8178 , n8215 );
xor ( n8217 , n8149 , n8216 );
and ( n8218 , n8004 , n8006 );
and ( n8219 , n8006 , n8060 );
and ( n8220 , n8004 , n8060 );
or ( n8221 , n8218 , n8219 , n8220 );
xor ( n8222 , n8217 , n8221 );
and ( n8223 , n8000 , n8061 );
and ( n8224 , n8062 , n8065 );
or ( n8225 , n8223 , n8224 );
xor ( n8226 , n8222 , n8225 );
buf ( n8227 , n8226 );
and ( n8228 , n8082 , n8093 );
and ( n8229 , n8093 , n8130 );
and ( n8230 , n8082 , n8130 );
or ( n8231 , n8228 , n8229 , n8230 );
buf ( n8232 , n850 );
buf ( n8233 , n8232 );
xor ( n8234 , n8231 , n8233 );
and ( n8235 , n8098 , n8112 );
and ( n8236 , n8112 , n8129 );
and ( n8237 , n8098 , n8129 );
or ( n8238 , n8235 , n8236 , n8237 );
and ( n8239 , n8116 , n6977 );
buf ( n8240 , n786 );
buf ( n8241 , n8240 );
and ( n8242 , n8241 , n6943 );
nor ( n8243 , n8239 , n8242 );
xnor ( n8244 , n8243 , n6974 );
not ( n8245 , n8111 );
buf ( n8246 , n818 );
buf ( n8247 , n8246 );
and ( n8248 , n8109 , n7935 );
not ( n8249 , n8248 );
and ( n8250 , n8247 , n8249 );
and ( n8251 , n8245 , n8250 );
xor ( n8252 , n8244 , n8251 );
and ( n8253 , n8102 , n8106 );
and ( n8254 , n8106 , n8111 );
and ( n8255 , n8102 , n8111 );
or ( n8256 , n8253 , n8254 , n8255 );
xor ( n8257 , n8252 , n8256 );
and ( n8258 , n8119 , n8123 );
and ( n8259 , n8123 , n8128 );
and ( n8260 , n8119 , n8128 );
or ( n8261 , n8258 , n8259 , n8260 );
xor ( n8262 , n8257 , n8261 );
xor ( n8263 , n8238 , n8262 );
and ( n8264 , n8086 , n8087 );
and ( n8265 , n8087 , n8092 );
and ( n8266 , n8086 , n8092 );
or ( n8267 , n8264 , n8265 , n8266 );
and ( n8268 , n7791 , n7098 );
and ( n8269 , n7966 , n7026 );
nor ( n8270 , n8268 , n8269 );
xnor ( n8271 , n8270 , n7093 );
and ( n8272 , n7333 , n7455 );
and ( n8273 , n7427 , n7344 );
nor ( n8274 , n8272 , n8273 );
xnor ( n8275 , n8274 , n7436 );
xor ( n8276 , n8271 , n8275 );
and ( n8277 , n7156 , n7674 );
and ( n8278 , n7241 , n7556 );
nor ( n8279 , n8277 , n8278 );
xnor ( n8280 , n8279 , n7680 );
xor ( n8281 , n8276 , n8280 );
xor ( n8282 , n8267 , n8281 );
and ( n8283 , n7545 , n7260 );
and ( n8284 , n7661 , n7167 );
nor ( n8285 , n8283 , n8284 );
xnor ( n8286 , n8285 , n7250 );
and ( n8287 , n7020 , n7948 );
and ( n8288 , n7084 , n7823 );
nor ( n8289 , n8287 , n8288 );
xnor ( n8290 , n8289 , n7938 );
xor ( n8291 , n8286 , n8290 );
xor ( n8292 , n8247 , n8109 );
not ( n8293 , n8110 );
and ( n8294 , n8292 , n8293 );
and ( n8295 , n6941 , n8294 );
and ( n8296 , n6980 , n8110 );
nor ( n8297 , n8295 , n8296 );
xnor ( n8298 , n8297 , n8250 );
xor ( n8299 , n8291 , n8298 );
xor ( n8300 , n8282 , n8299 );
xor ( n8301 , n8263 , n8300 );
xor ( n8302 , n8234 , n8301 );
and ( n8303 , n8075 , n8077 );
and ( n8304 , n8077 , n8131 );
and ( n8305 , n8075 , n8131 );
or ( n8306 , n8303 , n8304 , n8305 );
xor ( n8307 , n8302 , n8306 );
and ( n8308 , n8071 , n8132 );
and ( n8309 , n8133 , n8136 );
or ( n8310 , n8308 , n8309 );
xor ( n8311 , n8307 , n8310 );
buf ( n8312 , n8311 );
not ( n8313 , n831 );
and ( n8314 , n8313 , n8227 );
and ( n8315 , n8312 , n831 );
or ( n8316 , n8314 , n8315 );
and ( n8317 , n8153 , n8177 );
and ( n8318 , n8177 , n8215 );
and ( n8319 , n8153 , n8215 );
or ( n8320 , n8317 , n8318 , n8319 );
buf ( n8321 , n881 );
buf ( n8322 , n8321 );
xor ( n8323 , n8320 , n8322 );
and ( n8324 , n8182 , n8196 );
and ( n8325 , n8196 , n8214 );
and ( n8326 , n8182 , n8214 );
or ( n8327 , n8324 , n8325 , n8326 );
and ( n8328 , n8186 , n8190 );
and ( n8329 , n8190 , n8195 );
and ( n8330 , n8186 , n8195 );
or ( n8331 , n8328 , n8329 , n8330 );
and ( n8332 , n8201 , n8205 );
and ( n8333 , n8205 , n8213 );
and ( n8334 , n8201 , n8213 );
or ( n8335 , n8332 , n8333 , n8334 );
xor ( n8336 , n8331 , n8335 );
and ( n8337 , n8156 , n6957 );
buf ( n8338 , n785 );
buf ( n8339 , n8338 );
and ( n8340 , n8339 , n6934 );
nor ( n8341 , n8337 , n8340 );
xnor ( n8342 , n8341 , n6954 );
and ( n8343 , n7891 , n7063 );
and ( n8344 , n8045 , n7005 );
nor ( n8345 , n8343 , n8344 );
xnor ( n8346 , n8345 , n7058 );
xor ( n8347 , n8342 , n8346 );
buf ( n8348 , n817 );
buf ( n8349 , n8348 );
xor ( n8350 , n8349 , n8162 );
and ( n8351 , n6932 , n8350 );
xor ( n8352 , n8347 , n8351 );
xor ( n8353 , n8336 , n8352 );
xor ( n8354 , n8327 , n8353 );
and ( n8355 , n8167 , n8171 );
and ( n8356 , n8171 , n8176 );
and ( n8357 , n8167 , n8176 );
or ( n8358 , n8355 , n8356 , n8357 );
and ( n8359 , n7596 , n7215 );
and ( n8360 , n7730 , n7136 );
nor ( n8361 , n8359 , n8360 );
xnor ( n8362 , n8361 , n7205 );
and ( n8363 , n7372 , n7400 );
and ( n8364 , n7494 , n7303 );
nor ( n8365 , n8363 , n8364 );
xnor ( n8366 , n8365 , n7381 );
xor ( n8367 , n8362 , n8366 );
and ( n8368 , n7196 , n7609 );
and ( n8369 , n7292 , n7505 );
nor ( n8370 , n8368 , n8369 );
xnor ( n8371 , n8370 , n7615 );
xor ( n8372 , n8367 , n8371 );
xor ( n8373 , n8358 , n8372 );
and ( n8374 , n8159 , n8166 );
and ( n8375 , n7049 , n7873 );
and ( n8376 , n7125 , n7762 );
nor ( n8377 , n8375 , n8376 );
xnor ( n8378 , n8377 , n7863 );
xor ( n8379 , n8374 , n8378 );
and ( n8380 , n6960 , n8209 );
and ( n8381 , n6999 , n8039 );
nor ( n8382 , n8380 , n8381 );
xnor ( n8383 , n8382 , n8165 );
xor ( n8384 , n8379 , n8383 );
xor ( n8385 , n8373 , n8384 );
xor ( n8386 , n8354 , n8385 );
xor ( n8387 , n8323 , n8386 );
and ( n8388 , n8146 , n8148 );
and ( n8389 , n8148 , n8216 );
and ( n8390 , n8146 , n8216 );
or ( n8391 , n8388 , n8389 , n8390 );
xor ( n8392 , n8387 , n8391 );
and ( n8393 , n8217 , n8221 );
and ( n8394 , n8222 , n8225 );
or ( n8395 , n8393 , n8394 );
xor ( n8396 , n8392 , n8395 );
buf ( n8397 , n8396 );
and ( n8398 , n8238 , n8262 );
and ( n8399 , n8262 , n8300 );
and ( n8400 , n8238 , n8300 );
or ( n8401 , n8398 , n8399 , n8400 );
buf ( n8402 , n849 );
buf ( n8403 , n8402 );
xor ( n8404 , n8401 , n8403 );
and ( n8405 , n8267 , n8281 );
and ( n8406 , n8281 , n8299 );
and ( n8407 , n8267 , n8299 );
or ( n8408 , n8405 , n8406 , n8407 );
and ( n8409 , n8271 , n8275 );
and ( n8410 , n8275 , n8280 );
and ( n8411 , n8271 , n8280 );
or ( n8412 , n8409 , n8410 , n8411 );
and ( n8413 , n8286 , n8290 );
and ( n8414 , n8290 , n8298 );
and ( n8415 , n8286 , n8298 );
or ( n8416 , n8413 , n8414 , n8415 );
xor ( n8417 , n8412 , n8416 );
and ( n8418 , n8241 , n6977 );
buf ( n8419 , n785 );
buf ( n8420 , n8419 );
and ( n8421 , n8420 , n6943 );
nor ( n8422 , n8418 , n8421 );
xnor ( n8423 , n8422 , n6974 );
and ( n8424 , n7966 , n7098 );
and ( n8425 , n8116 , n7026 );
nor ( n8426 , n8424 , n8425 );
xnor ( n8427 , n8426 , n7093 );
xor ( n8428 , n8423 , n8427 );
buf ( n8429 , n817 );
buf ( n8430 , n8429 );
xor ( n8431 , n8430 , n8247 );
and ( n8432 , n6941 , n8431 );
xor ( n8433 , n8428 , n8432 );
xor ( n8434 , n8417 , n8433 );
xor ( n8435 , n8408 , n8434 );
and ( n8436 , n8252 , n8256 );
and ( n8437 , n8256 , n8261 );
and ( n8438 , n8252 , n8261 );
or ( n8439 , n8436 , n8437 , n8438 );
and ( n8440 , n7661 , n7260 );
and ( n8441 , n7791 , n7167 );
nor ( n8442 , n8440 , n8441 );
xnor ( n8443 , n8442 , n7250 );
and ( n8444 , n7427 , n7455 );
and ( n8445 , n7545 , n7344 );
nor ( n8446 , n8444 , n8445 );
xnor ( n8447 , n8446 , n7436 );
xor ( n8448 , n8443 , n8447 );
and ( n8449 , n7241 , n7674 );
and ( n8450 , n7333 , n7556 );
nor ( n8451 , n8449 , n8450 );
xnor ( n8452 , n8451 , n7680 );
xor ( n8453 , n8448 , n8452 );
xor ( n8454 , n8439 , n8453 );
and ( n8455 , n8244 , n8251 );
and ( n8456 , n7084 , n7948 );
and ( n8457 , n7156 , n7823 );
nor ( n8458 , n8456 , n8457 );
xnor ( n8459 , n8458 , n7938 );
xor ( n8460 , n8455 , n8459 );
and ( n8461 , n6980 , n8294 );
and ( n8462 , n7020 , n8110 );
nor ( n8463 , n8461 , n8462 );
xnor ( n8464 , n8463 , n8250 );
xor ( n8465 , n8460 , n8464 );
xor ( n8466 , n8454 , n8465 );
xor ( n8467 , n8435 , n8466 );
xor ( n8468 , n8404 , n8467 );
and ( n8469 , n8231 , n8233 );
and ( n8470 , n8233 , n8301 );
and ( n8471 , n8231 , n8301 );
or ( n8472 , n8469 , n8470 , n8471 );
xor ( n8473 , n8468 , n8472 );
and ( n8474 , n8302 , n8306 );
and ( n8475 , n8307 , n8310 );
or ( n8476 , n8474 , n8475 );
xor ( n8477 , n8473 , n8476 );
buf ( n8478 , n8477 );
not ( n8479 , n831 );
and ( n8480 , n8479 , n8397 );
and ( n8481 , n8478 , n831 );
or ( n8482 , n8480 , n8481 );
and ( n8483 , n8327 , n8353 );
and ( n8484 , n8353 , n8385 );
and ( n8485 , n8327 , n8385 );
or ( n8486 , n8483 , n8484 , n8485 );
buf ( n8487 , n880 );
buf ( n8488 , n8487 );
xor ( n8489 , n8486 , n8488 );
and ( n8490 , n8358 , n8372 );
and ( n8491 , n8372 , n8384 );
and ( n8492 , n8358 , n8384 );
or ( n8493 , n8490 , n8491 , n8492 );
and ( n8494 , n8362 , n8366 );
and ( n8495 , n8366 , n8371 );
and ( n8496 , n8362 , n8371 );
or ( n8497 , n8494 , n8495 , n8496 );
and ( n8498 , n8045 , n7063 );
and ( n8499 , n8156 , n7005 );
nor ( n8500 , n8498 , n8499 );
xnor ( n8501 , n8500 , n7058 );
and ( n8502 , n7494 , n7400 );
and ( n8503 , n7596 , n7303 );
nor ( n8504 , n8502 , n8503 );
xnor ( n8505 , n8504 , n7381 );
xor ( n8506 , n8501 , n8505 );
buf ( n8507 , n816 );
buf ( n8508 , n8507 );
xor ( n8509 , n8508 , n8349 );
not ( n8510 , n8350 );
and ( n8511 , n8509 , n8510 );
and ( n8512 , n6932 , n8511 );
and ( n8513 , n6960 , n8350 );
nor ( n8514 , n8512 , n8513 );
and ( n8515 , n8349 , n8162 );
not ( n8516 , n8515 );
and ( n8517 , n8508 , n8516 );
xnor ( n8518 , n8514 , n8517 );
xor ( n8519 , n8506 , n8518 );
xor ( n8520 , n8497 , n8519 );
and ( n8521 , n7730 , n7215 );
and ( n8522 , n7891 , n7136 );
nor ( n8523 , n8521 , n8522 );
xnor ( n8524 , n8523 , n7205 );
and ( n8525 , n7292 , n7609 );
and ( n8526 , n7372 , n7505 );
nor ( n8527 , n8525 , n8526 );
xnor ( n8528 , n8527 , n7615 );
xor ( n8529 , n8524 , n8528 );
and ( n8530 , n7125 , n7873 );
and ( n8531 , n7196 , n7762 );
nor ( n8532 , n8530 , n8531 );
xnor ( n8533 , n8532 , n7863 );
xor ( n8534 , n8529 , n8533 );
xor ( n8535 , n8520 , n8534 );
xor ( n8536 , n8493 , n8535 );
and ( n8537 , n8374 , n8378 );
and ( n8538 , n8378 , n8383 );
and ( n8539 , n8374 , n8383 );
or ( n8540 , n8537 , n8538 , n8539 );
and ( n8541 , n8331 , n8335 );
and ( n8542 , n8335 , n8352 );
and ( n8543 , n8331 , n8352 );
or ( n8544 , n8541 , n8542 , n8543 );
xor ( n8545 , n8540 , n8544 );
and ( n8546 , n8339 , n6957 );
buf ( n8547 , n784 );
buf ( n8548 , n8547 );
and ( n8549 , n8548 , n6934 );
nor ( n8550 , n8546 , n8549 );
xnor ( n8551 , n8550 , n6954 );
not ( n8552 , n8351 );
and ( n8553 , n8552 , n8517 );
xor ( n8554 , n8551 , n8553 );
and ( n8555 , n8342 , n8346 );
and ( n8556 , n8346 , n8351 );
and ( n8557 , n8342 , n8351 );
or ( n8558 , n8555 , n8556 , n8557 );
xor ( n8559 , n8554 , n8558 );
and ( n8560 , n6999 , n8209 );
and ( n8561 , n7049 , n8039 );
nor ( n8562 , n8560 , n8561 );
xnor ( n8563 , n8562 , n8165 );
xor ( n8564 , n8559 , n8563 );
xor ( n8565 , n8545 , n8564 );
xor ( n8566 , n8536 , n8565 );
xor ( n8567 , n8489 , n8566 );
and ( n8568 , n8320 , n8322 );
and ( n8569 , n8322 , n8386 );
and ( n8570 , n8320 , n8386 );
or ( n8571 , n8568 , n8569 , n8570 );
xor ( n8572 , n8567 , n8571 );
and ( n8573 , n8387 , n8391 );
and ( n8574 , n8392 , n8395 );
or ( n8575 , n8573 , n8574 );
xor ( n8576 , n8572 , n8575 );
buf ( n8577 , n8576 );
and ( n8578 , n8408 , n8434 );
and ( n8579 , n8434 , n8466 );
and ( n8580 , n8408 , n8466 );
or ( n8581 , n8578 , n8579 , n8580 );
buf ( n8582 , n848 );
buf ( n8583 , n8582 );
xor ( n8584 , n8581 , n8583 );
and ( n8585 , n8439 , n8453 );
and ( n8586 , n8453 , n8465 );
and ( n8587 , n8439 , n8465 );
or ( n8588 , n8585 , n8586 , n8587 );
and ( n8589 , n8443 , n8447 );
and ( n8590 , n8447 , n8452 );
and ( n8591 , n8443 , n8452 );
or ( n8592 , n8589 , n8590 , n8591 );
and ( n8593 , n8116 , n7098 );
and ( n8594 , n8241 , n7026 );
nor ( n8595 , n8593 , n8594 );
xnor ( n8596 , n8595 , n7093 );
and ( n8597 , n7545 , n7455 );
and ( n8598 , n7661 , n7344 );
nor ( n8599 , n8597 , n8598 );
xnor ( n8600 , n8599 , n7436 );
xor ( n8601 , n8596 , n8600 );
buf ( n8602 , n816 );
buf ( n8603 , n8602 );
xor ( n8604 , n8603 , n8430 );
not ( n8605 , n8431 );
and ( n8606 , n8604 , n8605 );
and ( n8607 , n6941 , n8606 );
and ( n8608 , n6980 , n8431 );
nor ( n8609 , n8607 , n8608 );
and ( n8610 , n8430 , n8247 );
not ( n8611 , n8610 );
and ( n8612 , n8603 , n8611 );
xnor ( n8613 , n8609 , n8612 );
xor ( n8614 , n8601 , n8613 );
xor ( n8615 , n8592 , n8614 );
and ( n8616 , n7791 , n7260 );
and ( n8617 , n7966 , n7167 );
nor ( n8618 , n8616 , n8617 );
xnor ( n8619 , n8618 , n7250 );
and ( n8620 , n7333 , n7674 );
and ( n8621 , n7427 , n7556 );
nor ( n8622 , n8620 , n8621 );
xnor ( n8623 , n8622 , n7680 );
xor ( n8624 , n8619 , n8623 );
and ( n8625 , n7156 , n7948 );
and ( n8626 , n7241 , n7823 );
nor ( n8627 , n8625 , n8626 );
xnor ( n8628 , n8627 , n7938 );
xor ( n8629 , n8624 , n8628 );
xor ( n8630 , n8615 , n8629 );
xor ( n8631 , n8588 , n8630 );
and ( n8632 , n8455 , n8459 );
and ( n8633 , n8459 , n8464 );
and ( n8634 , n8455 , n8464 );
or ( n8635 , n8632 , n8633 , n8634 );
and ( n8636 , n8412 , n8416 );
and ( n8637 , n8416 , n8433 );
and ( n8638 , n8412 , n8433 );
or ( n8639 , n8636 , n8637 , n8638 );
xor ( n8640 , n8635 , n8639 );
and ( n8641 , n8420 , n6977 );
buf ( n8642 , n784 );
buf ( n8643 , n8642 );
and ( n8644 , n8643 , n6943 );
nor ( n8645 , n8641 , n8644 );
xnor ( n8646 , n8645 , n6974 );
not ( n8647 , n8432 );
and ( n8648 , n8647 , n8612 );
xor ( n8649 , n8646 , n8648 );
and ( n8650 , n8423 , n8427 );
and ( n8651 , n8427 , n8432 );
and ( n8652 , n8423 , n8432 );
or ( n8653 , n8650 , n8651 , n8652 );
xor ( n8654 , n8649 , n8653 );
and ( n8655 , n7020 , n8294 );
and ( n8656 , n7084 , n8110 );
nor ( n8657 , n8655 , n8656 );
xnor ( n8658 , n8657 , n8250 );
xor ( n8659 , n8654 , n8658 );
xor ( n8660 , n8640 , n8659 );
xor ( n8661 , n8631 , n8660 );
xor ( n8662 , n8584 , n8661 );
and ( n8663 , n8401 , n8403 );
and ( n8664 , n8403 , n8467 );
and ( n8665 , n8401 , n8467 );
or ( n8666 , n8663 , n8664 , n8665 );
xor ( n8667 , n8662 , n8666 );
and ( n8668 , n8468 , n8472 );
and ( n8669 , n8473 , n8476 );
or ( n8670 , n8668 , n8669 );
xor ( n8671 , n8667 , n8670 );
buf ( n8672 , n8671 );
not ( n8673 , n831 );
and ( n8674 , n8673 , n8577 );
and ( n8675 , n8672 , n831 );
or ( n8676 , n8674 , n8675 );
and ( n8677 , n8493 , n8535 );
and ( n8678 , n8535 , n8565 );
and ( n8679 , n8493 , n8565 );
or ( n8680 , n8677 , n8678 , n8679 );
buf ( n8681 , n879 );
buf ( n8682 , n8681 );
xor ( n8683 , n8680 , n8682 );
and ( n8684 , n8540 , n8544 );
and ( n8685 , n8544 , n8564 );
and ( n8686 , n8540 , n8564 );
or ( n8687 , n8684 , n8685 , n8686 );
and ( n8688 , n8548 , n6957 );
buf ( n8689 , n783 );
buf ( n8690 , n8689 );
and ( n8691 , n8690 , n6934 );
nor ( n8692 , n8688 , n8691 );
xnor ( n8693 , n8692 , n6954 );
and ( n8694 , n8156 , n7063 );
and ( n8695 , n8339 , n7005 );
nor ( n8696 , n8694 , n8695 );
xnor ( n8697 , n8696 , n7058 );
xor ( n8698 , n8693 , n8697 );
buf ( n8699 , n815 );
buf ( n8700 , n8699 );
xor ( n8701 , n8700 , n8508 );
and ( n8702 , n6932 , n8701 );
xor ( n8703 , n8698 , n8702 );
and ( n8704 , n7891 , n7215 );
and ( n8705 , n8045 , n7136 );
nor ( n8706 , n8704 , n8705 );
xnor ( n8707 , n8706 , n7205 );
and ( n8708 , n7196 , n7873 );
and ( n8709 , n7292 , n7762 );
nor ( n8710 , n8708 , n8709 );
xnor ( n8711 , n8710 , n7863 );
xor ( n8712 , n8707 , n8711 );
and ( n8713 , n7049 , n8209 );
and ( n8714 , n7125 , n8039 );
nor ( n8715 , n8713 , n8714 );
xnor ( n8716 , n8715 , n8165 );
xor ( n8717 , n8712 , n8716 );
xor ( n8718 , n8703 , n8717 );
and ( n8719 , n7596 , n7400 );
and ( n8720 , n7730 , n7303 );
nor ( n8721 , n8719 , n8720 );
xnor ( n8722 , n8721 , n7381 );
and ( n8723 , n7372 , n7609 );
and ( n8724 , n7494 , n7505 );
nor ( n8725 , n8723 , n8724 );
xnor ( n8726 , n8725 , n7615 );
xor ( n8727 , n8722 , n8726 );
and ( n8728 , n6960 , n8511 );
and ( n8729 , n6999 , n8350 );
nor ( n8730 , n8728 , n8729 );
xnor ( n8731 , n8730 , n8517 );
xor ( n8732 , n8727 , n8731 );
xor ( n8733 , n8718 , n8732 );
xor ( n8734 , n8687 , n8733 );
and ( n8735 , n8554 , n8558 );
and ( n8736 , n8558 , n8563 );
and ( n8737 , n8554 , n8563 );
or ( n8738 , n8735 , n8736 , n8737 );
and ( n8739 , n8497 , n8519 );
and ( n8740 , n8519 , n8534 );
and ( n8741 , n8497 , n8534 );
or ( n8742 , n8739 , n8740 , n8741 );
xor ( n8743 , n8738 , n8742 );
and ( n8744 , n8501 , n8505 );
and ( n8745 , n8505 , n8518 );
and ( n8746 , n8501 , n8518 );
or ( n8747 , n8744 , n8745 , n8746 );
and ( n8748 , n8524 , n8528 );
and ( n8749 , n8528 , n8533 );
and ( n8750 , n8524 , n8533 );
or ( n8751 , n8748 , n8749 , n8750 );
xor ( n8752 , n8747 , n8751 );
and ( n8753 , n8551 , n8553 );
xor ( n8754 , n8752 , n8753 );
xor ( n8755 , n8743 , n8754 );
xor ( n8756 , n8734 , n8755 );
xor ( n8757 , n8683 , n8756 );
and ( n8758 , n8486 , n8488 );
and ( n8759 , n8488 , n8566 );
and ( n8760 , n8486 , n8566 );
or ( n8761 , n8758 , n8759 , n8760 );
xor ( n8762 , n8757 , n8761 );
and ( n8763 , n8567 , n8571 );
and ( n8764 , n8572 , n8575 );
or ( n8765 , n8763 , n8764 );
xor ( n8766 , n8762 , n8765 );
buf ( n8767 , n8766 );
and ( n8768 , n8588 , n8630 );
and ( n8769 , n8630 , n8660 );
and ( n8770 , n8588 , n8660 );
or ( n8771 , n8768 , n8769 , n8770 );
buf ( n8772 , n847 );
buf ( n8773 , n8772 );
xor ( n8774 , n8771 , n8773 );
and ( n8775 , n8635 , n8639 );
and ( n8776 , n8639 , n8659 );
and ( n8777 , n8635 , n8659 );
or ( n8778 , n8775 , n8776 , n8777 );
and ( n8779 , n8643 , n6977 );
buf ( n8780 , n783 );
buf ( n8781 , n8780 );
and ( n8782 , n8781 , n6943 );
nor ( n8783 , n8779 , n8782 );
xnor ( n8784 , n8783 , n6974 );
and ( n8785 , n8241 , n7098 );
and ( n8786 , n8420 , n7026 );
nor ( n8787 , n8785 , n8786 );
xnor ( n8788 , n8787 , n7093 );
xor ( n8789 , n8784 , n8788 );
buf ( n8790 , n815 );
buf ( n8791 , n8790 );
xor ( n8792 , n8791 , n8603 );
and ( n8793 , n6941 , n8792 );
xor ( n8794 , n8789 , n8793 );
and ( n8795 , n7966 , n7260 );
and ( n8796 , n8116 , n7167 );
nor ( n8797 , n8795 , n8796 );
xnor ( n8798 , n8797 , n7250 );
and ( n8799 , n7241 , n7948 );
and ( n8800 , n7333 , n7823 );
nor ( n8801 , n8799 , n8800 );
xnor ( n8802 , n8801 , n7938 );
xor ( n8803 , n8798 , n8802 );
and ( n8804 , n7084 , n8294 );
and ( n8805 , n7156 , n8110 );
nor ( n8806 , n8804 , n8805 );
xnor ( n8807 , n8806 , n8250 );
xor ( n8808 , n8803 , n8807 );
xor ( n8809 , n8794 , n8808 );
and ( n8810 , n7661 , n7455 );
and ( n8811 , n7791 , n7344 );
nor ( n8812 , n8810 , n8811 );
xnor ( n8813 , n8812 , n7436 );
and ( n8814 , n7427 , n7674 );
and ( n8815 , n7545 , n7556 );
nor ( n8816 , n8814 , n8815 );
xnor ( n8817 , n8816 , n7680 );
xor ( n8818 , n8813 , n8817 );
and ( n8819 , n6980 , n8606 );
and ( n8820 , n7020 , n8431 );
nor ( n8821 , n8819 , n8820 );
xnor ( n8822 , n8821 , n8612 );
xor ( n8823 , n8818 , n8822 );
xor ( n8824 , n8809 , n8823 );
xor ( n8825 , n8778 , n8824 );
and ( n8826 , n8649 , n8653 );
and ( n8827 , n8653 , n8658 );
and ( n8828 , n8649 , n8658 );
or ( n8829 , n8826 , n8827 , n8828 );
and ( n8830 , n8592 , n8614 );
and ( n8831 , n8614 , n8629 );
and ( n8832 , n8592 , n8629 );
or ( n8833 , n8830 , n8831 , n8832 );
xor ( n8834 , n8829 , n8833 );
and ( n8835 , n8596 , n8600 );
and ( n8836 , n8600 , n8613 );
and ( n8837 , n8596 , n8613 );
or ( n8838 , n8835 , n8836 , n8837 );
and ( n8839 , n8619 , n8623 );
and ( n8840 , n8623 , n8628 );
and ( n8841 , n8619 , n8628 );
or ( n8842 , n8839 , n8840 , n8841 );
xor ( n8843 , n8838 , n8842 );
and ( n8844 , n8646 , n8648 );
xor ( n8845 , n8843 , n8844 );
xor ( n8846 , n8834 , n8845 );
xor ( n8847 , n8825 , n8846 );
xor ( n8848 , n8774 , n8847 );
and ( n8849 , n8581 , n8583 );
and ( n8850 , n8583 , n8661 );
and ( n8851 , n8581 , n8661 );
or ( n8852 , n8849 , n8850 , n8851 );
xor ( n8853 , n8848 , n8852 );
and ( n8854 , n8662 , n8666 );
and ( n8855 , n8667 , n8670 );
or ( n8856 , n8854 , n8855 );
xor ( n8857 , n8853 , n8856 );
buf ( n8858 , n8857 );
not ( n8859 , n831 );
and ( n8860 , n8859 , n8767 );
and ( n8861 , n8858 , n831 );
or ( n8862 , n8860 , n8861 );
and ( n8863 , n8687 , n8733 );
and ( n8864 , n8733 , n8755 );
and ( n8865 , n8687 , n8755 );
or ( n8866 , n8863 , n8864 , n8865 );
buf ( n8867 , n878 );
buf ( n8868 , n8867 );
xor ( n8869 , n8866 , n8868 );
and ( n8870 , n8738 , n8742 );
and ( n8871 , n8742 , n8754 );
and ( n8872 , n8738 , n8754 );
or ( n8873 , n8870 , n8871 , n8872 );
and ( n8874 , n7730 , n7400 );
and ( n8875 , n7891 , n7303 );
nor ( n8876 , n8874 , n8875 );
xnor ( n8877 , n8876 , n7381 );
and ( n8878 , n6999 , n8511 );
and ( n8879 , n7049 , n8350 );
nor ( n8880 , n8878 , n8879 );
xnor ( n8881 , n8880 , n8517 );
xor ( n8882 , n8877 , n8881 );
buf ( n8883 , n814 );
buf ( n8884 , n8883 );
xor ( n8885 , n8884 , n8700 );
not ( n8886 , n8701 );
and ( n8887 , n8885 , n8886 );
and ( n8888 , n6932 , n8887 );
and ( n8889 , n6960 , n8701 );
nor ( n8890 , n8888 , n8889 );
and ( n8891 , n8700 , n8508 );
not ( n8892 , n8891 );
and ( n8893 , n8884 , n8892 );
xnor ( n8894 , n8890 , n8893 );
xor ( n8895 , n8882 , n8894 );
and ( n8896 , n8339 , n7063 );
and ( n8897 , n8548 , n7005 );
nor ( n8898 , n8896 , n8897 );
xnor ( n8899 , n8898 , n7058 );
and ( n8900 , n8045 , n7215 );
and ( n8901 , n8156 , n7136 );
nor ( n8902 , n8900 , n8901 );
xnor ( n8903 , n8902 , n7205 );
xor ( n8904 , n8899 , n8903 );
and ( n8905 , n7494 , n7609 );
and ( n8906 , n7596 , n7505 );
nor ( n8907 , n8905 , n8906 );
xnor ( n8908 , n8907 , n7615 );
xor ( n8909 , n8904 , n8908 );
xor ( n8910 , n8895 , n8909 );
and ( n8911 , n8690 , n6957 );
buf ( n8912 , n782 );
buf ( n8913 , n8912 );
and ( n8914 , n8913 , n6934 );
nor ( n8915 , n8911 , n8914 );
xnor ( n8916 , n8915 , n6954 );
not ( n8917 , n8702 );
and ( n8918 , n8917 , n8893 );
xor ( n8919 , n8916 , n8918 );
and ( n8920 , n7292 , n7873 );
and ( n8921 , n7372 , n7762 );
nor ( n8922 , n8920 , n8921 );
xnor ( n8923 , n8922 , n7863 );
xor ( n8924 , n8919 , n8923 );
and ( n8925 , n7125 , n8209 );
and ( n8926 , n7196 , n8039 );
nor ( n8927 , n8925 , n8926 );
xnor ( n8928 , n8927 , n8165 );
xor ( n8929 , n8924 , n8928 );
xor ( n8930 , n8910 , n8929 );
xor ( n8931 , n8873 , n8930 );
and ( n8932 , n8747 , n8751 );
and ( n8933 , n8751 , n8753 );
and ( n8934 , n8747 , n8753 );
or ( n8935 , n8932 , n8933 , n8934 );
and ( n8936 , n8703 , n8717 );
and ( n8937 , n8717 , n8732 );
and ( n8938 , n8703 , n8732 );
or ( n8939 , n8936 , n8937 , n8938 );
xor ( n8940 , n8935 , n8939 );
and ( n8941 , n8693 , n8697 );
and ( n8942 , n8697 , n8702 );
and ( n8943 , n8693 , n8702 );
or ( n8944 , n8941 , n8942 , n8943 );
and ( n8945 , n8707 , n8711 );
and ( n8946 , n8711 , n8716 );
and ( n8947 , n8707 , n8716 );
or ( n8948 , n8945 , n8946 , n8947 );
xor ( n8949 , n8944 , n8948 );
and ( n8950 , n8722 , n8726 );
and ( n8951 , n8726 , n8731 );
and ( n8952 , n8722 , n8731 );
or ( n8953 , n8950 , n8951 , n8952 );
xor ( n8954 , n8949 , n8953 );
xor ( n8955 , n8940 , n8954 );
xor ( n8956 , n8931 , n8955 );
xor ( n8957 , n8869 , n8956 );
and ( n8958 , n8680 , n8682 );
and ( n8959 , n8682 , n8756 );
and ( n8960 , n8680 , n8756 );
or ( n8961 , n8958 , n8959 , n8960 );
xor ( n8962 , n8957 , n8961 );
and ( n8963 , n8757 , n8761 );
and ( n8964 , n8762 , n8765 );
or ( n8965 , n8963 , n8964 );
xor ( n8966 , n8962 , n8965 );
buf ( n8967 , n8966 );
and ( n8968 , n8778 , n8824 );
and ( n8969 , n8824 , n8846 );
and ( n8970 , n8778 , n8846 );
or ( n8971 , n8968 , n8969 , n8970 );
buf ( n8972 , n846 );
buf ( n8973 , n8972 );
xor ( n8974 , n8971 , n8973 );
and ( n8975 , n8829 , n8833 );
and ( n8976 , n8833 , n8845 );
and ( n8977 , n8829 , n8845 );
or ( n8978 , n8975 , n8976 , n8977 );
and ( n8979 , n7791 , n7455 );
and ( n8980 , n7966 , n7344 );
nor ( n8981 , n8979 , n8980 );
xnor ( n8982 , n8981 , n7436 );
and ( n8983 , n7020 , n8606 );
and ( n8984 , n7084 , n8431 );
nor ( n8985 , n8983 , n8984 );
xnor ( n8986 , n8985 , n8612 );
xor ( n8987 , n8982 , n8986 );
buf ( n8988 , n814 );
buf ( n8989 , n8988 );
xor ( n8990 , n8989 , n8791 );
not ( n8991 , n8792 );
and ( n8992 , n8990 , n8991 );
and ( n8993 , n6941 , n8992 );
and ( n8994 , n6980 , n8792 );
nor ( n8995 , n8993 , n8994 );
and ( n8996 , n8791 , n8603 );
not ( n8997 , n8996 );
and ( n8998 , n8989 , n8997 );
xnor ( n8999 , n8995 , n8998 );
xor ( n9000 , n8987 , n8999 );
and ( n9001 , n8420 , n7098 );
and ( n9002 , n8643 , n7026 );
nor ( n9003 , n9001 , n9002 );
xnor ( n9004 , n9003 , n7093 );
and ( n9005 , n8116 , n7260 );
and ( n9006 , n8241 , n7167 );
nor ( n9007 , n9005 , n9006 );
xnor ( n9008 , n9007 , n7250 );
xor ( n9009 , n9004 , n9008 );
and ( n9010 , n7545 , n7674 );
and ( n9011 , n7661 , n7556 );
nor ( n9012 , n9010 , n9011 );
xnor ( n9013 , n9012 , n7680 );
xor ( n9014 , n9009 , n9013 );
xor ( n9015 , n9000 , n9014 );
and ( n9016 , n8781 , n6977 );
buf ( n9017 , n782 );
buf ( n9018 , n9017 );
and ( n9019 , n9018 , n6943 );
nor ( n9020 , n9016 , n9019 );
xnor ( n9021 , n9020 , n6974 );
not ( n9022 , n8793 );
and ( n9023 , n9022 , n8998 );
xor ( n9024 , n9021 , n9023 );
and ( n9025 , n7333 , n7948 );
and ( n9026 , n7427 , n7823 );
nor ( n9027 , n9025 , n9026 );
xnor ( n9028 , n9027 , n7938 );
xor ( n9029 , n9024 , n9028 );
and ( n9030 , n7156 , n8294 );
and ( n9031 , n7241 , n8110 );
nor ( n9032 , n9030 , n9031 );
xnor ( n9033 , n9032 , n8250 );
xor ( n9034 , n9029 , n9033 );
xor ( n9035 , n9015 , n9034 );
xor ( n9036 , n8978 , n9035 );
and ( n9037 , n8838 , n8842 );
and ( n9038 , n8842 , n8844 );
and ( n9039 , n8838 , n8844 );
or ( n9040 , n9037 , n9038 , n9039 );
and ( n9041 , n8794 , n8808 );
and ( n9042 , n8808 , n8823 );
and ( n9043 , n8794 , n8823 );
or ( n9044 , n9041 , n9042 , n9043 );
xor ( n9045 , n9040 , n9044 );
and ( n9046 , n8784 , n8788 );
and ( n9047 , n8788 , n8793 );
and ( n9048 , n8784 , n8793 );
or ( n9049 , n9046 , n9047 , n9048 );
and ( n9050 , n8798 , n8802 );
and ( n9051 , n8802 , n8807 );
and ( n9052 , n8798 , n8807 );
or ( n9053 , n9050 , n9051 , n9052 );
xor ( n9054 , n9049 , n9053 );
and ( n9055 , n8813 , n8817 );
and ( n9056 , n8817 , n8822 );
and ( n9057 , n8813 , n8822 );
or ( n9058 , n9055 , n9056 , n9057 );
xor ( n9059 , n9054 , n9058 );
xor ( n9060 , n9045 , n9059 );
xor ( n9061 , n9036 , n9060 );
xor ( n9062 , n8974 , n9061 );
and ( n9063 , n8771 , n8773 );
and ( n9064 , n8773 , n8847 );
and ( n9065 , n8771 , n8847 );
or ( n9066 , n9063 , n9064 , n9065 );
xor ( n9067 , n9062 , n9066 );
and ( n9068 , n8848 , n8852 );
and ( n9069 , n8853 , n8856 );
or ( n9070 , n9068 , n9069 );
xor ( n9071 , n9067 , n9070 );
buf ( n9072 , n9071 );
not ( n9073 , n831 );
and ( n9074 , n9073 , n8967 );
and ( n9075 , n9072 , n831 );
or ( n9076 , n9074 , n9075 );
and ( n9077 , n8866 , n8868 );
and ( n9078 , n8868 , n8956 );
and ( n9079 , n8866 , n8956 );
or ( n9080 , n9077 , n9078 , n9079 );
and ( n9081 , n8873 , n8930 );
and ( n9082 , n8930 , n8955 );
and ( n9083 , n8873 , n8955 );
or ( n9084 , n9081 , n9082 , n9083 );
buf ( n9085 , n877 );
buf ( n9086 , n9085 );
xor ( n9087 , n9084 , n9086 );
and ( n9088 , n8935 , n8939 );
and ( n9089 , n8939 , n8954 );
and ( n9090 , n8935 , n8954 );
or ( n9091 , n9088 , n9089 , n9090 );
and ( n9092 , n8919 , n8923 );
and ( n9093 , n8923 , n8928 );
and ( n9094 , n8919 , n8928 );
or ( n9095 , n9092 , n9093 , n9094 );
and ( n9096 , n8548 , n7063 );
and ( n9097 , n8690 , n7005 );
nor ( n9098 , n9096 , n9097 );
xnor ( n9099 , n9098 , n7058 );
and ( n9100 , n7049 , n8511 );
and ( n9101 , n7125 , n8350 );
nor ( n9102 , n9100 , n9101 );
xnor ( n9103 , n9102 , n8517 );
xor ( n9104 , n9099 , n9103 );
and ( n9105 , n6960 , n8887 );
and ( n9106 , n6999 , n8701 );
nor ( n9107 , n9105 , n9106 );
xnor ( n9108 , n9107 , n8893 );
xor ( n9109 , n9104 , n9108 );
xor ( n9110 , n9095 , n9109 );
and ( n9111 , n8877 , n8881 );
and ( n9112 , n8881 , n8894 );
and ( n9113 , n8877 , n8894 );
or ( n9114 , n9111 , n9112 , n9113 );
and ( n9115 , n8916 , n8918 );
xor ( n9116 , n9114 , n9115 );
and ( n9117 , n7196 , n8209 );
and ( n9118 , n7292 , n8039 );
nor ( n9119 , n9117 , n9118 );
xnor ( n9120 , n9119 , n8165 );
xor ( n9121 , n9116 , n9120 );
xor ( n9122 , n9110 , n9121 );
xor ( n9123 , n9091 , n9122 );
and ( n9124 , n8944 , n8948 );
and ( n9125 , n8948 , n8953 );
and ( n9126 , n8944 , n8953 );
or ( n9127 , n9124 , n9125 , n9126 );
and ( n9128 , n8895 , n8909 );
and ( n9129 , n8909 , n8929 );
and ( n9130 , n8895 , n8929 );
or ( n9131 , n9128 , n9129 , n9130 );
xor ( n9132 , n9127 , n9131 );
and ( n9133 , n8899 , n8903 );
and ( n9134 , n8903 , n8908 );
and ( n9135 , n8899 , n8908 );
or ( n9136 , n9133 , n9134 , n9135 );
and ( n9137 , n8913 , n6957 );
buf ( n9138 , n781 );
buf ( n9139 , n9138 );
and ( n9140 , n9139 , n6934 );
nor ( n9141 , n9137 , n9140 );
xnor ( n9142 , n9141 , n6954 );
and ( n9143 , n7891 , n7400 );
and ( n9144 , n8045 , n7303 );
nor ( n9145 , n9143 , n9144 );
xnor ( n9146 , n9145 , n7381 );
xor ( n9147 , n9142 , n9146 );
buf ( n9148 , n813 );
buf ( n9149 , n9148 );
xor ( n9150 , n9149 , n8884 );
and ( n9151 , n6932 , n9150 );
xor ( n9152 , n9147 , n9151 );
xor ( n9153 , n9136 , n9152 );
and ( n9154 , n8156 , n7215 );
and ( n9155 , n8339 , n7136 );
nor ( n9156 , n9154 , n9155 );
xnor ( n9157 , n9156 , n7205 );
and ( n9158 , n7596 , n7609 );
and ( n9159 , n7730 , n7505 );
nor ( n9160 , n9158 , n9159 );
xnor ( n9161 , n9160 , n7615 );
xor ( n9162 , n9157 , n9161 );
and ( n9163 , n7372 , n7873 );
and ( n9164 , n7494 , n7762 );
nor ( n9165 , n9163 , n9164 );
xnor ( n9166 , n9165 , n7863 );
xor ( n9167 , n9162 , n9166 );
xor ( n9168 , n9153 , n9167 );
xor ( n9169 , n9132 , n9168 );
xor ( n9170 , n9123 , n9169 );
xor ( n9171 , n9087 , n9170 );
xor ( n9172 , n9080 , n9171 );
and ( n9173 , n8957 , n8961 );
and ( n9174 , n8962 , n8965 );
or ( n9175 , n9173 , n9174 );
xor ( n9176 , n9172 , n9175 );
buf ( n9177 , n9176 );
and ( n9178 , n8971 , n8973 );
and ( n9179 , n8973 , n9061 );
and ( n9180 , n8971 , n9061 );
or ( n9181 , n9178 , n9179 , n9180 );
and ( n9182 , n8978 , n9035 );
and ( n9183 , n9035 , n9060 );
and ( n9184 , n8978 , n9060 );
or ( n9185 , n9182 , n9183 , n9184 );
buf ( n9186 , n845 );
buf ( n9187 , n9186 );
xor ( n9188 , n9185 , n9187 );
and ( n9189 , n9040 , n9044 );
and ( n9190 , n9044 , n9059 );
and ( n9191 , n9040 , n9059 );
or ( n9192 , n9189 , n9190 , n9191 );
and ( n9193 , n9024 , n9028 );
and ( n9194 , n9028 , n9033 );
and ( n9195 , n9024 , n9033 );
or ( n9196 , n9193 , n9194 , n9195 );
and ( n9197 , n8643 , n7098 );
and ( n9198 , n8781 , n7026 );
nor ( n9199 , n9197 , n9198 );
xnor ( n9200 , n9199 , n7093 );
and ( n9201 , n7084 , n8606 );
and ( n9202 , n7156 , n8431 );
nor ( n9203 , n9201 , n9202 );
xnor ( n9204 , n9203 , n8612 );
xor ( n9205 , n9200 , n9204 );
and ( n9206 , n6980 , n8992 );
and ( n9207 , n7020 , n8792 );
nor ( n9208 , n9206 , n9207 );
xnor ( n9209 , n9208 , n8998 );
xor ( n9210 , n9205 , n9209 );
xor ( n9211 , n9196 , n9210 );
and ( n9212 , n8982 , n8986 );
and ( n9213 , n8986 , n8999 );
and ( n9214 , n8982 , n8999 );
or ( n9215 , n9212 , n9213 , n9214 );
and ( n9216 , n9021 , n9023 );
xor ( n9217 , n9215 , n9216 );
and ( n9218 , n7241 , n8294 );
and ( n9219 , n7333 , n8110 );
nor ( n9220 , n9218 , n9219 );
xnor ( n9221 , n9220 , n8250 );
xor ( n9222 , n9217 , n9221 );
xor ( n9223 , n9211 , n9222 );
xor ( n9224 , n9192 , n9223 );
and ( n9225 , n9049 , n9053 );
and ( n9226 , n9053 , n9058 );
and ( n9227 , n9049 , n9058 );
or ( n9228 , n9225 , n9226 , n9227 );
and ( n9229 , n9000 , n9014 );
and ( n9230 , n9014 , n9034 );
and ( n9231 , n9000 , n9034 );
or ( n9232 , n9229 , n9230 , n9231 );
xor ( n9233 , n9228 , n9232 );
and ( n9234 , n9004 , n9008 );
and ( n9235 , n9008 , n9013 );
and ( n9236 , n9004 , n9013 );
or ( n9237 , n9234 , n9235 , n9236 );
and ( n9238 , n9018 , n6977 );
buf ( n9239 , n781 );
buf ( n9240 , n9239 );
and ( n9241 , n9240 , n6943 );
nor ( n9242 , n9238 , n9241 );
xnor ( n9243 , n9242 , n6974 );
and ( n9244 , n7966 , n7455 );
and ( n9245 , n8116 , n7344 );
nor ( n9246 , n9244 , n9245 );
xnor ( n9247 , n9246 , n7436 );
xor ( n9248 , n9243 , n9247 );
buf ( n9249 , n813 );
buf ( n9250 , n9249 );
xor ( n9251 , n9250 , n8989 );
and ( n9252 , n6941 , n9251 );
xor ( n9253 , n9248 , n9252 );
xor ( n9254 , n9237 , n9253 );
and ( n9255 , n8241 , n7260 );
and ( n9256 , n8420 , n7167 );
nor ( n9257 , n9255 , n9256 );
xnor ( n9258 , n9257 , n7250 );
and ( n9259 , n7661 , n7674 );
and ( n9260 , n7791 , n7556 );
nor ( n9261 , n9259 , n9260 );
xnor ( n9262 , n9261 , n7680 );
xor ( n9263 , n9258 , n9262 );
and ( n9264 , n7427 , n7948 );
and ( n9265 , n7545 , n7823 );
nor ( n9266 , n9264 , n9265 );
xnor ( n9267 , n9266 , n7938 );
xor ( n9268 , n9263 , n9267 );
xor ( n9269 , n9254 , n9268 );
xor ( n9270 , n9233 , n9269 );
xor ( n9271 , n9224 , n9270 );
xor ( n9272 , n9188 , n9271 );
xor ( n9273 , n9181 , n9272 );
and ( n9274 , n9062 , n9066 );
and ( n9275 , n9067 , n9070 );
or ( n9276 , n9274 , n9275 );
xor ( n9277 , n9273 , n9276 );
buf ( n9278 , n9277 );
not ( n9279 , n831 );
and ( n9280 , n9279 , n9177 );
and ( n9281 , n9278 , n831 );
or ( n9282 , n9280 , n9281 );
and ( n9283 , n9091 , n9122 );
and ( n9284 , n9122 , n9169 );
and ( n9285 , n9091 , n9169 );
or ( n9286 , n9283 , n9284 , n9285 );
buf ( n9287 , n876 );
buf ( n9288 , n9287 );
xor ( n9289 , n9286 , n9288 );
and ( n9290 , n9127 , n9131 );
and ( n9291 , n9131 , n9168 );
and ( n9292 , n9127 , n9168 );
or ( n9293 , n9290 , n9291 , n9292 );
and ( n9294 , n9114 , n9115 );
and ( n9295 , n9115 , n9120 );
and ( n9296 , n9114 , n9120 );
or ( n9297 , n9294 , n9295 , n9296 );
and ( n9298 , n8690 , n7063 );
and ( n9299 , n8913 , n7005 );
nor ( n9300 , n9298 , n9299 );
xnor ( n9301 , n9300 , n7058 );
and ( n9302 , n7730 , n7609 );
and ( n9303 , n7891 , n7505 );
nor ( n9304 , n9302 , n9303 );
xnor ( n9305 , n9304 , n7615 );
xor ( n9306 , n9301 , n9305 );
buf ( n9307 , n812 );
buf ( n9308 , n9307 );
xor ( n9309 , n9308 , n9149 );
not ( n9310 , n9150 );
and ( n9311 , n9309 , n9310 );
and ( n9312 , n6932 , n9311 );
and ( n9313 , n6960 , n9150 );
nor ( n9314 , n9312 , n9313 );
and ( n9315 , n9149 , n8884 );
not ( n9316 , n9315 );
and ( n9317 , n9308 , n9316 );
xnor ( n9318 , n9314 , n9317 );
xor ( n9319 , n9306 , n9318 );
xor ( n9320 , n9297 , n9319 );
and ( n9321 , n9139 , n6957 );
buf ( n9322 , n780 );
buf ( n9323 , n9322 );
and ( n9324 , n9323 , n6934 );
nor ( n9325 , n9321 , n9324 );
xnor ( n9326 , n9325 , n6954 );
not ( n9327 , n9151 );
and ( n9328 , n9327 , n9317 );
xor ( n9329 , n9326 , n9328 );
and ( n9330 , n9142 , n9146 );
and ( n9331 , n9146 , n9151 );
and ( n9332 , n9142 , n9151 );
or ( n9333 , n9330 , n9331 , n9332 );
xor ( n9334 , n9329 , n9333 );
and ( n9335 , n9099 , n9103 );
and ( n9336 , n9103 , n9108 );
and ( n9337 , n9099 , n9108 );
or ( n9338 , n9335 , n9336 , n9337 );
xor ( n9339 , n9334 , n9338 );
xor ( n9340 , n9320 , n9339 );
xor ( n9341 , n9293 , n9340 );
and ( n9342 , n9136 , n9152 );
and ( n9343 , n9152 , n9167 );
and ( n9344 , n9136 , n9167 );
or ( n9345 , n9342 , n9343 , n9344 );
and ( n9346 , n9095 , n9109 );
and ( n9347 , n9109 , n9121 );
and ( n9348 , n9095 , n9121 );
or ( n9349 , n9346 , n9347 , n9348 );
xor ( n9350 , n9345 , n9349 );
and ( n9351 , n9157 , n9161 );
and ( n9352 , n9161 , n9166 );
and ( n9353 , n9157 , n9166 );
or ( n9354 , n9351 , n9352 , n9353 );
and ( n9355 , n8045 , n7400 );
and ( n9356 , n8156 , n7303 );
nor ( n9357 , n9355 , n9356 );
xnor ( n9358 , n9357 , n7381 );
and ( n9359 , n7125 , n8511 );
and ( n9360 , n7196 , n8350 );
nor ( n9361 , n9359 , n9360 );
xnor ( n9362 , n9361 , n8517 );
xor ( n9363 , n9358 , n9362 );
and ( n9364 , n6999 , n8887 );
and ( n9365 , n7049 , n8701 );
nor ( n9366 , n9364 , n9365 );
xnor ( n9367 , n9366 , n8893 );
xor ( n9368 , n9363 , n9367 );
xor ( n9369 , n9354 , n9368 );
and ( n9370 , n8339 , n7215 );
and ( n9371 , n8548 , n7136 );
nor ( n9372 , n9370 , n9371 );
xnor ( n9373 , n9372 , n7205 );
and ( n9374 , n7494 , n7873 );
and ( n9375 , n7596 , n7762 );
nor ( n9376 , n9374 , n9375 );
xnor ( n9377 , n9376 , n7863 );
xor ( n9378 , n9373 , n9377 );
and ( n9379 , n7292 , n8209 );
and ( n9380 , n7372 , n8039 );
nor ( n9381 , n9379 , n9380 );
xnor ( n9382 , n9381 , n8165 );
xor ( n9383 , n9378 , n9382 );
xor ( n9384 , n9369 , n9383 );
xor ( n9385 , n9350 , n9384 );
xor ( n9386 , n9341 , n9385 );
xor ( n9387 , n9289 , n9386 );
and ( n9388 , n9084 , n9086 );
and ( n9389 , n9086 , n9170 );
and ( n9390 , n9084 , n9170 );
or ( n9391 , n9388 , n9389 , n9390 );
xor ( n9392 , n9387 , n9391 );
and ( n9393 , n9080 , n9171 );
and ( n9394 , n9172 , n9175 );
or ( n9395 , n9393 , n9394 );
xor ( n9396 , n9392 , n9395 );
buf ( n9397 , n9396 );
and ( n9398 , n9192 , n9223 );
and ( n9399 , n9223 , n9270 );
and ( n9400 , n9192 , n9270 );
or ( n9401 , n9398 , n9399 , n9400 );
buf ( n9402 , n844 );
buf ( n9403 , n9402 );
xor ( n9404 , n9401 , n9403 );
and ( n9405 , n9228 , n9232 );
and ( n9406 , n9232 , n9269 );
and ( n9407 , n9228 , n9269 );
or ( n9408 , n9405 , n9406 , n9407 );
and ( n9409 , n9215 , n9216 );
and ( n9410 , n9216 , n9221 );
and ( n9411 , n9215 , n9221 );
or ( n9412 , n9409 , n9410 , n9411 );
and ( n9413 , n8781 , n7098 );
and ( n9414 , n9018 , n7026 );
nor ( n9415 , n9413 , n9414 );
xnor ( n9416 , n9415 , n7093 );
and ( n9417 , n7791 , n7674 );
and ( n9418 , n7966 , n7556 );
nor ( n9419 , n9417 , n9418 );
xnor ( n9420 , n9419 , n7680 );
xor ( n9421 , n9416 , n9420 );
buf ( n9422 , n812 );
buf ( n9423 , n9422 );
xor ( n9424 , n9423 , n9250 );
not ( n9425 , n9251 );
and ( n9426 , n9424 , n9425 );
and ( n9427 , n6941 , n9426 );
and ( n9428 , n6980 , n9251 );
nor ( n9429 , n9427 , n9428 );
and ( n9430 , n9250 , n8989 );
not ( n9431 , n9430 );
and ( n9432 , n9423 , n9431 );
xnor ( n9433 , n9429 , n9432 );
xor ( n9434 , n9421 , n9433 );
xor ( n9435 , n9412 , n9434 );
and ( n9436 , n9240 , n6977 );
buf ( n9437 , n780 );
buf ( n9438 , n9437 );
and ( n9439 , n9438 , n6943 );
nor ( n9440 , n9436 , n9439 );
xnor ( n9441 , n9440 , n6974 );
not ( n9442 , n9252 );
and ( n9443 , n9442 , n9432 );
xor ( n9444 , n9441 , n9443 );
and ( n9445 , n9243 , n9247 );
and ( n9446 , n9247 , n9252 );
and ( n9447 , n9243 , n9252 );
or ( n9448 , n9445 , n9446 , n9447 );
xor ( n9449 , n9444 , n9448 );
and ( n9450 , n9200 , n9204 );
and ( n9451 , n9204 , n9209 );
and ( n9452 , n9200 , n9209 );
or ( n9453 , n9450 , n9451 , n9452 );
xor ( n9454 , n9449 , n9453 );
xor ( n9455 , n9435 , n9454 );
xor ( n9456 , n9408 , n9455 );
and ( n9457 , n9237 , n9253 );
and ( n9458 , n9253 , n9268 );
and ( n9459 , n9237 , n9268 );
or ( n9460 , n9457 , n9458 , n9459 );
and ( n9461 , n9196 , n9210 );
and ( n9462 , n9210 , n9222 );
and ( n9463 , n9196 , n9222 );
or ( n9464 , n9461 , n9462 , n9463 );
xor ( n9465 , n9460 , n9464 );
and ( n9466 , n9258 , n9262 );
and ( n9467 , n9262 , n9267 );
and ( n9468 , n9258 , n9267 );
or ( n9469 , n9466 , n9467 , n9468 );
and ( n9470 , n8116 , n7455 );
and ( n9471 , n8241 , n7344 );
nor ( n9472 , n9470 , n9471 );
xnor ( n9473 , n9472 , n7436 );
and ( n9474 , n7156 , n8606 );
and ( n9475 , n7241 , n8431 );
nor ( n9476 , n9474 , n9475 );
xnor ( n9477 , n9476 , n8612 );
xor ( n9478 , n9473 , n9477 );
and ( n9479 , n7020 , n8992 );
and ( n9480 , n7084 , n8792 );
nor ( n9481 , n9479 , n9480 );
xnor ( n9482 , n9481 , n8998 );
xor ( n9483 , n9478 , n9482 );
xor ( n9484 , n9469 , n9483 );
and ( n9485 , n8420 , n7260 );
and ( n9486 , n8643 , n7167 );
nor ( n9487 , n9485 , n9486 );
xnor ( n9488 , n9487 , n7250 );
and ( n9489 , n7545 , n7948 );
and ( n9490 , n7661 , n7823 );
nor ( n9491 , n9489 , n9490 );
xnor ( n9492 , n9491 , n7938 );
xor ( n9493 , n9488 , n9492 );
and ( n9494 , n7333 , n8294 );
and ( n9495 , n7427 , n8110 );
nor ( n9496 , n9494 , n9495 );
xnor ( n9497 , n9496 , n8250 );
xor ( n9498 , n9493 , n9497 );
xor ( n9499 , n9484 , n9498 );
xor ( n9500 , n9465 , n9499 );
xor ( n9501 , n9456 , n9500 );
xor ( n9502 , n9404 , n9501 );
and ( n9503 , n9185 , n9187 );
and ( n9504 , n9187 , n9271 );
and ( n9505 , n9185 , n9271 );
or ( n9506 , n9503 , n9504 , n9505 );
xor ( n9507 , n9502 , n9506 );
and ( n9508 , n9181 , n9272 );
and ( n9509 , n9273 , n9276 );
or ( n9510 , n9508 , n9509 );
xor ( n9511 , n9507 , n9510 );
buf ( n9512 , n9511 );
not ( n9513 , n831 );
and ( n9514 , n9513 , n9397 );
and ( n9515 , n9512 , n831 );
or ( n9516 , n9514 , n9515 );
and ( n9517 , n9293 , n9340 );
and ( n9518 , n9340 , n9385 );
and ( n9519 , n9293 , n9385 );
or ( n9520 , n9517 , n9518 , n9519 );
buf ( n9521 , n875 );
buf ( n9522 , n9521 );
xor ( n9523 , n9520 , n9522 );
and ( n9524 , n9297 , n9319 );
and ( n9525 , n9319 , n9339 );
and ( n9526 , n9297 , n9339 );
or ( n9527 , n9524 , n9525 , n9526 );
and ( n9528 , n9345 , n9349 );
and ( n9529 , n9349 , n9384 );
and ( n9530 , n9345 , n9384 );
or ( n9531 , n9528 , n9529 , n9530 );
xor ( n9532 , n9527 , n9531 );
and ( n9533 , n9358 , n9362 );
and ( n9534 , n9362 , n9367 );
and ( n9535 , n9358 , n9367 );
or ( n9536 , n9533 , n9534 , n9535 );
and ( n9537 , n9373 , n9377 );
and ( n9538 , n9377 , n9382 );
and ( n9539 , n9373 , n9382 );
or ( n9540 , n9537 , n9538 , n9539 );
xor ( n9541 , n9536 , n9540 );
and ( n9542 , n9301 , n9305 );
and ( n9543 , n9305 , n9318 );
and ( n9544 , n9301 , n9318 );
or ( n9545 , n9542 , n9543 , n9544 );
xor ( n9546 , n9541 , n9545 );
and ( n9547 , n9323 , n6957 );
buf ( n9548 , n779 );
buf ( n9549 , n9548 );
and ( n9550 , n9549 , n6934 );
nor ( n9551 , n9547 , n9550 );
xnor ( n9552 , n9551 , n6954 );
and ( n9553 , n8156 , n7400 );
and ( n9554 , n8339 , n7303 );
nor ( n9555 , n9553 , n9554 );
xnor ( n9556 , n9555 , n7381 );
xor ( n9557 , n9552 , n9556 );
buf ( n9558 , n811 );
buf ( n9559 , n9558 );
xor ( n9560 , n9559 , n9308 );
and ( n9561 , n6932 , n9560 );
xor ( n9562 , n9557 , n9561 );
and ( n9563 , n8913 , n7063 );
and ( n9564 , n9139 , n7005 );
nor ( n9565 , n9563 , n9564 );
xnor ( n9566 , n9565 , n7058 );
and ( n9567 , n7196 , n8511 );
and ( n9568 , n7292 , n8350 );
nor ( n9569 , n9567 , n9568 );
xnor ( n9570 , n9569 , n8517 );
xor ( n9571 , n9566 , n9570 );
and ( n9572 , n7049 , n8887 );
and ( n9573 , n7125 , n8701 );
nor ( n9574 , n9572 , n9573 );
xnor ( n9575 , n9574 , n8893 );
xor ( n9576 , n9571 , n9575 );
xor ( n9577 , n9562 , n9576 );
and ( n9578 , n8548 , n7215 );
and ( n9579 , n8690 , n7136 );
nor ( n9580 , n9578 , n9579 );
xnor ( n9581 , n9580 , n7205 );
and ( n9582 , n7891 , n7609 );
and ( n9583 , n8045 , n7505 );
nor ( n9584 , n9582 , n9583 );
xnor ( n9585 , n9584 , n7615 );
xor ( n9586 , n9581 , n9585 );
and ( n9587 , n6960 , n9311 );
and ( n9588 , n6999 , n9150 );
nor ( n9589 , n9587 , n9588 );
xnor ( n9590 , n9589 , n9317 );
xor ( n9591 , n9586 , n9590 );
xor ( n9592 , n9577 , n9591 );
xor ( n9593 , n9546 , n9592 );
and ( n9594 , n9329 , n9333 );
and ( n9595 , n9333 , n9338 );
and ( n9596 , n9329 , n9338 );
or ( n9597 , n9594 , n9595 , n9596 );
and ( n9598 , n9354 , n9368 );
and ( n9599 , n9368 , n9383 );
and ( n9600 , n9354 , n9383 );
or ( n9601 , n9598 , n9599 , n9600 );
xor ( n9602 , n9597 , n9601 );
and ( n9603 , n9326 , n9328 );
and ( n9604 , n7596 , n7873 );
and ( n9605 , n7730 , n7762 );
nor ( n9606 , n9604 , n9605 );
xnor ( n9607 , n9606 , n7863 );
xor ( n9608 , n9603 , n9607 );
and ( n9609 , n7372 , n8209 );
and ( n9610 , n7494 , n8039 );
nor ( n9611 , n9609 , n9610 );
xnor ( n9612 , n9611 , n8165 );
xor ( n9613 , n9608 , n9612 );
xor ( n9614 , n9602 , n9613 );
xor ( n9615 , n9593 , n9614 );
xor ( n9616 , n9532 , n9615 );
xor ( n9617 , n9523 , n9616 );
and ( n9618 , n9286 , n9288 );
and ( n9619 , n9288 , n9386 );
and ( n9620 , n9286 , n9386 );
or ( n9621 , n9618 , n9619 , n9620 );
xor ( n9622 , n9617 , n9621 );
and ( n9623 , n9387 , n9391 );
and ( n9624 , n9392 , n9395 );
or ( n9625 , n9623 , n9624 );
xor ( n9626 , n9622 , n9625 );
buf ( n9627 , n9626 );
and ( n9628 , n9408 , n9455 );
and ( n9629 , n9455 , n9500 );
and ( n9630 , n9408 , n9500 );
or ( n9631 , n9628 , n9629 , n9630 );
buf ( n9632 , n843 );
buf ( n9633 , n9632 );
xor ( n9634 , n9631 , n9633 );
and ( n9635 , n9412 , n9434 );
and ( n9636 , n9434 , n9454 );
and ( n9637 , n9412 , n9454 );
or ( n9638 , n9635 , n9636 , n9637 );
and ( n9639 , n9460 , n9464 );
and ( n9640 , n9464 , n9499 );
and ( n9641 , n9460 , n9499 );
or ( n9642 , n9639 , n9640 , n9641 );
xor ( n9643 , n9638 , n9642 );
and ( n9644 , n9473 , n9477 );
and ( n9645 , n9477 , n9482 );
and ( n9646 , n9473 , n9482 );
or ( n9647 , n9644 , n9645 , n9646 );
and ( n9648 , n9488 , n9492 );
and ( n9649 , n9492 , n9497 );
and ( n9650 , n9488 , n9497 );
or ( n9651 , n9648 , n9649 , n9650 );
xor ( n9652 , n9647 , n9651 );
and ( n9653 , n9416 , n9420 );
and ( n9654 , n9420 , n9433 );
and ( n9655 , n9416 , n9433 );
or ( n9656 , n9653 , n9654 , n9655 );
xor ( n9657 , n9652 , n9656 );
and ( n9658 , n9438 , n6977 );
buf ( n9659 , n779 );
buf ( n9660 , n9659 );
and ( n9661 , n9660 , n6943 );
nor ( n9662 , n9658 , n9661 );
xnor ( n9663 , n9662 , n6974 );
and ( n9664 , n8241 , n7455 );
and ( n9665 , n8420 , n7344 );
nor ( n9666 , n9664 , n9665 );
xnor ( n9667 , n9666 , n7436 );
xor ( n9668 , n9663 , n9667 );
buf ( n9669 , n811 );
buf ( n9670 , n9669 );
xor ( n9671 , n9670 , n9423 );
and ( n9672 , n6941 , n9671 );
xor ( n9673 , n9668 , n9672 );
and ( n9674 , n9018 , n7098 );
and ( n9675 , n9240 , n7026 );
nor ( n9676 , n9674 , n9675 );
xnor ( n9677 , n9676 , n7093 );
and ( n9678 , n7241 , n8606 );
and ( n9679 , n7333 , n8431 );
nor ( n9680 , n9678 , n9679 );
xnor ( n9681 , n9680 , n8612 );
xor ( n9682 , n9677 , n9681 );
and ( n9683 , n7084 , n8992 );
and ( n9684 , n7156 , n8792 );
nor ( n9685 , n9683 , n9684 );
xnor ( n9686 , n9685 , n8998 );
xor ( n9687 , n9682 , n9686 );
xor ( n9688 , n9673 , n9687 );
and ( n9689 , n8643 , n7260 );
and ( n9690 , n8781 , n7167 );
nor ( n9691 , n9689 , n9690 );
xnor ( n9692 , n9691 , n7250 );
and ( n9693 , n7966 , n7674 );
and ( n9694 , n8116 , n7556 );
nor ( n9695 , n9693 , n9694 );
xnor ( n9696 , n9695 , n7680 );
xor ( n9697 , n9692 , n9696 );
and ( n9698 , n6980 , n9426 );
and ( n9699 , n7020 , n9251 );
nor ( n9700 , n9698 , n9699 );
xnor ( n9701 , n9700 , n9432 );
xor ( n9702 , n9697 , n9701 );
xor ( n9703 , n9688 , n9702 );
xor ( n9704 , n9657 , n9703 );
and ( n9705 , n9444 , n9448 );
and ( n9706 , n9448 , n9453 );
and ( n9707 , n9444 , n9453 );
or ( n9708 , n9705 , n9706 , n9707 );
and ( n9709 , n9469 , n9483 );
and ( n9710 , n9483 , n9498 );
and ( n9711 , n9469 , n9498 );
or ( n9712 , n9709 , n9710 , n9711 );
xor ( n9713 , n9708 , n9712 );
and ( n9714 , n9441 , n9443 );
and ( n9715 , n7661 , n7948 );
and ( n9716 , n7791 , n7823 );
nor ( n9717 , n9715 , n9716 );
xnor ( n9718 , n9717 , n7938 );
xor ( n9719 , n9714 , n9718 );
and ( n9720 , n7427 , n8294 );
and ( n9721 , n7545 , n8110 );
nor ( n9722 , n9720 , n9721 );
xnor ( n9723 , n9722 , n8250 );
xor ( n9724 , n9719 , n9723 );
xor ( n9725 , n9713 , n9724 );
xor ( n9726 , n9704 , n9725 );
xor ( n9727 , n9643 , n9726 );
xor ( n9728 , n9634 , n9727 );
and ( n9729 , n9401 , n9403 );
and ( n9730 , n9403 , n9501 );
and ( n9731 , n9401 , n9501 );
or ( n9732 , n9729 , n9730 , n9731 );
xor ( n9733 , n9728 , n9732 );
and ( n9734 , n9502 , n9506 );
and ( n9735 , n9507 , n9510 );
or ( n9736 , n9734 , n9735 );
xor ( n9737 , n9733 , n9736 );
buf ( n9738 , n9737 );
not ( n9739 , n831 );
and ( n9740 , n9739 , n9627 );
and ( n9741 , n9738 , n831 );
or ( n9742 , n9740 , n9741 );
and ( n9743 , n9527 , n9531 );
and ( n9744 , n9531 , n9615 );
and ( n9745 , n9527 , n9615 );
or ( n9746 , n9743 , n9744 , n9745 );
buf ( n9747 , n874 );
buf ( n9748 , n9747 );
xor ( n9749 , n9746 , n9748 );
and ( n9750 , n9597 , n9601 );
and ( n9751 , n9601 , n9613 );
and ( n9752 , n9597 , n9613 );
or ( n9753 , n9750 , n9751 , n9752 );
and ( n9754 , n9546 , n9592 );
and ( n9755 , n9592 , n9614 );
and ( n9756 , n9546 , n9614 );
or ( n9757 , n9754 , n9755 , n9756 );
xor ( n9758 , n9753 , n9757 );
and ( n9759 , n9562 , n9576 );
and ( n9760 , n9576 , n9591 );
and ( n9761 , n9562 , n9591 );
or ( n9762 , n9759 , n9760 , n9761 );
and ( n9763 , n9603 , n9607 );
and ( n9764 , n9607 , n9612 );
and ( n9765 , n9603 , n9612 );
or ( n9766 , n9763 , n9764 , n9765 );
and ( n9767 , n8339 , n7400 );
and ( n9768 , n8548 , n7303 );
nor ( n9769 , n9767 , n9768 );
xnor ( n9770 , n9769 , n7381 );
and ( n9771 , n7292 , n8511 );
and ( n9772 , n7372 , n8350 );
nor ( n9773 , n9771 , n9772 );
xnor ( n9774 , n9773 , n8517 );
xor ( n9775 , n9770 , n9774 );
and ( n9776 , n7125 , n8887 );
and ( n9777 , n7196 , n8701 );
nor ( n9778 , n9776 , n9777 );
xnor ( n9779 , n9778 , n8893 );
xor ( n9780 , n9775 , n9779 );
xor ( n9781 , n9766 , n9780 );
and ( n9782 , n8045 , n7609 );
and ( n9783 , n8156 , n7505 );
nor ( n9784 , n9782 , n9783 );
xnor ( n9785 , n9784 , n7615 );
and ( n9786 , n6999 , n9311 );
and ( n9787 , n7049 , n9150 );
nor ( n9788 , n9786 , n9787 );
xnor ( n9789 , n9788 , n9317 );
xor ( n9790 , n9785 , n9789 );
buf ( n9791 , n810 );
buf ( n9792 , n9791 );
xor ( n9793 , n9792 , n9559 );
not ( n9794 , n9560 );
and ( n9795 , n9793 , n9794 );
and ( n9796 , n6932 , n9795 );
and ( n9797 , n6960 , n9560 );
nor ( n9798 , n9796 , n9797 );
and ( n9799 , n9559 , n9308 );
not ( n9800 , n9799 );
and ( n9801 , n9792 , n9800 );
xnor ( n9802 , n9798 , n9801 );
xor ( n9803 , n9790 , n9802 );
xor ( n9804 , n9781 , n9803 );
xor ( n9805 , n9762 , n9804 );
and ( n9806 , n9536 , n9540 );
and ( n9807 , n9540 , n9545 );
and ( n9808 , n9536 , n9545 );
or ( n9809 , n9806 , n9807 , n9808 );
and ( n9810 , n9139 , n7063 );
and ( n9811 , n9323 , n7005 );
nor ( n9812 , n9810 , n9811 );
xnor ( n9813 , n9812 , n7058 );
not ( n9814 , n9561 );
and ( n9815 , n9814 , n9801 );
xor ( n9816 , n9813 , n9815 );
and ( n9817 , n9566 , n9570 );
and ( n9818 , n9570 , n9575 );
and ( n9819 , n9566 , n9575 );
or ( n9820 , n9817 , n9818 , n9819 );
xor ( n9821 , n9816 , n9820 );
and ( n9822 , n7494 , n8209 );
and ( n9823 , n7596 , n8039 );
nor ( n9824 , n9822 , n9823 );
xnor ( n9825 , n9824 , n8165 );
xor ( n9826 , n9821 , n9825 );
xor ( n9827 , n9809 , n9826 );
and ( n9828 , n9552 , n9556 );
and ( n9829 , n9556 , n9561 );
and ( n9830 , n9552 , n9561 );
or ( n9831 , n9828 , n9829 , n9830 );
and ( n9832 , n9581 , n9585 );
and ( n9833 , n9585 , n9590 );
and ( n9834 , n9581 , n9590 );
or ( n9835 , n9832 , n9833 , n9834 );
xor ( n9836 , n9831 , n9835 );
and ( n9837 , n9549 , n6957 );
buf ( n9838 , n778 );
buf ( n9839 , n9838 );
and ( n9840 , n9839 , n6934 );
nor ( n9841 , n9837 , n9840 );
xnor ( n9842 , n9841 , n6954 );
and ( n9843 , n8690 , n7215 );
and ( n9844 , n8913 , n7136 );
nor ( n9845 , n9843 , n9844 );
xnor ( n9846 , n9845 , n7205 );
xor ( n9847 , n9842 , n9846 );
and ( n9848 , n7730 , n7873 );
and ( n9849 , n7891 , n7762 );
nor ( n9850 , n9848 , n9849 );
xnor ( n9851 , n9850 , n7863 );
xor ( n9852 , n9847 , n9851 );
xor ( n9853 , n9836 , n9852 );
xor ( n9854 , n9827 , n9853 );
xor ( n9855 , n9805 , n9854 );
xor ( n9856 , n9758 , n9855 );
xor ( n9857 , n9749 , n9856 );
and ( n9858 , n9520 , n9522 );
and ( n9859 , n9522 , n9616 );
and ( n9860 , n9520 , n9616 );
or ( n9861 , n9858 , n9859 , n9860 );
xor ( n9862 , n9857 , n9861 );
and ( n9863 , n9617 , n9621 );
and ( n9864 , n9622 , n9625 );
or ( n9865 , n9863 , n9864 );
xor ( n9866 , n9862 , n9865 );
buf ( n9867 , n9866 );
and ( n9868 , n9638 , n9642 );
and ( n9869 , n9642 , n9726 );
and ( n9870 , n9638 , n9726 );
or ( n9871 , n9868 , n9869 , n9870 );
buf ( n9872 , n842 );
buf ( n9873 , n9872 );
xor ( n9874 , n9871 , n9873 );
and ( n9875 , n9708 , n9712 );
and ( n9876 , n9712 , n9724 );
and ( n9877 , n9708 , n9724 );
or ( n9878 , n9875 , n9876 , n9877 );
and ( n9879 , n9657 , n9703 );
and ( n9880 , n9703 , n9725 );
and ( n9881 , n9657 , n9725 );
or ( n9882 , n9879 , n9880 , n9881 );
xor ( n9883 , n9878 , n9882 );
and ( n9884 , n9673 , n9687 );
and ( n9885 , n9687 , n9702 );
and ( n9886 , n9673 , n9702 );
or ( n9887 , n9884 , n9885 , n9886 );
and ( n9888 , n9714 , n9718 );
and ( n9889 , n9718 , n9723 );
and ( n9890 , n9714 , n9723 );
or ( n9891 , n9888 , n9889 , n9890 );
and ( n9892 , n8420 , n7455 );
and ( n9893 , n8643 , n7344 );
nor ( n9894 , n9892 , n9893 );
xnor ( n9895 , n9894 , n7436 );
and ( n9896 , n7333 , n8606 );
and ( n9897 , n7427 , n8431 );
nor ( n9898 , n9896 , n9897 );
xnor ( n9899 , n9898 , n8612 );
xor ( n9900 , n9895 , n9899 );
and ( n9901 , n7156 , n8992 );
and ( n9902 , n7241 , n8792 );
nor ( n9903 , n9901 , n9902 );
xnor ( n9904 , n9903 , n8998 );
xor ( n9905 , n9900 , n9904 );
xor ( n9906 , n9891 , n9905 );
and ( n9907 , n8116 , n7674 );
and ( n9908 , n8241 , n7556 );
nor ( n9909 , n9907 , n9908 );
xnor ( n9910 , n9909 , n7680 );
and ( n9911 , n7020 , n9426 );
and ( n9912 , n7084 , n9251 );
nor ( n9913 , n9911 , n9912 );
xnor ( n9914 , n9913 , n9432 );
xor ( n9915 , n9910 , n9914 );
buf ( n9916 , n810 );
buf ( n9917 , n9916 );
xor ( n9918 , n9917 , n9670 );
not ( n9919 , n9671 );
and ( n9920 , n9918 , n9919 );
and ( n9921 , n6941 , n9920 );
and ( n9922 , n6980 , n9671 );
nor ( n9923 , n9921 , n9922 );
and ( n9924 , n9670 , n9423 );
not ( n9925 , n9924 );
and ( n9926 , n9917 , n9925 );
xnor ( n9927 , n9923 , n9926 );
xor ( n9928 , n9915 , n9927 );
xor ( n9929 , n9906 , n9928 );
xor ( n9930 , n9887 , n9929 );
and ( n9931 , n9647 , n9651 );
and ( n9932 , n9651 , n9656 );
and ( n9933 , n9647 , n9656 );
or ( n9934 , n9931 , n9932 , n9933 );
and ( n9935 , n9240 , n7098 );
and ( n9936 , n9438 , n7026 );
nor ( n9937 , n9935 , n9936 );
xnor ( n9938 , n9937 , n7093 );
not ( n9939 , n9672 );
and ( n9940 , n9939 , n9926 );
xor ( n9941 , n9938 , n9940 );
and ( n9942 , n9677 , n9681 );
and ( n9943 , n9681 , n9686 );
and ( n9944 , n9677 , n9686 );
or ( n9945 , n9942 , n9943 , n9944 );
xor ( n9946 , n9941 , n9945 );
and ( n9947 , n7545 , n8294 );
and ( n9948 , n7661 , n8110 );
nor ( n9949 , n9947 , n9948 );
xnor ( n9950 , n9949 , n8250 );
xor ( n9951 , n9946 , n9950 );
xor ( n9952 , n9934 , n9951 );
and ( n9953 , n9663 , n9667 );
and ( n9954 , n9667 , n9672 );
and ( n9955 , n9663 , n9672 );
or ( n9956 , n9953 , n9954 , n9955 );
and ( n9957 , n9692 , n9696 );
and ( n9958 , n9696 , n9701 );
and ( n9959 , n9692 , n9701 );
or ( n9960 , n9957 , n9958 , n9959 );
xor ( n9961 , n9956 , n9960 );
and ( n9962 , n9660 , n6977 );
buf ( n9963 , n778 );
buf ( n9964 , n9963 );
and ( n9965 , n9964 , n6943 );
nor ( n9966 , n9962 , n9965 );
xnor ( n9967 , n9966 , n6974 );
and ( n9968 , n8781 , n7260 );
and ( n9969 , n9018 , n7167 );
nor ( n9970 , n9968 , n9969 );
xnor ( n9971 , n9970 , n7250 );
xor ( n9972 , n9967 , n9971 );
and ( n9973 , n7791 , n7948 );
and ( n9974 , n7966 , n7823 );
nor ( n9975 , n9973 , n9974 );
xnor ( n9976 , n9975 , n7938 );
xor ( n9977 , n9972 , n9976 );
xor ( n9978 , n9961 , n9977 );
xor ( n9979 , n9952 , n9978 );
xor ( n9980 , n9930 , n9979 );
xor ( n9981 , n9883 , n9980 );
xor ( n9982 , n9874 , n9981 );
and ( n9983 , n9631 , n9633 );
and ( n9984 , n9633 , n9727 );
and ( n9985 , n9631 , n9727 );
or ( n9986 , n9983 , n9984 , n9985 );
xor ( n9987 , n9982 , n9986 );
and ( n9988 , n9728 , n9732 );
and ( n9989 , n9733 , n9736 );
or ( n9990 , n9988 , n9989 );
xor ( n9991 , n9987 , n9990 );
buf ( n9992 , n9991 );
not ( n9993 , n831 );
and ( n9994 , n9993 , n9867 );
and ( n9995 , n9992 , n831 );
or ( n9996 , n9994 , n9995 );
and ( n9997 , n9753 , n9757 );
and ( n9998 , n9757 , n9855 );
and ( n9999 , n9753 , n9855 );
or ( n10000 , n9997 , n9998 , n9999 );
buf ( n10001 , n873 );
buf ( n10002 , n10001 );
xor ( n10003 , n10000 , n10002 );
and ( n10004 , n9762 , n9804 );
and ( n10005 , n9804 , n9854 );
and ( n10006 , n9762 , n9854 );
or ( n10007 , n10004 , n10005 , n10006 );
and ( n10008 , n9831 , n9835 );
and ( n10009 , n9835 , n9852 );
and ( n10010 , n9831 , n9852 );
or ( n10011 , n10008 , n10009 , n10010 );
and ( n10012 , n9766 , n9780 );
and ( n10013 , n9780 , n9803 );
and ( n10014 , n9766 , n9803 );
or ( n10015 , n10012 , n10013 , n10014 );
xor ( n10016 , n10011 , n10015 );
and ( n10017 , n9842 , n9846 );
and ( n10018 , n9846 , n9851 );
and ( n10019 , n9842 , n9851 );
or ( n10020 , n10017 , n10018 , n10019 );
and ( n10021 , n9785 , n9789 );
and ( n10022 , n9789 , n9802 );
and ( n10023 , n9785 , n9802 );
or ( n10024 , n10021 , n10022 , n10023 );
xor ( n10025 , n10020 , n10024 );
and ( n10026 , n9813 , n9815 );
xor ( n10027 , n10025 , n10026 );
xor ( n10028 , n10016 , n10027 );
xor ( n10029 , n10007 , n10028 );
and ( n10030 , n9809 , n9826 );
and ( n10031 , n9826 , n9853 );
and ( n10032 , n9809 , n9853 );
or ( n10033 , n10030 , n10031 , n10032 );
and ( n10034 , n9770 , n9774 );
and ( n10035 , n9774 , n9779 );
and ( n10036 , n9770 , n9779 );
or ( n10037 , n10034 , n10035 , n10036 );
and ( n10038 , n8156 , n7609 );
and ( n10039 , n8339 , n7505 );
nor ( n10040 , n10038 , n10039 );
xnor ( n10041 , n10040 , n7615 );
and ( n10042 , n7372 , n8511 );
and ( n10043 , n7494 , n8350 );
nor ( n10044 , n10042 , n10043 );
xnor ( n10045 , n10044 , n8517 );
xor ( n10046 , n10041 , n10045 );
and ( n10047 , n7196 , n8887 );
and ( n10048 , n7292 , n8701 );
nor ( n10049 , n10047 , n10048 );
xnor ( n10050 , n10049 , n8893 );
xor ( n10051 , n10046 , n10050 );
xor ( n10052 , n10037 , n10051 );
and ( n10053 , n8913 , n7215 );
and ( n10054 , n9139 , n7136 );
nor ( n10055 , n10053 , n10054 );
xnor ( n10056 , n10055 , n7205 );
and ( n10057 , n7891 , n7873 );
and ( n10058 , n8045 , n7762 );
nor ( n10059 , n10057 , n10058 );
xnor ( n10060 , n10059 , n7863 );
xor ( n10061 , n10056 , n10060 );
and ( n10062 , n7596 , n8209 );
and ( n10063 , n7730 , n8039 );
nor ( n10064 , n10062 , n10063 );
xnor ( n10065 , n10064 , n8165 );
xor ( n10066 , n10061 , n10065 );
xor ( n10067 , n10052 , n10066 );
xor ( n10068 , n10033 , n10067 );
and ( n10069 , n9816 , n9820 );
and ( n10070 , n9820 , n9825 );
and ( n10071 , n9816 , n9825 );
or ( n10072 , n10069 , n10070 , n10071 );
and ( n10073 , n9323 , n7063 );
and ( n10074 , n9549 , n7005 );
nor ( n10075 , n10073 , n10074 );
xnor ( n10076 , n10075 , n7058 );
and ( n10077 , n8548 , n7400 );
and ( n10078 , n8690 , n7303 );
nor ( n10079 , n10077 , n10078 );
xnor ( n10080 , n10079 , n7381 );
xor ( n10081 , n10076 , n10080 );
buf ( n10082 , n809 );
buf ( n10083 , n10082 );
xor ( n10084 , n10083 , n9792 );
and ( n10085 , n6932 , n10084 );
xor ( n10086 , n10081 , n10085 );
xor ( n10087 , n10072 , n10086 );
and ( n10088 , n9839 , n6957 );
buf ( n10089 , n777 );
buf ( n10090 , n10089 );
and ( n10091 , n10090 , n6934 );
nor ( n10092 , n10088 , n10091 );
xnor ( n10093 , n10092 , n6954 );
and ( n10094 , n7049 , n9311 );
and ( n10095 , n7125 , n9150 );
nor ( n10096 , n10094 , n10095 );
xnor ( n10097 , n10096 , n9317 );
xor ( n10098 , n10093 , n10097 );
and ( n10099 , n6960 , n9795 );
and ( n10100 , n6999 , n9560 );
nor ( n10101 , n10099 , n10100 );
xnor ( n10102 , n10101 , n9801 );
xor ( n10103 , n10098 , n10102 );
xor ( n10104 , n10087 , n10103 );
xor ( n10105 , n10068 , n10104 );
xor ( n10106 , n10029 , n10105 );
xor ( n10107 , n10003 , n10106 );
and ( n10108 , n9746 , n9748 );
and ( n10109 , n9748 , n9856 );
and ( n10110 , n9746 , n9856 );
or ( n10111 , n10108 , n10109 , n10110 );
xor ( n10112 , n10107 , n10111 );
and ( n10113 , n9857 , n9861 );
and ( n10114 , n9862 , n9865 );
or ( n10115 , n10113 , n10114 );
xor ( n10116 , n10112 , n10115 );
buf ( n10117 , n10116 );
and ( n10118 , n9878 , n9882 );
and ( n10119 , n9882 , n9980 );
and ( n10120 , n9878 , n9980 );
or ( n10121 , n10118 , n10119 , n10120 );
buf ( n10122 , n841 );
buf ( n10123 , n10122 );
xor ( n10124 , n10121 , n10123 );
and ( n10125 , n9887 , n9929 );
and ( n10126 , n9929 , n9979 );
and ( n10127 , n9887 , n9979 );
or ( n10128 , n10125 , n10126 , n10127 );
and ( n10129 , n9956 , n9960 );
and ( n10130 , n9960 , n9977 );
and ( n10131 , n9956 , n9977 );
or ( n10132 , n10129 , n10130 , n10131 );
and ( n10133 , n9891 , n9905 );
and ( n10134 , n9905 , n9928 );
and ( n10135 , n9891 , n9928 );
or ( n10136 , n10133 , n10134 , n10135 );
xor ( n10137 , n10132 , n10136 );
and ( n10138 , n9967 , n9971 );
and ( n10139 , n9971 , n9976 );
and ( n10140 , n9967 , n9976 );
or ( n10141 , n10138 , n10139 , n10140 );
and ( n10142 , n9910 , n9914 );
and ( n10143 , n9914 , n9927 );
and ( n10144 , n9910 , n9927 );
or ( n10145 , n10142 , n10143 , n10144 );
xor ( n10146 , n10141 , n10145 );
and ( n10147 , n9938 , n9940 );
xor ( n10148 , n10146 , n10147 );
xor ( n10149 , n10137 , n10148 );
xor ( n10150 , n10128 , n10149 );
and ( n10151 , n9934 , n9951 );
and ( n10152 , n9951 , n9978 );
and ( n10153 , n9934 , n9978 );
or ( n10154 , n10151 , n10152 , n10153 );
and ( n10155 , n9895 , n9899 );
and ( n10156 , n9899 , n9904 );
and ( n10157 , n9895 , n9904 );
or ( n10158 , n10155 , n10156 , n10157 );
and ( n10159 , n8241 , n7674 );
and ( n10160 , n8420 , n7556 );
nor ( n10161 , n10159 , n10160 );
xnor ( n10162 , n10161 , n7680 );
and ( n10163 , n7427 , n8606 );
and ( n10164 , n7545 , n8431 );
nor ( n10165 , n10163 , n10164 );
xnor ( n10166 , n10165 , n8612 );
xor ( n10167 , n10162 , n10166 );
and ( n10168 , n7241 , n8992 );
and ( n10169 , n7333 , n8792 );
nor ( n10170 , n10168 , n10169 );
xnor ( n10171 , n10170 , n8998 );
xor ( n10172 , n10167 , n10171 );
xor ( n10173 , n10158 , n10172 );
and ( n10174 , n9018 , n7260 );
and ( n10175 , n9240 , n7167 );
nor ( n10176 , n10174 , n10175 );
xnor ( n10177 , n10176 , n7250 );
and ( n10178 , n7966 , n7948 );
and ( n10179 , n8116 , n7823 );
nor ( n10180 , n10178 , n10179 );
xnor ( n10181 , n10180 , n7938 );
xor ( n10182 , n10177 , n10181 );
and ( n10183 , n7661 , n8294 );
and ( n10184 , n7791 , n8110 );
nor ( n10185 , n10183 , n10184 );
xnor ( n10186 , n10185 , n8250 );
xor ( n10187 , n10182 , n10186 );
xor ( n10188 , n10173 , n10187 );
xor ( n10189 , n10154 , n10188 );
and ( n10190 , n9941 , n9945 );
and ( n10191 , n9945 , n9950 );
and ( n10192 , n9941 , n9950 );
or ( n10193 , n10190 , n10191 , n10192 );
and ( n10194 , n9438 , n7098 );
and ( n10195 , n9660 , n7026 );
nor ( n10196 , n10194 , n10195 );
xnor ( n10197 , n10196 , n7093 );
and ( n10198 , n8643 , n7455 );
and ( n10199 , n8781 , n7344 );
nor ( n10200 , n10198 , n10199 );
xnor ( n10201 , n10200 , n7436 );
xor ( n10202 , n10197 , n10201 );
buf ( n10203 , n809 );
buf ( n10204 , n10203 );
xor ( n10205 , n10204 , n9917 );
and ( n10206 , n6941 , n10205 );
xor ( n10207 , n10202 , n10206 );
xor ( n10208 , n10193 , n10207 );
and ( n10209 , n9964 , n6977 );
buf ( n10210 , n777 );
buf ( n10211 , n10210 );
and ( n10212 , n10211 , n6943 );
nor ( n10213 , n10209 , n10212 );
xnor ( n10214 , n10213 , n6974 );
and ( n10215 , n7084 , n9426 );
and ( n10216 , n7156 , n9251 );
nor ( n10217 , n10215 , n10216 );
xnor ( n10218 , n10217 , n9432 );
xor ( n10219 , n10214 , n10218 );
and ( n10220 , n6980 , n9920 );
and ( n10221 , n7020 , n9671 );
nor ( n10222 , n10220 , n10221 );
xnor ( n10223 , n10222 , n9926 );
xor ( n10224 , n10219 , n10223 );
xor ( n10225 , n10208 , n10224 );
xor ( n10226 , n10189 , n10225 );
xor ( n10227 , n10150 , n10226 );
xor ( n10228 , n10124 , n10227 );
and ( n10229 , n9871 , n9873 );
and ( n10230 , n9873 , n9981 );
and ( n10231 , n9871 , n9981 );
or ( n10232 , n10229 , n10230 , n10231 );
xor ( n10233 , n10228 , n10232 );
and ( n10234 , n9982 , n9986 );
and ( n10235 , n9987 , n9990 );
or ( n10236 , n10234 , n10235 );
xor ( n10237 , n10233 , n10236 );
buf ( n10238 , n10237 );
not ( n10239 , n831 );
and ( n10240 , n10239 , n10117 );
and ( n10241 , n10238 , n831 );
or ( n10242 , n10240 , n10241 );
and ( n10243 , n10007 , n10028 );
and ( n10244 , n10028 , n10105 );
and ( n10245 , n10007 , n10105 );
or ( n10246 , n10243 , n10244 , n10245 );
buf ( n10247 , n872 );
buf ( n10248 , n10247 );
xor ( n10249 , n10246 , n10248 );
and ( n10250 , n10011 , n10015 );
and ( n10251 , n10015 , n10027 );
and ( n10252 , n10011 , n10027 );
or ( n10253 , n10250 , n10251 , n10252 );
and ( n10254 , n10033 , n10067 );
and ( n10255 , n10067 , n10104 );
and ( n10256 , n10033 , n10104 );
or ( n10257 , n10254 , n10255 , n10256 );
xor ( n10258 , n10253 , n10257 );
and ( n10259 , n10072 , n10086 );
and ( n10260 , n10086 , n10103 );
and ( n10261 , n10072 , n10103 );
or ( n10262 , n10259 , n10260 , n10261 );
and ( n10263 , n10020 , n10024 );
and ( n10264 , n10024 , n10026 );
and ( n10265 , n10020 , n10026 );
or ( n10266 , n10263 , n10264 , n10265 );
and ( n10267 , n8690 , n7400 );
and ( n10268 , n8913 , n7303 );
nor ( n10269 , n10267 , n10268 );
xnor ( n10270 , n10269 , n7381 );
and ( n10271 , n7494 , n8511 );
and ( n10272 , n7596 , n8350 );
nor ( n10273 , n10271 , n10272 );
xnor ( n10274 , n10273 , n8517 );
xor ( n10275 , n10270 , n10274 );
and ( n10276 , n7292 , n8887 );
and ( n10277 , n7372 , n8701 );
nor ( n10278 , n10276 , n10277 );
xnor ( n10279 , n10278 , n8893 );
xor ( n10280 , n10275 , n10279 );
xor ( n10281 , n10266 , n10280 );
and ( n10282 , n9549 , n7063 );
and ( n10283 , n9839 , n7005 );
nor ( n10284 , n10282 , n10283 );
xnor ( n10285 , n10284 , n7058 );
not ( n10286 , n10085 );
buf ( n10287 , n808 );
buf ( n10288 , n10287 );
and ( n10289 , n10083 , n9792 );
not ( n10290 , n10289 );
and ( n10291 , n10288 , n10290 );
and ( n10292 , n10286 , n10291 );
xor ( n10293 , n10285 , n10292 );
and ( n10294 , n8045 , n7873 );
and ( n10295 , n8156 , n7762 );
nor ( n10296 , n10294 , n10295 );
xnor ( n10297 , n10296 , n7863 );
xor ( n10298 , n10293 , n10297 );
and ( n10299 , n7730 , n8209 );
and ( n10300 , n7891 , n8039 );
nor ( n10301 , n10299 , n10300 );
xnor ( n10302 , n10301 , n8165 );
xor ( n10303 , n10298 , n10302 );
xor ( n10304 , n10281 , n10303 );
xor ( n10305 , n10262 , n10304 );
and ( n10306 , n10037 , n10051 );
and ( n10307 , n10051 , n10066 );
and ( n10308 , n10037 , n10066 );
or ( n10309 , n10306 , n10307 , n10308 );
and ( n10310 , n10056 , n10060 );
and ( n10311 , n10060 , n10065 );
and ( n10312 , n10056 , n10065 );
or ( n10313 , n10310 , n10311 , n10312 );
and ( n10314 , n10076 , n10080 );
and ( n10315 , n10080 , n10085 );
and ( n10316 , n10076 , n10085 );
or ( n10317 , n10314 , n10315 , n10316 );
xor ( n10318 , n10313 , n10317 );
and ( n10319 , n10093 , n10097 );
and ( n10320 , n10097 , n10102 );
and ( n10321 , n10093 , n10102 );
or ( n10322 , n10319 , n10320 , n10321 );
xor ( n10323 , n10318 , n10322 );
xor ( n10324 , n10309 , n10323 );
and ( n10325 , n10041 , n10045 );
and ( n10326 , n10045 , n10050 );
and ( n10327 , n10041 , n10050 );
or ( n10328 , n10325 , n10326 , n10327 );
and ( n10329 , n10090 , n6957 );
buf ( n10330 , n776 );
buf ( n10331 , n10330 );
and ( n10332 , n10331 , n6934 );
nor ( n10333 , n10329 , n10332 );
xnor ( n10334 , n10333 , n6954 );
and ( n10335 , n9139 , n7215 );
and ( n10336 , n9323 , n7136 );
nor ( n10337 , n10335 , n10336 );
xnor ( n10338 , n10337 , n7205 );
xor ( n10339 , n10334 , n10338 );
xor ( n10340 , n10288 , n10083 );
not ( n10341 , n10084 );
and ( n10342 , n10340 , n10341 );
and ( n10343 , n6932 , n10342 );
and ( n10344 , n6960 , n10084 );
nor ( n10345 , n10343 , n10344 );
xnor ( n10346 , n10345 , n10291 );
xor ( n10347 , n10339 , n10346 );
xor ( n10348 , n10328 , n10347 );
and ( n10349 , n8339 , n7609 );
and ( n10350 , n8548 , n7505 );
nor ( n10351 , n10349 , n10350 );
xnor ( n10352 , n10351 , n7615 );
and ( n10353 , n7125 , n9311 );
and ( n10354 , n7196 , n9150 );
nor ( n10355 , n10353 , n10354 );
xnor ( n10356 , n10355 , n9317 );
xor ( n10357 , n10352 , n10356 );
and ( n10358 , n6999 , n9795 );
and ( n10359 , n7049 , n9560 );
nor ( n10360 , n10358 , n10359 );
xnor ( n10361 , n10360 , n9801 );
xor ( n10362 , n10357 , n10361 );
xor ( n10363 , n10348 , n10362 );
xor ( n10364 , n10324 , n10363 );
xor ( n10365 , n10305 , n10364 );
xor ( n10366 , n10258 , n10365 );
xor ( n10367 , n10249 , n10366 );
and ( n10368 , n10000 , n10002 );
and ( n10369 , n10002 , n10106 );
and ( n10370 , n10000 , n10106 );
or ( n10371 , n10368 , n10369 , n10370 );
xor ( n10372 , n10367 , n10371 );
and ( n10373 , n10107 , n10111 );
and ( n10374 , n10112 , n10115 );
or ( n10375 , n10373 , n10374 );
xor ( n10376 , n10372 , n10375 );
buf ( n10377 , n10376 );
and ( n10378 , n10128 , n10149 );
and ( n10379 , n10149 , n10226 );
and ( n10380 , n10128 , n10226 );
or ( n10381 , n10378 , n10379 , n10380 );
buf ( n10382 , n840 );
buf ( n10383 , n10382 );
xor ( n10384 , n10381 , n10383 );
and ( n10385 , n10132 , n10136 );
and ( n10386 , n10136 , n10148 );
and ( n10387 , n10132 , n10148 );
or ( n10388 , n10385 , n10386 , n10387 );
and ( n10389 , n10154 , n10188 );
and ( n10390 , n10188 , n10225 );
and ( n10391 , n10154 , n10225 );
or ( n10392 , n10389 , n10390 , n10391 );
xor ( n10393 , n10388 , n10392 );
and ( n10394 , n10193 , n10207 );
and ( n10395 , n10207 , n10224 );
and ( n10396 , n10193 , n10224 );
or ( n10397 , n10394 , n10395 , n10396 );
and ( n10398 , n10141 , n10145 );
and ( n10399 , n10145 , n10147 );
and ( n10400 , n10141 , n10147 );
or ( n10401 , n10398 , n10399 , n10400 );
and ( n10402 , n8781 , n7455 );
and ( n10403 , n9018 , n7344 );
nor ( n10404 , n10402 , n10403 );
xnor ( n10405 , n10404 , n7436 );
and ( n10406 , n7545 , n8606 );
and ( n10407 , n7661 , n8431 );
nor ( n10408 , n10406 , n10407 );
xnor ( n10409 , n10408 , n8612 );
xor ( n10410 , n10405 , n10409 );
and ( n10411 , n7333 , n8992 );
and ( n10412 , n7427 , n8792 );
nor ( n10413 , n10411 , n10412 );
xnor ( n10414 , n10413 , n8998 );
xor ( n10415 , n10410 , n10414 );
xor ( n10416 , n10401 , n10415 );
and ( n10417 , n9660 , n7098 );
and ( n10418 , n9964 , n7026 );
nor ( n10419 , n10417 , n10418 );
xnor ( n10420 , n10419 , n7093 );
not ( n10421 , n10206 );
buf ( n10422 , n808 );
buf ( n10423 , n10422 );
and ( n10424 , n10204 , n9917 );
not ( n10425 , n10424 );
and ( n10426 , n10423 , n10425 );
and ( n10427 , n10421 , n10426 );
xor ( n10428 , n10420 , n10427 );
and ( n10429 , n8116 , n7948 );
and ( n10430 , n8241 , n7823 );
nor ( n10431 , n10429 , n10430 );
xnor ( n10432 , n10431 , n7938 );
xor ( n10433 , n10428 , n10432 );
and ( n10434 , n7791 , n8294 );
and ( n10435 , n7966 , n8110 );
nor ( n10436 , n10434 , n10435 );
xnor ( n10437 , n10436 , n8250 );
xor ( n10438 , n10433 , n10437 );
xor ( n10439 , n10416 , n10438 );
xor ( n10440 , n10397 , n10439 );
and ( n10441 , n10158 , n10172 );
and ( n10442 , n10172 , n10187 );
and ( n10443 , n10158 , n10187 );
or ( n10444 , n10441 , n10442 , n10443 );
and ( n10445 , n10177 , n10181 );
and ( n10446 , n10181 , n10186 );
and ( n10447 , n10177 , n10186 );
or ( n10448 , n10445 , n10446 , n10447 );
and ( n10449 , n10197 , n10201 );
and ( n10450 , n10201 , n10206 );
and ( n10451 , n10197 , n10206 );
or ( n10452 , n10449 , n10450 , n10451 );
xor ( n10453 , n10448 , n10452 );
and ( n10454 , n10214 , n10218 );
and ( n10455 , n10218 , n10223 );
and ( n10456 , n10214 , n10223 );
or ( n10457 , n10454 , n10455 , n10456 );
xor ( n10458 , n10453 , n10457 );
xor ( n10459 , n10444 , n10458 );
and ( n10460 , n10162 , n10166 );
and ( n10461 , n10166 , n10171 );
and ( n10462 , n10162 , n10171 );
or ( n10463 , n10460 , n10461 , n10462 );
and ( n10464 , n10211 , n6977 );
buf ( n10465 , n776 );
buf ( n10466 , n10465 );
and ( n10467 , n10466 , n6943 );
nor ( n10468 , n10464 , n10467 );
xnor ( n10469 , n10468 , n6974 );
and ( n10470 , n9240 , n7260 );
and ( n10471 , n9438 , n7167 );
nor ( n10472 , n10470 , n10471 );
xnor ( n10473 , n10472 , n7250 );
xor ( n10474 , n10469 , n10473 );
xor ( n10475 , n10423 , n10204 );
not ( n10476 , n10205 );
and ( n10477 , n10475 , n10476 );
and ( n10478 , n6941 , n10477 );
and ( n10479 , n6980 , n10205 );
nor ( n10480 , n10478 , n10479 );
xnor ( n10481 , n10480 , n10426 );
xor ( n10482 , n10474 , n10481 );
xor ( n10483 , n10463 , n10482 );
and ( n10484 , n8420 , n7674 );
and ( n10485 , n8643 , n7556 );
nor ( n10486 , n10484 , n10485 );
xnor ( n10487 , n10486 , n7680 );
and ( n10488 , n7156 , n9426 );
and ( n10489 , n7241 , n9251 );
nor ( n10490 , n10488 , n10489 );
xnor ( n10491 , n10490 , n9432 );
xor ( n10492 , n10487 , n10491 );
and ( n10493 , n7020 , n9920 );
and ( n10494 , n7084 , n9671 );
nor ( n10495 , n10493 , n10494 );
xnor ( n10496 , n10495 , n9926 );
xor ( n10497 , n10492 , n10496 );
xor ( n10498 , n10483 , n10497 );
xor ( n10499 , n10459 , n10498 );
xor ( n10500 , n10440 , n10499 );
xor ( n10501 , n10393 , n10500 );
xor ( n10502 , n10384 , n10501 );
and ( n10503 , n10121 , n10123 );
and ( n10504 , n10123 , n10227 );
and ( n10505 , n10121 , n10227 );
or ( n10506 , n10503 , n10504 , n10505 );
xor ( n10507 , n10502 , n10506 );
and ( n10508 , n10228 , n10232 );
and ( n10509 , n10233 , n10236 );
or ( n10510 , n10508 , n10509 );
xor ( n10511 , n10507 , n10510 );
buf ( n10512 , n10511 );
not ( n10513 , n831 );
and ( n10514 , n10513 , n10377 );
and ( n10515 , n10512 , n831 );
or ( n10516 , n10514 , n10515 );
and ( n10517 , n10253 , n10257 );
and ( n10518 , n10257 , n10365 );
and ( n10519 , n10253 , n10365 );
or ( n10520 , n10517 , n10518 , n10519 );
buf ( n10521 , n871 );
buf ( n10522 , n10521 );
xor ( n10523 , n10520 , n10522 );
and ( n10524 , n10262 , n10304 );
and ( n10525 , n10304 , n10364 );
and ( n10526 , n10262 , n10364 );
or ( n10527 , n10524 , n10525 , n10526 );
and ( n10528 , n10328 , n10347 );
and ( n10529 , n10347 , n10362 );
and ( n10530 , n10328 , n10362 );
or ( n10531 , n10528 , n10529 , n10530 );
and ( n10532 , n9839 , n7063 );
and ( n10533 , n10090 , n7005 );
nor ( n10534 , n10532 , n10533 );
xnor ( n10535 , n10534 , n7058 );
and ( n10536 , n8913 , n7400 );
and ( n10537 , n9139 , n7303 );
nor ( n10538 , n10536 , n10537 );
xnor ( n10539 , n10538 , n7381 );
xor ( n10540 , n10535 , n10539 );
buf ( n10541 , n807 );
buf ( n10542 , n10541 );
xor ( n10543 , n10542 , n10288 );
and ( n10544 , n6932 , n10543 );
xor ( n10545 , n10540 , n10544 );
and ( n10546 , n10331 , n6957 );
buf ( n10547 , n775 );
buf ( n10548 , n10547 );
and ( n10549 , n10548 , n6934 );
nor ( n10550 , n10546 , n10549 );
xnor ( n10551 , n10550 , n6954 );
and ( n10552 , n7196 , n9311 );
and ( n10553 , n7292 , n9150 );
nor ( n10554 , n10552 , n10553 );
xnor ( n10555 , n10554 , n9317 );
xor ( n10556 , n10551 , n10555 );
and ( n10557 , n7049 , n9795 );
and ( n10558 , n7125 , n9560 );
nor ( n10559 , n10557 , n10558 );
xnor ( n10560 , n10559 , n9801 );
xor ( n10561 , n10556 , n10560 );
xor ( n10562 , n10545 , n10561 );
and ( n10563 , n8548 , n7609 );
and ( n10564 , n8690 , n7505 );
nor ( n10565 , n10563 , n10564 );
xnor ( n10566 , n10565 , n7615 );
and ( n10567 , n7596 , n8511 );
and ( n10568 , n7730 , n8350 );
nor ( n10569 , n10567 , n10568 );
xnor ( n10570 , n10569 , n8517 );
xor ( n10571 , n10566 , n10570 );
and ( n10572 , n7372 , n8887 );
and ( n10573 , n7494 , n8701 );
nor ( n10574 , n10572 , n10573 );
xnor ( n10575 , n10574 , n8893 );
xor ( n10576 , n10571 , n10575 );
xor ( n10577 , n10562 , n10576 );
xor ( n10578 , n10531 , n10577 );
and ( n10579 , n10334 , n10338 );
and ( n10580 , n10338 , n10346 );
and ( n10581 , n10334 , n10346 );
or ( n10582 , n10579 , n10580 , n10581 );
and ( n10583 , n10270 , n10274 );
and ( n10584 , n10274 , n10279 );
and ( n10585 , n10270 , n10279 );
or ( n10586 , n10583 , n10584 , n10585 );
xor ( n10587 , n10582 , n10586 );
and ( n10588 , n9323 , n7215 );
and ( n10589 , n9549 , n7136 );
nor ( n10590 , n10588 , n10589 );
xnor ( n10591 , n10590 , n7205 );
and ( n10592 , n8156 , n7873 );
and ( n10593 , n8339 , n7762 );
nor ( n10594 , n10592 , n10593 );
xnor ( n10595 , n10594 , n7863 );
xor ( n10596 , n10591 , n10595 );
and ( n10597 , n6960 , n10342 );
and ( n10598 , n6999 , n10084 );
nor ( n10599 , n10597 , n10598 );
xnor ( n10600 , n10599 , n10291 );
xor ( n10601 , n10596 , n10600 );
xor ( n10602 , n10587 , n10601 );
xor ( n10603 , n10578 , n10602 );
xor ( n10604 , n10527 , n10603 );
and ( n10605 , n10266 , n10280 );
and ( n10606 , n10280 , n10303 );
and ( n10607 , n10266 , n10303 );
or ( n10608 , n10605 , n10606 , n10607 );
and ( n10609 , n10309 , n10323 );
and ( n10610 , n10323 , n10363 );
and ( n10611 , n10309 , n10363 );
or ( n10612 , n10609 , n10610 , n10611 );
xor ( n10613 , n10608 , n10612 );
and ( n10614 , n10313 , n10317 );
and ( n10615 , n10317 , n10322 );
and ( n10616 , n10313 , n10322 );
or ( n10617 , n10614 , n10615 , n10616 );
and ( n10618 , n10293 , n10297 );
and ( n10619 , n10297 , n10302 );
and ( n10620 , n10293 , n10302 );
or ( n10621 , n10618 , n10619 , n10620 );
xor ( n10622 , n10617 , n10621 );
and ( n10623 , n10352 , n10356 );
and ( n10624 , n10356 , n10361 );
and ( n10625 , n10352 , n10361 );
or ( n10626 , n10623 , n10624 , n10625 );
and ( n10627 , n10285 , n10292 );
xor ( n10628 , n10626 , n10627 );
and ( n10629 , n7891 , n8209 );
and ( n10630 , n8045 , n8039 );
nor ( n10631 , n10629 , n10630 );
xnor ( n10632 , n10631 , n8165 );
xor ( n10633 , n10628 , n10632 );
xor ( n10634 , n10622 , n10633 );
xor ( n10635 , n10613 , n10634 );
xor ( n10636 , n10604 , n10635 );
xor ( n10637 , n10523 , n10636 );
and ( n10638 , n10246 , n10248 );
and ( n10639 , n10248 , n10366 );
and ( n10640 , n10246 , n10366 );
or ( n10641 , n10638 , n10639 , n10640 );
xor ( n10642 , n10637 , n10641 );
and ( n10643 , n10367 , n10371 );
and ( n10644 , n10372 , n10375 );
or ( n10645 , n10643 , n10644 );
xor ( n10646 , n10642 , n10645 );
buf ( n10647 , n10646 );
and ( n10648 , n10388 , n10392 );
and ( n10649 , n10392 , n10500 );
and ( n10650 , n10388 , n10500 );
or ( n10651 , n10648 , n10649 , n10650 );
buf ( n10652 , n839 );
buf ( n10653 , n10652 );
xor ( n10654 , n10651 , n10653 );
and ( n10655 , n10397 , n10439 );
and ( n10656 , n10439 , n10499 );
and ( n10657 , n10397 , n10499 );
or ( n10658 , n10655 , n10656 , n10657 );
and ( n10659 , n10463 , n10482 );
and ( n10660 , n10482 , n10497 );
and ( n10661 , n10463 , n10497 );
or ( n10662 , n10659 , n10660 , n10661 );
and ( n10663 , n9964 , n7098 );
and ( n10664 , n10211 , n7026 );
nor ( n10665 , n10663 , n10664 );
xnor ( n10666 , n10665 , n7093 );
and ( n10667 , n9018 , n7455 );
and ( n10668 , n9240 , n7344 );
nor ( n10669 , n10667 , n10668 );
xnor ( n10670 , n10669 , n7436 );
xor ( n10671 , n10666 , n10670 );
buf ( n10672 , n807 );
buf ( n10673 , n10672 );
xor ( n10674 , n10673 , n10423 );
and ( n10675 , n6941 , n10674 );
xor ( n10676 , n10671 , n10675 );
and ( n10677 , n10466 , n6977 );
buf ( n10678 , n775 );
buf ( n10679 , n10678 );
and ( n10680 , n10679 , n6943 );
nor ( n10681 , n10677 , n10680 );
xnor ( n10682 , n10681 , n6974 );
and ( n10683 , n7241 , n9426 );
and ( n10684 , n7333 , n9251 );
nor ( n10685 , n10683 , n10684 );
xnor ( n10686 , n10685 , n9432 );
xor ( n10687 , n10682 , n10686 );
and ( n10688 , n7084 , n9920 );
and ( n10689 , n7156 , n9671 );
nor ( n10690 , n10688 , n10689 );
xnor ( n10691 , n10690 , n9926 );
xor ( n10692 , n10687 , n10691 );
xor ( n10693 , n10676 , n10692 );
and ( n10694 , n8643 , n7674 );
and ( n10695 , n8781 , n7556 );
nor ( n10696 , n10694 , n10695 );
xnor ( n10697 , n10696 , n7680 );
and ( n10698 , n7661 , n8606 );
and ( n10699 , n7791 , n8431 );
nor ( n10700 , n10698 , n10699 );
xnor ( n10701 , n10700 , n8612 );
xor ( n10702 , n10697 , n10701 );
and ( n10703 , n7427 , n8992 );
and ( n10704 , n7545 , n8792 );
nor ( n10705 , n10703 , n10704 );
xnor ( n10706 , n10705 , n8998 );
xor ( n10707 , n10702 , n10706 );
xor ( n10708 , n10693 , n10707 );
xor ( n10709 , n10662 , n10708 );
and ( n10710 , n10469 , n10473 );
and ( n10711 , n10473 , n10481 );
and ( n10712 , n10469 , n10481 );
or ( n10713 , n10710 , n10711 , n10712 );
and ( n10714 , n10405 , n10409 );
and ( n10715 , n10409 , n10414 );
and ( n10716 , n10405 , n10414 );
or ( n10717 , n10714 , n10715 , n10716 );
xor ( n10718 , n10713 , n10717 );
and ( n10719 , n9438 , n7260 );
and ( n10720 , n9660 , n7167 );
nor ( n10721 , n10719 , n10720 );
xnor ( n10722 , n10721 , n7250 );
and ( n10723 , n8241 , n7948 );
and ( n10724 , n8420 , n7823 );
nor ( n10725 , n10723 , n10724 );
xnor ( n10726 , n10725 , n7938 );
xor ( n10727 , n10722 , n10726 );
and ( n10728 , n6980 , n10477 );
and ( n10729 , n7020 , n10205 );
nor ( n10730 , n10728 , n10729 );
xnor ( n10731 , n10730 , n10426 );
xor ( n10732 , n10727 , n10731 );
xor ( n10733 , n10718 , n10732 );
xor ( n10734 , n10709 , n10733 );
xor ( n10735 , n10658 , n10734 );
and ( n10736 , n10401 , n10415 );
and ( n10737 , n10415 , n10438 );
and ( n10738 , n10401 , n10438 );
or ( n10739 , n10736 , n10737 , n10738 );
and ( n10740 , n10444 , n10458 );
and ( n10741 , n10458 , n10498 );
and ( n10742 , n10444 , n10498 );
or ( n10743 , n10740 , n10741 , n10742 );
xor ( n10744 , n10739 , n10743 );
and ( n10745 , n10448 , n10452 );
and ( n10746 , n10452 , n10457 );
and ( n10747 , n10448 , n10457 );
or ( n10748 , n10745 , n10746 , n10747 );
and ( n10749 , n10428 , n10432 );
and ( n10750 , n10432 , n10437 );
and ( n10751 , n10428 , n10437 );
or ( n10752 , n10749 , n10750 , n10751 );
xor ( n10753 , n10748 , n10752 );
and ( n10754 , n10487 , n10491 );
and ( n10755 , n10491 , n10496 );
and ( n10756 , n10487 , n10496 );
or ( n10757 , n10754 , n10755 , n10756 );
and ( n10758 , n10420 , n10427 );
xor ( n10759 , n10757 , n10758 );
and ( n10760 , n7966 , n8294 );
and ( n10761 , n8116 , n8110 );
nor ( n10762 , n10760 , n10761 );
xnor ( n10763 , n10762 , n8250 );
xor ( n10764 , n10759 , n10763 );
xor ( n10765 , n10753 , n10764 );
xor ( n10766 , n10744 , n10765 );
xor ( n10767 , n10735 , n10766 );
xor ( n10768 , n10654 , n10767 );
and ( n10769 , n10381 , n10383 );
and ( n10770 , n10383 , n10501 );
and ( n10771 , n10381 , n10501 );
or ( n10772 , n10769 , n10770 , n10771 );
xor ( n10773 , n10768 , n10772 );
and ( n10774 , n10502 , n10506 );
and ( n10775 , n10507 , n10510 );
or ( n10776 , n10774 , n10775 );
xor ( n10777 , n10773 , n10776 );
buf ( n10778 , n10777 );
not ( n10779 , n831 );
and ( n10780 , n10779 , n10647 );
and ( n10781 , n10778 , n831 );
or ( n10782 , n10780 , n10781 );
and ( n10783 , n10527 , n10603 );
and ( n10784 , n10603 , n10635 );
and ( n10785 , n10527 , n10635 );
or ( n10786 , n10783 , n10784 , n10785 );
buf ( n10787 , n870 );
buf ( n10788 , n10787 );
xor ( n10789 , n10786 , n10788 );
and ( n10790 , n10608 , n10612 );
and ( n10791 , n10612 , n10634 );
and ( n10792 , n10608 , n10634 );
or ( n10793 , n10790 , n10791 , n10792 );
and ( n10794 , n10582 , n10586 );
and ( n10795 , n10586 , n10601 );
and ( n10796 , n10582 , n10601 );
or ( n10797 , n10794 , n10795 , n10796 );
and ( n10798 , n10090 , n7063 );
and ( n10799 , n10331 , n7005 );
nor ( n10800 , n10798 , n10799 );
xnor ( n10801 , n10800 , n7058 );
not ( n10802 , n10544 );
buf ( n10803 , n806 );
buf ( n10804 , n10803 );
and ( n10805 , n10542 , n10288 );
not ( n10806 , n10805 );
and ( n10807 , n10804 , n10806 );
and ( n10808 , n10802 , n10807 );
xor ( n10809 , n10801 , n10808 );
and ( n10810 , n10551 , n10555 );
and ( n10811 , n10555 , n10560 );
and ( n10812 , n10551 , n10560 );
or ( n10813 , n10810 , n10811 , n10812 );
xor ( n10814 , n10809 , n10813 );
and ( n10815 , n10566 , n10570 );
and ( n10816 , n10570 , n10575 );
and ( n10817 , n10566 , n10575 );
or ( n10818 , n10815 , n10816 , n10817 );
xor ( n10819 , n10814 , n10818 );
xor ( n10820 , n10797 , n10819 );
and ( n10821 , n8690 , n7609 );
and ( n10822 , n8913 , n7505 );
nor ( n10823 , n10821 , n10822 );
xnor ( n10824 , n10823 , n7615 );
and ( n10825 , n7292 , n9311 );
and ( n10826 , n7372 , n9150 );
nor ( n10827 , n10825 , n10826 );
xnor ( n10828 , n10827 , n9317 );
xor ( n10829 , n10824 , n10828 );
and ( n10830 , n7125 , n9795 );
and ( n10831 , n7196 , n9560 );
nor ( n10832 , n10830 , n10831 );
xnor ( n10833 , n10832 , n9801 );
xor ( n10834 , n10829 , n10833 );
and ( n10835 , n10548 , n6957 );
buf ( n10836 , n774 );
buf ( n10837 , n10836 );
and ( n10838 , n10837 , n6934 );
nor ( n10839 , n10835 , n10838 );
xnor ( n10840 , n10839 , n6954 );
and ( n10841 , n8339 , n7873 );
and ( n10842 , n8548 , n7762 );
nor ( n10843 , n10841 , n10842 );
xnor ( n10844 , n10843 , n7863 );
xor ( n10845 , n10840 , n10844 );
and ( n10846 , n6999 , n10342 );
and ( n10847 , n7049 , n10084 );
nor ( n10848 , n10846 , n10847 );
xnor ( n10849 , n10848 , n10291 );
xor ( n10850 , n10845 , n10849 );
xor ( n10851 , n10834 , n10850 );
and ( n10852 , n9139 , n7400 );
and ( n10853 , n9323 , n7303 );
nor ( n10854 , n10852 , n10853 );
xnor ( n10855 , n10854 , n7381 );
and ( n10856 , n7730 , n8511 );
and ( n10857 , n7891 , n8350 );
nor ( n10858 , n10856 , n10857 );
xnor ( n10859 , n10858 , n8517 );
xor ( n10860 , n10855 , n10859 );
and ( n10861 , n7494 , n8887 );
and ( n10862 , n7596 , n8701 );
nor ( n10863 , n10861 , n10862 );
xnor ( n10864 , n10863 , n8893 );
xor ( n10865 , n10860 , n10864 );
xor ( n10866 , n10851 , n10865 );
xor ( n10867 , n10820 , n10866 );
xor ( n10868 , n10793 , n10867 );
and ( n10869 , n10617 , n10621 );
and ( n10870 , n10621 , n10633 );
and ( n10871 , n10617 , n10633 );
or ( n10872 , n10869 , n10870 , n10871 );
and ( n10873 , n10531 , n10577 );
and ( n10874 , n10577 , n10602 );
and ( n10875 , n10531 , n10602 );
or ( n10876 , n10873 , n10874 , n10875 );
xor ( n10877 , n10872 , n10876 );
and ( n10878 , n10626 , n10627 );
and ( n10879 , n10627 , n10632 );
and ( n10880 , n10626 , n10632 );
or ( n10881 , n10878 , n10879 , n10880 );
and ( n10882 , n10545 , n10561 );
and ( n10883 , n10561 , n10576 );
and ( n10884 , n10545 , n10576 );
or ( n10885 , n10882 , n10883 , n10884 );
xor ( n10886 , n10881 , n10885 );
and ( n10887 , n10535 , n10539 );
and ( n10888 , n10539 , n10544 );
and ( n10889 , n10535 , n10544 );
or ( n10890 , n10887 , n10888 , n10889 );
and ( n10891 , n10591 , n10595 );
and ( n10892 , n10595 , n10600 );
and ( n10893 , n10591 , n10600 );
or ( n10894 , n10891 , n10892 , n10893 );
xor ( n10895 , n10890 , n10894 );
and ( n10896 , n9549 , n7215 );
and ( n10897 , n9839 , n7136 );
nor ( n10898 , n10896 , n10897 );
xnor ( n10899 , n10898 , n7205 );
and ( n10900 , n8045 , n8209 );
and ( n10901 , n8156 , n8039 );
nor ( n10902 , n10900 , n10901 );
xnor ( n10903 , n10902 , n8165 );
xor ( n10904 , n10899 , n10903 );
xor ( n10905 , n10804 , n10542 );
not ( n10906 , n10543 );
and ( n10907 , n10905 , n10906 );
and ( n10908 , n6932 , n10907 );
and ( n10909 , n6960 , n10543 );
nor ( n10910 , n10908 , n10909 );
xnor ( n10911 , n10910 , n10807 );
xor ( n10912 , n10904 , n10911 );
xor ( n10913 , n10895 , n10912 );
xor ( n10914 , n10886 , n10913 );
xor ( n10915 , n10877 , n10914 );
xor ( n10916 , n10868 , n10915 );
xor ( n10917 , n10789 , n10916 );
and ( n10918 , n10520 , n10522 );
and ( n10919 , n10522 , n10636 );
and ( n10920 , n10520 , n10636 );
or ( n10921 , n10918 , n10919 , n10920 );
xor ( n10922 , n10917 , n10921 );
and ( n10923 , n10637 , n10641 );
and ( n10924 , n10642 , n10645 );
or ( n10925 , n10923 , n10924 );
xor ( n10926 , n10922 , n10925 );
buf ( n10927 , n10926 );
and ( n10928 , n10658 , n10734 );
and ( n10929 , n10734 , n10766 );
and ( n10930 , n10658 , n10766 );
or ( n10931 , n10928 , n10929 , n10930 );
buf ( n10932 , n838 );
buf ( n10933 , n10932 );
xor ( n10934 , n10931 , n10933 );
and ( n10935 , n10739 , n10743 );
and ( n10936 , n10743 , n10765 );
and ( n10937 , n10739 , n10765 );
or ( n10938 , n10935 , n10936 , n10937 );
and ( n10939 , n10713 , n10717 );
and ( n10940 , n10717 , n10732 );
and ( n10941 , n10713 , n10732 );
or ( n10942 , n10939 , n10940 , n10941 );
and ( n10943 , n10211 , n7098 );
and ( n10944 , n10466 , n7026 );
nor ( n10945 , n10943 , n10944 );
xnor ( n10946 , n10945 , n7093 );
not ( n10947 , n10675 );
buf ( n10948 , n806 );
buf ( n10949 , n10948 );
and ( n10950 , n10673 , n10423 );
not ( n10951 , n10950 );
and ( n10952 , n10949 , n10951 );
and ( n10953 , n10947 , n10952 );
xor ( n10954 , n10946 , n10953 );
and ( n10955 , n10682 , n10686 );
and ( n10956 , n10686 , n10691 );
and ( n10957 , n10682 , n10691 );
or ( n10958 , n10955 , n10956 , n10957 );
xor ( n10959 , n10954 , n10958 );
and ( n10960 , n10697 , n10701 );
and ( n10961 , n10701 , n10706 );
and ( n10962 , n10697 , n10706 );
or ( n10963 , n10960 , n10961 , n10962 );
xor ( n10964 , n10959 , n10963 );
xor ( n10965 , n10942 , n10964 );
and ( n10966 , n8781 , n7674 );
and ( n10967 , n9018 , n7556 );
nor ( n10968 , n10966 , n10967 );
xnor ( n10969 , n10968 , n7680 );
and ( n10970 , n7333 , n9426 );
and ( n10971 , n7427 , n9251 );
nor ( n10972 , n10970 , n10971 );
xnor ( n10973 , n10972 , n9432 );
xor ( n10974 , n10969 , n10973 );
and ( n10975 , n7156 , n9920 );
and ( n10976 , n7241 , n9671 );
nor ( n10977 , n10975 , n10976 );
xnor ( n10978 , n10977 , n9926 );
xor ( n10979 , n10974 , n10978 );
and ( n10980 , n10679 , n6977 );
buf ( n10981 , n774 );
buf ( n10982 , n10981 );
and ( n10983 , n10982 , n6943 );
nor ( n10984 , n10980 , n10983 );
xnor ( n10985 , n10984 , n6974 );
and ( n10986 , n8420 , n7948 );
and ( n10987 , n8643 , n7823 );
nor ( n10988 , n10986 , n10987 );
xnor ( n10989 , n10988 , n7938 );
xor ( n10990 , n10985 , n10989 );
and ( n10991 , n7020 , n10477 );
and ( n10992 , n7084 , n10205 );
nor ( n10993 , n10991 , n10992 );
xnor ( n10994 , n10993 , n10426 );
xor ( n10995 , n10990 , n10994 );
xor ( n10996 , n10979 , n10995 );
and ( n10997 , n9240 , n7455 );
and ( n10998 , n9438 , n7344 );
nor ( n10999 , n10997 , n10998 );
xnor ( n11000 , n10999 , n7436 );
and ( n11001 , n7791 , n8606 );
and ( n11002 , n7966 , n8431 );
nor ( n11003 , n11001 , n11002 );
xnor ( n11004 , n11003 , n8612 );
xor ( n11005 , n11000 , n11004 );
and ( n11006 , n7545 , n8992 );
and ( n11007 , n7661 , n8792 );
nor ( n11008 , n11006 , n11007 );
xnor ( n11009 , n11008 , n8998 );
xor ( n11010 , n11005 , n11009 );
xor ( n11011 , n10996 , n11010 );
xor ( n11012 , n10965 , n11011 );
xor ( n11013 , n10938 , n11012 );
and ( n11014 , n10748 , n10752 );
and ( n11015 , n10752 , n10764 );
and ( n11016 , n10748 , n10764 );
or ( n11017 , n11014 , n11015 , n11016 );
and ( n11018 , n10662 , n10708 );
and ( n11019 , n10708 , n10733 );
and ( n11020 , n10662 , n10733 );
or ( n11021 , n11018 , n11019 , n11020 );
xor ( n11022 , n11017 , n11021 );
and ( n11023 , n10757 , n10758 );
and ( n11024 , n10758 , n10763 );
and ( n11025 , n10757 , n10763 );
or ( n11026 , n11023 , n11024 , n11025 );
and ( n11027 , n10676 , n10692 );
and ( n11028 , n10692 , n10707 );
and ( n11029 , n10676 , n10707 );
or ( n11030 , n11027 , n11028 , n11029 );
xor ( n11031 , n11026 , n11030 );
and ( n11032 , n10666 , n10670 );
and ( n11033 , n10670 , n10675 );
and ( n11034 , n10666 , n10675 );
or ( n11035 , n11032 , n11033 , n11034 );
and ( n11036 , n10722 , n10726 );
and ( n11037 , n10726 , n10731 );
and ( n11038 , n10722 , n10731 );
or ( n11039 , n11036 , n11037 , n11038 );
xor ( n11040 , n11035 , n11039 );
and ( n11041 , n9660 , n7260 );
and ( n11042 , n9964 , n7167 );
nor ( n11043 , n11041 , n11042 );
xnor ( n11044 , n11043 , n7250 );
and ( n11045 , n8116 , n8294 );
and ( n11046 , n8241 , n8110 );
nor ( n11047 , n11045 , n11046 );
xnor ( n11048 , n11047 , n8250 );
xor ( n11049 , n11044 , n11048 );
xor ( n11050 , n10949 , n10673 );
not ( n11051 , n10674 );
and ( n11052 , n11050 , n11051 );
and ( n11053 , n6941 , n11052 );
and ( n11054 , n6980 , n10674 );
nor ( n11055 , n11053 , n11054 );
xnor ( n11056 , n11055 , n10952 );
xor ( n11057 , n11049 , n11056 );
xor ( n11058 , n11040 , n11057 );
xor ( n11059 , n11031 , n11058 );
xor ( n11060 , n11022 , n11059 );
xor ( n11061 , n11013 , n11060 );
xor ( n11062 , n10934 , n11061 );
and ( n11063 , n10651 , n10653 );
and ( n11064 , n10653 , n10767 );
and ( n11065 , n10651 , n10767 );
or ( n11066 , n11063 , n11064 , n11065 );
xor ( n11067 , n11062 , n11066 );
and ( n11068 , n10768 , n10772 );
and ( n11069 , n10773 , n10776 );
or ( n11070 , n11068 , n11069 );
xor ( n11071 , n11067 , n11070 );
buf ( n11072 , n11071 );
not ( n11073 , n831 );
and ( n11074 , n11073 , n10927 );
and ( n11075 , n11072 , n831 );
or ( n11076 , n11074 , n11075 );
and ( n11077 , n10793 , n10867 );
and ( n11078 , n10867 , n10915 );
and ( n11079 , n10793 , n10915 );
or ( n11080 , n11077 , n11078 , n11079 );
buf ( n11081 , n869 );
buf ( n11082 , n11081 );
xor ( n11083 , n11080 , n11082 );
and ( n11084 , n10872 , n10876 );
and ( n11085 , n10876 , n10914 );
and ( n11086 , n10872 , n10914 );
or ( n11087 , n11084 , n11085 , n11086 );
and ( n11088 , n10881 , n10885 );
and ( n11089 , n10885 , n10913 );
and ( n11090 , n10881 , n10913 );
or ( n11091 , n11088 , n11089 , n11090 );
and ( n11092 , n10797 , n10819 );
and ( n11093 , n10819 , n10866 );
and ( n11094 , n10797 , n10866 );
or ( n11095 , n11092 , n11093 , n11094 );
xor ( n11096 , n11091 , n11095 );
and ( n11097 , n10809 , n10813 );
and ( n11098 , n10813 , n10818 );
and ( n11099 , n10809 , n10818 );
or ( n11100 , n11097 , n11098 , n11099 );
and ( n11101 , n10890 , n10894 );
and ( n11102 , n10894 , n10912 );
and ( n11103 , n10890 , n10912 );
or ( n11104 , n11101 , n11102 , n11103 );
xor ( n11105 , n11100 , n11104 );
and ( n11106 , n10834 , n10850 );
and ( n11107 , n10850 , n10865 );
and ( n11108 , n10834 , n10865 );
or ( n11109 , n11106 , n11107 , n11108 );
xor ( n11110 , n11105 , n11109 );
xor ( n11111 , n11096 , n11110 );
xor ( n11112 , n11087 , n11111 );
and ( n11113 , n10824 , n10828 );
and ( n11114 , n10828 , n10833 );
and ( n11115 , n10824 , n10833 );
or ( n11116 , n11113 , n11114 , n11115 );
and ( n11117 , n10840 , n10844 );
and ( n11118 , n10844 , n10849 );
and ( n11119 , n10840 , n10849 );
or ( n11120 , n11117 , n11118 , n11119 );
xor ( n11121 , n11116 , n11120 );
and ( n11122 , n10855 , n10859 );
and ( n11123 , n10859 , n10864 );
and ( n11124 , n10855 , n10864 );
or ( n11125 , n11122 , n11123 , n11124 );
xor ( n11126 , n11121 , n11125 );
and ( n11127 , n10899 , n10903 );
and ( n11128 , n10903 , n10911 );
and ( n11129 , n10899 , n10911 );
or ( n11130 , n11127 , n11128 , n11129 );
and ( n11131 , n10837 , n6957 );
buf ( n11132 , n773 );
buf ( n11133 , n11132 );
and ( n11134 , n11133 , n6934 );
nor ( n11135 , n11131 , n11134 );
xnor ( n11136 , n11135 , n6954 );
and ( n11137 , n7372 , n9311 );
and ( n11138 , n7494 , n9150 );
nor ( n11139 , n11137 , n11138 );
xnor ( n11140 , n11139 , n9317 );
xor ( n11141 , n11136 , n11140 );
and ( n11142 , n7196 , n9795 );
and ( n11143 , n7292 , n9560 );
nor ( n11144 , n11142 , n11143 );
xnor ( n11145 , n11144 , n9801 );
xor ( n11146 , n11141 , n11145 );
xor ( n11147 , n11130 , n11146 );
and ( n11148 , n10331 , n7063 );
and ( n11149 , n10548 , n7005 );
nor ( n11150 , n11148 , n11149 );
xnor ( n11151 , n11150 , n7058 );
and ( n11152 , n9323 , n7400 );
and ( n11153 , n9549 , n7303 );
nor ( n11154 , n11152 , n11153 );
xnor ( n11155 , n11154 , n7381 );
xor ( n11156 , n11151 , n11155 );
buf ( n11157 , n805 );
buf ( n11158 , n11157 );
xor ( n11159 , n11158 , n10804 );
and ( n11160 , n6932 , n11159 );
xor ( n11161 , n11156 , n11160 );
xor ( n11162 , n11147 , n11161 );
xor ( n11163 , n11126 , n11162 );
and ( n11164 , n8548 , n7873 );
and ( n11165 , n8690 , n7762 );
nor ( n11166 , n11164 , n11165 );
xnor ( n11167 , n11166 , n7863 );
and ( n11168 , n7049 , n10342 );
and ( n11169 , n7125 , n10084 );
nor ( n11170 , n11168 , n11169 );
xnor ( n11171 , n11170 , n10291 );
xor ( n11172 , n11167 , n11171 );
and ( n11173 , n6960 , n10907 );
and ( n11174 , n6999 , n10543 );
nor ( n11175 , n11173 , n11174 );
xnor ( n11176 , n11175 , n10807 );
xor ( n11177 , n11172 , n11176 );
and ( n11178 , n8913 , n7609 );
and ( n11179 , n9139 , n7505 );
nor ( n11180 , n11178 , n11179 );
xnor ( n11181 , n11180 , n7615 );
and ( n11182 , n7891 , n8511 );
and ( n11183 , n8045 , n8350 );
nor ( n11184 , n11182 , n11183 );
xnor ( n11185 , n11184 , n8517 );
xor ( n11186 , n11181 , n11185 );
and ( n11187 , n7596 , n8887 );
and ( n11188 , n7730 , n8701 );
nor ( n11189 , n11187 , n11188 );
xnor ( n11190 , n11189 , n8893 );
xor ( n11191 , n11186 , n11190 );
xor ( n11192 , n11177 , n11191 );
and ( n11193 , n10801 , n10808 );
and ( n11194 , n9839 , n7215 );
and ( n11195 , n10090 , n7136 );
nor ( n11196 , n11194 , n11195 );
xnor ( n11197 , n11196 , n7205 );
xor ( n11198 , n11193 , n11197 );
and ( n11199 , n8156 , n8209 );
and ( n11200 , n8339 , n8039 );
nor ( n11201 , n11199 , n11200 );
xnor ( n11202 , n11201 , n8165 );
xor ( n11203 , n11198 , n11202 );
xor ( n11204 , n11192 , n11203 );
xor ( n11205 , n11163 , n11204 );
xor ( n11206 , n11112 , n11205 );
xor ( n11207 , n11083 , n11206 );
and ( n11208 , n10786 , n10788 );
and ( n11209 , n10788 , n10916 );
and ( n11210 , n10786 , n10916 );
or ( n11211 , n11208 , n11209 , n11210 );
xor ( n11212 , n11207 , n11211 );
and ( n11213 , n10917 , n10921 );
and ( n11214 , n10922 , n10925 );
or ( n11215 , n11213 , n11214 );
xor ( n11216 , n11212 , n11215 );
buf ( n11217 , n11216 );
and ( n11218 , n10938 , n11012 );
and ( n11219 , n11012 , n11060 );
and ( n11220 , n10938 , n11060 );
or ( n11221 , n11218 , n11219 , n11220 );
buf ( n11222 , n837 );
buf ( n11223 , n11222 );
xor ( n11224 , n11221 , n11223 );
and ( n11225 , n11017 , n11021 );
and ( n11226 , n11021 , n11059 );
and ( n11227 , n11017 , n11059 );
or ( n11228 , n11225 , n11226 , n11227 );
and ( n11229 , n11026 , n11030 );
and ( n11230 , n11030 , n11058 );
and ( n11231 , n11026 , n11058 );
or ( n11232 , n11229 , n11230 , n11231 );
and ( n11233 , n10942 , n10964 );
and ( n11234 , n10964 , n11011 );
and ( n11235 , n10942 , n11011 );
or ( n11236 , n11233 , n11234 , n11235 );
xor ( n11237 , n11232 , n11236 );
and ( n11238 , n10954 , n10958 );
and ( n11239 , n10958 , n10963 );
and ( n11240 , n10954 , n10963 );
or ( n11241 , n11238 , n11239 , n11240 );
and ( n11242 , n11035 , n11039 );
and ( n11243 , n11039 , n11057 );
and ( n11244 , n11035 , n11057 );
or ( n11245 , n11242 , n11243 , n11244 );
xor ( n11246 , n11241 , n11245 );
and ( n11247 , n10979 , n10995 );
and ( n11248 , n10995 , n11010 );
and ( n11249 , n10979 , n11010 );
or ( n11250 , n11247 , n11248 , n11249 );
xor ( n11251 , n11246 , n11250 );
xor ( n11252 , n11237 , n11251 );
xor ( n11253 , n11228 , n11252 );
and ( n11254 , n10969 , n10973 );
and ( n11255 , n10973 , n10978 );
and ( n11256 , n10969 , n10978 );
or ( n11257 , n11254 , n11255 , n11256 );
and ( n11258 , n10985 , n10989 );
and ( n11259 , n10989 , n10994 );
and ( n11260 , n10985 , n10994 );
or ( n11261 , n11258 , n11259 , n11260 );
xor ( n11262 , n11257 , n11261 );
and ( n11263 , n11000 , n11004 );
and ( n11264 , n11004 , n11009 );
and ( n11265 , n11000 , n11009 );
or ( n11266 , n11263 , n11264 , n11265 );
xor ( n11267 , n11262 , n11266 );
and ( n11268 , n11044 , n11048 );
and ( n11269 , n11048 , n11056 );
and ( n11270 , n11044 , n11056 );
or ( n11271 , n11268 , n11269 , n11270 );
and ( n11272 , n10982 , n6977 );
buf ( n11273 , n773 );
buf ( n11274 , n11273 );
and ( n11275 , n11274 , n6943 );
nor ( n11276 , n11272 , n11275 );
xnor ( n11277 , n11276 , n6974 );
and ( n11278 , n7427 , n9426 );
and ( n11279 , n7545 , n9251 );
nor ( n11280 , n11278 , n11279 );
xnor ( n11281 , n11280 , n9432 );
xor ( n11282 , n11277 , n11281 );
and ( n11283 , n7241 , n9920 );
and ( n11284 , n7333 , n9671 );
nor ( n11285 , n11283 , n11284 );
xnor ( n11286 , n11285 , n9926 );
xor ( n11287 , n11282 , n11286 );
xor ( n11288 , n11271 , n11287 );
and ( n11289 , n10466 , n7098 );
and ( n11290 , n10679 , n7026 );
nor ( n11291 , n11289 , n11290 );
xnor ( n11292 , n11291 , n7093 );
and ( n11293 , n9438 , n7455 );
and ( n11294 , n9660 , n7344 );
nor ( n11295 , n11293 , n11294 );
xnor ( n11296 , n11295 , n7436 );
xor ( n11297 , n11292 , n11296 );
buf ( n11298 , n805 );
buf ( n11299 , n11298 );
xor ( n11300 , n11299 , n10949 );
and ( n11301 , n6941 , n11300 );
xor ( n11302 , n11297 , n11301 );
xor ( n11303 , n11288 , n11302 );
xor ( n11304 , n11267 , n11303 );
and ( n11305 , n8643 , n7948 );
and ( n11306 , n8781 , n7823 );
nor ( n11307 , n11305 , n11306 );
xnor ( n11308 , n11307 , n7938 );
and ( n11309 , n7084 , n10477 );
and ( n11310 , n7156 , n10205 );
nor ( n11311 , n11309 , n11310 );
xnor ( n11312 , n11311 , n10426 );
xor ( n11313 , n11308 , n11312 );
and ( n11314 , n6980 , n11052 );
and ( n11315 , n7020 , n10674 );
nor ( n11316 , n11314 , n11315 );
xnor ( n11317 , n11316 , n10952 );
xor ( n11318 , n11313 , n11317 );
and ( n11319 , n9018 , n7674 );
and ( n11320 , n9240 , n7556 );
nor ( n11321 , n11319 , n11320 );
xnor ( n11322 , n11321 , n7680 );
and ( n11323 , n7966 , n8606 );
and ( n11324 , n8116 , n8431 );
nor ( n11325 , n11323 , n11324 );
xnor ( n11326 , n11325 , n8612 );
xor ( n11327 , n11322 , n11326 );
and ( n11328 , n7661 , n8992 );
and ( n11329 , n7791 , n8792 );
nor ( n11330 , n11328 , n11329 );
xnor ( n11331 , n11330 , n8998 );
xor ( n11332 , n11327 , n11331 );
xor ( n11333 , n11318 , n11332 );
and ( n11334 , n10946 , n10953 );
and ( n11335 , n9964 , n7260 );
and ( n11336 , n10211 , n7167 );
nor ( n11337 , n11335 , n11336 );
xnor ( n11338 , n11337 , n7250 );
xor ( n11339 , n11334 , n11338 );
and ( n11340 , n8241 , n8294 );
and ( n11341 , n8420 , n8110 );
nor ( n11342 , n11340 , n11341 );
xnor ( n11343 , n11342 , n8250 );
xor ( n11344 , n11339 , n11343 );
xor ( n11345 , n11333 , n11344 );
xor ( n11346 , n11304 , n11345 );
xor ( n11347 , n11253 , n11346 );
xor ( n11348 , n11224 , n11347 );
and ( n11349 , n10931 , n10933 );
and ( n11350 , n10933 , n11061 );
and ( n11351 , n10931 , n11061 );
or ( n11352 , n11349 , n11350 , n11351 );
xor ( n11353 , n11348 , n11352 );
and ( n11354 , n11062 , n11066 );
and ( n11355 , n11067 , n11070 );
or ( n11356 , n11354 , n11355 );
xor ( n11357 , n11353 , n11356 );
buf ( n11358 , n11357 );
not ( n11359 , n831 );
and ( n11360 , n11359 , n11217 );
and ( n11361 , n11358 , n831 );
or ( n11362 , n11360 , n11361 );
and ( n11363 , n11080 , n11082 );
and ( n11364 , n11082 , n11206 );
and ( n11365 , n11080 , n11206 );
or ( n11366 , n11363 , n11364 , n11365 );
and ( n11367 , n11087 , n11111 );
and ( n11368 , n11111 , n11205 );
and ( n11369 , n11087 , n11205 );
or ( n11370 , n11367 , n11368 , n11369 );
buf ( n11371 , n868 );
buf ( n11372 , n11371 );
xor ( n11373 , n11370 , n11372 );
and ( n11374 , n11091 , n11095 );
and ( n11375 , n11095 , n11110 );
and ( n11376 , n11091 , n11110 );
or ( n11377 , n11374 , n11375 , n11376 );
and ( n11378 , n11177 , n11191 );
and ( n11379 , n11191 , n11203 );
and ( n11380 , n11177 , n11203 );
or ( n11381 , n11378 , n11379 , n11380 );
and ( n11382 , n11133 , n6957 );
buf ( n11383 , n772 );
buf ( n11384 , n11383 );
and ( n11385 , n11384 , n6934 );
nor ( n11386 , n11382 , n11385 );
xnor ( n11387 , n11386 , n6954 );
and ( n11388 , n8690 , n7873 );
and ( n11389 , n8913 , n7762 );
nor ( n11390 , n11388 , n11389 );
xnor ( n11391 , n11390 , n7863 );
xor ( n11392 , n11387 , n11391 );
and ( n11393 , n7125 , n10342 );
and ( n11394 , n7196 , n10084 );
nor ( n11395 , n11393 , n11394 );
xnor ( n11396 , n11395 , n10291 );
xor ( n11397 , n11392 , n11396 );
and ( n11398 , n10090 , n7215 );
and ( n11399 , n10331 , n7136 );
nor ( n11400 , n11398 , n11399 );
xnor ( n11401 , n11400 , n7205 );
and ( n11402 , n6999 , n10907 );
and ( n11403 , n7049 , n10543 );
nor ( n11404 , n11402 , n11403 );
xnor ( n11405 , n11404 , n10807 );
xor ( n11406 , n11401 , n11405 );
buf ( n11407 , n804 );
buf ( n11408 , n11407 );
xor ( n11409 , n11408 , n11158 );
not ( n11410 , n11159 );
and ( n11411 , n11409 , n11410 );
and ( n11412 , n6932 , n11411 );
and ( n11413 , n6960 , n11159 );
nor ( n11414 , n11412 , n11413 );
and ( n11415 , n11158 , n10804 );
not ( n11416 , n11415 );
and ( n11417 , n11408 , n11416 );
xnor ( n11418 , n11414 , n11417 );
xor ( n11419 , n11406 , n11418 );
xor ( n11420 , n11397 , n11419 );
and ( n11421 , n9549 , n7400 );
and ( n11422 , n9839 , n7303 );
nor ( n11423 , n11421 , n11422 );
xnor ( n11424 , n11423 , n7381 );
and ( n11425 , n8045 , n8511 );
and ( n11426 , n8156 , n8350 );
nor ( n11427 , n11425 , n11426 );
xnor ( n11428 , n11427 , n8517 );
xor ( n11429 , n11424 , n11428 );
and ( n11430 , n7730 , n8887 );
and ( n11431 , n7891 , n8701 );
nor ( n11432 , n11430 , n11431 );
xnor ( n11433 , n11432 , n8893 );
xor ( n11434 , n11429 , n11433 );
xor ( n11435 , n11420 , n11434 );
xor ( n11436 , n11381 , n11435 );
and ( n11437 , n11193 , n11197 );
and ( n11438 , n11197 , n11202 );
and ( n11439 , n11193 , n11202 );
or ( n11440 , n11437 , n11438 , n11439 );
and ( n11441 , n9139 , n7609 );
and ( n11442 , n9323 , n7505 );
nor ( n11443 , n11441 , n11442 );
xnor ( n11444 , n11443 , n7615 );
and ( n11445 , n7494 , n9311 );
and ( n11446 , n7596 , n9150 );
nor ( n11447 , n11445 , n11446 );
xnor ( n11448 , n11447 , n9317 );
xor ( n11449 , n11444 , n11448 );
and ( n11450 , n7292 , n9795 );
and ( n11451 , n7372 , n9560 );
nor ( n11452 , n11450 , n11451 );
xnor ( n11453 , n11452 , n9801 );
xor ( n11454 , n11449 , n11453 );
xor ( n11455 , n11440 , n11454 );
and ( n11456 , n10548 , n7063 );
and ( n11457 , n10837 , n7005 );
nor ( n11458 , n11456 , n11457 );
xnor ( n11459 , n11458 , n7058 );
not ( n11460 , n11160 );
and ( n11461 , n11460 , n11417 );
xor ( n11462 , n11459 , n11461 );
and ( n11463 , n11151 , n11155 );
and ( n11464 , n11155 , n11160 );
and ( n11465 , n11151 , n11160 );
or ( n11466 , n11463 , n11464 , n11465 );
xor ( n11467 , n11462 , n11466 );
and ( n11468 , n8339 , n8209 );
and ( n11469 , n8548 , n8039 );
nor ( n11470 , n11468 , n11469 );
xnor ( n11471 , n11470 , n8165 );
xor ( n11472 , n11467 , n11471 );
xor ( n11473 , n11455 , n11472 );
xor ( n11474 , n11436 , n11473 );
xor ( n11475 , n11377 , n11474 );
and ( n11476 , n11100 , n11104 );
and ( n11477 , n11104 , n11109 );
and ( n11478 , n11100 , n11109 );
or ( n11479 , n11476 , n11477 , n11478 );
and ( n11480 , n11126 , n11162 );
and ( n11481 , n11162 , n11204 );
and ( n11482 , n11126 , n11204 );
or ( n11483 , n11480 , n11481 , n11482 );
xor ( n11484 , n11479 , n11483 );
and ( n11485 , n11116 , n11120 );
and ( n11486 , n11120 , n11125 );
and ( n11487 , n11116 , n11125 );
or ( n11488 , n11485 , n11486 , n11487 );
and ( n11489 , n11130 , n11146 );
and ( n11490 , n11146 , n11161 );
and ( n11491 , n11130 , n11161 );
or ( n11492 , n11489 , n11490 , n11491 );
xor ( n11493 , n11488 , n11492 );
and ( n11494 , n11136 , n11140 );
and ( n11495 , n11140 , n11145 );
and ( n11496 , n11136 , n11145 );
or ( n11497 , n11494 , n11495 , n11496 );
and ( n11498 , n11167 , n11171 );
and ( n11499 , n11171 , n11176 );
and ( n11500 , n11167 , n11176 );
or ( n11501 , n11498 , n11499 , n11500 );
xor ( n11502 , n11497 , n11501 );
and ( n11503 , n11181 , n11185 );
and ( n11504 , n11185 , n11190 );
and ( n11505 , n11181 , n11190 );
or ( n11506 , n11503 , n11504 , n11505 );
xor ( n11507 , n11502 , n11506 );
xor ( n11508 , n11493 , n11507 );
xor ( n11509 , n11484 , n11508 );
xor ( n11510 , n11475 , n11509 );
xor ( n11511 , n11373 , n11510 );
xor ( n11512 , n11366 , n11511 );
and ( n11513 , n11207 , n11211 );
and ( n11514 , n11212 , n11215 );
or ( n11515 , n11513 , n11514 );
xor ( n11516 , n11512 , n11515 );
buf ( n11517 , n11516 );
and ( n11518 , n11221 , n11223 );
and ( n11519 , n11223 , n11347 );
and ( n11520 , n11221 , n11347 );
or ( n11521 , n11518 , n11519 , n11520 );
and ( n11522 , n11228 , n11252 );
and ( n11523 , n11252 , n11346 );
and ( n11524 , n11228 , n11346 );
or ( n11525 , n11522 , n11523 , n11524 );
buf ( n11526 , n836 );
buf ( n11527 , n11526 );
xor ( n11528 , n11525 , n11527 );
and ( n11529 , n11232 , n11236 );
and ( n11530 , n11236 , n11251 );
and ( n11531 , n11232 , n11251 );
or ( n11532 , n11529 , n11530 , n11531 );
and ( n11533 , n11318 , n11332 );
and ( n11534 , n11332 , n11344 );
and ( n11535 , n11318 , n11344 );
or ( n11536 , n11533 , n11534 , n11535 );
and ( n11537 , n11274 , n6977 );
buf ( n11538 , n772 );
buf ( n11539 , n11538 );
and ( n11540 , n11539 , n6943 );
nor ( n11541 , n11537 , n11540 );
xnor ( n11542 , n11541 , n6974 );
and ( n11543 , n8781 , n7948 );
and ( n11544 , n9018 , n7823 );
nor ( n11545 , n11543 , n11544 );
xnor ( n11546 , n11545 , n7938 );
xor ( n11547 , n11542 , n11546 );
and ( n11548 , n7156 , n10477 );
and ( n11549 , n7241 , n10205 );
nor ( n11550 , n11548 , n11549 );
xnor ( n11551 , n11550 , n10426 );
xor ( n11552 , n11547 , n11551 );
and ( n11553 , n10211 , n7260 );
and ( n11554 , n10466 , n7167 );
nor ( n11555 , n11553 , n11554 );
xnor ( n11556 , n11555 , n7250 );
and ( n11557 , n7020 , n11052 );
and ( n11558 , n7084 , n10674 );
nor ( n11559 , n11557 , n11558 );
xnor ( n11560 , n11559 , n10952 );
xor ( n11561 , n11556 , n11560 );
buf ( n11562 , n804 );
buf ( n11563 , n11562 );
xor ( n11564 , n11563 , n11299 );
not ( n11565 , n11300 );
and ( n11566 , n11564 , n11565 );
and ( n11567 , n6941 , n11566 );
and ( n11568 , n6980 , n11300 );
nor ( n11569 , n11567 , n11568 );
and ( n11570 , n11299 , n10949 );
not ( n11571 , n11570 );
and ( n11572 , n11563 , n11571 );
xnor ( n11573 , n11569 , n11572 );
xor ( n11574 , n11561 , n11573 );
xor ( n11575 , n11552 , n11574 );
and ( n11576 , n9660 , n7455 );
and ( n11577 , n9964 , n7344 );
nor ( n11578 , n11576 , n11577 );
xnor ( n11579 , n11578 , n7436 );
and ( n11580 , n8116 , n8606 );
and ( n11581 , n8241 , n8431 );
nor ( n11582 , n11580 , n11581 );
xnor ( n11583 , n11582 , n8612 );
xor ( n11584 , n11579 , n11583 );
and ( n11585 , n7791 , n8992 );
and ( n11586 , n7966 , n8792 );
nor ( n11587 , n11585 , n11586 );
xnor ( n11588 , n11587 , n8998 );
xor ( n11589 , n11584 , n11588 );
xor ( n11590 , n11575 , n11589 );
xor ( n11591 , n11536 , n11590 );
and ( n11592 , n11334 , n11338 );
and ( n11593 , n11338 , n11343 );
and ( n11594 , n11334 , n11343 );
or ( n11595 , n11592 , n11593 , n11594 );
and ( n11596 , n9240 , n7674 );
and ( n11597 , n9438 , n7556 );
nor ( n11598 , n11596 , n11597 );
xnor ( n11599 , n11598 , n7680 );
and ( n11600 , n7545 , n9426 );
and ( n11601 , n7661 , n9251 );
nor ( n11602 , n11600 , n11601 );
xnor ( n11603 , n11602 , n9432 );
xor ( n11604 , n11599 , n11603 );
and ( n11605 , n7333 , n9920 );
and ( n11606 , n7427 , n9671 );
nor ( n11607 , n11605 , n11606 );
xnor ( n11608 , n11607 , n9926 );
xor ( n11609 , n11604 , n11608 );
xor ( n11610 , n11595 , n11609 );
and ( n11611 , n10679 , n7098 );
and ( n11612 , n10982 , n7026 );
nor ( n11613 , n11611 , n11612 );
xnor ( n11614 , n11613 , n7093 );
not ( n11615 , n11301 );
and ( n11616 , n11615 , n11572 );
xor ( n11617 , n11614 , n11616 );
and ( n11618 , n11292 , n11296 );
and ( n11619 , n11296 , n11301 );
and ( n11620 , n11292 , n11301 );
or ( n11621 , n11618 , n11619 , n11620 );
xor ( n11622 , n11617 , n11621 );
and ( n11623 , n8420 , n8294 );
and ( n11624 , n8643 , n8110 );
nor ( n11625 , n11623 , n11624 );
xnor ( n11626 , n11625 , n8250 );
xor ( n11627 , n11622 , n11626 );
xor ( n11628 , n11610 , n11627 );
xor ( n11629 , n11591 , n11628 );
xor ( n11630 , n11532 , n11629 );
and ( n11631 , n11241 , n11245 );
and ( n11632 , n11245 , n11250 );
and ( n11633 , n11241 , n11250 );
or ( n11634 , n11631 , n11632 , n11633 );
and ( n11635 , n11267 , n11303 );
and ( n11636 , n11303 , n11345 );
and ( n11637 , n11267 , n11345 );
or ( n11638 , n11635 , n11636 , n11637 );
xor ( n11639 , n11634 , n11638 );
and ( n11640 , n11257 , n11261 );
and ( n11641 , n11261 , n11266 );
and ( n11642 , n11257 , n11266 );
or ( n11643 , n11640 , n11641 , n11642 );
and ( n11644 , n11271 , n11287 );
and ( n11645 , n11287 , n11302 );
and ( n11646 , n11271 , n11302 );
or ( n11647 , n11644 , n11645 , n11646 );
xor ( n11648 , n11643 , n11647 );
and ( n11649 , n11277 , n11281 );
and ( n11650 , n11281 , n11286 );
and ( n11651 , n11277 , n11286 );
or ( n11652 , n11649 , n11650 , n11651 );
and ( n11653 , n11308 , n11312 );
and ( n11654 , n11312 , n11317 );
and ( n11655 , n11308 , n11317 );
or ( n11656 , n11653 , n11654 , n11655 );
xor ( n11657 , n11652 , n11656 );
and ( n11658 , n11322 , n11326 );
and ( n11659 , n11326 , n11331 );
and ( n11660 , n11322 , n11331 );
or ( n11661 , n11658 , n11659 , n11660 );
xor ( n11662 , n11657 , n11661 );
xor ( n11663 , n11648 , n11662 );
xor ( n11664 , n11639 , n11663 );
xor ( n11665 , n11630 , n11664 );
xor ( n11666 , n11528 , n11665 );
xor ( n11667 , n11521 , n11666 );
and ( n11668 , n11348 , n11352 );
and ( n11669 , n11353 , n11356 );
or ( n11670 , n11668 , n11669 );
xor ( n11671 , n11667 , n11670 );
buf ( n11672 , n11671 );
not ( n11673 , n831 );
and ( n11674 , n11673 , n11517 );
and ( n11675 , n11672 , n831 );
or ( n11676 , n11674 , n11675 );
and ( n11677 , n11377 , n11474 );
and ( n11678 , n11474 , n11509 );
and ( n11679 , n11377 , n11509 );
or ( n11680 , n11677 , n11678 , n11679 );
buf ( n11681 , n867 );
buf ( n11682 , n11681 );
xor ( n11683 , n11680 , n11682 );
and ( n11684 , n11479 , n11483 );
and ( n11685 , n11483 , n11508 );
and ( n11686 , n11479 , n11508 );
or ( n11687 , n11684 , n11685 , n11686 );
and ( n11688 , n11440 , n11454 );
and ( n11689 , n11454 , n11472 );
and ( n11690 , n11440 , n11472 );
or ( n11691 , n11688 , n11689 , n11690 );
and ( n11692 , n11488 , n11492 );
and ( n11693 , n11492 , n11507 );
and ( n11694 , n11488 , n11507 );
or ( n11695 , n11692 , n11693 , n11694 );
xor ( n11696 , n11691 , n11695 );
and ( n11697 , n11384 , n6957 );
buf ( n11698 , n771 );
buf ( n11699 , n11698 );
and ( n11700 , n11699 , n6934 );
nor ( n11701 , n11697 , n11700 );
xnor ( n11702 , n11701 , n6954 );
and ( n11703 , n7596 , n9311 );
and ( n11704 , n7730 , n9150 );
nor ( n11705 , n11703 , n11704 );
xnor ( n11706 , n11705 , n9317 );
xor ( n11707 , n11702 , n11706 );
and ( n11708 , n7372 , n9795 );
and ( n11709 , n7494 , n9560 );
nor ( n11710 , n11708 , n11709 );
xnor ( n11711 , n11710 , n9801 );
xor ( n11712 , n11707 , n11711 );
and ( n11713 , n10331 , n7215 );
and ( n11714 , n10548 , n7136 );
nor ( n11715 , n11713 , n11714 );
xnor ( n11716 , n11715 , n7205 );
and ( n11717 , n8548 , n8209 );
and ( n11718 , n8690 , n8039 );
nor ( n11719 , n11717 , n11718 );
xnor ( n11720 , n11719 , n8165 );
xor ( n11721 , n11716 , n11720 );
and ( n11722 , n6960 , n11411 );
and ( n11723 , n6999 , n11159 );
nor ( n11724 , n11722 , n11723 );
xnor ( n11725 , n11724 , n11417 );
xor ( n11726 , n11721 , n11725 );
xor ( n11727 , n11712 , n11726 );
and ( n11728 , n10837 , n7063 );
and ( n11729 , n11133 , n7005 );
nor ( n11730 , n11728 , n11729 );
xnor ( n11731 , n11730 , n7058 );
and ( n11732 , n9839 , n7400 );
and ( n11733 , n10090 , n7303 );
nor ( n11734 , n11732 , n11733 );
xnor ( n11735 , n11734 , n7381 );
xor ( n11736 , n11731 , n11735 );
buf ( n11737 , n803 );
buf ( n11738 , n11737 );
xor ( n11739 , n11738 , n11408 );
and ( n11740 , n6932 , n11739 );
xor ( n11741 , n11736 , n11740 );
xor ( n11742 , n11727 , n11741 );
xor ( n11743 , n11696 , n11742 );
xor ( n11744 , n11687 , n11743 );
and ( n11745 , n11381 , n11435 );
and ( n11746 , n11435 , n11473 );
and ( n11747 , n11381 , n11473 );
or ( n11748 , n11745 , n11746 , n11747 );
and ( n11749 , n11497 , n11501 );
and ( n11750 , n11501 , n11506 );
and ( n11751 , n11497 , n11506 );
or ( n11752 , n11749 , n11750 , n11751 );
and ( n11753 , n11462 , n11466 );
and ( n11754 , n11466 , n11471 );
and ( n11755 , n11462 , n11471 );
or ( n11756 , n11753 , n11754 , n11755 );
xor ( n11757 , n11752 , n11756 );
and ( n11758 , n8913 , n7873 );
and ( n11759 , n9139 , n7762 );
nor ( n11760 , n11758 , n11759 );
xnor ( n11761 , n11760 , n7863 );
and ( n11762 , n7196 , n10342 );
and ( n11763 , n7292 , n10084 );
nor ( n11764 , n11762 , n11763 );
xnor ( n11765 , n11764 , n10291 );
xor ( n11766 , n11761 , n11765 );
and ( n11767 , n7049 , n10907 );
and ( n11768 , n7125 , n10543 );
nor ( n11769 , n11767 , n11768 );
xnor ( n11770 , n11769 , n10807 );
xor ( n11771 , n11766 , n11770 );
xor ( n11772 , n11757 , n11771 );
xor ( n11773 , n11748 , n11772 );
and ( n11774 , n11397 , n11419 );
and ( n11775 , n11419 , n11434 );
and ( n11776 , n11397 , n11434 );
or ( n11777 , n11774 , n11775 , n11776 );
and ( n11778 , n11424 , n11428 );
and ( n11779 , n11428 , n11433 );
and ( n11780 , n11424 , n11433 );
or ( n11781 , n11778 , n11779 , n11780 );
and ( n11782 , n11444 , n11448 );
and ( n11783 , n11448 , n11453 );
and ( n11784 , n11444 , n11453 );
or ( n11785 , n11782 , n11783 , n11784 );
xor ( n11786 , n11781 , n11785 );
and ( n11787 , n11459 , n11461 );
xor ( n11788 , n11786 , n11787 );
xor ( n11789 , n11777 , n11788 );
and ( n11790 , n11387 , n11391 );
and ( n11791 , n11391 , n11396 );
and ( n11792 , n11387 , n11396 );
or ( n11793 , n11790 , n11791 , n11792 );
and ( n11794 , n11401 , n11405 );
and ( n11795 , n11405 , n11418 );
and ( n11796 , n11401 , n11418 );
or ( n11797 , n11794 , n11795 , n11796 );
xor ( n11798 , n11793 , n11797 );
and ( n11799 , n9323 , n7609 );
and ( n11800 , n9549 , n7505 );
nor ( n11801 , n11799 , n11800 );
xnor ( n11802 , n11801 , n7615 );
and ( n11803 , n8156 , n8511 );
and ( n11804 , n8339 , n8350 );
nor ( n11805 , n11803 , n11804 );
xnor ( n11806 , n11805 , n8517 );
xor ( n11807 , n11802 , n11806 );
and ( n11808 , n7891 , n8887 );
and ( n11809 , n8045 , n8701 );
nor ( n11810 , n11808 , n11809 );
xnor ( n11811 , n11810 , n8893 );
xor ( n11812 , n11807 , n11811 );
xor ( n11813 , n11798 , n11812 );
xor ( n11814 , n11789 , n11813 );
xor ( n11815 , n11773 , n11814 );
xor ( n11816 , n11744 , n11815 );
xor ( n11817 , n11683 , n11816 );
and ( n11818 , n11370 , n11372 );
and ( n11819 , n11372 , n11510 );
and ( n11820 , n11370 , n11510 );
or ( n11821 , n11818 , n11819 , n11820 );
xor ( n11822 , n11817 , n11821 );
and ( n11823 , n11366 , n11511 );
and ( n11824 , n11512 , n11515 );
or ( n11825 , n11823 , n11824 );
xor ( n11826 , n11822 , n11825 );
buf ( n11827 , n11826 );
and ( n11828 , n11532 , n11629 );
and ( n11829 , n11629 , n11664 );
and ( n11830 , n11532 , n11664 );
or ( n11831 , n11828 , n11829 , n11830 );
buf ( n11832 , n835 );
buf ( n11833 , n11832 );
xor ( n11834 , n11831 , n11833 );
and ( n11835 , n11634 , n11638 );
and ( n11836 , n11638 , n11663 );
and ( n11837 , n11634 , n11663 );
or ( n11838 , n11835 , n11836 , n11837 );
and ( n11839 , n11595 , n11609 );
and ( n11840 , n11609 , n11627 );
and ( n11841 , n11595 , n11627 );
or ( n11842 , n11839 , n11840 , n11841 );
and ( n11843 , n11643 , n11647 );
and ( n11844 , n11647 , n11662 );
and ( n11845 , n11643 , n11662 );
or ( n11846 , n11843 , n11844 , n11845 );
xor ( n11847 , n11842 , n11846 );
and ( n11848 , n11539 , n6977 );
buf ( n11849 , n771 );
buf ( n11850 , n11849 );
and ( n11851 , n11850 , n6943 );
nor ( n11852 , n11848 , n11851 );
xnor ( n11853 , n11852 , n6974 );
and ( n11854 , n7661 , n9426 );
and ( n11855 , n7791 , n9251 );
nor ( n11856 , n11854 , n11855 );
xnor ( n11857 , n11856 , n9432 );
xor ( n11858 , n11853 , n11857 );
and ( n11859 , n7427 , n9920 );
and ( n11860 , n7545 , n9671 );
nor ( n11861 , n11859 , n11860 );
xnor ( n11862 , n11861 , n9926 );
xor ( n11863 , n11858 , n11862 );
and ( n11864 , n10466 , n7260 );
and ( n11865 , n10679 , n7167 );
nor ( n11866 , n11864 , n11865 );
xnor ( n11867 , n11866 , n7250 );
and ( n11868 , n8643 , n8294 );
and ( n11869 , n8781 , n8110 );
nor ( n11870 , n11868 , n11869 );
xnor ( n11871 , n11870 , n8250 );
xor ( n11872 , n11867 , n11871 );
and ( n11873 , n6980 , n11566 );
and ( n11874 , n7020 , n11300 );
nor ( n11875 , n11873 , n11874 );
xnor ( n11876 , n11875 , n11572 );
xor ( n11877 , n11872 , n11876 );
xor ( n11878 , n11863 , n11877 );
and ( n11879 , n10982 , n7098 );
and ( n11880 , n11274 , n7026 );
nor ( n11881 , n11879 , n11880 );
xnor ( n11882 , n11881 , n7093 );
and ( n11883 , n9964 , n7455 );
and ( n11884 , n10211 , n7344 );
nor ( n11885 , n11883 , n11884 );
xnor ( n11886 , n11885 , n7436 );
xor ( n11887 , n11882 , n11886 );
buf ( n11888 , n803 );
buf ( n11889 , n11888 );
xor ( n11890 , n11889 , n11563 );
and ( n11891 , n6941 , n11890 );
xor ( n11892 , n11887 , n11891 );
xor ( n11893 , n11878 , n11892 );
xor ( n11894 , n11847 , n11893 );
xor ( n11895 , n11838 , n11894 );
and ( n11896 , n11536 , n11590 );
and ( n11897 , n11590 , n11628 );
and ( n11898 , n11536 , n11628 );
or ( n11899 , n11896 , n11897 , n11898 );
and ( n11900 , n11652 , n11656 );
and ( n11901 , n11656 , n11661 );
and ( n11902 , n11652 , n11661 );
or ( n11903 , n11900 , n11901 , n11902 );
and ( n11904 , n11617 , n11621 );
and ( n11905 , n11621 , n11626 );
and ( n11906 , n11617 , n11626 );
or ( n11907 , n11904 , n11905 , n11906 );
xor ( n11908 , n11903 , n11907 );
and ( n11909 , n9018 , n7948 );
and ( n11910 , n9240 , n7823 );
nor ( n11911 , n11909 , n11910 );
xnor ( n11912 , n11911 , n7938 );
and ( n11913 , n7241 , n10477 );
and ( n11914 , n7333 , n10205 );
nor ( n11915 , n11913 , n11914 );
xnor ( n11916 , n11915 , n10426 );
xor ( n11917 , n11912 , n11916 );
and ( n11918 , n7084 , n11052 );
and ( n11919 , n7156 , n10674 );
nor ( n11920 , n11918 , n11919 );
xnor ( n11921 , n11920 , n10952 );
xor ( n11922 , n11917 , n11921 );
xor ( n11923 , n11908 , n11922 );
xor ( n11924 , n11899 , n11923 );
and ( n11925 , n11552 , n11574 );
and ( n11926 , n11574 , n11589 );
and ( n11927 , n11552 , n11589 );
or ( n11928 , n11925 , n11926 , n11927 );
and ( n11929 , n11579 , n11583 );
and ( n11930 , n11583 , n11588 );
and ( n11931 , n11579 , n11588 );
or ( n11932 , n11929 , n11930 , n11931 );
and ( n11933 , n11599 , n11603 );
and ( n11934 , n11603 , n11608 );
and ( n11935 , n11599 , n11608 );
or ( n11936 , n11933 , n11934 , n11935 );
xor ( n11937 , n11932 , n11936 );
and ( n11938 , n11614 , n11616 );
xor ( n11939 , n11937 , n11938 );
xor ( n11940 , n11928 , n11939 );
and ( n11941 , n11542 , n11546 );
and ( n11942 , n11546 , n11551 );
and ( n11943 , n11542 , n11551 );
or ( n11944 , n11941 , n11942 , n11943 );
and ( n11945 , n11556 , n11560 );
and ( n11946 , n11560 , n11573 );
and ( n11947 , n11556 , n11573 );
or ( n11948 , n11945 , n11946 , n11947 );
xor ( n11949 , n11944 , n11948 );
and ( n11950 , n9438 , n7674 );
and ( n11951 , n9660 , n7556 );
nor ( n11952 , n11950 , n11951 );
xnor ( n11953 , n11952 , n7680 );
and ( n11954 , n8241 , n8606 );
and ( n11955 , n8420 , n8431 );
nor ( n11956 , n11954 , n11955 );
xnor ( n11957 , n11956 , n8612 );
xor ( n11958 , n11953 , n11957 );
and ( n11959 , n7966 , n8992 );
and ( n11960 , n8116 , n8792 );
nor ( n11961 , n11959 , n11960 );
xnor ( n11962 , n11961 , n8998 );
xor ( n11963 , n11958 , n11962 );
xor ( n11964 , n11949 , n11963 );
xor ( n11965 , n11940 , n11964 );
xor ( n11966 , n11924 , n11965 );
xor ( n11967 , n11895 , n11966 );
xor ( n11968 , n11834 , n11967 );
and ( n11969 , n11525 , n11527 );
and ( n11970 , n11527 , n11665 );
and ( n11971 , n11525 , n11665 );
or ( n11972 , n11969 , n11970 , n11971 );
xor ( n11973 , n11968 , n11972 );
and ( n11974 , n11521 , n11666 );
and ( n11975 , n11667 , n11670 );
or ( n11976 , n11974 , n11975 );
xor ( n11977 , n11973 , n11976 );
buf ( n11978 , n11977 );
not ( n11979 , n831 );
and ( n11980 , n11979 , n11827 );
and ( n11981 , n11978 , n831 );
or ( n11982 , n11980 , n11981 );
and ( n11983 , n11687 , n11743 );
and ( n11984 , n11743 , n11815 );
and ( n11985 , n11687 , n11815 );
or ( n11986 , n11983 , n11984 , n11985 );
buf ( n11987 , n866 );
buf ( n11988 , n11987 );
xor ( n11989 , n11986 , n11988 );
and ( n11990 , n11691 , n11695 );
and ( n11991 , n11695 , n11742 );
and ( n11992 , n11691 , n11742 );
or ( n11993 , n11990 , n11991 , n11992 );
and ( n11994 , n11748 , n11772 );
and ( n11995 , n11772 , n11814 );
and ( n11996 , n11748 , n11814 );
or ( n11997 , n11994 , n11995 , n11996 );
xor ( n11998 , n11993 , n11997 );
and ( n11999 , n11781 , n11785 );
and ( n12000 , n11785 , n11787 );
and ( n12001 , n11781 , n11787 );
or ( n12002 , n11999 , n12000 , n12001 );
and ( n12003 , n11712 , n11726 );
and ( n12004 , n11726 , n11741 );
and ( n12005 , n11712 , n11741 );
or ( n12006 , n12003 , n12004 , n12005 );
xor ( n12007 , n12002 , n12006 );
and ( n12008 , n11699 , n6957 );
buf ( n12009 , n770 );
buf ( n12010 , n12009 );
and ( n12011 , n12010 , n6934 );
nor ( n12012 , n12008 , n12011 );
xnor ( n12013 , n12012 , n6954 );
not ( n12014 , n11740 );
buf ( n12015 , n802 );
buf ( n12016 , n12015 );
and ( n12017 , n11738 , n11408 );
not ( n12018 , n12017 );
and ( n12019 , n12016 , n12018 );
and ( n12020 , n12014 , n12019 );
xor ( n12021 , n12013 , n12020 );
and ( n12022 , n6999 , n11411 );
and ( n12023 , n7049 , n11159 );
nor ( n12024 , n12022 , n12023 );
xnor ( n12025 , n12024 , n11417 );
xor ( n12026 , n12021 , n12025 );
xor ( n12027 , n12016 , n11738 );
not ( n12028 , n11739 );
and ( n12029 , n12027 , n12028 );
and ( n12030 , n6932 , n12029 );
and ( n12031 , n6960 , n11739 );
nor ( n12032 , n12030 , n12031 );
xnor ( n12033 , n12032 , n12019 );
xor ( n12034 , n12026 , n12033 );
xor ( n12035 , n12007 , n12034 );
and ( n12036 , n11793 , n11797 );
and ( n12037 , n11797 , n11812 );
and ( n12038 , n11793 , n11812 );
or ( n12039 , n12036 , n12037 , n12038 );
and ( n12040 , n11702 , n11706 );
and ( n12041 , n11706 , n11711 );
and ( n12042 , n11702 , n11711 );
or ( n12043 , n12040 , n12041 , n12042 );
and ( n12044 , n11731 , n11735 );
and ( n12045 , n11735 , n11740 );
and ( n12046 , n11731 , n11740 );
or ( n12047 , n12044 , n12045 , n12046 );
xor ( n12048 , n12043 , n12047 );
and ( n12049 , n11802 , n11806 );
and ( n12050 , n11806 , n11811 );
and ( n12051 , n11802 , n11811 );
or ( n12052 , n12049 , n12050 , n12051 );
xor ( n12053 , n12048 , n12052 );
xor ( n12054 , n12039 , n12053 );
and ( n12055 , n11716 , n11720 );
and ( n12056 , n11720 , n11725 );
and ( n12057 , n11716 , n11725 );
or ( n12058 , n12055 , n12056 , n12057 );
and ( n12059 , n11761 , n11765 );
and ( n12060 , n11765 , n11770 );
and ( n12061 , n11761 , n11770 );
or ( n12062 , n12059 , n12060 , n12061 );
xor ( n12063 , n12058 , n12062 );
and ( n12064 , n11133 , n7063 );
and ( n12065 , n11384 , n7005 );
nor ( n12066 , n12064 , n12065 );
xnor ( n12067 , n12066 , n7058 );
and ( n12068 , n10090 , n7400 );
and ( n12069 , n10331 , n7303 );
nor ( n12070 , n12068 , n12069 );
xnor ( n12071 , n12070 , n7381 );
xor ( n12072 , n12067 , n12071 );
and ( n12073 , n8339 , n8511 );
and ( n12074 , n8548 , n8350 );
nor ( n12075 , n12073 , n12074 );
xnor ( n12076 , n12075 , n8517 );
xor ( n12077 , n12072 , n12076 );
xor ( n12078 , n12063 , n12077 );
xor ( n12079 , n12054 , n12078 );
xor ( n12080 , n12035 , n12079 );
and ( n12081 , n11752 , n11756 );
and ( n12082 , n11756 , n11771 );
and ( n12083 , n11752 , n11771 );
or ( n12084 , n12081 , n12082 , n12083 );
and ( n12085 , n11777 , n11788 );
and ( n12086 , n11788 , n11813 );
and ( n12087 , n11777 , n11813 );
or ( n12088 , n12085 , n12086 , n12087 );
xor ( n12089 , n12084 , n12088 );
and ( n12090 , n9549 , n7609 );
and ( n12091 , n9839 , n7505 );
nor ( n12092 , n12090 , n12091 );
xnor ( n12093 , n12092 , n7615 );
and ( n12094 , n8045 , n8887 );
and ( n12095 , n8156 , n8701 );
nor ( n12096 , n12094 , n12095 );
xnor ( n12097 , n12096 , n8893 );
xor ( n12098 , n12093 , n12097 );
and ( n12099 , n7730 , n9311 );
and ( n12100 , n7891 , n9150 );
nor ( n12101 , n12099 , n12100 );
xnor ( n12102 , n12101 , n9317 );
xor ( n12103 , n12098 , n12102 );
and ( n12104 , n10548 , n7215 );
and ( n12105 , n10837 , n7136 );
nor ( n12106 , n12104 , n12105 );
xnor ( n12107 , n12106 , n7205 );
and ( n12108 , n9139 , n7873 );
and ( n12109 , n9323 , n7762 );
nor ( n12110 , n12108 , n12109 );
xnor ( n12111 , n12110 , n7863 );
xor ( n12112 , n12107 , n12111 );
and ( n12113 , n7494 , n9795 );
and ( n12114 , n7596 , n9560 );
nor ( n12115 , n12113 , n12114 );
xnor ( n12116 , n12115 , n9801 );
xor ( n12117 , n12112 , n12116 );
xor ( n12118 , n12103 , n12117 );
and ( n12119 , n8690 , n8209 );
and ( n12120 , n8913 , n8039 );
nor ( n12121 , n12119 , n12120 );
xnor ( n12122 , n12121 , n8165 );
and ( n12123 , n7292 , n10342 );
and ( n12124 , n7372 , n10084 );
nor ( n12125 , n12123 , n12124 );
xnor ( n12126 , n12125 , n10291 );
xor ( n12127 , n12122 , n12126 );
and ( n12128 , n7125 , n10907 );
and ( n12129 , n7196 , n10543 );
nor ( n12130 , n12128 , n12129 );
xnor ( n12131 , n12130 , n10807 );
xor ( n12132 , n12127 , n12131 );
xor ( n12133 , n12118 , n12132 );
xor ( n12134 , n12089 , n12133 );
xor ( n12135 , n12080 , n12134 );
xor ( n12136 , n11998 , n12135 );
xor ( n12137 , n11989 , n12136 );
and ( n12138 , n11680 , n11682 );
and ( n12139 , n11682 , n11816 );
and ( n12140 , n11680 , n11816 );
or ( n12141 , n12138 , n12139 , n12140 );
xor ( n12142 , n12137 , n12141 );
and ( n12143 , n11817 , n11821 );
and ( n12144 , n11822 , n11825 );
or ( n12145 , n12143 , n12144 );
xor ( n12146 , n12142 , n12145 );
buf ( n12147 , n12146 );
and ( n12148 , n11838 , n11894 );
and ( n12149 , n11894 , n11966 );
and ( n12150 , n11838 , n11966 );
or ( n12151 , n12148 , n12149 , n12150 );
buf ( n12152 , n834 );
buf ( n12153 , n12152 );
xor ( n12154 , n12151 , n12153 );
and ( n12155 , n11842 , n11846 );
and ( n12156 , n11846 , n11893 );
and ( n12157 , n11842 , n11893 );
or ( n12158 , n12155 , n12156 , n12157 );
and ( n12159 , n11899 , n11923 );
and ( n12160 , n11923 , n11965 );
and ( n12161 , n11899 , n11965 );
or ( n12162 , n12159 , n12160 , n12161 );
xor ( n12163 , n12158 , n12162 );
and ( n12164 , n11932 , n11936 );
and ( n12165 , n11936 , n11938 );
and ( n12166 , n11932 , n11938 );
or ( n12167 , n12164 , n12165 , n12166 );
and ( n12168 , n11863 , n11877 );
and ( n12169 , n11877 , n11892 );
and ( n12170 , n11863 , n11892 );
or ( n12171 , n12168 , n12169 , n12170 );
xor ( n12172 , n12167 , n12171 );
and ( n12173 , n11850 , n6977 );
buf ( n12174 , n770 );
buf ( n12175 , n12174 );
and ( n12176 , n12175 , n6943 );
nor ( n12177 , n12173 , n12176 );
xnor ( n12178 , n12177 , n6974 );
not ( n12179 , n11891 );
buf ( n12180 , n802 );
buf ( n12181 , n12180 );
and ( n12182 , n11889 , n11563 );
not ( n12183 , n12182 );
and ( n12184 , n12181 , n12183 );
and ( n12185 , n12179 , n12184 );
xor ( n12186 , n12178 , n12185 );
and ( n12187 , n7020 , n11566 );
and ( n12188 , n7084 , n11300 );
nor ( n12189 , n12187 , n12188 );
xnor ( n12190 , n12189 , n11572 );
xor ( n12191 , n12186 , n12190 );
xor ( n12192 , n12181 , n11889 );
not ( n12193 , n11890 );
and ( n12194 , n12192 , n12193 );
and ( n12195 , n6941 , n12194 );
and ( n12196 , n6980 , n11890 );
nor ( n12197 , n12195 , n12196 );
xnor ( n12198 , n12197 , n12184 );
xor ( n12199 , n12191 , n12198 );
xor ( n12200 , n12172 , n12199 );
and ( n12201 , n11944 , n11948 );
and ( n12202 , n11948 , n11963 );
and ( n12203 , n11944 , n11963 );
or ( n12204 , n12201 , n12202 , n12203 );
and ( n12205 , n11853 , n11857 );
and ( n12206 , n11857 , n11862 );
and ( n12207 , n11853 , n11862 );
or ( n12208 , n12205 , n12206 , n12207 );
and ( n12209 , n11882 , n11886 );
and ( n12210 , n11886 , n11891 );
and ( n12211 , n11882 , n11891 );
or ( n12212 , n12209 , n12210 , n12211 );
xor ( n12213 , n12208 , n12212 );
and ( n12214 , n11953 , n11957 );
and ( n12215 , n11957 , n11962 );
and ( n12216 , n11953 , n11962 );
or ( n12217 , n12214 , n12215 , n12216 );
xor ( n12218 , n12213 , n12217 );
xor ( n12219 , n12204 , n12218 );
and ( n12220 , n11867 , n11871 );
and ( n12221 , n11871 , n11876 );
and ( n12222 , n11867 , n11876 );
or ( n12223 , n12220 , n12221 , n12222 );
and ( n12224 , n11912 , n11916 );
and ( n12225 , n11916 , n11921 );
and ( n12226 , n11912 , n11921 );
or ( n12227 , n12224 , n12225 , n12226 );
xor ( n12228 , n12223 , n12227 );
and ( n12229 , n11274 , n7098 );
and ( n12230 , n11539 , n7026 );
nor ( n12231 , n12229 , n12230 );
xnor ( n12232 , n12231 , n7093 );
and ( n12233 , n10211 , n7455 );
and ( n12234 , n10466 , n7344 );
nor ( n12235 , n12233 , n12234 );
xnor ( n12236 , n12235 , n7436 );
xor ( n12237 , n12232 , n12236 );
and ( n12238 , n8420 , n8606 );
and ( n12239 , n8643 , n8431 );
nor ( n12240 , n12238 , n12239 );
xnor ( n12241 , n12240 , n8612 );
xor ( n12242 , n12237 , n12241 );
xor ( n12243 , n12228 , n12242 );
xor ( n12244 , n12219 , n12243 );
xor ( n12245 , n12200 , n12244 );
and ( n12246 , n11903 , n11907 );
and ( n12247 , n11907 , n11922 );
and ( n12248 , n11903 , n11922 );
or ( n12249 , n12246 , n12247 , n12248 );
and ( n12250 , n11928 , n11939 );
and ( n12251 , n11939 , n11964 );
and ( n12252 , n11928 , n11964 );
or ( n12253 , n12250 , n12251 , n12252 );
xor ( n12254 , n12249 , n12253 );
and ( n12255 , n9660 , n7674 );
and ( n12256 , n9964 , n7556 );
nor ( n12257 , n12255 , n12256 );
xnor ( n12258 , n12257 , n7680 );
and ( n12259 , n8116 , n8992 );
and ( n12260 , n8241 , n8792 );
nor ( n12261 , n12259 , n12260 );
xnor ( n12262 , n12261 , n8998 );
xor ( n12263 , n12258 , n12262 );
and ( n12264 , n7791 , n9426 );
and ( n12265 , n7966 , n9251 );
nor ( n12266 , n12264 , n12265 );
xnor ( n12267 , n12266 , n9432 );
xor ( n12268 , n12263 , n12267 );
and ( n12269 , n10679 , n7260 );
and ( n12270 , n10982 , n7167 );
nor ( n12271 , n12269 , n12270 );
xnor ( n12272 , n12271 , n7250 );
and ( n12273 , n9240 , n7948 );
and ( n12274 , n9438 , n7823 );
nor ( n12275 , n12273 , n12274 );
xnor ( n12276 , n12275 , n7938 );
xor ( n12277 , n12272 , n12276 );
and ( n12278 , n7545 , n9920 );
and ( n12279 , n7661 , n9671 );
nor ( n12280 , n12278 , n12279 );
xnor ( n12281 , n12280 , n9926 );
xor ( n12282 , n12277 , n12281 );
xor ( n12283 , n12268 , n12282 );
and ( n12284 , n8781 , n8294 );
and ( n12285 , n9018 , n8110 );
nor ( n12286 , n12284 , n12285 );
xnor ( n12287 , n12286 , n8250 );
and ( n12288 , n7333 , n10477 );
and ( n12289 , n7427 , n10205 );
nor ( n12290 , n12288 , n12289 );
xnor ( n12291 , n12290 , n10426 );
xor ( n12292 , n12287 , n12291 );
and ( n12293 , n7156 , n11052 );
and ( n12294 , n7241 , n10674 );
nor ( n12295 , n12293 , n12294 );
xnor ( n12296 , n12295 , n10952 );
xor ( n12297 , n12292 , n12296 );
xor ( n12298 , n12283 , n12297 );
xor ( n12299 , n12254 , n12298 );
xor ( n12300 , n12245 , n12299 );
xor ( n12301 , n12163 , n12300 );
xor ( n12302 , n12154 , n12301 );
and ( n12303 , n11831 , n11833 );
and ( n12304 , n11833 , n11967 );
and ( n12305 , n11831 , n11967 );
or ( n12306 , n12303 , n12304 , n12305 );
xor ( n12307 , n12302 , n12306 );
and ( n12308 , n11968 , n11972 );
and ( n12309 , n11973 , n11976 );
or ( n12310 , n12308 , n12309 );
xor ( n12311 , n12307 , n12310 );
buf ( n12312 , n12311 );
not ( n12313 , n831 );
and ( n12314 , n12313 , n12147 );
and ( n12315 , n12312 , n831 );
or ( n12316 , n12314 , n12315 );
and ( n12317 , n11993 , n11997 );
and ( n12318 , n11997 , n12135 );
and ( n12319 , n11993 , n12135 );
or ( n12320 , n12317 , n12318 , n12319 );
buf ( n12321 , n865 );
buf ( n12322 , n12321 );
xor ( n12323 , n12320 , n12322 );
and ( n12324 , n12035 , n12079 );
and ( n12325 , n12079 , n12134 );
and ( n12326 , n12035 , n12134 );
or ( n12327 , n12324 , n12325 , n12326 );
and ( n12328 , n12002 , n12006 );
and ( n12329 , n12006 , n12034 );
and ( n12330 , n12002 , n12034 );
or ( n12331 , n12328 , n12329 , n12330 );
and ( n12332 , n12039 , n12053 );
and ( n12333 , n12053 , n12078 );
and ( n12334 , n12039 , n12078 );
or ( n12335 , n12332 , n12333 , n12334 );
xor ( n12336 , n12331 , n12335 );
and ( n12337 , n12010 , n6957 );
buf ( n12338 , n769 );
buf ( n12339 , n12338 );
and ( n12340 , n12339 , n6934 );
nor ( n12341 , n12337 , n12340 );
xnor ( n12342 , n12341 , n6954 );
and ( n12343 , n11384 , n7063 );
and ( n12344 , n11699 , n7005 );
nor ( n12345 , n12343 , n12344 );
xnor ( n12346 , n12345 , n7058 );
xor ( n12347 , n12342 , n12346 );
buf ( n12348 , n801 );
buf ( n12349 , n12348 );
xor ( n12350 , n12349 , n12016 );
and ( n12351 , n6932 , n12350 );
xor ( n12352 , n12347 , n12351 );
and ( n12353 , n10837 , n7215 );
and ( n12354 , n11133 , n7136 );
nor ( n12355 , n12353 , n12354 );
xnor ( n12356 , n12355 , n7205 );
and ( n12357 , n9323 , n7873 );
and ( n12358 , n9549 , n7762 );
nor ( n12359 , n12357 , n12358 );
xnor ( n12360 , n12359 , n7863 );
xor ( n12361 , n12356 , n12360 );
and ( n12362 , n7372 , n10342 );
and ( n12363 , n7494 , n10084 );
nor ( n12364 , n12362 , n12363 );
xnor ( n12365 , n12364 , n10291 );
xor ( n12366 , n12361 , n12365 );
xor ( n12367 , n12352 , n12366 );
and ( n12368 , n8913 , n8209 );
and ( n12369 , n9139 , n8039 );
nor ( n12370 , n12368 , n12369 );
xnor ( n12371 , n12370 , n8165 );
and ( n12372 , n7196 , n10907 );
and ( n12373 , n7292 , n10543 );
nor ( n12374 , n12372 , n12373 );
xnor ( n12375 , n12374 , n10807 );
xor ( n12376 , n12371 , n12375 );
and ( n12377 , n7049 , n11411 );
and ( n12378 , n7125 , n11159 );
nor ( n12379 , n12377 , n12378 );
xnor ( n12380 , n12379 , n11417 );
xor ( n12381 , n12376 , n12380 );
xor ( n12382 , n12367 , n12381 );
xor ( n12383 , n12336 , n12382 );
xor ( n12384 , n12327 , n12383 );
and ( n12385 , n12084 , n12088 );
and ( n12386 , n12088 , n12133 );
and ( n12387 , n12084 , n12133 );
or ( n12388 , n12385 , n12386 , n12387 );
and ( n12389 , n12043 , n12047 );
and ( n12390 , n12047 , n12052 );
and ( n12391 , n12043 , n12052 );
or ( n12392 , n12389 , n12390 , n12391 );
and ( n12393 , n12103 , n12117 );
and ( n12394 , n12117 , n12132 );
and ( n12395 , n12103 , n12132 );
or ( n12396 , n12393 , n12394 , n12395 );
xor ( n12397 , n12392 , n12396 );
and ( n12398 , n12067 , n12071 );
and ( n12399 , n12071 , n12076 );
and ( n12400 , n12067 , n12076 );
or ( n12401 , n12398 , n12399 , n12400 );
and ( n12402 , n12013 , n12020 );
xor ( n12403 , n12401 , n12402 );
and ( n12404 , n6960 , n12029 );
and ( n12405 , n6999 , n11739 );
nor ( n12406 , n12404 , n12405 );
xnor ( n12407 , n12406 , n12019 );
xor ( n12408 , n12403 , n12407 );
xor ( n12409 , n12397 , n12408 );
xor ( n12410 , n12388 , n12409 );
and ( n12411 , n12058 , n12062 );
and ( n12412 , n12062 , n12077 );
and ( n12413 , n12058 , n12077 );
or ( n12414 , n12411 , n12412 , n12413 );
and ( n12415 , n12093 , n12097 );
and ( n12416 , n12097 , n12102 );
and ( n12417 , n12093 , n12102 );
or ( n12418 , n12415 , n12416 , n12417 );
and ( n12419 , n12107 , n12111 );
and ( n12420 , n12111 , n12116 );
and ( n12421 , n12107 , n12116 );
or ( n12422 , n12419 , n12420 , n12421 );
xor ( n12423 , n12418 , n12422 );
and ( n12424 , n12122 , n12126 );
and ( n12425 , n12126 , n12131 );
and ( n12426 , n12122 , n12131 );
or ( n12427 , n12424 , n12425 , n12426 );
xor ( n12428 , n12423 , n12427 );
xor ( n12429 , n12414 , n12428 );
and ( n12430 , n12021 , n12025 );
and ( n12431 , n12025 , n12033 );
and ( n12432 , n12021 , n12033 );
or ( n12433 , n12430 , n12431 , n12432 );
and ( n12434 , n9839 , n7609 );
and ( n12435 , n10090 , n7505 );
nor ( n12436 , n12434 , n12435 );
xnor ( n12437 , n12436 , n7615 );
and ( n12438 , n7891 , n9311 );
and ( n12439 , n8045 , n9150 );
nor ( n12440 , n12438 , n12439 );
xnor ( n12441 , n12440 , n9317 );
xor ( n12442 , n12437 , n12441 );
and ( n12443 , n7596 , n9795 );
and ( n12444 , n7730 , n9560 );
nor ( n12445 , n12443 , n12444 );
xnor ( n12446 , n12445 , n9801 );
xor ( n12447 , n12442 , n12446 );
xor ( n12448 , n12433 , n12447 );
and ( n12449 , n10331 , n7400 );
and ( n12450 , n10548 , n7303 );
nor ( n12451 , n12449 , n12450 );
xnor ( n12452 , n12451 , n7381 );
and ( n12453 , n8548 , n8511 );
and ( n12454 , n8690 , n8350 );
nor ( n12455 , n12453 , n12454 );
xnor ( n12456 , n12455 , n8517 );
xor ( n12457 , n12452 , n12456 );
and ( n12458 , n8156 , n8887 );
and ( n12459 , n8339 , n8701 );
nor ( n12460 , n12458 , n12459 );
xnor ( n12461 , n12460 , n8893 );
xor ( n12462 , n12457 , n12461 );
xor ( n12463 , n12448 , n12462 );
xor ( n12464 , n12429 , n12463 );
xor ( n12465 , n12410 , n12464 );
xor ( n12466 , n12384 , n12465 );
xor ( n12467 , n12323 , n12466 );
and ( n12468 , n11986 , n11988 );
and ( n12469 , n11988 , n12136 );
and ( n12470 , n11986 , n12136 );
or ( n12471 , n12468 , n12469 , n12470 );
xor ( n12472 , n12467 , n12471 );
and ( n12473 , n12137 , n12141 );
and ( n12474 , n12142 , n12145 );
or ( n12475 , n12473 , n12474 );
xor ( n12476 , n12472 , n12475 );
buf ( n12477 , n12476 );
and ( n12478 , n12158 , n12162 );
and ( n12479 , n12162 , n12300 );
and ( n12480 , n12158 , n12300 );
or ( n12481 , n12478 , n12479 , n12480 );
buf ( n12482 , n833 );
buf ( n12483 , n12482 );
xor ( n12484 , n12481 , n12483 );
and ( n12485 , n12200 , n12244 );
and ( n12486 , n12244 , n12299 );
and ( n12487 , n12200 , n12299 );
or ( n12488 , n12485 , n12486 , n12487 );
and ( n12489 , n12167 , n12171 );
and ( n12490 , n12171 , n12199 );
and ( n12491 , n12167 , n12199 );
or ( n12492 , n12489 , n12490 , n12491 );
and ( n12493 , n12204 , n12218 );
and ( n12494 , n12218 , n12243 );
and ( n12495 , n12204 , n12243 );
or ( n12496 , n12493 , n12494 , n12495 );
xor ( n12497 , n12492 , n12496 );
and ( n12498 , n12175 , n6977 );
buf ( n12499 , n769 );
buf ( n12500 , n12499 );
and ( n12501 , n12500 , n6943 );
nor ( n12502 , n12498 , n12501 );
xnor ( n12503 , n12502 , n6974 );
and ( n12504 , n11539 , n7098 );
and ( n12505 , n11850 , n7026 );
nor ( n12506 , n12504 , n12505 );
xnor ( n12507 , n12506 , n7093 );
xor ( n12508 , n12503 , n12507 );
buf ( n12509 , n801 );
buf ( n12510 , n12509 );
xor ( n12511 , n12510 , n12181 );
and ( n12512 , n6941 , n12511 );
xor ( n12513 , n12508 , n12512 );
and ( n12514 , n10982 , n7260 );
and ( n12515 , n11274 , n7167 );
nor ( n12516 , n12514 , n12515 );
xnor ( n12517 , n12516 , n7250 );
and ( n12518 , n9438 , n7948 );
and ( n12519 , n9660 , n7823 );
nor ( n12520 , n12518 , n12519 );
xnor ( n12521 , n12520 , n7938 );
xor ( n12522 , n12517 , n12521 );
and ( n12523 , n7427 , n10477 );
and ( n12524 , n7545 , n10205 );
nor ( n12525 , n12523 , n12524 );
xnor ( n12526 , n12525 , n10426 );
xor ( n12527 , n12522 , n12526 );
xor ( n12528 , n12513 , n12527 );
and ( n12529 , n9018 , n8294 );
and ( n12530 , n9240 , n8110 );
nor ( n12531 , n12529 , n12530 );
xnor ( n12532 , n12531 , n8250 );
and ( n12533 , n7241 , n11052 );
and ( n12534 , n7333 , n10674 );
nor ( n12535 , n12533 , n12534 );
xnor ( n12536 , n12535 , n10952 );
xor ( n12537 , n12532 , n12536 );
and ( n12538 , n7084 , n11566 );
and ( n12539 , n7156 , n11300 );
nor ( n12540 , n12538 , n12539 );
xnor ( n12541 , n12540 , n11572 );
xor ( n12542 , n12537 , n12541 );
xor ( n12543 , n12528 , n12542 );
xor ( n12544 , n12497 , n12543 );
xor ( n12545 , n12488 , n12544 );
and ( n12546 , n12249 , n12253 );
and ( n12547 , n12253 , n12298 );
and ( n12548 , n12249 , n12298 );
or ( n12549 , n12546 , n12547 , n12548 );
and ( n12550 , n12208 , n12212 );
and ( n12551 , n12212 , n12217 );
and ( n12552 , n12208 , n12217 );
or ( n12553 , n12550 , n12551 , n12552 );
and ( n12554 , n12268 , n12282 );
and ( n12555 , n12282 , n12297 );
and ( n12556 , n12268 , n12297 );
or ( n12557 , n12554 , n12555 , n12556 );
xor ( n12558 , n12553 , n12557 );
and ( n12559 , n12232 , n12236 );
and ( n12560 , n12236 , n12241 );
and ( n12561 , n12232 , n12241 );
or ( n12562 , n12559 , n12560 , n12561 );
and ( n12563 , n12178 , n12185 );
xor ( n12564 , n12562 , n12563 );
and ( n12565 , n6980 , n12194 );
and ( n12566 , n7020 , n11890 );
nor ( n12567 , n12565 , n12566 );
xnor ( n12568 , n12567 , n12184 );
xor ( n12569 , n12564 , n12568 );
xor ( n12570 , n12558 , n12569 );
xor ( n12571 , n12549 , n12570 );
and ( n12572 , n12223 , n12227 );
and ( n12573 , n12227 , n12242 );
and ( n12574 , n12223 , n12242 );
or ( n12575 , n12572 , n12573 , n12574 );
and ( n12576 , n12258 , n12262 );
and ( n12577 , n12262 , n12267 );
and ( n12578 , n12258 , n12267 );
or ( n12579 , n12576 , n12577 , n12578 );
and ( n12580 , n12272 , n12276 );
and ( n12581 , n12276 , n12281 );
and ( n12582 , n12272 , n12281 );
or ( n12583 , n12580 , n12581 , n12582 );
xor ( n12584 , n12579 , n12583 );
and ( n12585 , n12287 , n12291 );
and ( n12586 , n12291 , n12296 );
and ( n12587 , n12287 , n12296 );
or ( n12588 , n12585 , n12586 , n12587 );
xor ( n12589 , n12584 , n12588 );
xor ( n12590 , n12575 , n12589 );
and ( n12591 , n12186 , n12190 );
and ( n12592 , n12190 , n12198 );
and ( n12593 , n12186 , n12198 );
or ( n12594 , n12591 , n12592 , n12593 );
and ( n12595 , n9964 , n7674 );
and ( n12596 , n10211 , n7556 );
nor ( n12597 , n12595 , n12596 );
xnor ( n12598 , n12597 , n7680 );
and ( n12599 , n7966 , n9426 );
and ( n12600 , n8116 , n9251 );
nor ( n12601 , n12599 , n12600 );
xnor ( n12602 , n12601 , n9432 );
xor ( n12603 , n12598 , n12602 );
and ( n12604 , n7661 , n9920 );
and ( n12605 , n7791 , n9671 );
nor ( n12606 , n12604 , n12605 );
xnor ( n12607 , n12606 , n9926 );
xor ( n12608 , n12603 , n12607 );
xor ( n12609 , n12594 , n12608 );
and ( n12610 , n10466 , n7455 );
and ( n12611 , n10679 , n7344 );
nor ( n12612 , n12610 , n12611 );
xnor ( n12613 , n12612 , n7436 );
and ( n12614 , n8643 , n8606 );
and ( n12615 , n8781 , n8431 );
nor ( n12616 , n12614 , n12615 );
xnor ( n12617 , n12616 , n8612 );
xor ( n12618 , n12613 , n12617 );
and ( n12619 , n8241 , n8992 );
and ( n12620 , n8420 , n8792 );
nor ( n12621 , n12619 , n12620 );
xnor ( n12622 , n12621 , n8998 );
xor ( n12623 , n12618 , n12622 );
xor ( n12624 , n12609 , n12623 );
xor ( n12625 , n12590 , n12624 );
xor ( n12626 , n12571 , n12625 );
xor ( n12627 , n12545 , n12626 );
xor ( n12628 , n12484 , n12627 );
and ( n12629 , n12151 , n12153 );
and ( n12630 , n12153 , n12301 );
and ( n12631 , n12151 , n12301 );
or ( n12632 , n12629 , n12630 , n12631 );
xor ( n12633 , n12628 , n12632 );
and ( n12634 , n12302 , n12306 );
and ( n12635 , n12307 , n12310 );
or ( n12636 , n12634 , n12635 );
xor ( n12637 , n12633 , n12636 );
buf ( n12638 , n12637 );
not ( n12639 , n831 );
and ( n12640 , n12639 , n12477 );
and ( n12641 , n12638 , n831 );
or ( n12642 , n12640 , n12641 );
and ( n12643 , n12327 , n12383 );
and ( n12644 , n12383 , n12465 );
and ( n12645 , n12327 , n12465 );
or ( n12646 , n12643 , n12644 , n12645 );
buf ( n12647 , n864 );
buf ( n12648 , n12647 );
xor ( n12649 , n12646 , n12648 );
and ( n12650 , n12388 , n12409 );
and ( n12651 , n12409 , n12464 );
and ( n12652 , n12388 , n12464 );
or ( n12653 , n12650 , n12651 , n12652 );
and ( n12654 , n12392 , n12396 );
and ( n12655 , n12396 , n12408 );
and ( n12656 , n12392 , n12408 );
or ( n12657 , n12654 , n12655 , n12656 );
and ( n12658 , n12414 , n12428 );
and ( n12659 , n12428 , n12463 );
and ( n12660 , n12414 , n12463 );
or ( n12661 , n12658 , n12659 , n12660 );
xor ( n12662 , n12657 , n12661 );
and ( n12663 , n12418 , n12422 );
and ( n12664 , n12422 , n12427 );
and ( n12665 , n12418 , n12427 );
or ( n12666 , n12663 , n12664 , n12665 );
and ( n12667 , n9549 , n7873 );
and ( n12668 , n9839 , n7762 );
nor ( n12669 , n12667 , n12668 );
xnor ( n12670 , n12669 , n7863 );
and ( n12671 , n7494 , n10342 );
and ( n12672 , n7596 , n10084 );
nor ( n12673 , n12671 , n12672 );
xnor ( n12674 , n12673 , n10291 );
xor ( n12675 , n12670 , n12674 );
and ( n12676 , n7292 , n10907 );
and ( n12677 , n7372 , n10543 );
nor ( n12678 , n12676 , n12677 );
xnor ( n12679 , n12678 , n10807 );
xor ( n12680 , n12675 , n12679 );
xor ( n12681 , n12666 , n12680 );
and ( n12682 , n11133 , n7215 );
and ( n12683 , n11384 , n7136 );
nor ( n12684 , n12682 , n12683 );
xnor ( n12685 , n12684 , n7205 );
and ( n12686 , n8045 , n9311 );
and ( n12687 , n8156 , n9150 );
nor ( n12688 , n12686 , n12687 );
xnor ( n12689 , n12688 , n9317 );
xor ( n12690 , n12685 , n12689 );
and ( n12691 , n7730 , n9795 );
and ( n12692 , n7891 , n9560 );
nor ( n12693 , n12691 , n12692 );
xnor ( n12694 , n12693 , n9801 );
xor ( n12695 , n12690 , n12694 );
xor ( n12696 , n12681 , n12695 );
xor ( n12697 , n12662 , n12696 );
xor ( n12698 , n12653 , n12697 );
and ( n12699 , n12331 , n12335 );
and ( n12700 , n12335 , n12382 );
and ( n12701 , n12331 , n12382 );
or ( n12702 , n12699 , n12700 , n12701 );
and ( n12703 , n12401 , n12402 );
and ( n12704 , n12402 , n12407 );
and ( n12705 , n12401 , n12407 );
or ( n12706 , n12703 , n12704 , n12705 );
and ( n12707 , n12356 , n12360 );
and ( n12708 , n12360 , n12365 );
and ( n12709 , n12356 , n12365 );
or ( n12710 , n12707 , n12708 , n12709 );
and ( n12711 , n12371 , n12375 );
and ( n12712 , n12375 , n12380 );
and ( n12713 , n12371 , n12380 );
or ( n12714 , n12711 , n12712 , n12713 );
xor ( n12715 , n12710 , n12714 );
and ( n12716 , n12437 , n12441 );
and ( n12717 , n12441 , n12446 );
and ( n12718 , n12437 , n12446 );
or ( n12719 , n12716 , n12717 , n12718 );
xor ( n12720 , n12715 , n12719 );
xor ( n12721 , n12706 , n12720 );
and ( n12722 , n12339 , n6957 );
buf ( n12723 , n768 );
buf ( n12724 , n12723 );
and ( n12725 , n12724 , n6934 );
nor ( n12726 , n12722 , n12725 );
xnor ( n12727 , n12726 , n6954 );
not ( n12728 , n12351 );
buf ( n12729 , n800 );
buf ( n12730 , n12729 );
and ( n12731 , n12349 , n12016 );
not ( n12732 , n12731 );
and ( n12733 , n12730 , n12732 );
and ( n12734 , n12728 , n12733 );
xor ( n12735 , n12727 , n12734 );
and ( n12736 , n12342 , n12346 );
and ( n12737 , n12346 , n12351 );
and ( n12738 , n12342 , n12351 );
or ( n12739 , n12736 , n12737 , n12738 );
xor ( n12740 , n12735 , n12739 );
and ( n12741 , n12452 , n12456 );
and ( n12742 , n12456 , n12461 );
and ( n12743 , n12452 , n12461 );
or ( n12744 , n12741 , n12742 , n12743 );
xor ( n12745 , n12740 , n12744 );
xor ( n12746 , n12721 , n12745 );
xor ( n12747 , n12702 , n12746 );
and ( n12748 , n12352 , n12366 );
and ( n12749 , n12366 , n12381 );
and ( n12750 , n12352 , n12381 );
or ( n12751 , n12748 , n12749 , n12750 );
and ( n12752 , n12433 , n12447 );
and ( n12753 , n12447 , n12462 );
and ( n12754 , n12433 , n12462 );
or ( n12755 , n12752 , n12753 , n12754 );
xor ( n12756 , n12751 , n12755 );
and ( n12757 , n9139 , n8209 );
and ( n12758 , n9323 , n8039 );
nor ( n12759 , n12757 , n12758 );
xnor ( n12760 , n12759 , n8165 );
and ( n12761 , n7125 , n11411 );
and ( n12762 , n7196 , n11159 );
nor ( n12763 , n12761 , n12762 );
xnor ( n12764 , n12763 , n11417 );
xor ( n12765 , n12760 , n12764 );
and ( n12766 , n6999 , n12029 );
and ( n12767 , n7049 , n11739 );
nor ( n12768 , n12766 , n12767 );
xnor ( n12769 , n12768 , n12019 );
xor ( n12770 , n12765 , n12769 );
and ( n12771 , n11699 , n7063 );
and ( n12772 , n12010 , n7005 );
nor ( n12773 , n12771 , n12772 );
xnor ( n12774 , n12773 , n7058 );
and ( n12775 , n10548 , n7400 );
and ( n12776 , n10837 , n7303 );
nor ( n12777 , n12775 , n12776 );
xnor ( n12778 , n12777 , n7381 );
xor ( n12779 , n12774 , n12778 );
xor ( n12780 , n12730 , n12349 );
not ( n12781 , n12350 );
and ( n12782 , n12780 , n12781 );
and ( n12783 , n6932 , n12782 );
and ( n12784 , n6960 , n12350 );
nor ( n12785 , n12783 , n12784 );
xnor ( n12786 , n12785 , n12733 );
xor ( n12787 , n12779 , n12786 );
xor ( n12788 , n12770 , n12787 );
and ( n12789 , n10090 , n7609 );
and ( n12790 , n10331 , n7505 );
nor ( n12791 , n12789 , n12790 );
xnor ( n12792 , n12791 , n7615 );
and ( n12793 , n8690 , n8511 );
and ( n12794 , n8913 , n8350 );
nor ( n12795 , n12793 , n12794 );
xnor ( n12796 , n12795 , n8517 );
xor ( n12797 , n12792 , n12796 );
and ( n12798 , n8339 , n8887 );
and ( n12799 , n8548 , n8701 );
nor ( n12800 , n12798 , n12799 );
xnor ( n12801 , n12800 , n8893 );
xor ( n12802 , n12797 , n12801 );
xor ( n12803 , n12788 , n12802 );
xor ( n12804 , n12756 , n12803 );
xor ( n12805 , n12747 , n12804 );
xor ( n12806 , n12698 , n12805 );
xor ( n12807 , n12649 , n12806 );
and ( n12808 , n12320 , n12322 );
and ( n12809 , n12322 , n12466 );
and ( n12810 , n12320 , n12466 );
or ( n12811 , n12808 , n12809 , n12810 );
xor ( n12812 , n12807 , n12811 );
and ( n12813 , n12467 , n12471 );
and ( n12814 , n12472 , n12475 );
or ( n12815 , n12813 , n12814 );
xor ( n12816 , n12812 , n12815 );
buf ( n12817 , n12816 );
and ( n12818 , n12488 , n12544 );
and ( n12819 , n12544 , n12626 );
and ( n12820 , n12488 , n12626 );
or ( n12821 , n12818 , n12819 , n12820 );
buf ( n12822 , n832 );
buf ( n12823 , n12822 );
xor ( n12824 , n12821 , n12823 );
and ( n12825 , n12549 , n12570 );
and ( n12826 , n12570 , n12625 );
and ( n12827 , n12549 , n12625 );
or ( n12828 , n12825 , n12826 , n12827 );
and ( n12829 , n12553 , n12557 );
and ( n12830 , n12557 , n12569 );
and ( n12831 , n12553 , n12569 );
or ( n12832 , n12829 , n12830 , n12831 );
and ( n12833 , n12575 , n12589 );
and ( n12834 , n12589 , n12624 );
and ( n12835 , n12575 , n12624 );
or ( n12836 , n12833 , n12834 , n12835 );
xor ( n12837 , n12832 , n12836 );
and ( n12838 , n12579 , n12583 );
and ( n12839 , n12583 , n12588 );
and ( n12840 , n12579 , n12588 );
or ( n12841 , n12838 , n12839 , n12840 );
and ( n12842 , n9660 , n7948 );
and ( n12843 , n9964 , n7823 );
nor ( n12844 , n12842 , n12843 );
xnor ( n12845 , n12844 , n7938 );
and ( n12846 , n7545 , n10477 );
and ( n12847 , n7661 , n10205 );
nor ( n12848 , n12846 , n12847 );
xnor ( n12849 , n12848 , n10426 );
xor ( n12850 , n12845 , n12849 );
and ( n12851 , n7333 , n11052 );
and ( n12852 , n7427 , n10674 );
nor ( n12853 , n12851 , n12852 );
xnor ( n12854 , n12853 , n10952 );
xor ( n12855 , n12850 , n12854 );
xor ( n12856 , n12841 , n12855 );
and ( n12857 , n11274 , n7260 );
and ( n12858 , n11539 , n7167 );
nor ( n12859 , n12857 , n12858 );
xnor ( n12860 , n12859 , n7250 );
and ( n12861 , n8116 , n9426 );
and ( n12862 , n8241 , n9251 );
nor ( n12863 , n12861 , n12862 );
xnor ( n12864 , n12863 , n9432 );
xor ( n12865 , n12860 , n12864 );
and ( n12866 , n7791 , n9920 );
and ( n12867 , n7966 , n9671 );
nor ( n12868 , n12866 , n12867 );
xnor ( n12869 , n12868 , n9926 );
xor ( n12870 , n12865 , n12869 );
xor ( n12871 , n12856 , n12870 );
xor ( n12872 , n12837 , n12871 );
xor ( n12873 , n12828 , n12872 );
and ( n12874 , n12492 , n12496 );
and ( n12875 , n12496 , n12543 );
and ( n12876 , n12492 , n12543 );
or ( n12877 , n12874 , n12875 , n12876 );
and ( n12878 , n12562 , n12563 );
and ( n12879 , n12563 , n12568 );
and ( n12880 , n12562 , n12568 );
or ( n12881 , n12878 , n12879 , n12880 );
and ( n12882 , n12517 , n12521 );
and ( n12883 , n12521 , n12526 );
and ( n12884 , n12517 , n12526 );
or ( n12885 , n12882 , n12883 , n12884 );
and ( n12886 , n12532 , n12536 );
and ( n12887 , n12536 , n12541 );
and ( n12888 , n12532 , n12541 );
or ( n12889 , n12886 , n12887 , n12888 );
xor ( n12890 , n12885 , n12889 );
and ( n12891 , n12598 , n12602 );
and ( n12892 , n12602 , n12607 );
and ( n12893 , n12598 , n12607 );
or ( n12894 , n12891 , n12892 , n12893 );
xor ( n12895 , n12890 , n12894 );
xor ( n12896 , n12881 , n12895 );
and ( n12897 , n12500 , n6977 );
buf ( n12898 , n768 );
buf ( n12899 , n12898 );
and ( n12900 , n12899 , n6943 );
nor ( n12901 , n12897 , n12900 );
xnor ( n12902 , n12901 , n6974 );
not ( n12903 , n12512 );
buf ( n12904 , n800 );
buf ( n12905 , n12904 );
and ( n12906 , n12510 , n12181 );
not ( n12907 , n12906 );
and ( n12908 , n12905 , n12907 );
and ( n12909 , n12903 , n12908 );
xor ( n12910 , n12902 , n12909 );
and ( n12911 , n12503 , n12507 );
and ( n12912 , n12507 , n12512 );
and ( n12913 , n12503 , n12512 );
or ( n12914 , n12911 , n12912 , n12913 );
xor ( n12915 , n12910 , n12914 );
and ( n12916 , n12613 , n12617 );
and ( n12917 , n12617 , n12622 );
and ( n12918 , n12613 , n12622 );
or ( n12919 , n12916 , n12917 , n12918 );
xor ( n12920 , n12915 , n12919 );
xor ( n12921 , n12896 , n12920 );
xor ( n12922 , n12877 , n12921 );
and ( n12923 , n12513 , n12527 );
and ( n12924 , n12527 , n12542 );
and ( n12925 , n12513 , n12542 );
or ( n12926 , n12923 , n12924 , n12925 );
and ( n12927 , n12594 , n12608 );
and ( n12928 , n12608 , n12623 );
and ( n12929 , n12594 , n12623 );
or ( n12930 , n12927 , n12928 , n12929 );
xor ( n12931 , n12926 , n12930 );
and ( n12932 , n9240 , n8294 );
and ( n12933 , n9438 , n8110 );
nor ( n12934 , n12932 , n12933 );
xnor ( n12935 , n12934 , n8250 );
and ( n12936 , n7156 , n11566 );
and ( n12937 , n7241 , n11300 );
nor ( n12938 , n12936 , n12937 );
xnor ( n12939 , n12938 , n11572 );
xor ( n12940 , n12935 , n12939 );
and ( n12941 , n7020 , n12194 );
and ( n12942 , n7084 , n11890 );
nor ( n12943 , n12941 , n12942 );
xnor ( n12944 , n12943 , n12184 );
xor ( n12945 , n12940 , n12944 );
and ( n12946 , n11850 , n7098 );
and ( n12947 , n12175 , n7026 );
nor ( n12948 , n12946 , n12947 );
xnor ( n12949 , n12948 , n7093 );
and ( n12950 , n10679 , n7455 );
and ( n12951 , n10982 , n7344 );
nor ( n12952 , n12950 , n12951 );
xnor ( n12953 , n12952 , n7436 );
xor ( n12954 , n12949 , n12953 );
xor ( n12955 , n12905 , n12510 );
not ( n12956 , n12511 );
and ( n12957 , n12955 , n12956 );
and ( n12958 , n6941 , n12957 );
and ( n12959 , n6980 , n12511 );
nor ( n12960 , n12958 , n12959 );
xnor ( n12961 , n12960 , n12908 );
xor ( n12962 , n12954 , n12961 );
xor ( n12963 , n12945 , n12962 );
and ( n12964 , n10211 , n7674 );
and ( n12965 , n10466 , n7556 );
nor ( n12966 , n12964 , n12965 );
xnor ( n12967 , n12966 , n7680 );
and ( n12968 , n8781 , n8606 );
and ( n12969 , n9018 , n8431 );
nor ( n12970 , n12968 , n12969 );
xnor ( n12971 , n12970 , n8612 );
xor ( n12972 , n12967 , n12971 );
and ( n12973 , n8420 , n8992 );
and ( n12974 , n8643 , n8792 );
nor ( n12975 , n12973 , n12974 );
xnor ( n12976 , n12975 , n8998 );
xor ( n12977 , n12972 , n12976 );
xor ( n12978 , n12963 , n12977 );
xor ( n12979 , n12931 , n12978 );
xor ( n12980 , n12922 , n12979 );
xor ( n12981 , n12873 , n12980 );
xor ( n12982 , n12824 , n12981 );
and ( n12983 , n12481 , n12483 );
and ( n12984 , n12483 , n12627 );
and ( n12985 , n12481 , n12627 );
or ( n12986 , n12983 , n12984 , n12985 );
xor ( n12987 , n12982 , n12986 );
and ( n12988 , n12628 , n12632 );
and ( n12989 , n12633 , n12636 );
or ( n12990 , n12988 , n12989 );
xor ( n12991 , n12987 , n12990 );
buf ( n12992 , n12991 );
not ( n12993 , n831 );
and ( n12994 , n12993 , n12817 );
and ( n12995 , n12992 , n831 );
or ( n12996 , n12994 , n12995 );
and ( n12997 , n12646 , n12648 );
and ( n12998 , n12648 , n12806 );
and ( n12999 , n12646 , n12806 );
or ( n13000 , n12997 , n12998 , n12999 );
and ( n13001 , n12653 , n12697 );
and ( n13002 , n12697 , n12805 );
and ( n13003 , n12653 , n12805 );
or ( n13004 , n13001 , n13002 , n13003 );
and ( n13005 , n12657 , n12661 );
and ( n13006 , n12661 , n12696 );
and ( n13007 , n12657 , n12696 );
or ( n13008 , n13005 , n13006 , n13007 );
and ( n13009 , n12702 , n12746 );
and ( n13010 , n12746 , n12804 );
and ( n13011 , n12702 , n12804 );
or ( n13012 , n13009 , n13010 , n13011 );
xor ( n13013 , n13008 , n13012 );
and ( n13014 , n12735 , n12739 );
and ( n13015 , n12739 , n12744 );
and ( n13016 , n12735 , n12744 );
or ( n13017 , n13014 , n13015 , n13016 );
and ( n13018 , n12770 , n12787 );
and ( n13019 , n12787 , n12802 );
and ( n13020 , n12770 , n12802 );
or ( n13021 , n13018 , n13019 , n13020 );
xor ( n13022 , n13017 , n13021 );
and ( n13023 , n12670 , n12674 );
and ( n13024 , n12674 , n12679 );
and ( n13025 , n12670 , n12679 );
or ( n13026 , n13023 , n13024 , n13025 );
and ( n13027 , n12760 , n12764 );
and ( n13028 , n12764 , n12769 );
and ( n13029 , n12760 , n12769 );
or ( n13030 , n13027 , n13028 , n13029 );
xor ( n13031 , n13026 , n13030 );
and ( n13032 , n12724 , n6957 );
not ( n13033 , n13032 );
xnor ( n13034 , n13033 , n6954 );
and ( n13035 , n12010 , n7063 );
and ( n13036 , n12339 , n7005 );
nor ( n13037 , n13035 , n13036 );
xnor ( n13038 , n13037 , n7058 );
xor ( n13039 , n13034 , n13038 );
and ( n13040 , n6932 , n12730 );
xor ( n13041 , n13039 , n13040 );
xor ( n13042 , n13031 , n13041 );
xor ( n13043 , n13022 , n13042 );
and ( n13044 , n12666 , n12680 );
and ( n13045 , n12680 , n12695 );
and ( n13046 , n12666 , n12695 );
or ( n13047 , n13044 , n13045 , n13046 );
and ( n13048 , n12685 , n12689 );
and ( n13049 , n12689 , n12694 );
and ( n13050 , n12685 , n12694 );
or ( n13051 , n13048 , n13049 , n13050 );
and ( n13052 , n12774 , n12778 );
and ( n13053 , n12778 , n12786 );
and ( n13054 , n12774 , n12786 );
or ( n13055 , n13052 , n13053 , n13054 );
xor ( n13056 , n13051 , n13055 );
and ( n13057 , n12792 , n12796 );
and ( n13058 , n12796 , n12801 );
and ( n13059 , n12792 , n12801 );
or ( n13060 , n13057 , n13058 , n13059 );
xor ( n13061 , n13056 , n13060 );
xor ( n13062 , n13047 , n13061 );
and ( n13063 , n10331 , n7609 );
and ( n13064 , n10548 , n7505 );
nor ( n13065 , n13063 , n13064 );
xnor ( n13066 , n13065 , n7615 );
and ( n13067 , n8548 , n8887 );
and ( n13068 , n8690 , n8701 );
nor ( n13069 , n13067 , n13068 );
xnor ( n13070 , n13069 , n8893 );
xor ( n13071 , n13066 , n13070 );
and ( n13072 , n8156 , n9311 );
and ( n13073 , n8339 , n9150 );
nor ( n13074 , n13072 , n13073 );
xnor ( n13075 , n13074 , n9317 );
xor ( n13076 , n13071 , n13075 );
and ( n13077 , n11384 , n7215 );
and ( n13078 , n11699 , n7136 );
nor ( n13079 , n13077 , n13078 );
xnor ( n13080 , n13079 , n7205 );
and ( n13081 , n9839 , n7873 );
and ( n13082 , n10090 , n7762 );
nor ( n13083 , n13081 , n13082 );
xnor ( n13084 , n13083 , n7863 );
xor ( n13085 , n13080 , n13084 );
and ( n13086 , n7891 , n9795 );
and ( n13087 , n8045 , n9560 );
nor ( n13088 , n13086 , n13087 );
xnor ( n13089 , n13088 , n9801 );
xor ( n13090 , n13085 , n13089 );
xor ( n13091 , n13076 , n13090 );
and ( n13092 , n9323 , n8209 );
and ( n13093 , n9549 , n8039 );
nor ( n13094 , n13092 , n13093 );
xnor ( n13095 , n13094 , n8165 );
and ( n13096 , n7596 , n10342 );
and ( n13097 , n7730 , n10084 );
nor ( n13098 , n13096 , n13097 );
xnor ( n13099 , n13098 , n10291 );
xor ( n13100 , n13095 , n13099 );
and ( n13101 , n7372 , n10907 );
and ( n13102 , n7494 , n10543 );
nor ( n13103 , n13101 , n13102 );
xnor ( n13104 , n13103 , n10807 );
xor ( n13105 , n13100 , n13104 );
xor ( n13106 , n13091 , n13105 );
xor ( n13107 , n13062 , n13106 );
xor ( n13108 , n13043 , n13107 );
and ( n13109 , n12706 , n12720 );
and ( n13110 , n12720 , n12745 );
and ( n13111 , n12706 , n12745 );
or ( n13112 , n13109 , n13110 , n13111 );
and ( n13113 , n12751 , n12755 );
and ( n13114 , n12755 , n12803 );
and ( n13115 , n12751 , n12803 );
or ( n13116 , n13113 , n13114 , n13115 );
xor ( n13117 , n13112 , n13116 );
and ( n13118 , n12710 , n12714 );
and ( n13119 , n12714 , n12719 );
and ( n13120 , n12710 , n12719 );
or ( n13121 , n13118 , n13119 , n13120 );
and ( n13122 , n10837 , n7400 );
and ( n13123 , n11133 , n7303 );
nor ( n13124 , n13122 , n13123 );
xnor ( n13125 , n13124 , n7381 );
and ( n13126 , n8913 , n8511 );
and ( n13127 , n9139 , n8350 );
nor ( n13128 , n13126 , n13127 );
xnor ( n13129 , n13128 , n8517 );
xor ( n13130 , n13125 , n13129 );
and ( n13131 , n6960 , n12782 );
and ( n13132 , n6999 , n12350 );
nor ( n13133 , n13131 , n13132 );
xnor ( n13134 , n13133 , n12733 );
xor ( n13135 , n13130 , n13134 );
xor ( n13136 , n13121 , n13135 );
and ( n13137 , n12727 , n12734 );
and ( n13138 , n7196 , n11411 );
and ( n13139 , n7292 , n11159 );
nor ( n13140 , n13138 , n13139 );
xnor ( n13141 , n13140 , n11417 );
xor ( n13142 , n13137 , n13141 );
and ( n13143 , n7049 , n12029 );
and ( n13144 , n7125 , n11739 );
nor ( n13145 , n13143 , n13144 );
xnor ( n13146 , n13145 , n12019 );
xor ( n13147 , n13142 , n13146 );
xor ( n13148 , n13136 , n13147 );
xor ( n13149 , n13117 , n13148 );
xor ( n13150 , n13108 , n13149 );
xor ( n13151 , n13013 , n13150 );
xor ( n13152 , n13004 , n13151 );
xor ( n13153 , n13000 , n13152 );
and ( n13154 , n12807 , n12811 );
and ( n13155 , n12812 , n12815 );
or ( n13156 , n13154 , n13155 );
xor ( n13157 , n13153 , n13156 );
buf ( n13158 , n13157 );
and ( n13159 , n12821 , n12823 );
and ( n13160 , n12823 , n12981 );
and ( n13161 , n12821 , n12981 );
or ( n13162 , n13159 , n13160 , n13161 );
and ( n13163 , n12828 , n12872 );
and ( n13164 , n12872 , n12980 );
and ( n13165 , n12828 , n12980 );
or ( n13166 , n13163 , n13164 , n13165 );
and ( n13167 , n12832 , n12836 );
and ( n13168 , n12836 , n12871 );
and ( n13169 , n12832 , n12871 );
or ( n13170 , n13167 , n13168 , n13169 );
and ( n13171 , n12877 , n12921 );
and ( n13172 , n12921 , n12979 );
and ( n13173 , n12877 , n12979 );
or ( n13174 , n13171 , n13172 , n13173 );
xor ( n13175 , n13170 , n13174 );
and ( n13176 , n12910 , n12914 );
and ( n13177 , n12914 , n12919 );
and ( n13178 , n12910 , n12919 );
or ( n13179 , n13176 , n13177 , n13178 );
and ( n13180 , n12945 , n12962 );
and ( n13181 , n12962 , n12977 );
and ( n13182 , n12945 , n12977 );
or ( n13183 , n13180 , n13181 , n13182 );
xor ( n13184 , n13179 , n13183 );
and ( n13185 , n12845 , n12849 );
and ( n13186 , n12849 , n12854 );
and ( n13187 , n12845 , n12854 );
or ( n13188 , n13185 , n13186 , n13187 );
and ( n13189 , n12935 , n12939 );
and ( n13190 , n12939 , n12944 );
and ( n13191 , n12935 , n12944 );
or ( n13192 , n13189 , n13190 , n13191 );
xor ( n13193 , n13188 , n13192 );
and ( n13194 , n12899 , n6977 );
not ( n13195 , n13194 );
xnor ( n13196 , n13195 , n6974 );
and ( n13197 , n12175 , n7098 );
and ( n13198 , n12500 , n7026 );
nor ( n13199 , n13197 , n13198 );
xnor ( n13200 , n13199 , n7093 );
xor ( n13201 , n13196 , n13200 );
and ( n13202 , n6941 , n12905 );
xor ( n13203 , n13201 , n13202 );
xor ( n13204 , n13193 , n13203 );
xor ( n13205 , n13184 , n13204 );
and ( n13206 , n12841 , n12855 );
and ( n13207 , n12855 , n12870 );
and ( n13208 , n12841 , n12870 );
or ( n13209 , n13206 , n13207 , n13208 );
and ( n13210 , n12860 , n12864 );
and ( n13211 , n12864 , n12869 );
and ( n13212 , n12860 , n12869 );
or ( n13213 , n13210 , n13211 , n13212 );
and ( n13214 , n12949 , n12953 );
and ( n13215 , n12953 , n12961 );
and ( n13216 , n12949 , n12961 );
or ( n13217 , n13214 , n13215 , n13216 );
xor ( n13218 , n13213 , n13217 );
and ( n13219 , n12967 , n12971 );
and ( n13220 , n12971 , n12976 );
and ( n13221 , n12967 , n12976 );
or ( n13222 , n13219 , n13220 , n13221 );
xor ( n13223 , n13218 , n13222 );
xor ( n13224 , n13209 , n13223 );
and ( n13225 , n10466 , n7674 );
and ( n13226 , n10679 , n7556 );
nor ( n13227 , n13225 , n13226 );
xnor ( n13228 , n13227 , n7680 );
and ( n13229 , n8643 , n8992 );
and ( n13230 , n8781 , n8792 );
nor ( n13231 , n13229 , n13230 );
xnor ( n13232 , n13231 , n8998 );
xor ( n13233 , n13228 , n13232 );
and ( n13234 , n8241 , n9426 );
and ( n13235 , n8420 , n9251 );
nor ( n13236 , n13234 , n13235 );
xnor ( n13237 , n13236 , n9432 );
xor ( n13238 , n13233 , n13237 );
and ( n13239 , n11539 , n7260 );
and ( n13240 , n11850 , n7167 );
nor ( n13241 , n13239 , n13240 );
xnor ( n13242 , n13241 , n7250 );
and ( n13243 , n9964 , n7948 );
and ( n13244 , n10211 , n7823 );
nor ( n13245 , n13243 , n13244 );
xnor ( n13246 , n13245 , n7938 );
xor ( n13247 , n13242 , n13246 );
and ( n13248 , n7966 , n9920 );
and ( n13249 , n8116 , n9671 );
nor ( n13250 , n13248 , n13249 );
xnor ( n13251 , n13250 , n9926 );
xor ( n13252 , n13247 , n13251 );
xor ( n13253 , n13238 , n13252 );
and ( n13254 , n9438 , n8294 );
and ( n13255 , n9660 , n8110 );
nor ( n13256 , n13254 , n13255 );
xnor ( n13257 , n13256 , n8250 );
and ( n13258 , n7661 , n10477 );
and ( n13259 , n7791 , n10205 );
nor ( n13260 , n13258 , n13259 );
xnor ( n13261 , n13260 , n10426 );
xor ( n13262 , n13257 , n13261 );
and ( n13263 , n7427 , n11052 );
and ( n13264 , n7545 , n10674 );
nor ( n13265 , n13263 , n13264 );
xnor ( n13266 , n13265 , n10952 );
xor ( n13267 , n13262 , n13266 );
xor ( n13268 , n13253 , n13267 );
xor ( n13269 , n13224 , n13268 );
xor ( n13270 , n13205 , n13269 );
and ( n13271 , n12881 , n12895 );
and ( n13272 , n12895 , n12920 );
and ( n13273 , n12881 , n12920 );
or ( n13274 , n13271 , n13272 , n13273 );
and ( n13275 , n12926 , n12930 );
and ( n13276 , n12930 , n12978 );
and ( n13277 , n12926 , n12978 );
or ( n13278 , n13275 , n13276 , n13277 );
xor ( n13279 , n13274 , n13278 );
and ( n13280 , n12885 , n12889 );
and ( n13281 , n12889 , n12894 );
and ( n13282 , n12885 , n12894 );
or ( n13283 , n13280 , n13281 , n13282 );
and ( n13284 , n10982 , n7455 );
and ( n13285 , n11274 , n7344 );
nor ( n13286 , n13284 , n13285 );
xnor ( n13287 , n13286 , n7436 );
and ( n13288 , n9018 , n8606 );
and ( n13289 , n9240 , n8431 );
nor ( n13290 , n13288 , n13289 );
xnor ( n13291 , n13290 , n8612 );
xor ( n13292 , n13287 , n13291 );
and ( n13293 , n6980 , n12957 );
and ( n13294 , n7020 , n12511 );
nor ( n13295 , n13293 , n13294 );
xnor ( n13296 , n13295 , n12908 );
xor ( n13297 , n13292 , n13296 );
xor ( n13298 , n13283 , n13297 );
and ( n13299 , n12902 , n12909 );
and ( n13300 , n7241 , n11566 );
and ( n13301 , n7333 , n11300 );
nor ( n13302 , n13300 , n13301 );
xnor ( n13303 , n13302 , n11572 );
xor ( n13304 , n13299 , n13303 );
and ( n13305 , n7084 , n12194 );
and ( n13306 , n7156 , n11890 );
nor ( n13307 , n13305 , n13306 );
xnor ( n13308 , n13307 , n12184 );
xor ( n13309 , n13304 , n13308 );
xor ( n13310 , n13298 , n13309 );
xor ( n13311 , n13279 , n13310 );
xor ( n13312 , n13270 , n13311 );
xor ( n13313 , n13175 , n13312 );
xor ( n13314 , n13166 , n13313 );
xor ( n13315 , n13162 , n13314 );
and ( n13316 , n12982 , n12986 );
and ( n13317 , n12987 , n12990 );
or ( n13318 , n13316 , n13317 );
xor ( n13319 , n13315 , n13318 );
buf ( n13320 , n13319 );
not ( n13321 , n831 );
and ( n13322 , n13321 , n13158 );
and ( n13323 , n13320 , n831 );
or ( n13324 , n13322 , n13323 );
and ( n13325 , n13000 , n13152 );
and ( n13326 , n13008 , n13012 );
and ( n13327 , n13012 , n13150 );
and ( n13328 , n13008 , n13150 );
or ( n13329 , n13326 , n13327 , n13328 );
and ( n13330 , n13043 , n13107 );
and ( n13331 , n13107 , n13149 );
and ( n13332 , n13043 , n13149 );
or ( n13333 , n13330 , n13331 , n13332 );
and ( n13334 , n13017 , n13021 );
and ( n13335 , n13021 , n13042 );
and ( n13336 , n13017 , n13042 );
or ( n13337 , n13334 , n13335 , n13336 );
and ( n13338 , n13051 , n13055 );
and ( n13339 , n13055 , n13060 );
and ( n13340 , n13051 , n13060 );
or ( n13341 , n13338 , n13339 , n13340 );
and ( n13342 , n13137 , n13141 );
and ( n13343 , n13141 , n13146 );
and ( n13344 , n13137 , n13146 );
or ( n13345 , n13342 , n13343 , n13344 );
xor ( n13346 , n13341 , n13345 );
and ( n13347 , n13026 , n13030 );
and ( n13348 , n13030 , n13041 );
and ( n13349 , n13026 , n13041 );
or ( n13350 , n13347 , n13348 , n13349 );
xor ( n13351 , n13346 , n13350 );
xor ( n13352 , n13337 , n13351 );
and ( n13353 , n13076 , n13090 );
and ( n13354 , n13090 , n13105 );
and ( n13355 , n13076 , n13105 );
or ( n13356 , n13353 , n13354 , n13355 );
and ( n13357 , n13066 , n13070 );
and ( n13358 , n13070 , n13075 );
and ( n13359 , n13066 , n13075 );
or ( n13360 , n13357 , n13358 , n13359 );
and ( n13361 , n13095 , n13099 );
and ( n13362 , n13099 , n13104 );
and ( n13363 , n13095 , n13104 );
or ( n13364 , n13361 , n13362 , n13363 );
xor ( n13365 , n13360 , n13364 );
and ( n13366 , n13125 , n13129 );
and ( n13367 , n13129 , n13134 );
and ( n13368 , n13125 , n13134 );
or ( n13369 , n13366 , n13367 , n13368 );
xor ( n13370 , n13365 , n13369 );
xor ( n13371 , n13356 , n13370 );
and ( n13372 , n13034 , n13038 );
and ( n13373 , n13038 , n13040 );
and ( n13374 , n13034 , n13040 );
or ( n13375 , n13372 , n13373 , n13374 );
xor ( n13376 , n13375 , n6954 );
and ( n13377 , n7125 , n12029 );
and ( n13378 , n7196 , n11739 );
nor ( n13379 , n13377 , n13378 );
xnor ( n13380 , n13379 , n12019 );
xor ( n13381 , n13376 , n13380 );
xor ( n13382 , n13371 , n13381 );
xor ( n13383 , n13352 , n13382 );
xor ( n13384 , n13333 , n13383 );
and ( n13385 , n13047 , n13061 );
and ( n13386 , n13061 , n13106 );
and ( n13387 , n13047 , n13106 );
or ( n13388 , n13385 , n13386 , n13387 );
and ( n13389 , n13112 , n13116 );
and ( n13390 , n13116 , n13148 );
and ( n13391 , n13112 , n13148 );
or ( n13392 , n13389 , n13390 , n13391 );
xor ( n13393 , n13388 , n13392 );
and ( n13394 , n13121 , n13135 );
and ( n13395 , n13135 , n13147 );
and ( n13396 , n13121 , n13147 );
or ( n13397 , n13394 , n13395 , n13396 );
and ( n13398 , n11699 , n7215 );
and ( n13399 , n12010 , n7136 );
nor ( n13400 , n13398 , n13399 );
xnor ( n13401 , n13400 , n7205 );
and ( n13402 , n10090 , n7873 );
and ( n13403 , n10331 , n7762 );
nor ( n13404 , n13402 , n13403 );
xnor ( n13405 , n13404 , n7863 );
xor ( n13406 , n13401 , n13405 );
and ( n13407 , n7730 , n10342 );
and ( n13408 , n7891 , n10084 );
nor ( n13409 , n13407 , n13408 );
xnor ( n13410 , n13409 , n10291 );
xor ( n13411 , n13406 , n13410 );
and ( n13412 , n10548 , n7609 );
and ( n13413 , n10837 , n7505 );
nor ( n13414 , n13412 , n13413 );
xnor ( n13415 , n13414 , n7615 );
and ( n13416 , n8339 , n9311 );
and ( n13417 , n8548 , n9150 );
nor ( n13418 , n13416 , n13417 );
xnor ( n13419 , n13418 , n9317 );
xor ( n13420 , n13415 , n13419 );
and ( n13421 , n8045 , n9795 );
and ( n13422 , n8156 , n9560 );
nor ( n13423 , n13421 , n13422 );
xnor ( n13424 , n13423 , n9801 );
xor ( n13425 , n13420 , n13424 );
xor ( n13426 , n13411 , n13425 );
and ( n13427 , n12339 , n7063 );
and ( n13428 , n12724 , n7005 );
nor ( n13429 , n13427 , n13428 );
xnor ( n13430 , n13429 , n7058 );
and ( n13431 , n11133 , n7400 );
and ( n13432 , n11384 , n7303 );
nor ( n13433 , n13431 , n13432 );
xnor ( n13434 , n13433 , n7381 );
xor ( n13435 , n13430 , n13434 );
and ( n13436 , n8690 , n8887 );
and ( n13437 , n8913 , n8701 );
nor ( n13438 , n13436 , n13437 );
xnor ( n13439 , n13438 , n8893 );
xor ( n13440 , n13435 , n13439 );
xor ( n13441 , n13426 , n13440 );
xor ( n13442 , n13397 , n13441 );
and ( n13443 , n13080 , n13084 );
and ( n13444 , n13084 , n13089 );
and ( n13445 , n13080 , n13089 );
or ( n13446 , n13443 , n13444 , n13445 );
and ( n13447 , n9549 , n8209 );
and ( n13448 , n9839 , n8039 );
nor ( n13449 , n13447 , n13448 );
xnor ( n13450 , n13449 , n8165 );
and ( n13451 , n7494 , n10907 );
and ( n13452 , n7596 , n10543 );
nor ( n13453 , n13451 , n13452 );
xnor ( n13454 , n13453 , n10807 );
xor ( n13455 , n13450 , n13454 );
and ( n13456 , n7292 , n11411 );
and ( n13457 , n7372 , n11159 );
nor ( n13458 , n13456 , n13457 );
xnor ( n13459 , n13458 , n11417 );
xor ( n13460 , n13455 , n13459 );
xor ( n13461 , n13446 , n13460 );
and ( n13462 , n9139 , n8511 );
and ( n13463 , n9323 , n8350 );
nor ( n13464 , n13462 , n13463 );
xnor ( n13465 , n13464 , n8517 );
and ( n13466 , n6999 , n12782 );
and ( n13467 , n7049 , n12350 );
nor ( n13468 , n13466 , n13467 );
xnor ( n13469 , n13468 , n12733 );
xor ( n13470 , n13465 , n13469 );
and ( n13471 , n6960 , n12730 );
xor ( n13472 , n13470 , n13471 );
xor ( n13473 , n13461 , n13472 );
xor ( n13474 , n13442 , n13473 );
xor ( n13475 , n13393 , n13474 );
xor ( n13476 , n13384 , n13475 );
xor ( n13477 , n13329 , n13476 );
and ( n13478 , n13004 , n13151 );
xor ( n13479 , n13477 , n13478 );
xor ( n13480 , n13325 , n13479 );
and ( n13481 , n13153 , n13156 );
xor ( n13482 , n13480 , n13481 );
buf ( n13483 , n13482 );
and ( n13484 , n13162 , n13314 );
and ( n13485 , n13170 , n13174 );
and ( n13486 , n13174 , n13312 );
and ( n13487 , n13170 , n13312 );
or ( n13488 , n13485 , n13486 , n13487 );
and ( n13489 , n13205 , n13269 );
and ( n13490 , n13269 , n13311 );
and ( n13491 , n13205 , n13311 );
or ( n13492 , n13489 , n13490 , n13491 );
and ( n13493 , n13179 , n13183 );
and ( n13494 , n13183 , n13204 );
and ( n13495 , n13179 , n13204 );
or ( n13496 , n13493 , n13494 , n13495 );
and ( n13497 , n13213 , n13217 );
and ( n13498 , n13217 , n13222 );
and ( n13499 , n13213 , n13222 );
or ( n13500 , n13497 , n13498 , n13499 );
and ( n13501 , n13299 , n13303 );
and ( n13502 , n13303 , n13308 );
and ( n13503 , n13299 , n13308 );
or ( n13504 , n13501 , n13502 , n13503 );
xor ( n13505 , n13500 , n13504 );
and ( n13506 , n13188 , n13192 );
and ( n13507 , n13192 , n13203 );
and ( n13508 , n13188 , n13203 );
or ( n13509 , n13506 , n13507 , n13508 );
xor ( n13510 , n13505 , n13509 );
xor ( n13511 , n13496 , n13510 );
and ( n13512 , n13238 , n13252 );
and ( n13513 , n13252 , n13267 );
and ( n13514 , n13238 , n13267 );
or ( n13515 , n13512 , n13513 , n13514 );
and ( n13516 , n13228 , n13232 );
and ( n13517 , n13232 , n13237 );
and ( n13518 , n13228 , n13237 );
or ( n13519 , n13516 , n13517 , n13518 );
and ( n13520 , n13257 , n13261 );
and ( n13521 , n13261 , n13266 );
and ( n13522 , n13257 , n13266 );
or ( n13523 , n13520 , n13521 , n13522 );
xor ( n13524 , n13519 , n13523 );
and ( n13525 , n13287 , n13291 );
and ( n13526 , n13291 , n13296 );
and ( n13527 , n13287 , n13296 );
or ( n13528 , n13525 , n13526 , n13527 );
xor ( n13529 , n13524 , n13528 );
xor ( n13530 , n13515 , n13529 );
and ( n13531 , n13196 , n13200 );
and ( n13532 , n13200 , n13202 );
and ( n13533 , n13196 , n13202 );
or ( n13534 , n13531 , n13532 , n13533 );
xor ( n13535 , n13534 , n6974 );
and ( n13536 , n7156 , n12194 );
and ( n13537 , n7241 , n11890 );
nor ( n13538 , n13536 , n13537 );
xnor ( n13539 , n13538 , n12184 );
xor ( n13540 , n13535 , n13539 );
xor ( n13541 , n13530 , n13540 );
xor ( n13542 , n13511 , n13541 );
xor ( n13543 , n13492 , n13542 );
and ( n13544 , n13209 , n13223 );
and ( n13545 , n13223 , n13268 );
and ( n13546 , n13209 , n13268 );
or ( n13547 , n13544 , n13545 , n13546 );
and ( n13548 , n13274 , n13278 );
and ( n13549 , n13278 , n13310 );
and ( n13550 , n13274 , n13310 );
or ( n13551 , n13548 , n13549 , n13550 );
xor ( n13552 , n13547 , n13551 );
and ( n13553 , n13283 , n13297 );
and ( n13554 , n13297 , n13309 );
and ( n13555 , n13283 , n13309 );
or ( n13556 , n13553 , n13554 , n13555 );
and ( n13557 , n11850 , n7260 );
and ( n13558 , n12175 , n7167 );
nor ( n13559 , n13557 , n13558 );
xnor ( n13560 , n13559 , n7250 );
and ( n13561 , n10211 , n7948 );
and ( n13562 , n10466 , n7823 );
nor ( n13563 , n13561 , n13562 );
xnor ( n13564 , n13563 , n7938 );
xor ( n13565 , n13560 , n13564 );
and ( n13566 , n7791 , n10477 );
and ( n13567 , n7966 , n10205 );
nor ( n13568 , n13566 , n13567 );
xnor ( n13569 , n13568 , n10426 );
xor ( n13570 , n13565 , n13569 );
and ( n13571 , n10679 , n7674 );
and ( n13572 , n10982 , n7556 );
nor ( n13573 , n13571 , n13572 );
xnor ( n13574 , n13573 , n7680 );
and ( n13575 , n8420 , n9426 );
and ( n13576 , n8643 , n9251 );
nor ( n13577 , n13575 , n13576 );
xnor ( n13578 , n13577 , n9432 );
xor ( n13579 , n13574 , n13578 );
and ( n13580 , n8116 , n9920 );
and ( n13581 , n8241 , n9671 );
nor ( n13582 , n13580 , n13581 );
xnor ( n13583 , n13582 , n9926 );
xor ( n13584 , n13579 , n13583 );
xor ( n13585 , n13570 , n13584 );
and ( n13586 , n12500 , n7098 );
and ( n13587 , n12899 , n7026 );
nor ( n13588 , n13586 , n13587 );
xnor ( n13589 , n13588 , n7093 );
and ( n13590 , n11274 , n7455 );
and ( n13591 , n11539 , n7344 );
nor ( n13592 , n13590 , n13591 );
xnor ( n13593 , n13592 , n7436 );
xor ( n13594 , n13589 , n13593 );
and ( n13595 , n8781 , n8992 );
and ( n13596 , n9018 , n8792 );
nor ( n13597 , n13595 , n13596 );
xnor ( n13598 , n13597 , n8998 );
xor ( n13599 , n13594 , n13598 );
xor ( n13600 , n13585 , n13599 );
xor ( n13601 , n13556 , n13600 );
and ( n13602 , n13242 , n13246 );
and ( n13603 , n13246 , n13251 );
and ( n13604 , n13242 , n13251 );
or ( n13605 , n13602 , n13603 , n13604 );
and ( n13606 , n9660 , n8294 );
and ( n13607 , n9964 , n8110 );
nor ( n13608 , n13606 , n13607 );
xnor ( n13609 , n13608 , n8250 );
and ( n13610 , n7545 , n11052 );
and ( n13611 , n7661 , n10674 );
nor ( n13612 , n13610 , n13611 );
xnor ( n13613 , n13612 , n10952 );
xor ( n13614 , n13609 , n13613 );
and ( n13615 , n7333 , n11566 );
and ( n13616 , n7427 , n11300 );
nor ( n13617 , n13615 , n13616 );
xnor ( n13618 , n13617 , n11572 );
xor ( n13619 , n13614 , n13618 );
xor ( n13620 , n13605 , n13619 );
and ( n13621 , n9240 , n8606 );
and ( n13622 , n9438 , n8431 );
nor ( n13623 , n13621 , n13622 );
xnor ( n13624 , n13623 , n8612 );
and ( n13625 , n7020 , n12957 );
and ( n13626 , n7084 , n12511 );
nor ( n13627 , n13625 , n13626 );
xnor ( n13628 , n13627 , n12908 );
xor ( n13629 , n13624 , n13628 );
and ( n13630 , n6980 , n12905 );
xor ( n13631 , n13629 , n13630 );
xor ( n13632 , n13620 , n13631 );
xor ( n13633 , n13601 , n13632 );
xor ( n13634 , n13552 , n13633 );
xor ( n13635 , n13543 , n13634 );
xor ( n13636 , n13488 , n13635 );
and ( n13637 , n13166 , n13313 );
xor ( n13638 , n13636 , n13637 );
xor ( n13639 , n13484 , n13638 );
and ( n13640 , n13315 , n13318 );
xor ( n13641 , n13639 , n13640 );
buf ( n13642 , n13641 );
not ( n13643 , n831 );
and ( n13644 , n13643 , n13483 );
and ( n13645 , n13642 , n831 );
or ( n13646 , n13644 , n13645 );
and ( n13647 , n13477 , n13478 );
and ( n13648 , n13333 , n13383 );
and ( n13649 , n13383 , n13475 );
and ( n13650 , n13333 , n13475 );
or ( n13651 , n13648 , n13649 , n13650 );
and ( n13652 , n13388 , n13392 );
and ( n13653 , n13392 , n13474 );
and ( n13654 , n13388 , n13474 );
or ( n13655 , n13652 , n13653 , n13654 );
and ( n13656 , n13341 , n13345 );
and ( n13657 , n13345 , n13350 );
and ( n13658 , n13341 , n13350 );
or ( n13659 , n13656 , n13657 , n13658 );
and ( n13660 , n13360 , n13364 );
and ( n13661 , n13364 , n13369 );
and ( n13662 , n13360 , n13369 );
or ( n13663 , n13660 , n13661 , n13662 );
and ( n13664 , n13375 , n6954 );
and ( n13665 , n6954 , n13380 );
and ( n13666 , n13375 , n13380 );
or ( n13667 , n13664 , n13665 , n13666 );
xor ( n13668 , n13663 , n13667 );
and ( n13669 , n13401 , n13405 );
and ( n13670 , n13405 , n13410 );
and ( n13671 , n13401 , n13410 );
or ( n13672 , n13669 , n13670 , n13671 );
and ( n13673 , n13415 , n13419 );
and ( n13674 , n13419 , n13424 );
and ( n13675 , n13415 , n13424 );
or ( n13676 , n13673 , n13674 , n13675 );
xor ( n13677 , n13672 , n13676 );
and ( n13678 , n13430 , n13434 );
and ( n13679 , n13434 , n13439 );
and ( n13680 , n13430 , n13439 );
or ( n13681 , n13678 , n13679 , n13680 );
xor ( n13682 , n13677 , n13681 );
xor ( n13683 , n13668 , n13682 );
xor ( n13684 , n13659 , n13683 );
and ( n13685 , n13411 , n13425 );
and ( n13686 , n13425 , n13440 );
and ( n13687 , n13411 , n13440 );
or ( n13688 , n13685 , n13686 , n13687 );
and ( n13689 , n13446 , n13460 );
and ( n13690 , n13460 , n13472 );
and ( n13691 , n13446 , n13472 );
or ( n13692 , n13689 , n13690 , n13691 );
xor ( n13693 , n13688 , n13692 );
and ( n13694 , n13465 , n13469 );
and ( n13695 , n13469 , n13471 );
and ( n13696 , n13465 , n13471 );
or ( n13697 , n13694 , n13695 , n13696 );
not ( n13698 , n6954 );
buf ( n13699 , n13698 );
xor ( n13700 , n13697 , n13699 );
and ( n13701 , n12724 , n7063 );
not ( n13702 , n13701 );
xnor ( n13703 , n13702 , n7058 );
not ( n13704 , n13703 );
xor ( n13705 , n13700 , n13704 );
xor ( n13706 , n13693 , n13705 );
xor ( n13707 , n13684 , n13706 );
xor ( n13708 , n13655 , n13707 );
and ( n13709 , n13397 , n13441 );
and ( n13710 , n13441 , n13473 );
and ( n13711 , n13397 , n13473 );
or ( n13712 , n13709 , n13710 , n13711 );
and ( n13713 , n13337 , n13351 );
and ( n13714 , n13351 , n13382 );
and ( n13715 , n13337 , n13382 );
or ( n13716 , n13713 , n13714 , n13715 );
xor ( n13717 , n13712 , n13716 );
and ( n13718 , n13356 , n13370 );
and ( n13719 , n13370 , n13381 );
and ( n13720 , n13356 , n13381 );
or ( n13721 , n13718 , n13719 , n13720 );
and ( n13722 , n13450 , n13454 );
and ( n13723 , n13454 , n13459 );
and ( n13724 , n13450 , n13459 );
or ( n13725 , n13722 , n13723 , n13724 );
and ( n13726 , n9323 , n8511 );
and ( n13727 , n9549 , n8350 );
nor ( n13728 , n13726 , n13727 );
xnor ( n13729 , n13728 , n8517 );
and ( n13730 , n7196 , n12029 );
and ( n13731 , n7292 , n11739 );
nor ( n13732 , n13730 , n13731 );
xnor ( n13733 , n13732 , n12019 );
xor ( n13734 , n13729 , n13733 );
and ( n13735 , n7049 , n12782 );
and ( n13736 , n7125 , n12350 );
nor ( n13737 , n13735 , n13736 );
xnor ( n13738 , n13737 , n12733 );
xor ( n13739 , n13734 , n13738 );
xor ( n13740 , n13725 , n13739 );
and ( n13741 , n10331 , n7873 );
and ( n13742 , n10548 , n7762 );
nor ( n13743 , n13741 , n13742 );
xnor ( n13744 , n13743 , n7863 );
and ( n13745 , n8913 , n8887 );
and ( n13746 , n9139 , n8701 );
nor ( n13747 , n13745 , n13746 );
xnor ( n13748 , n13747 , n8893 );
xor ( n13749 , n13744 , n13748 );
and ( n13750 , n8548 , n9311 );
and ( n13751 , n8690 , n9150 );
nor ( n13752 , n13750 , n13751 );
xnor ( n13753 , n13752 , n9317 );
xor ( n13754 , n13749 , n13753 );
xor ( n13755 , n13740 , n13754 );
xor ( n13756 , n13721 , n13755 );
and ( n13757 , n12010 , n7215 );
and ( n13758 , n12339 , n7136 );
nor ( n13759 , n13757 , n13758 );
xnor ( n13760 , n13759 , n7205 );
and ( n13761 , n10837 , n7609 );
and ( n13762 , n11133 , n7505 );
nor ( n13763 , n13761 , n13762 );
xnor ( n13764 , n13763 , n7615 );
xor ( n13765 , n13760 , n13764 );
and ( n13766 , n6999 , n12730 );
xor ( n13767 , n13765 , n13766 );
and ( n13768 , n9839 , n8209 );
and ( n13769 , n10090 , n8039 );
nor ( n13770 , n13768 , n13769 );
xnor ( n13771 , n13770 , n8165 );
and ( n13772 , n7596 , n10907 );
and ( n13773 , n7730 , n10543 );
nor ( n13774 , n13772 , n13773 );
xnor ( n13775 , n13774 , n10807 );
xor ( n13776 , n13771 , n13775 );
and ( n13777 , n7372 , n11411 );
and ( n13778 , n7494 , n11159 );
nor ( n13779 , n13777 , n13778 );
xnor ( n13780 , n13779 , n11417 );
xor ( n13781 , n13776 , n13780 );
xor ( n13782 , n13767 , n13781 );
and ( n13783 , n11384 , n7400 );
and ( n13784 , n11699 , n7303 );
nor ( n13785 , n13783 , n13784 );
xnor ( n13786 , n13785 , n7381 );
and ( n13787 , n8156 , n9795 );
and ( n13788 , n8339 , n9560 );
nor ( n13789 , n13787 , n13788 );
xnor ( n13790 , n13789 , n9801 );
xor ( n13791 , n13786 , n13790 );
and ( n13792 , n7891 , n10342 );
and ( n13793 , n8045 , n10084 );
nor ( n13794 , n13792 , n13793 );
xnor ( n13795 , n13794 , n10291 );
xor ( n13796 , n13791 , n13795 );
xor ( n13797 , n13782 , n13796 );
xor ( n13798 , n13756 , n13797 );
xor ( n13799 , n13717 , n13798 );
xor ( n13800 , n13708 , n13799 );
xor ( n13801 , n13651 , n13800 );
and ( n13802 , n13329 , n13476 );
xor ( n13803 , n13801 , n13802 );
xor ( n13804 , n13647 , n13803 );
and ( n13805 , n13325 , n13479 );
and ( n13806 , n13480 , n13481 );
or ( n13807 , n13805 , n13806 );
xor ( n13808 , n13804 , n13807 );
buf ( n13809 , n13808 );
and ( n13810 , n13636 , n13637 );
and ( n13811 , n13492 , n13542 );
and ( n13812 , n13542 , n13634 );
and ( n13813 , n13492 , n13634 );
or ( n13814 , n13811 , n13812 , n13813 );
and ( n13815 , n13547 , n13551 );
and ( n13816 , n13551 , n13633 );
and ( n13817 , n13547 , n13633 );
or ( n13818 , n13815 , n13816 , n13817 );
and ( n13819 , n13500 , n13504 );
and ( n13820 , n13504 , n13509 );
and ( n13821 , n13500 , n13509 );
or ( n13822 , n13819 , n13820 , n13821 );
and ( n13823 , n13519 , n13523 );
and ( n13824 , n13523 , n13528 );
and ( n13825 , n13519 , n13528 );
or ( n13826 , n13823 , n13824 , n13825 );
and ( n13827 , n13534 , n6974 );
and ( n13828 , n6974 , n13539 );
and ( n13829 , n13534 , n13539 );
or ( n13830 , n13827 , n13828 , n13829 );
xor ( n13831 , n13826 , n13830 );
and ( n13832 , n13560 , n13564 );
and ( n13833 , n13564 , n13569 );
and ( n13834 , n13560 , n13569 );
or ( n13835 , n13832 , n13833 , n13834 );
and ( n13836 , n13574 , n13578 );
and ( n13837 , n13578 , n13583 );
and ( n13838 , n13574 , n13583 );
or ( n13839 , n13836 , n13837 , n13838 );
xor ( n13840 , n13835 , n13839 );
and ( n13841 , n13589 , n13593 );
and ( n13842 , n13593 , n13598 );
and ( n13843 , n13589 , n13598 );
or ( n13844 , n13841 , n13842 , n13843 );
xor ( n13845 , n13840 , n13844 );
xor ( n13846 , n13831 , n13845 );
xor ( n13847 , n13822 , n13846 );
and ( n13848 , n13570 , n13584 );
and ( n13849 , n13584 , n13599 );
and ( n13850 , n13570 , n13599 );
or ( n13851 , n13848 , n13849 , n13850 );
and ( n13852 , n13605 , n13619 );
and ( n13853 , n13619 , n13631 );
and ( n13854 , n13605 , n13631 );
or ( n13855 , n13852 , n13853 , n13854 );
xor ( n13856 , n13851 , n13855 );
and ( n13857 , n13624 , n13628 );
and ( n13858 , n13628 , n13630 );
and ( n13859 , n13624 , n13630 );
or ( n13860 , n13857 , n13858 , n13859 );
not ( n13861 , n6974 );
buf ( n13862 , n13861 );
xor ( n13863 , n13860 , n13862 );
and ( n13864 , n12899 , n7098 );
not ( n13865 , n13864 );
xnor ( n13866 , n13865 , n7093 );
not ( n13867 , n13866 );
xor ( n13868 , n13863 , n13867 );
xor ( n13869 , n13856 , n13868 );
xor ( n13870 , n13847 , n13869 );
xor ( n13871 , n13818 , n13870 );
and ( n13872 , n13556 , n13600 );
and ( n13873 , n13600 , n13632 );
and ( n13874 , n13556 , n13632 );
or ( n13875 , n13872 , n13873 , n13874 );
and ( n13876 , n13496 , n13510 );
and ( n13877 , n13510 , n13541 );
and ( n13878 , n13496 , n13541 );
or ( n13879 , n13876 , n13877 , n13878 );
xor ( n13880 , n13875 , n13879 );
and ( n13881 , n13515 , n13529 );
and ( n13882 , n13529 , n13540 );
and ( n13883 , n13515 , n13540 );
or ( n13884 , n13881 , n13882 , n13883 );
and ( n13885 , n13609 , n13613 );
and ( n13886 , n13613 , n13618 );
and ( n13887 , n13609 , n13618 );
or ( n13888 , n13885 , n13886 , n13887 );
and ( n13889 , n9438 , n8606 );
and ( n13890 , n9660 , n8431 );
nor ( n13891 , n13889 , n13890 );
xnor ( n13892 , n13891 , n8612 );
and ( n13893 , n7241 , n12194 );
and ( n13894 , n7333 , n11890 );
nor ( n13895 , n13893 , n13894 );
xnor ( n13896 , n13895 , n12184 );
xor ( n13897 , n13892 , n13896 );
and ( n13898 , n7084 , n12957 );
and ( n13899 , n7156 , n12511 );
nor ( n13900 , n13898 , n13899 );
xnor ( n13901 , n13900 , n12908 );
xor ( n13902 , n13897 , n13901 );
xor ( n13903 , n13888 , n13902 );
and ( n13904 , n10466 , n7948 );
and ( n13905 , n10679 , n7823 );
nor ( n13906 , n13904 , n13905 );
xnor ( n13907 , n13906 , n7938 );
and ( n13908 , n9018 , n8992 );
and ( n13909 , n9240 , n8792 );
nor ( n13910 , n13908 , n13909 );
xnor ( n13911 , n13910 , n8998 );
xor ( n13912 , n13907 , n13911 );
and ( n13913 , n8643 , n9426 );
and ( n13914 , n8781 , n9251 );
nor ( n13915 , n13913 , n13914 );
xnor ( n13916 , n13915 , n9432 );
xor ( n13917 , n13912 , n13916 );
xor ( n13918 , n13903 , n13917 );
xor ( n13919 , n13884 , n13918 );
and ( n13920 , n12175 , n7260 );
and ( n13921 , n12500 , n7167 );
nor ( n13922 , n13920 , n13921 );
xnor ( n13923 , n13922 , n7250 );
and ( n13924 , n10982 , n7674 );
and ( n13925 , n11274 , n7556 );
nor ( n13926 , n13924 , n13925 );
xnor ( n13927 , n13926 , n7680 );
xor ( n13928 , n13923 , n13927 );
and ( n13929 , n7020 , n12905 );
xor ( n13930 , n13928 , n13929 );
and ( n13931 , n9964 , n8294 );
and ( n13932 , n10211 , n8110 );
nor ( n13933 , n13931 , n13932 );
xnor ( n13934 , n13933 , n8250 );
and ( n13935 , n7661 , n11052 );
and ( n13936 , n7791 , n10674 );
nor ( n13937 , n13935 , n13936 );
xnor ( n13938 , n13937 , n10952 );
xor ( n13939 , n13934 , n13938 );
and ( n13940 , n7427 , n11566 );
and ( n13941 , n7545 , n11300 );
nor ( n13942 , n13940 , n13941 );
xnor ( n13943 , n13942 , n11572 );
xor ( n13944 , n13939 , n13943 );
xor ( n13945 , n13930 , n13944 );
and ( n13946 , n11539 , n7455 );
and ( n13947 , n11850 , n7344 );
nor ( n13948 , n13946 , n13947 );
xnor ( n13949 , n13948 , n7436 );
and ( n13950 , n8241 , n9920 );
and ( n13951 , n8420 , n9671 );
nor ( n13952 , n13950 , n13951 );
xnor ( n13953 , n13952 , n9926 );
xor ( n13954 , n13949 , n13953 );
and ( n13955 , n7966 , n10477 );
and ( n13956 , n8116 , n10205 );
nor ( n13957 , n13955 , n13956 );
xnor ( n13958 , n13957 , n10426 );
xor ( n13959 , n13954 , n13958 );
xor ( n13960 , n13945 , n13959 );
xor ( n13961 , n13919 , n13960 );
xor ( n13962 , n13880 , n13961 );
xor ( n13963 , n13871 , n13962 );
xor ( n13964 , n13814 , n13963 );
and ( n13965 , n13488 , n13635 );
xor ( n13966 , n13964 , n13965 );
xor ( n13967 , n13810 , n13966 );
and ( n13968 , n13484 , n13638 );
and ( n13969 , n13639 , n13640 );
or ( n13970 , n13968 , n13969 );
xor ( n13971 , n13967 , n13970 );
buf ( n13972 , n13971 );
not ( n13973 , n831 );
and ( n13974 , n13973 , n13809 );
and ( n13975 , n13972 , n831 );
or ( n13976 , n13974 , n13975 );
and ( n13977 , n13801 , n13802 );
and ( n13978 , n13651 , n13800 );
and ( n13979 , n13655 , n13707 );
and ( n13980 , n13707 , n13799 );
and ( n13981 , n13655 , n13799 );
or ( n13982 , n13979 , n13980 , n13981 );
and ( n13983 , n13712 , n13716 );
and ( n13984 , n13716 , n13798 );
and ( n13985 , n13712 , n13798 );
or ( n13986 , n13983 , n13984 , n13985 );
and ( n13987 , n13663 , n13667 );
and ( n13988 , n13667 , n13682 );
and ( n13989 , n13663 , n13682 );
or ( n13990 , n13987 , n13988 , n13989 );
and ( n13991 , n13688 , n13692 );
and ( n13992 , n13692 , n13705 );
and ( n13993 , n13688 , n13705 );
or ( n13994 , n13991 , n13992 , n13993 );
xor ( n13995 , n13990 , n13994 );
and ( n13996 , n13725 , n13739 );
and ( n13997 , n13739 , n13754 );
and ( n13998 , n13725 , n13754 );
or ( n13999 , n13996 , n13997 , n13998 );
and ( n14000 , n13767 , n13781 );
and ( n14001 , n13781 , n13796 );
and ( n14002 , n13767 , n13796 );
or ( n14003 , n14000 , n14001 , n14002 );
xor ( n14004 , n13999 , n14003 );
and ( n14005 , n13744 , n13748 );
and ( n14006 , n13748 , n13753 );
and ( n14007 , n13744 , n13753 );
or ( n14008 , n14005 , n14006 , n14007 );
and ( n14009 , n13771 , n13775 );
and ( n14010 , n13775 , n13780 );
and ( n14011 , n13771 , n13780 );
or ( n14012 , n14009 , n14010 , n14011 );
xor ( n14013 , n14008 , n14012 );
and ( n14014 , n13786 , n13790 );
and ( n14015 , n13790 , n13795 );
and ( n14016 , n13786 , n13795 );
or ( n14017 , n14014 , n14015 , n14016 );
xor ( n14018 , n14013 , n14017 );
xor ( n14019 , n14004 , n14018 );
xor ( n14020 , n13995 , n14019 );
xor ( n14021 , n13986 , n14020 );
and ( n14022 , n13721 , n13755 );
and ( n14023 , n13755 , n13797 );
and ( n14024 , n13721 , n13797 );
or ( n14025 , n14022 , n14023 , n14024 );
and ( n14026 , n13659 , n13683 );
and ( n14027 , n13683 , n13706 );
and ( n14028 , n13659 , n13706 );
or ( n14029 , n14026 , n14027 , n14028 );
xor ( n14030 , n14025 , n14029 );
and ( n14031 , n13729 , n13733 );
and ( n14032 , n13733 , n13738 );
and ( n14033 , n13729 , n13738 );
or ( n14034 , n14031 , n14032 , n14033 );
and ( n14035 , n9139 , n8887 );
and ( n14036 , n9323 , n8701 );
nor ( n14037 , n14035 , n14036 );
xnor ( n14038 , n14037 , n8893 );
and ( n14039 , n8690 , n9311 );
and ( n14040 , n8913 , n9150 );
nor ( n14041 , n14039 , n14040 );
xnor ( n14042 , n14041 , n9317 );
xor ( n14043 , n14038 , n14042 );
and ( n14044 , n7049 , n12730 );
xor ( n14045 , n14043 , n14044 );
xor ( n14046 , n14034 , n14045 );
not ( n14047 , n7058 );
and ( n14048 , n12339 , n7215 );
and ( n14049 , n12724 , n7136 );
nor ( n14050 , n14048 , n14049 );
xnor ( n14051 , n14050 , n7205 );
xor ( n14052 , n14047 , n14051 );
and ( n14053 , n11133 , n7609 );
and ( n14054 , n11384 , n7505 );
nor ( n14055 , n14053 , n14054 );
xnor ( n14056 , n14055 , n7615 );
xor ( n14057 , n14052 , n14056 );
xor ( n14058 , n14046 , n14057 );
and ( n14059 , n11699 , n7400 );
and ( n14060 , n12010 , n7303 );
nor ( n14061 , n14059 , n14060 );
xnor ( n14062 , n14061 , n7381 );
and ( n14063 , n10090 , n8209 );
and ( n14064 , n10331 , n8039 );
nor ( n14065 , n14063 , n14064 );
xnor ( n14066 , n14065 , n8165 );
xor ( n14067 , n14062 , n14066 );
and ( n14068 , n7730 , n10907 );
and ( n14069 , n7891 , n10543 );
nor ( n14070 , n14068 , n14069 );
xnor ( n14071 , n14070 , n10807 );
xor ( n14072 , n14067 , n14071 );
and ( n14073 , n10548 , n7873 );
and ( n14074 , n10837 , n7762 );
nor ( n14075 , n14073 , n14074 );
xnor ( n14076 , n14075 , n7863 );
and ( n14077 , n8339 , n9795 );
and ( n14078 , n8548 , n9560 );
nor ( n14079 , n14077 , n14078 );
xnor ( n14080 , n14079 , n9801 );
xor ( n14081 , n14076 , n14080 );
and ( n14082 , n8045 , n10342 );
and ( n14083 , n8156 , n10084 );
nor ( n14084 , n14082 , n14083 );
xnor ( n14085 , n14084 , n10291 );
xor ( n14086 , n14081 , n14085 );
xor ( n14087 , n14072 , n14086 );
and ( n14088 , n9549 , n8511 );
and ( n14089 , n9839 , n8350 );
nor ( n14090 , n14088 , n14089 );
xnor ( n14091 , n14090 , n8517 );
and ( n14092 , n7494 , n11411 );
and ( n14093 , n7596 , n11159 );
nor ( n14094 , n14092 , n14093 );
xnor ( n14095 , n14094 , n11417 );
xor ( n14096 , n14091 , n14095 );
and ( n14097 , n7292 , n12029 );
and ( n14098 , n7372 , n11739 );
nor ( n14099 , n14097 , n14098 );
xnor ( n14100 , n14099 , n12019 );
xor ( n14101 , n14096 , n14100 );
xor ( n14102 , n14087 , n14101 );
xor ( n14103 , n14058 , n14102 );
and ( n14104 , n13672 , n13676 );
and ( n14105 , n13676 , n13681 );
and ( n14106 , n13672 , n13681 );
or ( n14107 , n14104 , n14105 , n14106 );
and ( n14108 , n13697 , n13699 );
and ( n14109 , n13699 , n13704 );
and ( n14110 , n13697 , n13704 );
or ( n14111 , n14108 , n14109 , n14110 );
xor ( n14112 , n14107 , n14111 );
and ( n14113 , n13760 , n13764 );
and ( n14114 , n13764 , n13766 );
and ( n14115 , n13760 , n13766 );
or ( n14116 , n14113 , n14114 , n14115 );
buf ( n14117 , n13703 );
xor ( n14118 , n14116 , n14117 );
and ( n14119 , n7125 , n12782 );
and ( n14120 , n7196 , n12350 );
nor ( n14121 , n14119 , n14120 );
xnor ( n14122 , n14121 , n12733 );
xor ( n14123 , n14118 , n14122 );
xor ( n14124 , n14112 , n14123 );
xor ( n14125 , n14103 , n14124 );
xor ( n14126 , n14030 , n14125 );
xor ( n14127 , n14021 , n14126 );
xor ( n14128 , n13982 , n14127 );
xor ( n14129 , n13978 , n14128 );
xor ( n14130 , n13977 , n14129 );
and ( n14131 , n13647 , n13803 );
and ( n14132 , n13804 , n13807 );
or ( n14133 , n14131 , n14132 );
xor ( n14134 , n14130 , n14133 );
buf ( n14135 , n14134 );
and ( n14136 , n13964 , n13965 );
and ( n14137 , n13814 , n13963 );
and ( n14138 , n13818 , n13870 );
and ( n14139 , n13870 , n13962 );
and ( n14140 , n13818 , n13962 );
or ( n14141 , n14138 , n14139 , n14140 );
and ( n14142 , n13875 , n13879 );
and ( n14143 , n13879 , n13961 );
and ( n14144 , n13875 , n13961 );
or ( n14145 , n14142 , n14143 , n14144 );
and ( n14146 , n13826 , n13830 );
and ( n14147 , n13830 , n13845 );
and ( n14148 , n13826 , n13845 );
or ( n14149 , n14146 , n14147 , n14148 );
and ( n14150 , n13851 , n13855 );
and ( n14151 , n13855 , n13868 );
and ( n14152 , n13851 , n13868 );
or ( n14153 , n14150 , n14151 , n14152 );
xor ( n14154 , n14149 , n14153 );
and ( n14155 , n13888 , n13902 );
and ( n14156 , n13902 , n13917 );
and ( n14157 , n13888 , n13917 );
or ( n14158 , n14155 , n14156 , n14157 );
and ( n14159 , n13930 , n13944 );
and ( n14160 , n13944 , n13959 );
and ( n14161 , n13930 , n13959 );
or ( n14162 , n14159 , n14160 , n14161 );
xor ( n14163 , n14158 , n14162 );
and ( n14164 , n13907 , n13911 );
and ( n14165 , n13911 , n13916 );
and ( n14166 , n13907 , n13916 );
or ( n14167 , n14164 , n14165 , n14166 );
and ( n14168 , n13934 , n13938 );
and ( n14169 , n13938 , n13943 );
and ( n14170 , n13934 , n13943 );
or ( n14171 , n14168 , n14169 , n14170 );
xor ( n14172 , n14167 , n14171 );
and ( n14173 , n13949 , n13953 );
and ( n14174 , n13953 , n13958 );
and ( n14175 , n13949 , n13958 );
or ( n14176 , n14173 , n14174 , n14175 );
xor ( n14177 , n14172 , n14176 );
xor ( n14178 , n14163 , n14177 );
xor ( n14179 , n14154 , n14178 );
xor ( n14180 , n14145 , n14179 );
and ( n14181 , n13884 , n13918 );
and ( n14182 , n13918 , n13960 );
and ( n14183 , n13884 , n13960 );
or ( n14184 , n14181 , n14182 , n14183 );
and ( n14185 , n13822 , n13846 );
and ( n14186 , n13846 , n13869 );
and ( n14187 , n13822 , n13869 );
or ( n14188 , n14185 , n14186 , n14187 );
xor ( n14189 , n14184 , n14188 );
and ( n14190 , n13892 , n13896 );
and ( n14191 , n13896 , n13901 );
and ( n14192 , n13892 , n13901 );
or ( n14193 , n14190 , n14191 , n14192 );
and ( n14194 , n9240 , n8992 );
and ( n14195 , n9438 , n8792 );
nor ( n14196 , n14194 , n14195 );
xnor ( n14197 , n14196 , n8998 );
and ( n14198 , n8781 , n9426 );
and ( n14199 , n9018 , n9251 );
nor ( n14200 , n14198 , n14199 );
xnor ( n14201 , n14200 , n9432 );
xor ( n14202 , n14197 , n14201 );
and ( n14203 , n7084 , n12905 );
xor ( n14204 , n14202 , n14203 );
xor ( n14205 , n14193 , n14204 );
not ( n14206 , n7093 );
and ( n14207 , n12500 , n7260 );
and ( n14208 , n12899 , n7167 );
nor ( n14209 , n14207 , n14208 );
xnor ( n14210 , n14209 , n7250 );
xor ( n14211 , n14206 , n14210 );
and ( n14212 , n11274 , n7674 );
and ( n14213 , n11539 , n7556 );
nor ( n14214 , n14212 , n14213 );
xnor ( n14215 , n14214 , n7680 );
xor ( n14216 , n14211 , n14215 );
xor ( n14217 , n14205 , n14216 );
and ( n14218 , n11850 , n7455 );
and ( n14219 , n12175 , n7344 );
nor ( n14220 , n14218 , n14219 );
xnor ( n14221 , n14220 , n7436 );
and ( n14222 , n10211 , n8294 );
and ( n14223 , n10466 , n8110 );
nor ( n14224 , n14222 , n14223 );
xnor ( n14225 , n14224 , n8250 );
xor ( n14226 , n14221 , n14225 );
and ( n14227 , n7791 , n11052 );
and ( n14228 , n7966 , n10674 );
nor ( n14229 , n14227 , n14228 );
xnor ( n14230 , n14229 , n10952 );
xor ( n14231 , n14226 , n14230 );
and ( n14232 , n10679 , n7948 );
and ( n14233 , n10982 , n7823 );
nor ( n14234 , n14232 , n14233 );
xnor ( n14235 , n14234 , n7938 );
and ( n14236 , n8420 , n9920 );
and ( n14237 , n8643 , n9671 );
nor ( n14238 , n14236 , n14237 );
xnor ( n14239 , n14238 , n9926 );
xor ( n14240 , n14235 , n14239 );
and ( n14241 , n8116 , n10477 );
and ( n14242 , n8241 , n10205 );
nor ( n14243 , n14241 , n14242 );
xnor ( n14244 , n14243 , n10426 );
xor ( n14245 , n14240 , n14244 );
xor ( n14246 , n14231 , n14245 );
and ( n14247 , n9660 , n8606 );
and ( n14248 , n9964 , n8431 );
nor ( n14249 , n14247 , n14248 );
xnor ( n14250 , n14249 , n8612 );
and ( n14251 , n7545 , n11566 );
and ( n14252 , n7661 , n11300 );
nor ( n14253 , n14251 , n14252 );
xnor ( n14254 , n14253 , n11572 );
xor ( n14255 , n14250 , n14254 );
and ( n14256 , n7333 , n12194 );
and ( n14257 , n7427 , n11890 );
nor ( n14258 , n14256 , n14257 );
xnor ( n14259 , n14258 , n12184 );
xor ( n14260 , n14255 , n14259 );
xor ( n14261 , n14246 , n14260 );
xor ( n14262 , n14217 , n14261 );
and ( n14263 , n13835 , n13839 );
and ( n14264 , n13839 , n13844 );
and ( n14265 , n13835 , n13844 );
or ( n14266 , n14263 , n14264 , n14265 );
and ( n14267 , n13860 , n13862 );
and ( n14268 , n13862 , n13867 );
and ( n14269 , n13860 , n13867 );
or ( n14270 , n14267 , n14268 , n14269 );
xor ( n14271 , n14266 , n14270 );
and ( n14272 , n13923 , n13927 );
and ( n14273 , n13927 , n13929 );
and ( n14274 , n13923 , n13929 );
or ( n14275 , n14272 , n14273 , n14274 );
buf ( n14276 , n13866 );
xor ( n14277 , n14275 , n14276 );
and ( n14278 , n7156 , n12957 );
and ( n14279 , n7241 , n12511 );
nor ( n14280 , n14278 , n14279 );
xnor ( n14281 , n14280 , n12908 );
xor ( n14282 , n14277 , n14281 );
xor ( n14283 , n14271 , n14282 );
xor ( n14284 , n14262 , n14283 );
xor ( n14285 , n14189 , n14284 );
xor ( n14286 , n14180 , n14285 );
xor ( n14287 , n14141 , n14286 );
xor ( n14288 , n14137 , n14287 );
xor ( n14289 , n14136 , n14288 );
and ( n14290 , n13810 , n13966 );
and ( n14291 , n13967 , n13970 );
or ( n14292 , n14290 , n14291 );
xor ( n14293 , n14289 , n14292 );
buf ( n14294 , n14293 );
not ( n14295 , n831 );
and ( n14296 , n14295 , n14135 );
and ( n14297 , n14294 , n831 );
or ( n14298 , n14296 , n14297 );
and ( n14299 , n13978 , n14128 );
and ( n14300 , n13986 , n14020 );
and ( n14301 , n14020 , n14126 );
and ( n14302 , n13986 , n14126 );
or ( n14303 , n14300 , n14301 , n14302 );
and ( n14304 , n14025 , n14029 );
and ( n14305 , n14029 , n14125 );
and ( n14306 , n14025 , n14125 );
or ( n14307 , n14304 , n14305 , n14306 );
and ( n14308 , n13999 , n14003 );
and ( n14309 , n14003 , n14018 );
and ( n14310 , n13999 , n14018 );
or ( n14311 , n14308 , n14309 , n14310 );
and ( n14312 , n14008 , n14012 );
and ( n14313 , n14012 , n14017 );
and ( n14314 , n14008 , n14017 );
or ( n14315 , n14312 , n14313 , n14314 );
and ( n14316 , n14116 , n14117 );
and ( n14317 , n14117 , n14122 );
and ( n14318 , n14116 , n14122 );
or ( n14319 , n14316 , n14317 , n14318 );
xor ( n14320 , n14315 , n14319 );
and ( n14321 , n12724 , n7215 );
not ( n14322 , n14321 );
xnor ( n14323 , n14322 , n7205 );
not ( n14324 , n14323 );
and ( n14325 , n7196 , n12782 );
and ( n14326 , n7292 , n12350 );
nor ( n14327 , n14325 , n14326 );
xnor ( n14328 , n14327 , n12733 );
xor ( n14329 , n14324 , n14328 );
and ( n14330 , n7125 , n12730 );
xor ( n14331 , n14329 , n14330 );
xor ( n14332 , n14320 , n14331 );
xor ( n14333 , n14311 , n14332 );
and ( n14334 , n14034 , n14045 );
and ( n14335 , n14045 , n14057 );
and ( n14336 , n14034 , n14057 );
or ( n14337 , n14334 , n14335 , n14336 );
and ( n14338 , n14038 , n14042 );
and ( n14339 , n14042 , n14044 );
and ( n14340 , n14038 , n14044 );
or ( n14341 , n14338 , n14339 , n14340 );
and ( n14342 , n14047 , n14051 );
and ( n14343 , n14051 , n14056 );
and ( n14344 , n14047 , n14056 );
or ( n14345 , n14342 , n14343 , n14344 );
xor ( n14346 , n14341 , n14345 );
and ( n14347 , n14076 , n14080 );
and ( n14348 , n14080 , n14085 );
and ( n14349 , n14076 , n14085 );
or ( n14350 , n14347 , n14348 , n14349 );
xor ( n14351 , n14346 , n14350 );
xor ( n14352 , n14337 , n14351 );
and ( n14353 , n14062 , n14066 );
and ( n14354 , n14066 , n14071 );
and ( n14355 , n14062 , n14071 );
or ( n14356 , n14353 , n14354 , n14355 );
and ( n14357 , n14091 , n14095 );
and ( n14358 , n14095 , n14100 );
and ( n14359 , n14091 , n14100 );
or ( n14360 , n14357 , n14358 , n14359 );
xor ( n14361 , n14356 , n14360 );
and ( n14362 , n12010 , n7400 );
and ( n14363 , n12339 , n7303 );
nor ( n14364 , n14362 , n14363 );
xnor ( n14365 , n14364 , n7381 );
and ( n14366 , n10837 , n7873 );
and ( n14367 , n11133 , n7762 );
nor ( n14368 , n14366 , n14367 );
xnor ( n14369 , n14368 , n7863 );
xor ( n14370 , n14365 , n14369 );
and ( n14371 , n8913 , n9311 );
and ( n14372 , n9139 , n9150 );
nor ( n14373 , n14371 , n14372 );
xnor ( n14374 , n14373 , n9317 );
xor ( n14375 , n14370 , n14374 );
xor ( n14376 , n14361 , n14375 );
xor ( n14377 , n14352 , n14376 );
xor ( n14378 , n14333 , n14377 );
xor ( n14379 , n14307 , n14378 );
and ( n14380 , n13990 , n13994 );
and ( n14381 , n13994 , n14019 );
and ( n14382 , n13990 , n14019 );
or ( n14383 , n14380 , n14381 , n14382 );
and ( n14384 , n14058 , n14102 );
and ( n14385 , n14102 , n14124 );
and ( n14386 , n14058 , n14124 );
or ( n14387 , n14384 , n14385 , n14386 );
xor ( n14388 , n14383 , n14387 );
and ( n14389 , n14072 , n14086 );
and ( n14390 , n14086 , n14101 );
and ( n14391 , n14072 , n14101 );
or ( n14392 , n14389 , n14390 , n14391 );
and ( n14393 , n14107 , n14111 );
and ( n14394 , n14111 , n14123 );
and ( n14395 , n14107 , n14123 );
or ( n14396 , n14393 , n14394 , n14395 );
xor ( n14397 , n14392 , n14396 );
and ( n14398 , n9323 , n8887 );
and ( n14399 , n9549 , n8701 );
nor ( n14400 , n14398 , n14399 );
xnor ( n14401 , n14400 , n8893 );
and ( n14402 , n7596 , n11411 );
and ( n14403 , n7730 , n11159 );
nor ( n14404 , n14402 , n14403 );
xnor ( n14405 , n14404 , n11417 );
xor ( n14406 , n14401 , n14405 );
and ( n14407 , n7372 , n12029 );
and ( n14408 , n7494 , n11739 );
nor ( n14409 , n14407 , n14408 );
xnor ( n14410 , n14409 , n12019 );
xor ( n14411 , n14406 , n14410 );
and ( n14412 , n10331 , n8209 );
and ( n14413 , n10548 , n8039 );
nor ( n14414 , n14412 , n14413 );
xnor ( n14415 , n14414 , n8165 );
and ( n14416 , n8548 , n9795 );
and ( n14417 , n8690 , n9560 );
nor ( n14418 , n14416 , n14417 );
xnor ( n14419 , n14418 , n9801 );
xor ( n14420 , n14415 , n14419 );
and ( n14421 , n8156 , n10342 );
and ( n14422 , n8339 , n10084 );
nor ( n14423 , n14421 , n14422 );
xnor ( n14424 , n14423 , n10291 );
xor ( n14425 , n14420 , n14424 );
xor ( n14426 , n14411 , n14425 );
and ( n14427 , n11384 , n7609 );
and ( n14428 , n11699 , n7505 );
nor ( n14429 , n14427 , n14428 );
xnor ( n14430 , n14429 , n7615 );
and ( n14431 , n9839 , n8511 );
and ( n14432 , n10090 , n8350 );
nor ( n14433 , n14431 , n14432 );
xnor ( n14434 , n14433 , n8517 );
xor ( n14435 , n14430 , n14434 );
and ( n14436 , n7891 , n10907 );
and ( n14437 , n8045 , n10543 );
nor ( n14438 , n14436 , n14437 );
xnor ( n14439 , n14438 , n10807 );
xor ( n14440 , n14435 , n14439 );
xor ( n14441 , n14426 , n14440 );
xor ( n14442 , n14397 , n14441 );
xor ( n14443 , n14388 , n14442 );
xor ( n14444 , n14379 , n14443 );
xor ( n14445 , n14303 , n14444 );
and ( n14446 , n13982 , n14127 );
xor ( n14447 , n14445 , n14446 );
xor ( n14448 , n14299 , n14447 );
and ( n14449 , n13977 , n14129 );
and ( n14450 , n14130 , n14133 );
or ( n14451 , n14449 , n14450 );
xor ( n14452 , n14448 , n14451 );
buf ( n14453 , n14452 );
and ( n14454 , n14137 , n14287 );
and ( n14455 , n14145 , n14179 );
and ( n14456 , n14179 , n14285 );
and ( n14457 , n14145 , n14285 );
or ( n14458 , n14455 , n14456 , n14457 );
and ( n14459 , n14184 , n14188 );
and ( n14460 , n14188 , n14284 );
and ( n14461 , n14184 , n14284 );
or ( n14462 , n14459 , n14460 , n14461 );
and ( n14463 , n14158 , n14162 );
and ( n14464 , n14162 , n14177 );
and ( n14465 , n14158 , n14177 );
or ( n14466 , n14463 , n14464 , n14465 );
and ( n14467 , n14167 , n14171 );
and ( n14468 , n14171 , n14176 );
and ( n14469 , n14167 , n14176 );
or ( n14470 , n14467 , n14468 , n14469 );
and ( n14471 , n14275 , n14276 );
and ( n14472 , n14276 , n14281 );
and ( n14473 , n14275 , n14281 );
or ( n14474 , n14471 , n14472 , n14473 );
xor ( n14475 , n14470 , n14474 );
and ( n14476 , n12899 , n7260 );
not ( n14477 , n14476 );
xnor ( n14478 , n14477 , n7250 );
not ( n14479 , n14478 );
and ( n14480 , n7241 , n12957 );
and ( n14481 , n7333 , n12511 );
nor ( n14482 , n14480 , n14481 );
xnor ( n14483 , n14482 , n12908 );
xor ( n14484 , n14479 , n14483 );
and ( n14485 , n7156 , n12905 );
xor ( n14486 , n14484 , n14485 );
xor ( n14487 , n14475 , n14486 );
xor ( n14488 , n14466 , n14487 );
and ( n14489 , n14193 , n14204 );
and ( n14490 , n14204 , n14216 );
and ( n14491 , n14193 , n14216 );
or ( n14492 , n14489 , n14490 , n14491 );
and ( n14493 , n14197 , n14201 );
and ( n14494 , n14201 , n14203 );
and ( n14495 , n14197 , n14203 );
or ( n14496 , n14493 , n14494 , n14495 );
and ( n14497 , n14206 , n14210 );
and ( n14498 , n14210 , n14215 );
and ( n14499 , n14206 , n14215 );
or ( n14500 , n14497 , n14498 , n14499 );
xor ( n14501 , n14496 , n14500 );
and ( n14502 , n14235 , n14239 );
and ( n14503 , n14239 , n14244 );
and ( n14504 , n14235 , n14244 );
or ( n14505 , n14502 , n14503 , n14504 );
xor ( n14506 , n14501 , n14505 );
xor ( n14507 , n14492 , n14506 );
and ( n14508 , n14221 , n14225 );
and ( n14509 , n14225 , n14230 );
and ( n14510 , n14221 , n14230 );
or ( n14511 , n14508 , n14509 , n14510 );
and ( n14512 , n14250 , n14254 );
and ( n14513 , n14254 , n14259 );
and ( n14514 , n14250 , n14259 );
or ( n14515 , n14512 , n14513 , n14514 );
xor ( n14516 , n14511 , n14515 );
and ( n14517 , n12175 , n7455 );
and ( n14518 , n12500 , n7344 );
nor ( n14519 , n14517 , n14518 );
xnor ( n14520 , n14519 , n7436 );
and ( n14521 , n10982 , n7948 );
and ( n14522 , n11274 , n7823 );
nor ( n14523 , n14521 , n14522 );
xnor ( n14524 , n14523 , n7938 );
xor ( n14525 , n14520 , n14524 );
and ( n14526 , n9018 , n9426 );
and ( n14527 , n9240 , n9251 );
nor ( n14528 , n14526 , n14527 );
xnor ( n14529 , n14528 , n9432 );
xor ( n14530 , n14525 , n14529 );
xor ( n14531 , n14516 , n14530 );
xor ( n14532 , n14507 , n14531 );
xor ( n14533 , n14488 , n14532 );
xor ( n14534 , n14462 , n14533 );
and ( n14535 , n14149 , n14153 );
and ( n14536 , n14153 , n14178 );
and ( n14537 , n14149 , n14178 );
or ( n14538 , n14535 , n14536 , n14537 );
and ( n14539 , n14217 , n14261 );
and ( n14540 , n14261 , n14283 );
and ( n14541 , n14217 , n14283 );
or ( n14542 , n14539 , n14540 , n14541 );
xor ( n14543 , n14538 , n14542 );
and ( n14544 , n14231 , n14245 );
and ( n14545 , n14245 , n14260 );
and ( n14546 , n14231 , n14260 );
or ( n14547 , n14544 , n14545 , n14546 );
and ( n14548 , n14266 , n14270 );
and ( n14549 , n14270 , n14282 );
and ( n14550 , n14266 , n14282 );
or ( n14551 , n14548 , n14549 , n14550 );
xor ( n14552 , n14547 , n14551 );
and ( n14553 , n9438 , n8992 );
and ( n14554 , n9660 , n8792 );
nor ( n14555 , n14553 , n14554 );
xnor ( n14556 , n14555 , n8998 );
and ( n14557 , n7661 , n11566 );
and ( n14558 , n7791 , n11300 );
nor ( n14559 , n14557 , n14558 );
xnor ( n14560 , n14559 , n11572 );
xor ( n14561 , n14556 , n14560 );
and ( n14562 , n7427 , n12194 );
and ( n14563 , n7545 , n11890 );
nor ( n14564 , n14562 , n14563 );
xnor ( n14565 , n14564 , n12184 );
xor ( n14566 , n14561 , n14565 );
and ( n14567 , n10466 , n8294 );
and ( n14568 , n10679 , n8110 );
nor ( n14569 , n14567 , n14568 );
xnor ( n14570 , n14569 , n8250 );
and ( n14571 , n8643 , n9920 );
and ( n14572 , n8781 , n9671 );
nor ( n14573 , n14571 , n14572 );
xnor ( n14574 , n14573 , n9926 );
xor ( n14575 , n14570 , n14574 );
and ( n14576 , n8241 , n10477 );
and ( n14577 , n8420 , n10205 );
nor ( n14578 , n14576 , n14577 );
xnor ( n14579 , n14578 , n10426 );
xor ( n14580 , n14575 , n14579 );
xor ( n14581 , n14566 , n14580 );
and ( n14582 , n11539 , n7674 );
and ( n14583 , n11850 , n7556 );
nor ( n14584 , n14582 , n14583 );
xnor ( n14585 , n14584 , n7680 );
and ( n14586 , n9964 , n8606 );
and ( n14587 , n10211 , n8431 );
nor ( n14588 , n14586 , n14587 );
xnor ( n14589 , n14588 , n8612 );
xor ( n14590 , n14585 , n14589 );
and ( n14591 , n7966 , n11052 );
and ( n14592 , n8116 , n10674 );
nor ( n14593 , n14591 , n14592 );
xnor ( n14594 , n14593 , n10952 );
xor ( n14595 , n14590 , n14594 );
xor ( n14596 , n14581 , n14595 );
xor ( n14597 , n14552 , n14596 );
xor ( n14598 , n14543 , n14597 );
xor ( n14599 , n14534 , n14598 );
xor ( n14600 , n14458 , n14599 );
and ( n14601 , n14141 , n14286 );
xor ( n14602 , n14600 , n14601 );
xor ( n14603 , n14454 , n14602 );
and ( n14604 , n14136 , n14288 );
and ( n14605 , n14289 , n14292 );
or ( n14606 , n14604 , n14605 );
xor ( n14607 , n14603 , n14606 );
buf ( n14608 , n14607 );
not ( n14609 , n831 );
and ( n14610 , n14609 , n14453 );
and ( n14611 , n14608 , n831 );
or ( n14612 , n14610 , n14611 );
and ( n14613 , n14445 , n14446 );
and ( n14614 , n14307 , n14378 );
and ( n14615 , n14378 , n14443 );
and ( n14616 , n14307 , n14443 );
or ( n14617 , n14614 , n14615 , n14616 );
and ( n14618 , n14383 , n14387 );
and ( n14619 , n14387 , n14442 );
and ( n14620 , n14383 , n14442 );
or ( n14621 , n14618 , n14619 , n14620 );
and ( n14622 , n14315 , n14319 );
and ( n14623 , n14319 , n14331 );
and ( n14624 , n14315 , n14331 );
or ( n14625 , n14622 , n14623 , n14624 );
and ( n14626 , n14337 , n14351 );
and ( n14627 , n14351 , n14376 );
and ( n14628 , n14337 , n14376 );
or ( n14629 , n14626 , n14627 , n14628 );
xor ( n14630 , n14625 , n14629 );
and ( n14631 , n14356 , n14360 );
and ( n14632 , n14360 , n14375 );
and ( n14633 , n14356 , n14375 );
or ( n14634 , n14631 , n14632 , n14633 );
and ( n14635 , n14365 , n14369 );
and ( n14636 , n14369 , n14374 );
and ( n14637 , n14365 , n14374 );
or ( n14638 , n14635 , n14636 , n14637 );
and ( n14639 , n14415 , n14419 );
and ( n14640 , n14419 , n14424 );
and ( n14641 , n14415 , n14424 );
or ( n14642 , n14639 , n14640 , n14641 );
xor ( n14643 , n14638 , n14642 );
buf ( n14644 , n14323 );
xor ( n14645 , n14643 , n14644 );
xor ( n14646 , n14634 , n14645 );
and ( n14647 , n14401 , n14405 );
and ( n14648 , n14405 , n14410 );
and ( n14649 , n14401 , n14410 );
or ( n14650 , n14647 , n14648 , n14649 );
and ( n14651 , n14430 , n14434 );
and ( n14652 , n14434 , n14439 );
and ( n14653 , n14430 , n14439 );
or ( n14654 , n14651 , n14652 , n14653 );
xor ( n14655 , n14650 , n14654 );
and ( n14656 , n10548 , n8209 );
and ( n14657 , n10837 , n8039 );
nor ( n14658 , n14656 , n14657 );
xnor ( n14659 , n14658 , n8165 );
and ( n14660 , n9139 , n9311 );
and ( n14661 , n9323 , n9150 );
nor ( n14662 , n14660 , n14661 );
xnor ( n14663 , n14662 , n9317 );
xor ( n14664 , n14659 , n14663 );
and ( n14665 , n8690 , n9795 );
and ( n14666 , n8913 , n9560 );
nor ( n14667 , n14665 , n14666 );
xnor ( n14668 , n14667 , n9801 );
xor ( n14669 , n14664 , n14668 );
xor ( n14670 , n14655 , n14669 );
xor ( n14671 , n14646 , n14670 );
xor ( n14672 , n14630 , n14671 );
xor ( n14673 , n14621 , n14672 );
and ( n14674 , n14392 , n14396 );
and ( n14675 , n14396 , n14441 );
and ( n14676 , n14392 , n14441 );
or ( n14677 , n14674 , n14675 , n14676 );
and ( n14678 , n14311 , n14332 );
and ( n14679 , n14332 , n14377 );
and ( n14680 , n14311 , n14377 );
or ( n14681 , n14678 , n14679 , n14680 );
xor ( n14682 , n14677 , n14681 );
and ( n14683 , n14411 , n14425 );
and ( n14684 , n14425 , n14440 );
and ( n14685 , n14411 , n14440 );
or ( n14686 , n14683 , n14684 , n14685 );
and ( n14687 , n10090 , n8511 );
and ( n14688 , n10331 , n8350 );
nor ( n14689 , n14687 , n14688 );
xnor ( n14690 , n14689 , n8517 );
and ( n14691 , n7730 , n11411 );
and ( n14692 , n7891 , n11159 );
nor ( n14693 , n14691 , n14692 );
xnor ( n14694 , n14693 , n11417 );
xor ( n14695 , n14690 , n14694 );
and ( n14696 , n7494 , n12029 );
and ( n14697 , n7596 , n11739 );
nor ( n14698 , n14696 , n14697 );
xnor ( n14699 , n14698 , n12019 );
xor ( n14700 , n14695 , n14699 );
and ( n14701 , n9549 , n8887 );
and ( n14702 , n9839 , n8701 );
nor ( n14703 , n14701 , n14702 );
xnor ( n14704 , n14703 , n8893 );
and ( n14705 , n7292 , n12782 );
and ( n14706 , n7372 , n12350 );
nor ( n14707 , n14705 , n14706 );
xnor ( n14708 , n14707 , n12733 );
xor ( n14709 , n14704 , n14708 );
and ( n14710 , n7196 , n12730 );
xor ( n14711 , n14709 , n14710 );
xor ( n14712 , n14700 , n14711 );
not ( n14713 , n7205 );
and ( n14714 , n12339 , n7400 );
and ( n14715 , n12724 , n7303 );
nor ( n14716 , n14714 , n14715 );
xnor ( n14717 , n14716 , n7381 );
xor ( n14718 , n14713 , n14717 );
and ( n14719 , n11133 , n7873 );
and ( n14720 , n11384 , n7762 );
nor ( n14721 , n14719 , n14720 );
xnor ( n14722 , n14721 , n7863 );
xor ( n14723 , n14718 , n14722 );
xor ( n14724 , n14712 , n14723 );
xor ( n14725 , n14686 , n14724 );
and ( n14726 , n14341 , n14345 );
and ( n14727 , n14345 , n14350 );
and ( n14728 , n14341 , n14350 );
or ( n14729 , n14726 , n14727 , n14728 );
and ( n14730 , n14324 , n14328 );
and ( n14731 , n14328 , n14330 );
and ( n14732 , n14324 , n14330 );
or ( n14733 , n14730 , n14731 , n14732 );
xor ( n14734 , n14729 , n14733 );
and ( n14735 , n11699 , n7609 );
and ( n14736 , n12010 , n7505 );
nor ( n14737 , n14735 , n14736 );
xnor ( n14738 , n14737 , n7615 );
and ( n14739 , n8339 , n10342 );
and ( n14740 , n8548 , n10084 );
nor ( n14741 , n14739 , n14740 );
xnor ( n14742 , n14741 , n10291 );
xor ( n14743 , n14738 , n14742 );
and ( n14744 , n8045 , n10907 );
and ( n14745 , n8156 , n10543 );
nor ( n14746 , n14744 , n14745 );
xnor ( n14747 , n14746 , n10807 );
xor ( n14748 , n14743 , n14747 );
xor ( n14749 , n14734 , n14748 );
xor ( n14750 , n14725 , n14749 );
xor ( n14751 , n14682 , n14750 );
xor ( n14752 , n14673 , n14751 );
xor ( n14753 , n14617 , n14752 );
and ( n14754 , n14303 , n14444 );
xor ( n14755 , n14753 , n14754 );
xor ( n14756 , n14613 , n14755 );
and ( n14757 , n14299 , n14447 );
and ( n14758 , n14448 , n14451 );
or ( n14759 , n14757 , n14758 );
xor ( n14760 , n14756 , n14759 );
buf ( n14761 , n14760 );
and ( n14762 , n14600 , n14601 );
and ( n14763 , n14462 , n14533 );
and ( n14764 , n14533 , n14598 );
and ( n14765 , n14462 , n14598 );
or ( n14766 , n14763 , n14764 , n14765 );
and ( n14767 , n14538 , n14542 );
and ( n14768 , n14542 , n14597 );
and ( n14769 , n14538 , n14597 );
or ( n14770 , n14767 , n14768 , n14769 );
and ( n14771 , n14470 , n14474 );
and ( n14772 , n14474 , n14486 );
and ( n14773 , n14470 , n14486 );
or ( n14774 , n14771 , n14772 , n14773 );
and ( n14775 , n14492 , n14506 );
and ( n14776 , n14506 , n14531 );
and ( n14777 , n14492 , n14531 );
or ( n14778 , n14775 , n14776 , n14777 );
xor ( n14779 , n14774 , n14778 );
and ( n14780 , n14511 , n14515 );
and ( n14781 , n14515 , n14530 );
and ( n14782 , n14511 , n14530 );
or ( n14783 , n14780 , n14781 , n14782 );
and ( n14784 , n14520 , n14524 );
and ( n14785 , n14524 , n14529 );
and ( n14786 , n14520 , n14529 );
or ( n14787 , n14784 , n14785 , n14786 );
and ( n14788 , n14570 , n14574 );
and ( n14789 , n14574 , n14579 );
and ( n14790 , n14570 , n14579 );
or ( n14791 , n14788 , n14789 , n14790 );
xor ( n14792 , n14787 , n14791 );
buf ( n14793 , n14478 );
xor ( n14794 , n14792 , n14793 );
xor ( n14795 , n14783 , n14794 );
and ( n14796 , n14556 , n14560 );
and ( n14797 , n14560 , n14565 );
and ( n14798 , n14556 , n14565 );
or ( n14799 , n14796 , n14797 , n14798 );
and ( n14800 , n14585 , n14589 );
and ( n14801 , n14589 , n14594 );
and ( n14802 , n14585 , n14594 );
or ( n14803 , n14800 , n14801 , n14802 );
xor ( n14804 , n14799 , n14803 );
and ( n14805 , n10679 , n8294 );
and ( n14806 , n10982 , n8110 );
nor ( n14807 , n14805 , n14806 );
xnor ( n14808 , n14807 , n8250 );
and ( n14809 , n9240 , n9426 );
and ( n14810 , n9438 , n9251 );
nor ( n14811 , n14809 , n14810 );
xnor ( n14812 , n14811 , n9432 );
xor ( n14813 , n14808 , n14812 );
and ( n14814 , n8781 , n9920 );
and ( n14815 , n9018 , n9671 );
nor ( n14816 , n14814 , n14815 );
xnor ( n14817 , n14816 , n9926 );
xor ( n14818 , n14813 , n14817 );
xor ( n14819 , n14804 , n14818 );
xor ( n14820 , n14795 , n14819 );
xor ( n14821 , n14779 , n14820 );
xor ( n14822 , n14770 , n14821 );
and ( n14823 , n14547 , n14551 );
and ( n14824 , n14551 , n14596 );
and ( n14825 , n14547 , n14596 );
or ( n14826 , n14823 , n14824 , n14825 );
and ( n14827 , n14466 , n14487 );
and ( n14828 , n14487 , n14532 );
and ( n14829 , n14466 , n14532 );
or ( n14830 , n14827 , n14828 , n14829 );
xor ( n14831 , n14826 , n14830 );
and ( n14832 , n14566 , n14580 );
and ( n14833 , n14580 , n14595 );
and ( n14834 , n14566 , n14595 );
or ( n14835 , n14832 , n14833 , n14834 );
and ( n14836 , n10211 , n8606 );
and ( n14837 , n10466 , n8431 );
nor ( n14838 , n14836 , n14837 );
xnor ( n14839 , n14838 , n8612 );
and ( n14840 , n7791 , n11566 );
and ( n14841 , n7966 , n11300 );
nor ( n14842 , n14840 , n14841 );
xnor ( n14843 , n14842 , n11572 );
xor ( n14844 , n14839 , n14843 );
and ( n14845 , n7545 , n12194 );
and ( n14846 , n7661 , n11890 );
nor ( n14847 , n14845 , n14846 );
xnor ( n14848 , n14847 , n12184 );
xor ( n14849 , n14844 , n14848 );
and ( n14850 , n9660 , n8992 );
and ( n14851 , n9964 , n8792 );
nor ( n14852 , n14850 , n14851 );
xnor ( n14853 , n14852 , n8998 );
and ( n14854 , n7333 , n12957 );
and ( n14855 , n7427 , n12511 );
nor ( n14856 , n14854 , n14855 );
xnor ( n14857 , n14856 , n12908 );
xor ( n14858 , n14853 , n14857 );
and ( n14859 , n7241 , n12905 );
xor ( n14860 , n14858 , n14859 );
xor ( n14861 , n14849 , n14860 );
not ( n14862 , n7250 );
and ( n14863 , n12500 , n7455 );
and ( n14864 , n12899 , n7344 );
nor ( n14865 , n14863 , n14864 );
xnor ( n14866 , n14865 , n7436 );
xor ( n14867 , n14862 , n14866 );
and ( n14868 , n11274 , n7948 );
and ( n14869 , n11539 , n7823 );
nor ( n14870 , n14868 , n14869 );
xnor ( n14871 , n14870 , n7938 );
xor ( n14872 , n14867 , n14871 );
xor ( n14873 , n14861 , n14872 );
xor ( n14874 , n14835 , n14873 );
and ( n14875 , n14496 , n14500 );
and ( n14876 , n14500 , n14505 );
and ( n14877 , n14496 , n14505 );
or ( n14878 , n14875 , n14876 , n14877 );
and ( n14879 , n14479 , n14483 );
and ( n14880 , n14483 , n14485 );
and ( n14881 , n14479 , n14485 );
or ( n14882 , n14879 , n14880 , n14881 );
xor ( n14883 , n14878 , n14882 );
and ( n14884 , n11850 , n7674 );
and ( n14885 , n12175 , n7556 );
nor ( n14886 , n14884 , n14885 );
xnor ( n14887 , n14886 , n7680 );
and ( n14888 , n8420 , n10477 );
and ( n14889 , n8643 , n10205 );
nor ( n14890 , n14888 , n14889 );
xnor ( n14891 , n14890 , n10426 );
xor ( n14892 , n14887 , n14891 );
and ( n14893 , n8116 , n11052 );
and ( n14894 , n8241 , n10674 );
nor ( n14895 , n14893 , n14894 );
xnor ( n14896 , n14895 , n10952 );
xor ( n14897 , n14892 , n14896 );
xor ( n14898 , n14883 , n14897 );
xor ( n14899 , n14874 , n14898 );
xor ( n14900 , n14831 , n14899 );
xor ( n14901 , n14822 , n14900 );
xor ( n14902 , n14766 , n14901 );
and ( n14903 , n14458 , n14599 );
xor ( n14904 , n14902 , n14903 );
xor ( n14905 , n14762 , n14904 );
and ( n14906 , n14454 , n14602 );
and ( n14907 , n14603 , n14606 );
or ( n14908 , n14906 , n14907 );
xor ( n14909 , n14905 , n14908 );
buf ( n14910 , n14909 );
not ( n14911 , n831 );
and ( n14912 , n14911 , n14761 );
and ( n14913 , n14910 , n831 );
or ( n14914 , n14912 , n14913 );
and ( n14915 , n14753 , n14754 );
and ( n14916 , n14621 , n14672 );
and ( n14917 , n14672 , n14751 );
and ( n14918 , n14621 , n14751 );
or ( n14919 , n14916 , n14917 , n14918 );
and ( n14920 , n14625 , n14629 );
and ( n14921 , n14629 , n14671 );
and ( n14922 , n14625 , n14671 );
or ( n14923 , n14920 , n14921 , n14922 );
and ( n14924 , n14677 , n14681 );
and ( n14925 , n14681 , n14750 );
and ( n14926 , n14677 , n14750 );
or ( n14927 , n14924 , n14925 , n14926 );
xor ( n14928 , n14923 , n14927 );
and ( n14929 , n14686 , n14724 );
and ( n14930 , n14724 , n14749 );
and ( n14931 , n14686 , n14749 );
or ( n14932 , n14929 , n14930 , n14931 );
and ( n14933 , n14700 , n14711 );
and ( n14934 , n14711 , n14723 );
and ( n14935 , n14700 , n14723 );
or ( n14936 , n14933 , n14934 , n14935 );
and ( n14937 , n14729 , n14733 );
and ( n14938 , n14733 , n14748 );
and ( n14939 , n14729 , n14748 );
or ( n14940 , n14937 , n14938 , n14939 );
xor ( n14941 , n14936 , n14940 );
and ( n14942 , n14704 , n14708 );
and ( n14943 , n14708 , n14710 );
and ( n14944 , n14704 , n14710 );
or ( n14945 , n14942 , n14943 , n14944 );
and ( n14946 , n10837 , n8209 );
and ( n14947 , n11133 , n8039 );
nor ( n14948 , n14946 , n14947 );
xnor ( n14949 , n14948 , n8165 );
and ( n14950 , n8913 , n9795 );
and ( n14951 , n9139 , n9560 );
nor ( n14952 , n14950 , n14951 );
xnor ( n14953 , n14952 , n9801 );
xor ( n14954 , n14949 , n14953 );
and ( n14955 , n8548 , n10342 );
and ( n14956 , n8690 , n10084 );
nor ( n14957 , n14955 , n14956 );
xnor ( n14958 , n14957 , n10291 );
xor ( n14959 , n14954 , n14958 );
xor ( n14960 , n14945 , n14959 );
and ( n14961 , n11384 , n7873 );
and ( n14962 , n11699 , n7762 );
nor ( n14963 , n14961 , n14962 );
xnor ( n14964 , n14963 , n7863 );
and ( n14965 , n7372 , n12782 );
and ( n14966 , n7494 , n12350 );
nor ( n14967 , n14965 , n14966 );
xnor ( n14968 , n14967 , n12733 );
xor ( n14969 , n14964 , n14968 );
and ( n14970 , n7292 , n12730 );
xor ( n14971 , n14969 , n14970 );
xor ( n14972 , n14960 , n14971 );
xor ( n14973 , n14941 , n14972 );
xor ( n14974 , n14932 , n14973 );
and ( n14975 , n14634 , n14645 );
and ( n14976 , n14645 , n14670 );
and ( n14977 , n14634 , n14670 );
or ( n14978 , n14975 , n14976 , n14977 );
and ( n14979 , n12724 , n7400 );
not ( n14980 , n14979 );
xnor ( n14981 , n14980 , n7381 );
and ( n14982 , n9839 , n8887 );
and ( n14983 , n10090 , n8701 );
nor ( n14984 , n14982 , n14983 );
xnor ( n14985 , n14984 , n8893 );
xor ( n14986 , n14981 , n14985 );
and ( n14987 , n7596 , n12029 );
and ( n14988 , n7730 , n11739 );
nor ( n14989 , n14987 , n14988 );
xnor ( n14990 , n14989 , n12019 );
xor ( n14991 , n14986 , n14990 );
and ( n14992 , n10331 , n8511 );
and ( n14993 , n10548 , n8350 );
nor ( n14994 , n14992 , n14993 );
xnor ( n14995 , n14994 , n8517 );
and ( n14996 , n8156 , n10907 );
and ( n14997 , n8339 , n10543 );
nor ( n14998 , n14996 , n14997 );
xnor ( n14999 , n14998 , n10807 );
xor ( n15000 , n14995 , n14999 );
and ( n15001 , n7891 , n11411 );
and ( n15002 , n8045 , n11159 );
nor ( n15003 , n15001 , n15002 );
xnor ( n15004 , n15003 , n11417 );
xor ( n15005 , n15000 , n15004 );
xor ( n15006 , n14991 , n15005 );
and ( n15007 , n14690 , n14694 );
and ( n15008 , n14694 , n14699 );
and ( n15009 , n14690 , n14699 );
or ( n15010 , n15007 , n15008 , n15009 );
and ( n15011 , n12010 , n7609 );
and ( n15012 , n12339 , n7505 );
nor ( n15013 , n15011 , n15012 );
xnor ( n15014 , n15013 , n7615 );
not ( n15015 , n15014 );
xor ( n15016 , n15010 , n15015 );
and ( n15017 , n9323 , n9311 );
and ( n15018 , n9549 , n9150 );
nor ( n15019 , n15017 , n15018 );
xnor ( n15020 , n15019 , n9317 );
xor ( n15021 , n15016 , n15020 );
xor ( n15022 , n15006 , n15021 );
xor ( n15023 , n14978 , n15022 );
and ( n15024 , n14638 , n14642 );
and ( n15025 , n14642 , n14644 );
and ( n15026 , n14638 , n14644 );
or ( n15027 , n15024 , n15025 , n15026 );
and ( n15028 , n14650 , n14654 );
and ( n15029 , n14654 , n14669 );
and ( n15030 , n14650 , n14669 );
or ( n15031 , n15028 , n15029 , n15030 );
xor ( n15032 , n15027 , n15031 );
and ( n15033 , n14659 , n14663 );
and ( n15034 , n14663 , n14668 );
and ( n15035 , n14659 , n14668 );
or ( n15036 , n15033 , n15034 , n15035 );
and ( n15037 , n14713 , n14717 );
and ( n15038 , n14717 , n14722 );
and ( n15039 , n14713 , n14722 );
or ( n15040 , n15037 , n15038 , n15039 );
xor ( n15041 , n15036 , n15040 );
and ( n15042 , n14738 , n14742 );
and ( n15043 , n14742 , n14747 );
and ( n15044 , n14738 , n14747 );
or ( n15045 , n15042 , n15043 , n15044 );
xor ( n15046 , n15041 , n15045 );
xor ( n15047 , n15032 , n15046 );
xor ( n15048 , n15023 , n15047 );
xor ( n15049 , n14974 , n15048 );
xor ( n15050 , n14928 , n15049 );
xor ( n15051 , n14919 , n15050 );
and ( n15052 , n14617 , n14752 );
xor ( n15053 , n15051 , n15052 );
xor ( n15054 , n14915 , n15053 );
and ( n15055 , n14613 , n14755 );
and ( n15056 , n14756 , n14759 );
or ( n15057 , n15055 , n15056 );
xor ( n15058 , n15054 , n15057 );
buf ( n15059 , n15058 );
and ( n15060 , n14902 , n14903 );
and ( n15061 , n14770 , n14821 );
and ( n15062 , n14821 , n14900 );
and ( n15063 , n14770 , n14900 );
or ( n15064 , n15061 , n15062 , n15063 );
and ( n15065 , n14774 , n14778 );
and ( n15066 , n14778 , n14820 );
and ( n15067 , n14774 , n14820 );
or ( n15068 , n15065 , n15066 , n15067 );
and ( n15069 , n14826 , n14830 );
and ( n15070 , n14830 , n14899 );
and ( n15071 , n14826 , n14899 );
or ( n15072 , n15069 , n15070 , n15071 );
xor ( n15073 , n15068 , n15072 );
and ( n15074 , n14835 , n14873 );
and ( n15075 , n14873 , n14898 );
and ( n15076 , n14835 , n14898 );
or ( n15077 , n15074 , n15075 , n15076 );
and ( n15078 , n14849 , n14860 );
and ( n15079 , n14860 , n14872 );
and ( n15080 , n14849 , n14872 );
or ( n15081 , n15078 , n15079 , n15080 );
and ( n15082 , n14878 , n14882 );
and ( n15083 , n14882 , n14897 );
and ( n15084 , n14878 , n14897 );
or ( n15085 , n15082 , n15083 , n15084 );
xor ( n15086 , n15081 , n15085 );
and ( n15087 , n14853 , n14857 );
and ( n15088 , n14857 , n14859 );
and ( n15089 , n14853 , n14859 );
or ( n15090 , n15087 , n15088 , n15089 );
and ( n15091 , n10982 , n8294 );
and ( n15092 , n11274 , n8110 );
nor ( n15093 , n15091 , n15092 );
xnor ( n15094 , n15093 , n8250 );
and ( n15095 , n9018 , n9920 );
and ( n15096 , n9240 , n9671 );
nor ( n15097 , n15095 , n15096 );
xnor ( n15098 , n15097 , n9926 );
xor ( n15099 , n15094 , n15098 );
and ( n15100 , n8643 , n10477 );
and ( n15101 , n8781 , n10205 );
nor ( n15102 , n15100 , n15101 );
xnor ( n15103 , n15102 , n10426 );
xor ( n15104 , n15099 , n15103 );
xor ( n15105 , n15090 , n15104 );
and ( n15106 , n11539 , n7948 );
and ( n15107 , n11850 , n7823 );
nor ( n15108 , n15106 , n15107 );
xnor ( n15109 , n15108 , n7938 );
and ( n15110 , n7427 , n12957 );
and ( n15111 , n7545 , n12511 );
nor ( n15112 , n15110 , n15111 );
xnor ( n15113 , n15112 , n12908 );
xor ( n15114 , n15109 , n15113 );
and ( n15115 , n7333 , n12905 );
xor ( n15116 , n15114 , n15115 );
xor ( n15117 , n15105 , n15116 );
xor ( n15118 , n15086 , n15117 );
xor ( n15119 , n15077 , n15118 );
and ( n15120 , n14783 , n14794 );
and ( n15121 , n14794 , n14819 );
and ( n15122 , n14783 , n14819 );
or ( n15123 , n15120 , n15121 , n15122 );
and ( n15124 , n12899 , n7455 );
not ( n15125 , n15124 );
xnor ( n15126 , n15125 , n7436 );
and ( n15127 , n9964 , n8992 );
and ( n15128 , n10211 , n8792 );
nor ( n15129 , n15127 , n15128 );
xnor ( n15130 , n15129 , n8998 );
xor ( n15131 , n15126 , n15130 );
and ( n15132 , n7661 , n12194 );
and ( n15133 , n7791 , n11890 );
nor ( n15134 , n15132 , n15133 );
xnor ( n15135 , n15134 , n12184 );
xor ( n15136 , n15131 , n15135 );
and ( n15137 , n10466 , n8606 );
and ( n15138 , n10679 , n8431 );
nor ( n15139 , n15137 , n15138 );
xnor ( n15140 , n15139 , n8612 );
and ( n15141 , n8241 , n11052 );
and ( n15142 , n8420 , n10674 );
nor ( n15143 , n15141 , n15142 );
xnor ( n15144 , n15143 , n10952 );
xor ( n15145 , n15140 , n15144 );
and ( n15146 , n7966 , n11566 );
and ( n15147 , n8116 , n11300 );
nor ( n15148 , n15146 , n15147 );
xnor ( n15149 , n15148 , n11572 );
xor ( n15150 , n15145 , n15149 );
xor ( n15151 , n15136 , n15150 );
and ( n15152 , n14839 , n14843 );
and ( n15153 , n14843 , n14848 );
and ( n15154 , n14839 , n14848 );
or ( n15155 , n15152 , n15153 , n15154 );
and ( n15156 , n12175 , n7674 );
and ( n15157 , n12500 , n7556 );
nor ( n15158 , n15156 , n15157 );
xnor ( n15159 , n15158 , n7680 );
not ( n15160 , n15159 );
xor ( n15161 , n15155 , n15160 );
and ( n15162 , n9438 , n9426 );
and ( n15163 , n9660 , n9251 );
nor ( n15164 , n15162 , n15163 );
xnor ( n15165 , n15164 , n9432 );
xor ( n15166 , n15161 , n15165 );
xor ( n15167 , n15151 , n15166 );
xor ( n15168 , n15123 , n15167 );
and ( n15169 , n14787 , n14791 );
and ( n15170 , n14791 , n14793 );
and ( n15171 , n14787 , n14793 );
or ( n15172 , n15169 , n15170 , n15171 );
and ( n15173 , n14799 , n14803 );
and ( n15174 , n14803 , n14818 );
and ( n15175 , n14799 , n14818 );
or ( n15176 , n15173 , n15174 , n15175 );
xor ( n15177 , n15172 , n15176 );
and ( n15178 , n14808 , n14812 );
and ( n15179 , n14812 , n14817 );
and ( n15180 , n14808 , n14817 );
or ( n15181 , n15178 , n15179 , n15180 );
and ( n15182 , n14862 , n14866 );
and ( n15183 , n14866 , n14871 );
and ( n15184 , n14862 , n14871 );
or ( n15185 , n15182 , n15183 , n15184 );
xor ( n15186 , n15181 , n15185 );
and ( n15187 , n14887 , n14891 );
and ( n15188 , n14891 , n14896 );
and ( n15189 , n14887 , n14896 );
or ( n15190 , n15187 , n15188 , n15189 );
xor ( n15191 , n15186 , n15190 );
xor ( n15192 , n15177 , n15191 );
xor ( n15193 , n15168 , n15192 );
xor ( n15194 , n15119 , n15193 );
xor ( n15195 , n15073 , n15194 );
xor ( n15196 , n15064 , n15195 );
and ( n15197 , n14766 , n14901 );
xor ( n15198 , n15196 , n15197 );
xor ( n15199 , n15060 , n15198 );
and ( n15200 , n14762 , n14904 );
and ( n15201 , n14905 , n14908 );
or ( n15202 , n15200 , n15201 );
xor ( n15203 , n15199 , n15202 );
buf ( n15204 , n15203 );
not ( n15205 , n831 );
and ( n15206 , n15205 , n15059 );
and ( n15207 , n15204 , n831 );
or ( n15208 , n15206 , n15207 );
and ( n15209 , n15051 , n15052 );
and ( n15210 , n14923 , n14927 );
and ( n15211 , n14927 , n15049 );
and ( n15212 , n14923 , n15049 );
or ( n15213 , n15210 , n15211 , n15212 );
and ( n15214 , n14978 , n15022 );
and ( n15215 , n15022 , n15047 );
and ( n15216 , n14978 , n15047 );
or ( n15217 , n15214 , n15215 , n15216 );
and ( n15218 , n14932 , n14973 );
and ( n15219 , n14973 , n15048 );
and ( n15220 , n14932 , n15048 );
or ( n15221 , n15218 , n15219 , n15220 );
xor ( n15222 , n15217 , n15221 );
and ( n15223 , n14936 , n14940 );
and ( n15224 , n14940 , n14972 );
and ( n15225 , n14936 , n14972 );
or ( n15226 , n15223 , n15224 , n15225 );
and ( n15227 , n14991 , n15005 );
and ( n15228 , n15005 , n15021 );
and ( n15229 , n14991 , n15021 );
or ( n15230 , n15227 , n15228 , n15229 );
and ( n15231 , n15027 , n15031 );
and ( n15232 , n15031 , n15046 );
and ( n15233 , n15027 , n15046 );
or ( n15234 , n15231 , n15232 , n15233 );
xor ( n15235 , n15230 , n15234 );
and ( n15236 , n15036 , n15040 );
and ( n15237 , n15040 , n15045 );
and ( n15238 , n15036 , n15045 );
or ( n15239 , n15236 , n15237 , n15238 );
and ( n15240 , n15010 , n15015 );
and ( n15241 , n15015 , n15020 );
and ( n15242 , n15010 , n15020 );
or ( n15243 , n15240 , n15241 , n15242 );
xor ( n15244 , n15239 , n15243 );
and ( n15245 , n14949 , n14953 );
and ( n15246 , n14953 , n14958 );
and ( n15247 , n14949 , n14958 );
or ( n15248 , n15245 , n15246 , n15247 );
and ( n15249 , n14981 , n14985 );
and ( n15250 , n14985 , n14990 );
and ( n15251 , n14981 , n14990 );
or ( n15252 , n15249 , n15250 , n15251 );
xor ( n15253 , n15248 , n15252 );
and ( n15254 , n14995 , n14999 );
and ( n15255 , n14999 , n15004 );
and ( n15256 , n14995 , n15004 );
or ( n15257 , n15254 , n15255 , n15256 );
xor ( n15258 , n15253 , n15257 );
xor ( n15259 , n15244 , n15258 );
xor ( n15260 , n15235 , n15259 );
xor ( n15261 , n15226 , n15260 );
and ( n15262 , n14945 , n14959 );
and ( n15263 , n14959 , n14971 );
and ( n15264 , n14945 , n14971 );
or ( n15265 , n15262 , n15263 , n15264 );
and ( n15266 , n14964 , n14968 );
and ( n15267 , n14968 , n14970 );
and ( n15268 , n14964 , n14970 );
or ( n15269 , n15266 , n15267 , n15268 );
and ( n15270 , n10548 , n8511 );
and ( n15271 , n10837 , n8350 );
nor ( n15272 , n15270 , n15271 );
xnor ( n15273 , n15272 , n8517 );
and ( n15274 , n9139 , n9795 );
and ( n15275 , n9323 , n9560 );
nor ( n15276 , n15274 , n15275 );
xnor ( n15277 , n15276 , n9801 );
xor ( n15278 , n15273 , n15277 );
and ( n15279 , n8690 , n10342 );
and ( n15280 , n8913 , n10084 );
nor ( n15281 , n15279 , n15280 );
xnor ( n15282 , n15281 , n10291 );
xor ( n15283 , n15278 , n15282 );
xor ( n15284 , n15269 , n15283 );
not ( n15285 , n7381 );
and ( n15286 , n12339 , n7609 );
and ( n15287 , n12724 , n7505 );
nor ( n15288 , n15286 , n15287 );
xnor ( n15289 , n15288 , n7615 );
xor ( n15290 , n15285 , n15289 );
and ( n15291 , n11133 , n8209 );
and ( n15292 , n11384 , n8039 );
nor ( n15293 , n15291 , n15292 );
xnor ( n15294 , n15293 , n8165 );
xor ( n15295 , n15290 , n15294 );
xor ( n15296 , n15284 , n15295 );
xor ( n15297 , n15265 , n15296 );
and ( n15298 , n10090 , n8887 );
and ( n15299 , n10331 , n8701 );
nor ( n15300 , n15298 , n15299 );
xnor ( n15301 , n15300 , n8893 );
and ( n15302 , n7730 , n12029 );
and ( n15303 , n7891 , n11739 );
nor ( n15304 , n15302 , n15303 );
xnor ( n15305 , n15304 , n12019 );
xor ( n15306 , n15301 , n15305 );
and ( n15307 , n7494 , n12782 );
and ( n15308 , n7596 , n12350 );
nor ( n15309 , n15307 , n15308 );
xnor ( n15310 , n15309 , n12733 );
xor ( n15311 , n15306 , n15310 );
and ( n15312 , n11699 , n7873 );
and ( n15313 , n12010 , n7762 );
nor ( n15314 , n15312 , n15313 );
xnor ( n15315 , n15314 , n7863 );
and ( n15316 , n8339 , n10907 );
and ( n15317 , n8548 , n10543 );
nor ( n15318 , n15316 , n15317 );
xnor ( n15319 , n15318 , n10807 );
xor ( n15320 , n15315 , n15319 );
and ( n15321 , n8045 , n11411 );
and ( n15322 , n8156 , n11159 );
nor ( n15323 , n15321 , n15322 );
xnor ( n15324 , n15323 , n11417 );
xor ( n15325 , n15320 , n15324 );
xor ( n15326 , n15311 , n15325 );
buf ( n15327 , n15014 );
and ( n15328 , n9549 , n9311 );
and ( n15329 , n9839 , n9150 );
nor ( n15330 , n15328 , n15329 );
xnor ( n15331 , n15330 , n9317 );
xor ( n15332 , n15327 , n15331 );
and ( n15333 , n7372 , n12730 );
xor ( n15334 , n15332 , n15333 );
xor ( n15335 , n15326 , n15334 );
xor ( n15336 , n15297 , n15335 );
xor ( n15337 , n15261 , n15336 );
xor ( n15338 , n15222 , n15337 );
xor ( n15339 , n15213 , n15338 );
and ( n15340 , n14919 , n15050 );
xor ( n15341 , n15339 , n15340 );
xor ( n15342 , n15209 , n15341 );
and ( n15343 , n14915 , n15053 );
and ( n15344 , n15054 , n15057 );
or ( n15345 , n15343 , n15344 );
xor ( n15346 , n15342 , n15345 );
buf ( n15347 , n15346 );
and ( n15348 , n15196 , n15197 );
and ( n15349 , n15068 , n15072 );
and ( n15350 , n15072 , n15194 );
and ( n15351 , n15068 , n15194 );
or ( n15352 , n15349 , n15350 , n15351 );
and ( n15353 , n15123 , n15167 );
and ( n15354 , n15167 , n15192 );
and ( n15355 , n15123 , n15192 );
or ( n15356 , n15353 , n15354 , n15355 );
and ( n15357 , n15077 , n15118 );
and ( n15358 , n15118 , n15193 );
and ( n15359 , n15077 , n15193 );
or ( n15360 , n15357 , n15358 , n15359 );
xor ( n15361 , n15356 , n15360 );
and ( n15362 , n15081 , n15085 );
and ( n15363 , n15085 , n15117 );
and ( n15364 , n15081 , n15117 );
or ( n15365 , n15362 , n15363 , n15364 );
and ( n15366 , n15136 , n15150 );
and ( n15367 , n15150 , n15166 );
and ( n15368 , n15136 , n15166 );
or ( n15369 , n15366 , n15367 , n15368 );
and ( n15370 , n15172 , n15176 );
and ( n15371 , n15176 , n15191 );
and ( n15372 , n15172 , n15191 );
or ( n15373 , n15370 , n15371 , n15372 );
xor ( n15374 , n15369 , n15373 );
and ( n15375 , n15181 , n15185 );
and ( n15376 , n15185 , n15190 );
and ( n15377 , n15181 , n15190 );
or ( n15378 , n15375 , n15376 , n15377 );
and ( n15379 , n15155 , n15160 );
and ( n15380 , n15160 , n15165 );
and ( n15381 , n15155 , n15165 );
or ( n15382 , n15379 , n15380 , n15381 );
xor ( n15383 , n15378 , n15382 );
and ( n15384 , n15094 , n15098 );
and ( n15385 , n15098 , n15103 );
and ( n15386 , n15094 , n15103 );
or ( n15387 , n15384 , n15385 , n15386 );
and ( n15388 , n15126 , n15130 );
and ( n15389 , n15130 , n15135 );
and ( n15390 , n15126 , n15135 );
or ( n15391 , n15388 , n15389 , n15390 );
xor ( n15392 , n15387 , n15391 );
and ( n15393 , n15140 , n15144 );
and ( n15394 , n15144 , n15149 );
and ( n15395 , n15140 , n15149 );
or ( n15396 , n15393 , n15394 , n15395 );
xor ( n15397 , n15392 , n15396 );
xor ( n15398 , n15383 , n15397 );
xor ( n15399 , n15374 , n15398 );
xor ( n15400 , n15365 , n15399 );
and ( n15401 , n15090 , n15104 );
and ( n15402 , n15104 , n15116 );
and ( n15403 , n15090 , n15116 );
or ( n15404 , n15401 , n15402 , n15403 );
and ( n15405 , n15109 , n15113 );
and ( n15406 , n15113 , n15115 );
and ( n15407 , n15109 , n15115 );
or ( n15408 , n15405 , n15406 , n15407 );
and ( n15409 , n10679 , n8606 );
and ( n15410 , n10982 , n8431 );
nor ( n15411 , n15409 , n15410 );
xnor ( n15412 , n15411 , n8612 );
and ( n15413 , n9240 , n9920 );
and ( n15414 , n9438 , n9671 );
nor ( n15415 , n15413 , n15414 );
xnor ( n15416 , n15415 , n9926 );
xor ( n15417 , n15412 , n15416 );
and ( n15418 , n8781 , n10477 );
and ( n15419 , n9018 , n10205 );
nor ( n15420 , n15418 , n15419 );
xnor ( n15421 , n15420 , n10426 );
xor ( n15422 , n15417 , n15421 );
xor ( n15423 , n15408 , n15422 );
not ( n15424 , n7436 );
and ( n15425 , n12500 , n7674 );
and ( n15426 , n12899 , n7556 );
nor ( n15427 , n15425 , n15426 );
xnor ( n15428 , n15427 , n7680 );
xor ( n15429 , n15424 , n15428 );
and ( n15430 , n11274 , n8294 );
and ( n15431 , n11539 , n8110 );
nor ( n15432 , n15430 , n15431 );
xnor ( n15433 , n15432 , n8250 );
xor ( n15434 , n15429 , n15433 );
xor ( n15435 , n15423 , n15434 );
xor ( n15436 , n15404 , n15435 );
and ( n15437 , n10211 , n8992 );
and ( n15438 , n10466 , n8792 );
nor ( n15439 , n15437 , n15438 );
xnor ( n15440 , n15439 , n8998 );
and ( n15441 , n7791 , n12194 );
and ( n15442 , n7966 , n11890 );
nor ( n15443 , n15441 , n15442 );
xnor ( n15444 , n15443 , n12184 );
xor ( n15445 , n15440 , n15444 );
and ( n15446 , n7545 , n12957 );
and ( n15447 , n7661 , n12511 );
nor ( n15448 , n15446 , n15447 );
xnor ( n15449 , n15448 , n12908 );
xor ( n15450 , n15445 , n15449 );
and ( n15451 , n11850 , n7948 );
and ( n15452 , n12175 , n7823 );
nor ( n15453 , n15451 , n15452 );
xnor ( n15454 , n15453 , n7938 );
and ( n15455 , n8420 , n11052 );
and ( n15456 , n8643 , n10674 );
nor ( n15457 , n15455 , n15456 );
xnor ( n15458 , n15457 , n10952 );
xor ( n15459 , n15454 , n15458 );
and ( n15460 , n8116 , n11566 );
and ( n15461 , n8241 , n11300 );
nor ( n15462 , n15460 , n15461 );
xnor ( n15463 , n15462 , n11572 );
xor ( n15464 , n15459 , n15463 );
xor ( n15465 , n15450 , n15464 );
buf ( n15466 , n15159 );
and ( n15467 , n9660 , n9426 );
and ( n15468 , n9964 , n9251 );
nor ( n15469 , n15467 , n15468 );
xnor ( n15470 , n15469 , n9432 );
xor ( n15471 , n15466 , n15470 );
and ( n15472 , n7427 , n12905 );
xor ( n15473 , n15471 , n15472 );
xor ( n15474 , n15465 , n15473 );
xor ( n15475 , n15436 , n15474 );
xor ( n15476 , n15400 , n15475 );
xor ( n15477 , n15361 , n15476 );
xor ( n15478 , n15352 , n15477 );
and ( n15479 , n15064 , n15195 );
xor ( n15480 , n15478 , n15479 );
xor ( n15481 , n15348 , n15480 );
and ( n15482 , n15060 , n15198 );
and ( n15483 , n15199 , n15202 );
or ( n15484 , n15482 , n15483 );
xor ( n15485 , n15481 , n15484 );
buf ( n15486 , n15485 );
not ( n15487 , n831 );
and ( n15488 , n15487 , n15347 );
and ( n15489 , n15486 , n831 );
or ( n15490 , n15488 , n15489 );
and ( n15491 , n15339 , n15340 );
and ( n15492 , n15217 , n15221 );
and ( n15493 , n15221 , n15337 );
and ( n15494 , n15217 , n15337 );
or ( n15495 , n15492 , n15493 , n15494 );
and ( n15496 , n15226 , n15260 );
and ( n15497 , n15260 , n15336 );
and ( n15498 , n15226 , n15336 );
or ( n15499 , n15496 , n15497 , n15498 );
and ( n15500 , n15239 , n15243 );
and ( n15501 , n15243 , n15258 );
and ( n15502 , n15239 , n15258 );
or ( n15503 , n15500 , n15501 , n15502 );
and ( n15504 , n12724 , n7609 );
not ( n15505 , n15504 );
xnor ( n15506 , n15505 , n7615 );
and ( n15507 , n9839 , n9311 );
and ( n15508 , n10090 , n9150 );
nor ( n15509 , n15507 , n15508 );
xnor ( n15510 , n15509 , n9317 );
xor ( n15511 , n15506 , n15510 );
and ( n15512 , n7596 , n12782 );
and ( n15513 , n7730 , n12350 );
nor ( n15514 , n15512 , n15513 );
xnor ( n15515 , n15514 , n12733 );
xor ( n15516 , n15511 , n15515 );
and ( n15517 , n10837 , n8511 );
and ( n15518 , n11133 , n8350 );
nor ( n15519 , n15517 , n15518 );
xnor ( n15520 , n15519 , n8517 );
and ( n15521 , n8913 , n10342 );
and ( n15522 , n9139 , n10084 );
nor ( n15523 , n15521 , n15522 );
xnor ( n15524 , n15523 , n10291 );
xor ( n15525 , n15520 , n15524 );
and ( n15526 , n8548 , n10907 );
and ( n15527 , n8690 , n10543 );
nor ( n15528 , n15526 , n15527 );
xnor ( n15529 , n15528 , n10807 );
xor ( n15530 , n15525 , n15529 );
xor ( n15531 , n15516 , n15530 );
and ( n15532 , n10331 , n8887 );
and ( n15533 , n10548 , n8701 );
nor ( n15534 , n15532 , n15533 );
xnor ( n15535 , n15534 , n8893 );
and ( n15536 , n8156 , n11411 );
and ( n15537 , n8339 , n11159 );
nor ( n15538 , n15536 , n15537 );
xnor ( n15539 , n15538 , n11417 );
xor ( n15540 , n15535 , n15539 );
and ( n15541 , n7891 , n12029 );
and ( n15542 , n8045 , n11739 );
nor ( n15543 , n15541 , n15542 );
xnor ( n15544 , n15543 , n12019 );
xor ( n15545 , n15540 , n15544 );
xor ( n15546 , n15531 , n15545 );
xor ( n15547 , n15503 , n15546 );
and ( n15548 , n15248 , n15252 );
and ( n15549 , n15252 , n15257 );
and ( n15550 , n15248 , n15257 );
or ( n15551 , n15548 , n15549 , n15550 );
and ( n15552 , n15327 , n15331 );
and ( n15553 , n15331 , n15333 );
and ( n15554 , n15327 , n15333 );
or ( n15555 , n15552 , n15553 , n15554 );
xor ( n15556 , n15551 , n15555 );
and ( n15557 , n15273 , n15277 );
and ( n15558 , n15277 , n15282 );
and ( n15559 , n15273 , n15282 );
or ( n15560 , n15557 , n15558 , n15559 );
and ( n15561 , n15315 , n15319 );
and ( n15562 , n15319 , n15324 );
and ( n15563 , n15315 , n15324 );
or ( n15564 , n15561 , n15562 , n15563 );
xor ( n15565 , n15560 , n15564 );
and ( n15566 , n12010 , n7873 );
and ( n15567 , n12339 , n7762 );
nor ( n15568 , n15566 , n15567 );
xnor ( n15569 , n15568 , n7863 );
not ( n15570 , n15569 );
xor ( n15571 , n15565 , n15570 );
xor ( n15572 , n15556 , n15571 );
xor ( n15573 , n15547 , n15572 );
xor ( n15574 , n15499 , n15573 );
and ( n15575 , n15230 , n15234 );
and ( n15576 , n15234 , n15259 );
and ( n15577 , n15230 , n15259 );
or ( n15578 , n15575 , n15576 , n15577 );
and ( n15579 , n15265 , n15296 );
and ( n15580 , n15296 , n15335 );
and ( n15581 , n15265 , n15335 );
or ( n15582 , n15579 , n15580 , n15581 );
xor ( n15583 , n15578 , n15582 );
and ( n15584 , n15269 , n15283 );
and ( n15585 , n15283 , n15295 );
and ( n15586 , n15269 , n15295 );
or ( n15587 , n15584 , n15585 , n15586 );
and ( n15588 , n15311 , n15325 );
and ( n15589 , n15325 , n15334 );
and ( n15590 , n15311 , n15334 );
or ( n15591 , n15588 , n15589 , n15590 );
xor ( n15592 , n15587 , n15591 );
and ( n15593 , n15285 , n15289 );
and ( n15594 , n15289 , n15294 );
and ( n15595 , n15285 , n15294 );
or ( n15596 , n15593 , n15594 , n15595 );
and ( n15597 , n15301 , n15305 );
and ( n15598 , n15305 , n15310 );
and ( n15599 , n15301 , n15310 );
or ( n15600 , n15597 , n15598 , n15599 );
xor ( n15601 , n15596 , n15600 );
and ( n15602 , n11384 , n8209 );
and ( n15603 , n11699 , n8039 );
nor ( n15604 , n15602 , n15603 );
xnor ( n15605 , n15604 , n8165 );
and ( n15606 , n9323 , n9795 );
and ( n15607 , n9549 , n9560 );
nor ( n15608 , n15606 , n15607 );
xnor ( n15609 , n15608 , n9801 );
xor ( n15610 , n15605 , n15609 );
and ( n15611 , n7494 , n12730 );
xor ( n15612 , n15610 , n15611 );
xor ( n15613 , n15601 , n15612 );
xor ( n15614 , n15592 , n15613 );
xor ( n15615 , n15583 , n15614 );
xor ( n15616 , n15574 , n15615 );
xor ( n15617 , n15495 , n15616 );
and ( n15618 , n15213 , n15338 );
xor ( n15619 , n15617 , n15618 );
xor ( n15620 , n15491 , n15619 );
and ( n15621 , n15209 , n15341 );
and ( n15622 , n15342 , n15345 );
or ( n15623 , n15621 , n15622 );
xor ( n15624 , n15620 , n15623 );
buf ( n15625 , n15624 );
and ( n15626 , n15478 , n15479 );
and ( n15627 , n15356 , n15360 );
and ( n15628 , n15360 , n15476 );
and ( n15629 , n15356 , n15476 );
or ( n15630 , n15627 , n15628 , n15629 );
and ( n15631 , n15365 , n15399 );
and ( n15632 , n15399 , n15475 );
and ( n15633 , n15365 , n15475 );
or ( n15634 , n15631 , n15632 , n15633 );
and ( n15635 , n15378 , n15382 );
and ( n15636 , n15382 , n15397 );
and ( n15637 , n15378 , n15397 );
or ( n15638 , n15635 , n15636 , n15637 );
and ( n15639 , n12899 , n7674 );
not ( n15640 , n15639 );
xnor ( n15641 , n15640 , n7680 );
and ( n15642 , n9964 , n9426 );
and ( n15643 , n10211 , n9251 );
nor ( n15644 , n15642 , n15643 );
xnor ( n15645 , n15644 , n9432 );
xor ( n15646 , n15641 , n15645 );
and ( n15647 , n7661 , n12957 );
and ( n15648 , n7791 , n12511 );
nor ( n15649 , n15647 , n15648 );
xnor ( n15650 , n15649 , n12908 );
xor ( n15651 , n15646 , n15650 );
and ( n15652 , n10982 , n8606 );
and ( n15653 , n11274 , n8431 );
nor ( n15654 , n15652 , n15653 );
xnor ( n15655 , n15654 , n8612 );
and ( n15656 , n9018 , n10477 );
and ( n15657 , n9240 , n10205 );
nor ( n15658 , n15656 , n15657 );
xnor ( n15659 , n15658 , n10426 );
xor ( n15660 , n15655 , n15659 );
and ( n15661 , n8643 , n11052 );
and ( n15662 , n8781 , n10674 );
nor ( n15663 , n15661 , n15662 );
xnor ( n15664 , n15663 , n10952 );
xor ( n15665 , n15660 , n15664 );
xor ( n15666 , n15651 , n15665 );
and ( n15667 , n10466 , n8992 );
and ( n15668 , n10679 , n8792 );
nor ( n15669 , n15667 , n15668 );
xnor ( n15670 , n15669 , n8998 );
and ( n15671 , n8241 , n11566 );
and ( n15672 , n8420 , n11300 );
nor ( n15673 , n15671 , n15672 );
xnor ( n15674 , n15673 , n11572 );
xor ( n15675 , n15670 , n15674 );
and ( n15676 , n7966 , n12194 );
and ( n15677 , n8116 , n11890 );
nor ( n15678 , n15676 , n15677 );
xnor ( n15679 , n15678 , n12184 );
xor ( n15680 , n15675 , n15679 );
xor ( n15681 , n15666 , n15680 );
xor ( n15682 , n15638 , n15681 );
and ( n15683 , n15387 , n15391 );
and ( n15684 , n15391 , n15396 );
and ( n15685 , n15387 , n15396 );
or ( n15686 , n15683 , n15684 , n15685 );
and ( n15687 , n15466 , n15470 );
and ( n15688 , n15470 , n15472 );
and ( n15689 , n15466 , n15472 );
or ( n15690 , n15687 , n15688 , n15689 );
xor ( n15691 , n15686 , n15690 );
and ( n15692 , n15412 , n15416 );
and ( n15693 , n15416 , n15421 );
and ( n15694 , n15412 , n15421 );
or ( n15695 , n15692 , n15693 , n15694 );
and ( n15696 , n15454 , n15458 );
and ( n15697 , n15458 , n15463 );
and ( n15698 , n15454 , n15463 );
or ( n15699 , n15696 , n15697 , n15698 );
xor ( n15700 , n15695 , n15699 );
and ( n15701 , n12175 , n7948 );
and ( n15702 , n12500 , n7823 );
nor ( n15703 , n15701 , n15702 );
xnor ( n15704 , n15703 , n7938 );
not ( n15705 , n15704 );
xor ( n15706 , n15700 , n15705 );
xor ( n15707 , n15691 , n15706 );
xor ( n15708 , n15682 , n15707 );
xor ( n15709 , n15634 , n15708 );
and ( n15710 , n15369 , n15373 );
and ( n15711 , n15373 , n15398 );
and ( n15712 , n15369 , n15398 );
or ( n15713 , n15710 , n15711 , n15712 );
and ( n15714 , n15404 , n15435 );
and ( n15715 , n15435 , n15474 );
and ( n15716 , n15404 , n15474 );
or ( n15717 , n15714 , n15715 , n15716 );
xor ( n15718 , n15713 , n15717 );
and ( n15719 , n15408 , n15422 );
and ( n15720 , n15422 , n15434 );
and ( n15721 , n15408 , n15434 );
or ( n15722 , n15719 , n15720 , n15721 );
and ( n15723 , n15450 , n15464 );
and ( n15724 , n15464 , n15473 );
and ( n15725 , n15450 , n15473 );
or ( n15726 , n15723 , n15724 , n15725 );
xor ( n15727 , n15722 , n15726 );
and ( n15728 , n15424 , n15428 );
and ( n15729 , n15428 , n15433 );
and ( n15730 , n15424 , n15433 );
or ( n15731 , n15728 , n15729 , n15730 );
and ( n15732 , n15440 , n15444 );
and ( n15733 , n15444 , n15449 );
and ( n15734 , n15440 , n15449 );
or ( n15735 , n15732 , n15733 , n15734 );
xor ( n15736 , n15731 , n15735 );
and ( n15737 , n11539 , n8294 );
and ( n15738 , n11850 , n8110 );
nor ( n15739 , n15737 , n15738 );
xnor ( n15740 , n15739 , n8250 );
and ( n15741 , n9438 , n9920 );
and ( n15742 , n9660 , n9671 );
nor ( n15743 , n15741 , n15742 );
xnor ( n15744 , n15743 , n9926 );
xor ( n15745 , n15740 , n15744 );
and ( n15746 , n7545 , n12905 );
xor ( n15747 , n15745 , n15746 );
xor ( n15748 , n15736 , n15747 );
xor ( n15749 , n15727 , n15748 );
xor ( n15750 , n15718 , n15749 );
xor ( n15751 , n15709 , n15750 );
xor ( n15752 , n15630 , n15751 );
and ( n15753 , n15352 , n15477 );
xor ( n15754 , n15752 , n15753 );
xor ( n15755 , n15626 , n15754 );
and ( n15756 , n15348 , n15480 );
and ( n15757 , n15481 , n15484 );
or ( n15758 , n15756 , n15757 );
xor ( n15759 , n15755 , n15758 );
buf ( n15760 , n15759 );
not ( n15761 , n831 );
and ( n15762 , n15761 , n15625 );
and ( n15763 , n15760 , n831 );
or ( n15764 , n15762 , n15763 );
and ( n15765 , n15499 , n15573 );
and ( n15766 , n15573 , n15615 );
and ( n15767 , n15499 , n15615 );
or ( n15768 , n15765 , n15766 , n15767 );
and ( n15769 , n15578 , n15582 );
and ( n15770 , n15582 , n15614 );
and ( n15771 , n15578 , n15614 );
or ( n15772 , n15769 , n15770 , n15771 );
and ( n15773 , n15551 , n15555 );
and ( n15774 , n15555 , n15571 );
and ( n15775 , n15551 , n15571 );
or ( n15776 , n15773 , n15774 , n15775 );
and ( n15777 , n11699 , n8209 );
and ( n15778 , n12010 , n8039 );
nor ( n15779 , n15777 , n15778 );
xnor ( n15780 , n15779 , n8165 );
and ( n15781 , n8339 , n11411 );
and ( n15782 , n8548 , n11159 );
nor ( n15783 , n15781 , n15782 );
xnor ( n15784 , n15783 , n11417 );
xor ( n15785 , n15780 , n15784 );
and ( n15786 , n8045 , n12029 );
and ( n15787 , n8156 , n11739 );
nor ( n15788 , n15786 , n15787 );
xnor ( n15789 , n15788 , n12019 );
xor ( n15790 , n15785 , n15789 );
not ( n15791 , n7615 );
and ( n15792 , n12339 , n7873 );
and ( n15793 , n12724 , n7762 );
nor ( n15794 , n15792 , n15793 );
xnor ( n15795 , n15794 , n7863 );
xor ( n15796 , n15791 , n15795 );
and ( n15797 , n11133 , n8511 );
and ( n15798 , n11384 , n8350 );
nor ( n15799 , n15797 , n15798 );
xnor ( n15800 , n15799 , n8517 );
xor ( n15801 , n15796 , n15800 );
xor ( n15802 , n15790 , n15801 );
and ( n15803 , n10548 , n8887 );
and ( n15804 , n10837 , n8701 );
nor ( n15805 , n15803 , n15804 );
xnor ( n15806 , n15805 , n8893 );
and ( n15807 , n9139 , n10342 );
and ( n15808 , n9323 , n10084 );
nor ( n15809 , n15807 , n15808 );
xnor ( n15810 , n15809 , n10291 );
xor ( n15811 , n15806 , n15810 );
and ( n15812 , n8690 , n10907 );
and ( n15813 , n8913 , n10543 );
nor ( n15814 , n15812 , n15813 );
xnor ( n15815 , n15814 , n10807 );
xor ( n15816 , n15811 , n15815 );
xor ( n15817 , n15802 , n15816 );
xor ( n15818 , n15776 , n15817 );
and ( n15819 , n15560 , n15564 );
and ( n15820 , n15564 , n15570 );
and ( n15821 , n15560 , n15570 );
or ( n15822 , n15819 , n15820 , n15821 );
and ( n15823 , n10090 , n9311 );
and ( n15824 , n10331 , n9150 );
nor ( n15825 , n15823 , n15824 );
xnor ( n15826 , n15825 , n9317 );
and ( n15827 , n7730 , n12782 );
and ( n15828 , n7891 , n12350 );
nor ( n15829 , n15827 , n15828 );
xnor ( n15830 , n15829 , n12733 );
xor ( n15831 , n15826 , n15830 );
and ( n15832 , n7596 , n12730 );
xor ( n15833 , n15831 , n15832 );
xor ( n15834 , n15822 , n15833 );
and ( n15835 , n15535 , n15539 );
and ( n15836 , n15539 , n15544 );
and ( n15837 , n15535 , n15544 );
or ( n15838 , n15835 , n15836 , n15837 );
buf ( n15839 , n15569 );
xor ( n15840 , n15838 , n15839 );
and ( n15841 , n9549 , n9795 );
and ( n15842 , n9839 , n9560 );
nor ( n15843 , n15841 , n15842 );
xnor ( n15844 , n15843 , n9801 );
xor ( n15845 , n15840 , n15844 );
xor ( n15846 , n15834 , n15845 );
xor ( n15847 , n15818 , n15846 );
xor ( n15848 , n15772 , n15847 );
and ( n15849 , n15503 , n15546 );
and ( n15850 , n15546 , n15572 );
and ( n15851 , n15503 , n15572 );
or ( n15852 , n15849 , n15850 , n15851 );
and ( n15853 , n15587 , n15591 );
and ( n15854 , n15591 , n15613 );
and ( n15855 , n15587 , n15613 );
or ( n15856 , n15853 , n15854 , n15855 );
xor ( n15857 , n15852 , n15856 );
and ( n15858 , n15516 , n15530 );
and ( n15859 , n15530 , n15545 );
and ( n15860 , n15516 , n15545 );
or ( n15861 , n15858 , n15859 , n15860 );
and ( n15862 , n15596 , n15600 );
and ( n15863 , n15600 , n15612 );
and ( n15864 , n15596 , n15612 );
or ( n15865 , n15862 , n15863 , n15864 );
xor ( n15866 , n15861 , n15865 );
and ( n15867 , n15506 , n15510 );
and ( n15868 , n15510 , n15515 );
and ( n15869 , n15506 , n15515 );
or ( n15870 , n15867 , n15868 , n15869 );
and ( n15871 , n15520 , n15524 );
and ( n15872 , n15524 , n15529 );
and ( n15873 , n15520 , n15529 );
or ( n15874 , n15871 , n15872 , n15873 );
xor ( n15875 , n15870 , n15874 );
and ( n15876 , n15605 , n15609 );
and ( n15877 , n15609 , n15611 );
and ( n15878 , n15605 , n15611 );
or ( n15879 , n15876 , n15877 , n15878 );
xor ( n15880 , n15875 , n15879 );
xor ( n15881 , n15866 , n15880 );
xor ( n15882 , n15857 , n15881 );
xor ( n15883 , n15848 , n15882 );
xor ( n15884 , n15768 , n15883 );
and ( n15885 , n15495 , n15616 );
xor ( n15886 , n15884 , n15885 );
and ( n15887 , n15617 , n15618 );
xor ( n15888 , n15886 , n15887 );
and ( n15889 , n15491 , n15619 );
and ( n15890 , n15620 , n15623 );
or ( n15891 , n15889 , n15890 );
xor ( n15892 , n15888 , n15891 );
buf ( n15893 , n15892 );
and ( n15894 , n15634 , n15708 );
and ( n15895 , n15708 , n15750 );
and ( n15896 , n15634 , n15750 );
or ( n15897 , n15894 , n15895 , n15896 );
and ( n15898 , n15713 , n15717 );
and ( n15899 , n15717 , n15749 );
and ( n15900 , n15713 , n15749 );
or ( n15901 , n15898 , n15899 , n15900 );
and ( n15902 , n15686 , n15690 );
and ( n15903 , n15690 , n15706 );
and ( n15904 , n15686 , n15706 );
or ( n15905 , n15902 , n15903 , n15904 );
and ( n15906 , n11850 , n8294 );
and ( n15907 , n12175 , n8110 );
nor ( n15908 , n15906 , n15907 );
xnor ( n15909 , n15908 , n8250 );
and ( n15910 , n8420 , n11566 );
and ( n15911 , n8643 , n11300 );
nor ( n15912 , n15910 , n15911 );
xnor ( n15913 , n15912 , n11572 );
xor ( n15914 , n15909 , n15913 );
and ( n15915 , n8116 , n12194 );
and ( n15916 , n8241 , n11890 );
nor ( n15917 , n15915 , n15916 );
xnor ( n15918 , n15917 , n12184 );
xor ( n15919 , n15914 , n15918 );
not ( n15920 , n7680 );
and ( n15921 , n12500 , n7948 );
and ( n15922 , n12899 , n7823 );
nor ( n15923 , n15921 , n15922 );
xnor ( n15924 , n15923 , n7938 );
xor ( n15925 , n15920 , n15924 );
and ( n15926 , n11274 , n8606 );
and ( n15927 , n11539 , n8431 );
nor ( n15928 , n15926 , n15927 );
xnor ( n15929 , n15928 , n8612 );
xor ( n15930 , n15925 , n15929 );
xor ( n15931 , n15919 , n15930 );
and ( n15932 , n10679 , n8992 );
and ( n15933 , n10982 , n8792 );
nor ( n15934 , n15932 , n15933 );
xnor ( n15935 , n15934 , n8998 );
and ( n15936 , n9240 , n10477 );
and ( n15937 , n9438 , n10205 );
nor ( n15938 , n15936 , n15937 );
xnor ( n15939 , n15938 , n10426 );
xor ( n15940 , n15935 , n15939 );
and ( n15941 , n8781 , n11052 );
and ( n15942 , n9018 , n10674 );
nor ( n15943 , n15941 , n15942 );
xnor ( n15944 , n15943 , n10952 );
xor ( n15945 , n15940 , n15944 );
xor ( n15946 , n15931 , n15945 );
xor ( n15947 , n15905 , n15946 );
and ( n15948 , n15695 , n15699 );
and ( n15949 , n15699 , n15705 );
and ( n15950 , n15695 , n15705 );
or ( n15951 , n15948 , n15949 , n15950 );
and ( n15952 , n10211 , n9426 );
and ( n15953 , n10466 , n9251 );
nor ( n15954 , n15952 , n15953 );
xnor ( n15955 , n15954 , n9432 );
and ( n15956 , n7791 , n12957 );
and ( n15957 , n7966 , n12511 );
nor ( n15958 , n15956 , n15957 );
xnor ( n15959 , n15958 , n12908 );
xor ( n15960 , n15955 , n15959 );
and ( n15961 , n7661 , n12905 );
xor ( n15962 , n15960 , n15961 );
xor ( n15963 , n15951 , n15962 );
and ( n15964 , n15670 , n15674 );
and ( n15965 , n15674 , n15679 );
and ( n15966 , n15670 , n15679 );
or ( n15967 , n15964 , n15965 , n15966 );
buf ( n15968 , n15704 );
xor ( n15969 , n15967 , n15968 );
and ( n15970 , n9660 , n9920 );
and ( n15971 , n9964 , n9671 );
nor ( n15972 , n15970 , n15971 );
xnor ( n15973 , n15972 , n9926 );
xor ( n15974 , n15969 , n15973 );
xor ( n15975 , n15963 , n15974 );
xor ( n15976 , n15947 , n15975 );
xor ( n15977 , n15901 , n15976 );
and ( n15978 , n15638 , n15681 );
and ( n15979 , n15681 , n15707 );
and ( n15980 , n15638 , n15707 );
or ( n15981 , n15978 , n15979 , n15980 );
and ( n15982 , n15722 , n15726 );
and ( n15983 , n15726 , n15748 );
and ( n15984 , n15722 , n15748 );
or ( n15985 , n15982 , n15983 , n15984 );
xor ( n15986 , n15981 , n15985 );
and ( n15987 , n15651 , n15665 );
and ( n15988 , n15665 , n15680 );
and ( n15989 , n15651 , n15680 );
or ( n15990 , n15987 , n15988 , n15989 );
and ( n15991 , n15731 , n15735 );
and ( n15992 , n15735 , n15747 );
and ( n15993 , n15731 , n15747 );
or ( n15994 , n15991 , n15992 , n15993 );
xor ( n15995 , n15990 , n15994 );
and ( n15996 , n15641 , n15645 );
and ( n15997 , n15645 , n15650 );
and ( n15998 , n15641 , n15650 );
or ( n15999 , n15996 , n15997 , n15998 );
and ( n16000 , n15655 , n15659 );
and ( n16001 , n15659 , n15664 );
and ( n16002 , n15655 , n15664 );
or ( n16003 , n16000 , n16001 , n16002 );
xor ( n16004 , n15999 , n16003 );
and ( n16005 , n15740 , n15744 );
and ( n16006 , n15744 , n15746 );
and ( n16007 , n15740 , n15746 );
or ( n16008 , n16005 , n16006 , n16007 );
xor ( n16009 , n16004 , n16008 );
xor ( n16010 , n15995 , n16009 );
xor ( n16011 , n15986 , n16010 );
xor ( n16012 , n15977 , n16011 );
xor ( n16013 , n15897 , n16012 );
and ( n16014 , n15630 , n15751 );
xor ( n16015 , n16013 , n16014 );
and ( n16016 , n15752 , n15753 );
xor ( n16017 , n16015 , n16016 );
and ( n16018 , n15626 , n15754 );
and ( n16019 , n15755 , n15758 );
or ( n16020 , n16018 , n16019 );
xor ( n16021 , n16017 , n16020 );
buf ( n16022 , n16021 );
not ( n16023 , n831 );
and ( n16024 , n16023 , n15893 );
and ( n16025 , n16022 , n831 );
or ( n16026 , n16024 , n16025 );
and ( n16027 , n15884 , n15885 );
and ( n16028 , n15772 , n15847 );
and ( n16029 , n15847 , n15882 );
and ( n16030 , n15772 , n15882 );
or ( n16031 , n16028 , n16029 , n16030 );
and ( n16032 , n15852 , n15856 );
and ( n16033 , n15856 , n15881 );
and ( n16034 , n15852 , n15881 );
or ( n16035 , n16032 , n16033 , n16034 );
and ( n16036 , n15822 , n15833 );
and ( n16037 , n15833 , n15845 );
and ( n16038 , n15822 , n15845 );
or ( n16039 , n16036 , n16037 , n16038 );
and ( n16040 , n15806 , n15810 );
and ( n16041 , n15810 , n15815 );
and ( n16042 , n15806 , n15815 );
or ( n16043 , n16040 , n16041 , n16042 );
and ( n16044 , n12724 , n7873 );
not ( n16045 , n16044 );
xnor ( n16046 , n16045 , n7863 );
and ( n16047 , n11384 , n8511 );
and ( n16048 , n11699 , n8350 );
nor ( n16049 , n16047 , n16048 );
xnor ( n16050 , n16049 , n8517 );
xor ( n16051 , n16046 , n16050 );
and ( n16052 , n7730 , n12730 );
xor ( n16053 , n16051 , n16052 );
xor ( n16054 , n16043 , n16053 );
and ( n16055 , n10837 , n8887 );
and ( n16056 , n11133 , n8701 );
nor ( n16057 , n16055 , n16056 );
xnor ( n16058 , n16057 , n8893 );
and ( n16059 , n8913 , n10907 );
and ( n16060 , n9139 , n10543 );
nor ( n16061 , n16059 , n16060 );
xnor ( n16062 , n16061 , n10807 );
xor ( n16063 , n16058 , n16062 );
and ( n16064 , n8548 , n11411 );
and ( n16065 , n8690 , n11159 );
nor ( n16066 , n16064 , n16065 );
xnor ( n16067 , n16066 , n11417 );
xor ( n16068 , n16063 , n16067 );
xor ( n16069 , n16054 , n16068 );
xor ( n16070 , n16039 , n16069 );
and ( n16071 , n15870 , n15874 );
and ( n16072 , n15874 , n15879 );
and ( n16073 , n15870 , n15879 );
or ( n16074 , n16071 , n16072 , n16073 );
and ( n16075 , n10331 , n9311 );
and ( n16076 , n10548 , n9150 );
nor ( n16077 , n16075 , n16076 );
xnor ( n16078 , n16077 , n9317 );
and ( n16079 , n8156 , n12029 );
and ( n16080 , n8339 , n11739 );
nor ( n16081 , n16079 , n16080 );
xnor ( n16082 , n16081 , n12019 );
xor ( n16083 , n16078 , n16082 );
and ( n16084 , n7891 , n12782 );
and ( n16085 , n8045 , n12350 );
nor ( n16086 , n16084 , n16085 );
xnor ( n16087 , n16086 , n12733 );
xor ( n16088 , n16083 , n16087 );
xor ( n16089 , n16074 , n16088 );
and ( n16090 , n12010 , n8209 );
and ( n16091 , n12339 , n8039 );
nor ( n16092 , n16090 , n16091 );
xnor ( n16093 , n16092 , n8165 );
not ( n16094 , n16093 );
and ( n16095 , n9839 , n9795 );
and ( n16096 , n10090 , n9560 );
nor ( n16097 , n16095 , n16096 );
xnor ( n16098 , n16097 , n9801 );
xor ( n16099 , n16094 , n16098 );
and ( n16100 , n9323 , n10342 );
and ( n16101 , n9549 , n10084 );
nor ( n16102 , n16100 , n16101 );
xnor ( n16103 , n16102 , n10291 );
xor ( n16104 , n16099 , n16103 );
xor ( n16105 , n16089 , n16104 );
xor ( n16106 , n16070 , n16105 );
xor ( n16107 , n16035 , n16106 );
and ( n16108 , n15861 , n15865 );
and ( n16109 , n15865 , n15880 );
and ( n16110 , n15861 , n15880 );
or ( n16111 , n16108 , n16109 , n16110 );
and ( n16112 , n15776 , n15817 );
and ( n16113 , n15817 , n15846 );
and ( n16114 , n15776 , n15846 );
or ( n16115 , n16112 , n16113 , n16114 );
xor ( n16116 , n16111 , n16115 );
and ( n16117 , n15838 , n15839 );
and ( n16118 , n15839 , n15844 );
and ( n16119 , n15838 , n15844 );
or ( n16120 , n16117 , n16118 , n16119 );
and ( n16121 , n15790 , n15801 );
and ( n16122 , n15801 , n15816 );
and ( n16123 , n15790 , n15816 );
or ( n16124 , n16121 , n16122 , n16123 );
xor ( n16125 , n16120 , n16124 );
and ( n16126 , n15780 , n15784 );
and ( n16127 , n15784 , n15789 );
and ( n16128 , n15780 , n15789 );
or ( n16129 , n16126 , n16127 , n16128 );
and ( n16130 , n15791 , n15795 );
and ( n16131 , n15795 , n15800 );
and ( n16132 , n15791 , n15800 );
or ( n16133 , n16130 , n16131 , n16132 );
xor ( n16134 , n16129 , n16133 );
and ( n16135 , n15826 , n15830 );
and ( n16136 , n15830 , n15832 );
and ( n16137 , n15826 , n15832 );
or ( n16138 , n16135 , n16136 , n16137 );
xor ( n16139 , n16134 , n16138 );
xor ( n16140 , n16125 , n16139 );
xor ( n16141 , n16116 , n16140 );
xor ( n16142 , n16107 , n16141 );
xor ( n16143 , n16031 , n16142 );
and ( n16144 , n15768 , n15883 );
xor ( n16145 , n16143 , n16144 );
xor ( n16146 , n16027 , n16145 );
and ( n16147 , n15886 , n15887 );
and ( n16148 , n15888 , n15891 );
or ( n16149 , n16147 , n16148 );
xor ( n16150 , n16146 , n16149 );
buf ( n16151 , n16150 );
and ( n16152 , n16013 , n16014 );
and ( n16153 , n15901 , n15976 );
and ( n16154 , n15976 , n16011 );
and ( n16155 , n15901 , n16011 );
or ( n16156 , n16153 , n16154 , n16155 );
and ( n16157 , n15981 , n15985 );
and ( n16158 , n15985 , n16010 );
and ( n16159 , n15981 , n16010 );
or ( n16160 , n16157 , n16158 , n16159 );
and ( n16161 , n15951 , n15962 );
and ( n16162 , n15962 , n15974 );
and ( n16163 , n15951 , n15974 );
or ( n16164 , n16161 , n16162 , n16163 );
and ( n16165 , n15935 , n15939 );
and ( n16166 , n15939 , n15944 );
and ( n16167 , n15935 , n15944 );
or ( n16168 , n16165 , n16166 , n16167 );
and ( n16169 , n12899 , n7948 );
not ( n16170 , n16169 );
xnor ( n16171 , n16170 , n7938 );
and ( n16172 , n11539 , n8606 );
and ( n16173 , n11850 , n8431 );
nor ( n16174 , n16172 , n16173 );
xnor ( n16175 , n16174 , n8612 );
xor ( n16176 , n16171 , n16175 );
and ( n16177 , n7791 , n12905 );
xor ( n16178 , n16176 , n16177 );
xor ( n16179 , n16168 , n16178 );
and ( n16180 , n10982 , n8992 );
and ( n16181 , n11274 , n8792 );
nor ( n16182 , n16180 , n16181 );
xnor ( n16183 , n16182 , n8998 );
and ( n16184 , n9018 , n11052 );
and ( n16185 , n9240 , n10674 );
nor ( n16186 , n16184 , n16185 );
xnor ( n16187 , n16186 , n10952 );
xor ( n16188 , n16183 , n16187 );
and ( n16189 , n8643 , n11566 );
and ( n16190 , n8781 , n11300 );
nor ( n16191 , n16189 , n16190 );
xnor ( n16192 , n16191 , n11572 );
xor ( n16193 , n16188 , n16192 );
xor ( n16194 , n16179 , n16193 );
xor ( n16195 , n16164 , n16194 );
and ( n16196 , n15999 , n16003 );
and ( n16197 , n16003 , n16008 );
and ( n16198 , n15999 , n16008 );
or ( n16199 , n16196 , n16197 , n16198 );
and ( n16200 , n10466 , n9426 );
and ( n16201 , n10679 , n9251 );
nor ( n16202 , n16200 , n16201 );
xnor ( n16203 , n16202 , n9432 );
and ( n16204 , n8241 , n12194 );
and ( n16205 , n8420 , n11890 );
nor ( n16206 , n16204 , n16205 );
xnor ( n16207 , n16206 , n12184 );
xor ( n16208 , n16203 , n16207 );
and ( n16209 , n7966 , n12957 );
and ( n16210 , n8116 , n12511 );
nor ( n16211 , n16209 , n16210 );
xnor ( n16212 , n16211 , n12908 );
xor ( n16213 , n16208 , n16212 );
xor ( n16214 , n16199 , n16213 );
and ( n16215 , n12175 , n8294 );
and ( n16216 , n12500 , n8110 );
nor ( n16217 , n16215 , n16216 );
xnor ( n16218 , n16217 , n8250 );
not ( n16219 , n16218 );
and ( n16220 , n9964 , n9920 );
and ( n16221 , n10211 , n9671 );
nor ( n16222 , n16220 , n16221 );
xnor ( n16223 , n16222 , n9926 );
xor ( n16224 , n16219 , n16223 );
and ( n16225 , n9438 , n10477 );
and ( n16226 , n9660 , n10205 );
nor ( n16227 , n16225 , n16226 );
xnor ( n16228 , n16227 , n10426 );
xor ( n16229 , n16224 , n16228 );
xor ( n16230 , n16214 , n16229 );
xor ( n16231 , n16195 , n16230 );
xor ( n16232 , n16160 , n16231 );
and ( n16233 , n15990 , n15994 );
and ( n16234 , n15994 , n16009 );
and ( n16235 , n15990 , n16009 );
or ( n16236 , n16233 , n16234 , n16235 );
and ( n16237 , n15905 , n15946 );
and ( n16238 , n15946 , n15975 );
and ( n16239 , n15905 , n15975 );
or ( n16240 , n16237 , n16238 , n16239 );
xor ( n16241 , n16236 , n16240 );
and ( n16242 , n15967 , n15968 );
and ( n16243 , n15968 , n15973 );
and ( n16244 , n15967 , n15973 );
or ( n16245 , n16242 , n16243 , n16244 );
and ( n16246 , n15919 , n15930 );
and ( n16247 , n15930 , n15945 );
and ( n16248 , n15919 , n15945 );
or ( n16249 , n16246 , n16247 , n16248 );
xor ( n16250 , n16245 , n16249 );
and ( n16251 , n15909 , n15913 );
and ( n16252 , n15913 , n15918 );
and ( n16253 , n15909 , n15918 );
or ( n16254 , n16251 , n16252 , n16253 );
and ( n16255 , n15920 , n15924 );
and ( n16256 , n15924 , n15929 );
and ( n16257 , n15920 , n15929 );
or ( n16258 , n16255 , n16256 , n16257 );
xor ( n16259 , n16254 , n16258 );
and ( n16260 , n15955 , n15959 );
and ( n16261 , n15959 , n15961 );
and ( n16262 , n15955 , n15961 );
or ( n16263 , n16260 , n16261 , n16262 );
xor ( n16264 , n16259 , n16263 );
xor ( n16265 , n16250 , n16264 );
xor ( n16266 , n16241 , n16265 );
xor ( n16267 , n16232 , n16266 );
xor ( n16268 , n16156 , n16267 );
and ( n16269 , n15897 , n16012 );
xor ( n16270 , n16268 , n16269 );
xor ( n16271 , n16152 , n16270 );
and ( n16272 , n16015 , n16016 );
and ( n16273 , n16017 , n16020 );
or ( n16274 , n16272 , n16273 );
xor ( n16275 , n16271 , n16274 );
buf ( n16276 , n16275 );
not ( n16277 , n831 );
and ( n16278 , n16277 , n16151 );
and ( n16279 , n16276 , n831 );
or ( n16280 , n16278 , n16279 );
and ( n16281 , n16143 , n16144 );
and ( n16282 , n16035 , n16106 );
and ( n16283 , n16106 , n16141 );
and ( n16284 , n16035 , n16141 );
or ( n16285 , n16282 , n16283 , n16284 );
and ( n16286 , n16111 , n16115 );
and ( n16287 , n16115 , n16140 );
and ( n16288 , n16111 , n16140 );
or ( n16289 , n16286 , n16287 , n16288 );
and ( n16290 , n16074 , n16088 );
and ( n16291 , n16088 , n16104 );
and ( n16292 , n16074 , n16104 );
or ( n16293 , n16290 , n16291 , n16292 );
and ( n16294 , n16094 , n16098 );
and ( n16295 , n16098 , n16103 );
and ( n16296 , n16094 , n16103 );
or ( n16297 , n16294 , n16295 , n16296 );
not ( n16298 , n7863 );
and ( n16299 , n12339 , n8209 );
and ( n16300 , n12724 , n8039 );
nor ( n16301 , n16299 , n16300 );
xnor ( n16302 , n16301 , n8165 );
xor ( n16303 , n16298 , n16302 );
and ( n16304 , n11133 , n8887 );
and ( n16305 , n11384 , n8701 );
nor ( n16306 , n16304 , n16305 );
xnor ( n16307 , n16306 , n8893 );
xor ( n16308 , n16303 , n16307 );
xor ( n16309 , n16297 , n16308 );
and ( n16310 , n10548 , n9311 );
and ( n16311 , n10837 , n9150 );
nor ( n16312 , n16310 , n16311 );
xnor ( n16313 , n16312 , n9317 );
and ( n16314 , n9139 , n10907 );
and ( n16315 , n9323 , n10543 );
nor ( n16316 , n16314 , n16315 );
xnor ( n16317 , n16316 , n10807 );
xor ( n16318 , n16313 , n16317 );
and ( n16319 , n8690 , n11411 );
and ( n16320 , n8913 , n11159 );
nor ( n16321 , n16319 , n16320 );
xnor ( n16322 , n16321 , n11417 );
xor ( n16323 , n16318 , n16322 );
xor ( n16324 , n16309 , n16323 );
xor ( n16325 , n16293 , n16324 );
and ( n16326 , n16078 , n16082 );
and ( n16327 , n16082 , n16087 );
and ( n16328 , n16078 , n16087 );
or ( n16329 , n16326 , n16327 , n16328 );
and ( n16330 , n10090 , n9795 );
and ( n16331 , n10331 , n9560 );
nor ( n16332 , n16330 , n16331 );
xnor ( n16333 , n16332 , n9801 );
and ( n16334 , n9549 , n10342 );
and ( n16335 , n9839 , n10084 );
nor ( n16336 , n16334 , n16335 );
xnor ( n16337 , n16336 , n10291 );
xor ( n16338 , n16333 , n16337 );
and ( n16339 , n7891 , n12730 );
xor ( n16340 , n16338 , n16339 );
xor ( n16341 , n16329 , n16340 );
and ( n16342 , n11699 , n8511 );
and ( n16343 , n12010 , n8350 );
nor ( n16344 , n16342 , n16343 );
xnor ( n16345 , n16344 , n8517 );
and ( n16346 , n8339 , n12029 );
and ( n16347 , n8548 , n11739 );
nor ( n16348 , n16346 , n16347 );
xnor ( n16349 , n16348 , n12019 );
xor ( n16350 , n16345 , n16349 );
and ( n16351 , n8045 , n12782 );
and ( n16352 , n8156 , n12350 );
nor ( n16353 , n16351 , n16352 );
xnor ( n16354 , n16353 , n12733 );
xor ( n16355 , n16350 , n16354 );
xor ( n16356 , n16341 , n16355 );
xor ( n16357 , n16325 , n16356 );
xor ( n16358 , n16289 , n16357 );
and ( n16359 , n16120 , n16124 );
and ( n16360 , n16124 , n16139 );
and ( n16361 , n16120 , n16139 );
or ( n16362 , n16359 , n16360 , n16361 );
and ( n16363 , n16039 , n16069 );
and ( n16364 , n16069 , n16105 );
and ( n16365 , n16039 , n16105 );
or ( n16366 , n16363 , n16364 , n16365 );
xor ( n16367 , n16362 , n16366 );
and ( n16368 , n16129 , n16133 );
and ( n16369 , n16133 , n16138 );
and ( n16370 , n16129 , n16138 );
or ( n16371 , n16368 , n16369 , n16370 );
and ( n16372 , n16043 , n16053 );
and ( n16373 , n16053 , n16068 );
and ( n16374 , n16043 , n16068 );
or ( n16375 , n16372 , n16373 , n16374 );
xor ( n16376 , n16371 , n16375 );
and ( n16377 , n16046 , n16050 );
and ( n16378 , n16050 , n16052 );
and ( n16379 , n16046 , n16052 );
or ( n16380 , n16377 , n16378 , n16379 );
and ( n16381 , n16058 , n16062 );
and ( n16382 , n16062 , n16067 );
and ( n16383 , n16058 , n16067 );
or ( n16384 , n16381 , n16382 , n16383 );
xor ( n16385 , n16380 , n16384 );
buf ( n16386 , n16093 );
xor ( n16387 , n16385 , n16386 );
xor ( n16388 , n16376 , n16387 );
xor ( n16389 , n16367 , n16388 );
xor ( n16390 , n16358 , n16389 );
xor ( n16391 , n16285 , n16390 );
and ( n16392 , n16031 , n16142 );
xor ( n16393 , n16391 , n16392 );
xor ( n16394 , n16281 , n16393 );
and ( n16395 , n16027 , n16145 );
and ( n16396 , n16146 , n16149 );
or ( n16397 , n16395 , n16396 );
xor ( n16398 , n16394 , n16397 );
buf ( n16399 , n16398 );
and ( n16400 , n16268 , n16269 );
and ( n16401 , n16160 , n16231 );
and ( n16402 , n16231 , n16266 );
and ( n16403 , n16160 , n16266 );
or ( n16404 , n16401 , n16402 , n16403 );
and ( n16405 , n16236 , n16240 );
and ( n16406 , n16240 , n16265 );
and ( n16407 , n16236 , n16265 );
or ( n16408 , n16405 , n16406 , n16407 );
and ( n16409 , n16199 , n16213 );
and ( n16410 , n16213 , n16229 );
and ( n16411 , n16199 , n16229 );
or ( n16412 , n16409 , n16410 , n16411 );
and ( n16413 , n16219 , n16223 );
and ( n16414 , n16223 , n16228 );
and ( n16415 , n16219 , n16228 );
or ( n16416 , n16413 , n16414 , n16415 );
not ( n16417 , n7938 );
and ( n16418 , n12500 , n8294 );
and ( n16419 , n12899 , n8110 );
nor ( n16420 , n16418 , n16419 );
xnor ( n16421 , n16420 , n8250 );
xor ( n16422 , n16417 , n16421 );
and ( n16423 , n11274 , n8992 );
and ( n16424 , n11539 , n8792 );
nor ( n16425 , n16423 , n16424 );
xnor ( n16426 , n16425 , n8998 );
xor ( n16427 , n16422 , n16426 );
xor ( n16428 , n16416 , n16427 );
and ( n16429 , n10679 , n9426 );
and ( n16430 , n10982 , n9251 );
nor ( n16431 , n16429 , n16430 );
xnor ( n16432 , n16431 , n9432 );
and ( n16433 , n9240 , n11052 );
and ( n16434 , n9438 , n10674 );
nor ( n16435 , n16433 , n16434 );
xnor ( n16436 , n16435 , n10952 );
xor ( n16437 , n16432 , n16436 );
and ( n16438 , n8781 , n11566 );
and ( n16439 , n9018 , n11300 );
nor ( n16440 , n16438 , n16439 );
xnor ( n16441 , n16440 , n11572 );
xor ( n16442 , n16437 , n16441 );
xor ( n16443 , n16428 , n16442 );
xor ( n16444 , n16412 , n16443 );
and ( n16445 , n16203 , n16207 );
and ( n16446 , n16207 , n16212 );
and ( n16447 , n16203 , n16212 );
or ( n16448 , n16445 , n16446 , n16447 );
and ( n16449 , n10211 , n9920 );
and ( n16450 , n10466 , n9671 );
nor ( n16451 , n16449 , n16450 );
xnor ( n16452 , n16451 , n9926 );
and ( n16453 , n9660 , n10477 );
and ( n16454 , n9964 , n10205 );
nor ( n16455 , n16453 , n16454 );
xnor ( n16456 , n16455 , n10426 );
xor ( n16457 , n16452 , n16456 );
and ( n16458 , n7966 , n12905 );
xor ( n16459 , n16457 , n16458 );
xor ( n16460 , n16448 , n16459 );
and ( n16461 , n11850 , n8606 );
and ( n16462 , n12175 , n8431 );
nor ( n16463 , n16461 , n16462 );
xnor ( n16464 , n16463 , n8612 );
and ( n16465 , n8420 , n12194 );
and ( n16466 , n8643 , n11890 );
nor ( n16467 , n16465 , n16466 );
xnor ( n16468 , n16467 , n12184 );
xor ( n16469 , n16464 , n16468 );
and ( n16470 , n8116 , n12957 );
and ( n16471 , n8241 , n12511 );
nor ( n16472 , n16470 , n16471 );
xnor ( n16473 , n16472 , n12908 );
xor ( n16474 , n16469 , n16473 );
xor ( n16475 , n16460 , n16474 );
xor ( n16476 , n16444 , n16475 );
xor ( n16477 , n16408 , n16476 );
and ( n16478 , n16245 , n16249 );
and ( n16479 , n16249 , n16264 );
and ( n16480 , n16245 , n16264 );
or ( n16481 , n16478 , n16479 , n16480 );
and ( n16482 , n16164 , n16194 );
and ( n16483 , n16194 , n16230 );
and ( n16484 , n16164 , n16230 );
or ( n16485 , n16482 , n16483 , n16484 );
xor ( n16486 , n16481 , n16485 );
and ( n16487 , n16254 , n16258 );
and ( n16488 , n16258 , n16263 );
and ( n16489 , n16254 , n16263 );
or ( n16490 , n16487 , n16488 , n16489 );
and ( n16491 , n16168 , n16178 );
and ( n16492 , n16178 , n16193 );
and ( n16493 , n16168 , n16193 );
or ( n16494 , n16491 , n16492 , n16493 );
xor ( n16495 , n16490 , n16494 );
and ( n16496 , n16171 , n16175 );
and ( n16497 , n16175 , n16177 );
and ( n16498 , n16171 , n16177 );
or ( n16499 , n16496 , n16497 , n16498 );
and ( n16500 , n16183 , n16187 );
and ( n16501 , n16187 , n16192 );
and ( n16502 , n16183 , n16192 );
or ( n16503 , n16500 , n16501 , n16502 );
xor ( n16504 , n16499 , n16503 );
buf ( n16505 , n16218 );
xor ( n16506 , n16504 , n16505 );
xor ( n16507 , n16495 , n16506 );
xor ( n16508 , n16486 , n16507 );
xor ( n16509 , n16477 , n16508 );
xor ( n16510 , n16404 , n16509 );
and ( n16511 , n16156 , n16267 );
xor ( n16512 , n16510 , n16511 );
xor ( n16513 , n16400 , n16512 );
and ( n16514 , n16152 , n16270 );
and ( n16515 , n16271 , n16274 );
or ( n16516 , n16514 , n16515 );
xor ( n16517 , n16513 , n16516 );
buf ( n16518 , n16517 );
not ( n16519 , n831 );
and ( n16520 , n16519 , n16399 );
and ( n16521 , n16518 , n831 );
or ( n16522 , n16520 , n16521 );
and ( n16523 , n16391 , n16392 );
and ( n16524 , n16289 , n16357 );
and ( n16525 , n16357 , n16389 );
and ( n16526 , n16289 , n16389 );
or ( n16527 , n16524 , n16525 , n16526 );
and ( n16528 , n16362 , n16366 );
and ( n16529 , n16366 , n16388 );
and ( n16530 , n16362 , n16388 );
or ( n16531 , n16528 , n16529 , n16530 );
and ( n16532 , n16297 , n16308 );
and ( n16533 , n16308 , n16323 );
and ( n16534 , n16297 , n16323 );
or ( n16535 , n16532 , n16533 , n16534 );
and ( n16536 , n16329 , n16340 );
and ( n16537 , n16340 , n16355 );
and ( n16538 , n16329 , n16355 );
or ( n16539 , n16536 , n16537 , n16538 );
xor ( n16540 , n16535 , n16539 );
and ( n16541 , n10331 , n9795 );
and ( n16542 , n10548 , n9560 );
nor ( n16543 , n16541 , n16542 );
xnor ( n16544 , n16543 , n9801 );
and ( n16545 , n8156 , n12782 );
and ( n16546 , n8339 , n12350 );
nor ( n16547 , n16545 , n16546 );
xnor ( n16548 , n16547 , n12733 );
xor ( n16549 , n16544 , n16548 );
and ( n16550 , n8045 , n12730 );
xor ( n16551 , n16549 , n16550 );
and ( n16552 , n10837 , n9311 );
and ( n16553 , n11133 , n9150 );
nor ( n16554 , n16552 , n16553 );
xnor ( n16555 , n16554 , n9317 );
and ( n16556 , n8913 , n11411 );
and ( n16557 , n9139 , n11159 );
nor ( n16558 , n16556 , n16557 );
xnor ( n16559 , n16558 , n11417 );
xor ( n16560 , n16555 , n16559 );
and ( n16561 , n8548 , n12029 );
and ( n16562 , n8690 , n11739 );
nor ( n16563 , n16561 , n16562 );
xnor ( n16564 , n16563 , n12019 );
xor ( n16565 , n16560 , n16564 );
xor ( n16566 , n16551 , n16565 );
and ( n16567 , n12724 , n8209 );
not ( n16568 , n16567 );
xnor ( n16569 , n16568 , n8165 );
and ( n16570 , n11384 , n8887 );
and ( n16571 , n11699 , n8701 );
nor ( n16572 , n16570 , n16571 );
xnor ( n16573 , n16572 , n8893 );
xor ( n16574 , n16569 , n16573 );
and ( n16575 , n9839 , n10342 );
and ( n16576 , n10090 , n10084 );
nor ( n16577 , n16575 , n16576 );
xnor ( n16578 , n16577 , n10291 );
xor ( n16579 , n16574 , n16578 );
xor ( n16580 , n16566 , n16579 );
xor ( n16581 , n16540 , n16580 );
xor ( n16582 , n16531 , n16581 );
and ( n16583 , n16371 , n16375 );
and ( n16584 , n16375 , n16387 );
and ( n16585 , n16371 , n16387 );
or ( n16586 , n16583 , n16584 , n16585 );
and ( n16587 , n16293 , n16324 );
and ( n16588 , n16324 , n16356 );
and ( n16589 , n16293 , n16356 );
or ( n16590 , n16587 , n16588 , n16589 );
xor ( n16591 , n16586 , n16590 );
and ( n16592 , n16380 , n16384 );
and ( n16593 , n16384 , n16386 );
and ( n16594 , n16380 , n16386 );
or ( n16595 , n16592 , n16593 , n16594 );
and ( n16596 , n16298 , n16302 );
and ( n16597 , n16302 , n16307 );
and ( n16598 , n16298 , n16307 );
or ( n16599 , n16596 , n16597 , n16598 );
and ( n16600 , n16313 , n16317 );
and ( n16601 , n16317 , n16322 );
and ( n16602 , n16313 , n16322 );
or ( n16603 , n16600 , n16601 , n16602 );
xor ( n16604 , n16599 , n16603 );
and ( n16605 , n16333 , n16337 );
and ( n16606 , n16337 , n16339 );
and ( n16607 , n16333 , n16339 );
or ( n16608 , n16605 , n16606 , n16607 );
xor ( n16609 , n16604 , n16608 );
xor ( n16610 , n16595 , n16609 );
and ( n16611 , n16345 , n16349 );
and ( n16612 , n16349 , n16354 );
and ( n16613 , n16345 , n16354 );
or ( n16614 , n16611 , n16612 , n16613 );
and ( n16615 , n12010 , n8511 );
and ( n16616 , n12339 , n8350 );
nor ( n16617 , n16615 , n16616 );
xnor ( n16618 , n16617 , n8517 );
not ( n16619 , n16618 );
xor ( n16620 , n16614 , n16619 );
and ( n16621 , n9323 , n10907 );
and ( n16622 , n9549 , n10543 );
nor ( n16623 , n16621 , n16622 );
xnor ( n16624 , n16623 , n10807 );
xor ( n16625 , n16620 , n16624 );
xor ( n16626 , n16610 , n16625 );
xor ( n16627 , n16591 , n16626 );
xor ( n16628 , n16582 , n16627 );
xor ( n16629 , n16527 , n16628 );
and ( n16630 , n16285 , n16390 );
xor ( n16631 , n16629 , n16630 );
xor ( n16632 , n16523 , n16631 );
and ( n16633 , n16281 , n16393 );
and ( n16634 , n16394 , n16397 );
or ( n16635 , n16633 , n16634 );
xor ( n16636 , n16632 , n16635 );
buf ( n16637 , n16636 );
and ( n16638 , n16510 , n16511 );
and ( n16639 , n16408 , n16476 );
and ( n16640 , n16476 , n16508 );
and ( n16641 , n16408 , n16508 );
or ( n16642 , n16639 , n16640 , n16641 );
and ( n16643 , n16481 , n16485 );
and ( n16644 , n16485 , n16507 );
and ( n16645 , n16481 , n16507 );
or ( n16646 , n16643 , n16644 , n16645 );
and ( n16647 , n16416 , n16427 );
and ( n16648 , n16427 , n16442 );
and ( n16649 , n16416 , n16442 );
or ( n16650 , n16647 , n16648 , n16649 );
and ( n16651 , n16448 , n16459 );
and ( n16652 , n16459 , n16474 );
and ( n16653 , n16448 , n16474 );
or ( n16654 , n16651 , n16652 , n16653 );
xor ( n16655 , n16650 , n16654 );
and ( n16656 , n10466 , n9920 );
and ( n16657 , n10679 , n9671 );
nor ( n16658 , n16656 , n16657 );
xnor ( n16659 , n16658 , n9926 );
and ( n16660 , n8241 , n12957 );
and ( n16661 , n8420 , n12511 );
nor ( n16662 , n16660 , n16661 );
xnor ( n16663 , n16662 , n12908 );
xor ( n16664 , n16659 , n16663 );
and ( n16665 , n8116 , n12905 );
xor ( n16666 , n16664 , n16665 );
and ( n16667 , n10982 , n9426 );
and ( n16668 , n11274 , n9251 );
nor ( n16669 , n16667 , n16668 );
xnor ( n16670 , n16669 , n9432 );
and ( n16671 , n9018 , n11566 );
and ( n16672 , n9240 , n11300 );
nor ( n16673 , n16671 , n16672 );
xnor ( n16674 , n16673 , n11572 );
xor ( n16675 , n16670 , n16674 );
and ( n16676 , n8643 , n12194 );
and ( n16677 , n8781 , n11890 );
nor ( n16678 , n16676 , n16677 );
xnor ( n16679 , n16678 , n12184 );
xor ( n16680 , n16675 , n16679 );
xor ( n16681 , n16666 , n16680 );
and ( n16682 , n12899 , n8294 );
not ( n16683 , n16682 );
xnor ( n16684 , n16683 , n8250 );
and ( n16685 , n11539 , n8992 );
and ( n16686 , n11850 , n8792 );
nor ( n16687 , n16685 , n16686 );
xnor ( n16688 , n16687 , n8998 );
xor ( n16689 , n16684 , n16688 );
and ( n16690 , n9964 , n10477 );
and ( n16691 , n10211 , n10205 );
nor ( n16692 , n16690 , n16691 );
xnor ( n16693 , n16692 , n10426 );
xor ( n16694 , n16689 , n16693 );
xor ( n16695 , n16681 , n16694 );
xor ( n16696 , n16655 , n16695 );
xor ( n16697 , n16646 , n16696 );
and ( n16698 , n16490 , n16494 );
and ( n16699 , n16494 , n16506 );
and ( n16700 , n16490 , n16506 );
or ( n16701 , n16698 , n16699 , n16700 );
and ( n16702 , n16412 , n16443 );
and ( n16703 , n16443 , n16475 );
and ( n16704 , n16412 , n16475 );
or ( n16705 , n16702 , n16703 , n16704 );
xor ( n16706 , n16701 , n16705 );
and ( n16707 , n16499 , n16503 );
and ( n16708 , n16503 , n16505 );
and ( n16709 , n16499 , n16505 );
or ( n16710 , n16707 , n16708 , n16709 );
and ( n16711 , n16417 , n16421 );
and ( n16712 , n16421 , n16426 );
and ( n16713 , n16417 , n16426 );
or ( n16714 , n16711 , n16712 , n16713 );
and ( n16715 , n16432 , n16436 );
and ( n16716 , n16436 , n16441 );
and ( n16717 , n16432 , n16441 );
or ( n16718 , n16715 , n16716 , n16717 );
xor ( n16719 , n16714 , n16718 );
and ( n16720 , n16452 , n16456 );
and ( n16721 , n16456 , n16458 );
and ( n16722 , n16452 , n16458 );
or ( n16723 , n16720 , n16721 , n16722 );
xor ( n16724 , n16719 , n16723 );
xor ( n16725 , n16710 , n16724 );
and ( n16726 , n16464 , n16468 );
and ( n16727 , n16468 , n16473 );
and ( n16728 , n16464 , n16473 );
or ( n16729 , n16726 , n16727 , n16728 );
and ( n16730 , n12175 , n8606 );
and ( n16731 , n12500 , n8431 );
nor ( n16732 , n16730 , n16731 );
xnor ( n16733 , n16732 , n8612 );
not ( n16734 , n16733 );
xor ( n16735 , n16729 , n16734 );
and ( n16736 , n9438 , n11052 );
and ( n16737 , n9660 , n10674 );
nor ( n16738 , n16736 , n16737 );
xnor ( n16739 , n16738 , n10952 );
xor ( n16740 , n16735 , n16739 );
xor ( n16741 , n16725 , n16740 );
xor ( n16742 , n16706 , n16741 );
xor ( n16743 , n16697 , n16742 );
xor ( n16744 , n16642 , n16743 );
and ( n16745 , n16404 , n16509 );
xor ( n16746 , n16744 , n16745 );
xor ( n16747 , n16638 , n16746 );
and ( n16748 , n16400 , n16512 );
and ( n16749 , n16513 , n16516 );
or ( n16750 , n16748 , n16749 );
xor ( n16751 , n16747 , n16750 );
buf ( n16752 , n16751 );
not ( n16753 , n831 );
and ( n16754 , n16753 , n16637 );
and ( n16755 , n16752 , n831 );
or ( n16756 , n16754 , n16755 );
and ( n16757 , n16629 , n16630 );
and ( n16758 , n16531 , n16581 );
and ( n16759 , n16581 , n16627 );
and ( n16760 , n16531 , n16627 );
or ( n16761 , n16758 , n16759 , n16760 );
and ( n16762 , n16535 , n16539 );
and ( n16763 , n16539 , n16580 );
and ( n16764 , n16535 , n16580 );
or ( n16765 , n16762 , n16763 , n16764 );
and ( n16766 , n16586 , n16590 );
and ( n16767 , n16590 , n16626 );
and ( n16768 , n16586 , n16626 );
or ( n16769 , n16766 , n16767 , n16768 );
xor ( n16770 , n16765 , n16769 );
and ( n16771 , n16595 , n16609 );
and ( n16772 , n16609 , n16625 );
and ( n16773 , n16595 , n16625 );
or ( n16774 , n16771 , n16772 , n16773 );
and ( n16775 , n16599 , n16603 );
and ( n16776 , n16603 , n16608 );
and ( n16777 , n16599 , n16608 );
or ( n16778 , n16775 , n16776 , n16777 );
and ( n16779 , n16614 , n16619 );
and ( n16780 , n16619 , n16624 );
and ( n16781 , n16614 , n16624 );
or ( n16782 , n16779 , n16780 , n16781 );
xor ( n16783 , n16778 , n16782 );
buf ( n16784 , n16618 );
and ( n16785 , n10090 , n10342 );
and ( n16786 , n10331 , n10084 );
nor ( n16787 , n16785 , n16786 );
xnor ( n16788 , n16787 , n10291 );
xor ( n16789 , n16784 , n16788 );
and ( n16790 , n9549 , n10907 );
and ( n16791 , n9839 , n10543 );
nor ( n16792 , n16790 , n16791 );
xnor ( n16793 , n16792 , n10807 );
xor ( n16794 , n16789 , n16793 );
xor ( n16795 , n16783 , n16794 );
xor ( n16796 , n16774 , n16795 );
and ( n16797 , n16551 , n16565 );
and ( n16798 , n16565 , n16579 );
and ( n16799 , n16551 , n16579 );
or ( n16800 , n16797 , n16798 , n16799 );
and ( n16801 , n16544 , n16548 );
and ( n16802 , n16548 , n16550 );
and ( n16803 , n16544 , n16550 );
or ( n16804 , n16801 , n16802 , n16803 );
and ( n16805 , n16555 , n16559 );
and ( n16806 , n16559 , n16564 );
and ( n16807 , n16555 , n16564 );
or ( n16808 , n16805 , n16806 , n16807 );
xor ( n16809 , n16804 , n16808 );
and ( n16810 , n16569 , n16573 );
and ( n16811 , n16573 , n16578 );
and ( n16812 , n16569 , n16578 );
or ( n16813 , n16810 , n16811 , n16812 );
xor ( n16814 , n16809 , n16813 );
xor ( n16815 , n16800 , n16814 );
and ( n16816 , n11699 , n8887 );
and ( n16817 , n12010 , n8701 );
nor ( n16818 , n16816 , n16817 );
xnor ( n16819 , n16818 , n8893 );
and ( n16820 , n8339 , n12782 );
and ( n16821 , n8548 , n12350 );
nor ( n16822 , n16820 , n16821 );
xnor ( n16823 , n16822 , n12733 );
xor ( n16824 , n16819 , n16823 );
and ( n16825 , n8156 , n12730 );
xor ( n16826 , n16824 , n16825 );
not ( n16827 , n8165 );
and ( n16828 , n12339 , n8511 );
and ( n16829 , n12724 , n8350 );
nor ( n16830 , n16828 , n16829 );
xnor ( n16831 , n16830 , n8517 );
xor ( n16832 , n16827 , n16831 );
and ( n16833 , n11133 , n9311 );
and ( n16834 , n11384 , n9150 );
nor ( n16835 , n16833 , n16834 );
xnor ( n16836 , n16835 , n9317 );
xor ( n16837 , n16832 , n16836 );
xor ( n16838 , n16826 , n16837 );
and ( n16839 , n10548 , n9795 );
and ( n16840 , n10837 , n9560 );
nor ( n16841 , n16839 , n16840 );
xnor ( n16842 , n16841 , n9801 );
and ( n16843 , n9139 , n11411 );
and ( n16844 , n9323 , n11159 );
nor ( n16845 , n16843 , n16844 );
xnor ( n16846 , n16845 , n11417 );
xor ( n16847 , n16842 , n16846 );
and ( n16848 , n8690 , n12029 );
and ( n16849 , n8913 , n11739 );
nor ( n16850 , n16848 , n16849 );
xnor ( n16851 , n16850 , n12019 );
xor ( n16852 , n16847 , n16851 );
xor ( n16853 , n16838 , n16852 );
xor ( n16854 , n16815 , n16853 );
xor ( n16855 , n16796 , n16854 );
xor ( n16856 , n16770 , n16855 );
xor ( n16857 , n16761 , n16856 );
and ( n16858 , n16527 , n16628 );
xor ( n16859 , n16857 , n16858 );
xor ( n16860 , n16757 , n16859 );
and ( n16861 , n16523 , n16631 );
and ( n16862 , n16632 , n16635 );
or ( n16863 , n16861 , n16862 );
xor ( n16864 , n16860 , n16863 );
buf ( n16865 , n16864 );
and ( n16866 , n16744 , n16745 );
and ( n16867 , n16646 , n16696 );
and ( n16868 , n16696 , n16742 );
and ( n16869 , n16646 , n16742 );
or ( n16870 , n16867 , n16868 , n16869 );
and ( n16871 , n16650 , n16654 );
and ( n16872 , n16654 , n16695 );
and ( n16873 , n16650 , n16695 );
or ( n16874 , n16871 , n16872 , n16873 );
and ( n16875 , n16701 , n16705 );
and ( n16876 , n16705 , n16741 );
and ( n16877 , n16701 , n16741 );
or ( n16878 , n16875 , n16876 , n16877 );
xor ( n16879 , n16874 , n16878 );
and ( n16880 , n16710 , n16724 );
and ( n16881 , n16724 , n16740 );
and ( n16882 , n16710 , n16740 );
or ( n16883 , n16880 , n16881 , n16882 );
and ( n16884 , n16714 , n16718 );
and ( n16885 , n16718 , n16723 );
and ( n16886 , n16714 , n16723 );
or ( n16887 , n16884 , n16885 , n16886 );
and ( n16888 , n16729 , n16734 );
and ( n16889 , n16734 , n16739 );
and ( n16890 , n16729 , n16739 );
or ( n16891 , n16888 , n16889 , n16890 );
xor ( n16892 , n16887 , n16891 );
buf ( n16893 , n16733 );
and ( n16894 , n10211 , n10477 );
and ( n16895 , n10466 , n10205 );
nor ( n16896 , n16894 , n16895 );
xnor ( n16897 , n16896 , n10426 );
xor ( n16898 , n16893 , n16897 );
and ( n16899 , n9660 , n11052 );
and ( n16900 , n9964 , n10674 );
nor ( n16901 , n16899 , n16900 );
xnor ( n16902 , n16901 , n10952 );
xor ( n16903 , n16898 , n16902 );
xor ( n16904 , n16892 , n16903 );
xor ( n16905 , n16883 , n16904 );
and ( n16906 , n16666 , n16680 );
and ( n16907 , n16680 , n16694 );
and ( n16908 , n16666 , n16694 );
or ( n16909 , n16906 , n16907 , n16908 );
and ( n16910 , n16659 , n16663 );
and ( n16911 , n16663 , n16665 );
and ( n16912 , n16659 , n16665 );
or ( n16913 , n16910 , n16911 , n16912 );
and ( n16914 , n16670 , n16674 );
and ( n16915 , n16674 , n16679 );
and ( n16916 , n16670 , n16679 );
or ( n16917 , n16914 , n16915 , n16916 );
xor ( n16918 , n16913 , n16917 );
and ( n16919 , n16684 , n16688 );
and ( n16920 , n16688 , n16693 );
and ( n16921 , n16684 , n16693 );
or ( n16922 , n16919 , n16920 , n16921 );
xor ( n16923 , n16918 , n16922 );
xor ( n16924 , n16909 , n16923 );
and ( n16925 , n11850 , n8992 );
and ( n16926 , n12175 , n8792 );
nor ( n16927 , n16925 , n16926 );
xnor ( n16928 , n16927 , n8998 );
and ( n16929 , n8420 , n12957 );
and ( n16930 , n8643 , n12511 );
nor ( n16931 , n16929 , n16930 );
xnor ( n16932 , n16931 , n12908 );
xor ( n16933 , n16928 , n16932 );
and ( n16934 , n8241 , n12905 );
xor ( n16935 , n16933 , n16934 );
not ( n16936 , n8250 );
and ( n16937 , n12500 , n8606 );
and ( n16938 , n12899 , n8431 );
nor ( n16939 , n16937 , n16938 );
xnor ( n16940 , n16939 , n8612 );
xor ( n16941 , n16936 , n16940 );
and ( n16942 , n11274 , n9426 );
and ( n16943 , n11539 , n9251 );
nor ( n16944 , n16942 , n16943 );
xnor ( n16945 , n16944 , n9432 );
xor ( n16946 , n16941 , n16945 );
xor ( n16947 , n16935 , n16946 );
and ( n16948 , n10679 , n9920 );
and ( n16949 , n10982 , n9671 );
nor ( n16950 , n16948 , n16949 );
xnor ( n16951 , n16950 , n9926 );
and ( n16952 , n9240 , n11566 );
and ( n16953 , n9438 , n11300 );
nor ( n16954 , n16952 , n16953 );
xnor ( n16955 , n16954 , n11572 );
xor ( n16956 , n16951 , n16955 );
and ( n16957 , n8781 , n12194 );
and ( n16958 , n9018 , n11890 );
nor ( n16959 , n16957 , n16958 );
xnor ( n16960 , n16959 , n12184 );
xor ( n16961 , n16956 , n16960 );
xor ( n16962 , n16947 , n16961 );
xor ( n16963 , n16924 , n16962 );
xor ( n16964 , n16905 , n16963 );
xor ( n16965 , n16879 , n16964 );
xor ( n16966 , n16870 , n16965 );
and ( n16967 , n16642 , n16743 );
xor ( n16968 , n16966 , n16967 );
xor ( n16969 , n16866 , n16968 );
and ( n16970 , n16638 , n16746 );
and ( n16971 , n16747 , n16750 );
or ( n16972 , n16970 , n16971 );
xor ( n16973 , n16969 , n16972 );
buf ( n16974 , n16973 );
not ( n16975 , n831 );
and ( n16976 , n16975 , n16865 );
and ( n16977 , n16974 , n831 );
or ( n16978 , n16976 , n16977 );
and ( n16979 , n16857 , n16858 );
and ( n16980 , n16765 , n16769 );
and ( n16981 , n16769 , n16855 );
and ( n16982 , n16765 , n16855 );
or ( n16983 , n16980 , n16981 , n16982 );
and ( n16984 , n16774 , n16795 );
and ( n16985 , n16795 , n16854 );
and ( n16986 , n16774 , n16854 );
or ( n16987 , n16984 , n16985 , n16986 );
and ( n16988 , n16826 , n16837 );
and ( n16989 , n16837 , n16852 );
and ( n16990 , n16826 , n16852 );
or ( n16991 , n16988 , n16989 , n16990 );
and ( n16992 , n16827 , n16831 );
and ( n16993 , n16831 , n16836 );
and ( n16994 , n16827 , n16836 );
or ( n16995 , n16992 , n16993 , n16994 );
and ( n16996 , n16842 , n16846 );
and ( n16997 , n16846 , n16851 );
and ( n16998 , n16842 , n16851 );
or ( n16999 , n16996 , n16997 , n16998 );
xor ( n17000 , n16995 , n16999 );
and ( n17001 , n12724 , n8511 );
not ( n17002 , n17001 );
xnor ( n17003 , n17002 , n8517 );
not ( n17004 , n17003 );
xor ( n17005 , n17000 , n17004 );
xor ( n17006 , n16991 , n17005 );
and ( n17007 , n16819 , n16823 );
and ( n17008 , n16823 , n16825 );
and ( n17009 , n16819 , n16825 );
or ( n17010 , n17007 , n17008 , n17009 );
and ( n17011 , n10837 , n9795 );
and ( n17012 , n11133 , n9560 );
nor ( n17013 , n17011 , n17012 );
xnor ( n17014 , n17013 , n9801 );
and ( n17015 , n8913 , n12029 );
and ( n17016 , n9139 , n11739 );
nor ( n17017 , n17015 , n17016 );
xnor ( n17018 , n17017 , n12019 );
xor ( n17019 , n17014 , n17018 );
and ( n17020 , n8548 , n12782 );
and ( n17021 , n8690 , n12350 );
nor ( n17022 , n17020 , n17021 );
xnor ( n17023 , n17022 , n12733 );
xor ( n17024 , n17019 , n17023 );
xor ( n17025 , n17010 , n17024 );
and ( n17026 , n12010 , n8887 );
and ( n17027 , n12339 , n8701 );
nor ( n17028 , n17026 , n17027 );
xnor ( n17029 , n17028 , n8893 );
and ( n17030 , n10331 , n10342 );
and ( n17031 , n10548 , n10084 );
nor ( n17032 , n17030 , n17031 );
xnor ( n17033 , n17032 , n10291 );
xor ( n17034 , n17029 , n17033 );
and ( n17035 , n8339 , n12730 );
xor ( n17036 , n17034 , n17035 );
xor ( n17037 , n17025 , n17036 );
xor ( n17038 , n17006 , n17037 );
xor ( n17039 , n16987 , n17038 );
and ( n17040 , n16778 , n16782 );
and ( n17041 , n16782 , n16794 );
and ( n17042 , n16778 , n16794 );
or ( n17043 , n17040 , n17041 , n17042 );
and ( n17044 , n16800 , n16814 );
and ( n17045 , n16814 , n16853 );
and ( n17046 , n16800 , n16853 );
or ( n17047 , n17044 , n17045 , n17046 );
xor ( n17048 , n17043 , n17047 );
and ( n17049 , n16804 , n16808 );
and ( n17050 , n16808 , n16813 );
and ( n17051 , n16804 , n16813 );
or ( n17052 , n17049 , n17050 , n17051 );
and ( n17053 , n16784 , n16788 );
and ( n17054 , n16788 , n16793 );
and ( n17055 , n16784 , n16793 );
or ( n17056 , n17053 , n17054 , n17055 );
xor ( n17057 , n17052 , n17056 );
and ( n17058 , n11384 , n9311 );
and ( n17059 , n11699 , n9150 );
nor ( n17060 , n17058 , n17059 );
xnor ( n17061 , n17060 , n9317 );
and ( n17062 , n9839 , n10907 );
and ( n17063 , n10090 , n10543 );
nor ( n17064 , n17062 , n17063 );
xnor ( n17065 , n17064 , n10807 );
xor ( n17066 , n17061 , n17065 );
and ( n17067 , n9323 , n11411 );
and ( n17068 , n9549 , n11159 );
nor ( n17069 , n17067 , n17068 );
xnor ( n17070 , n17069 , n11417 );
xor ( n17071 , n17066 , n17070 );
xor ( n17072 , n17057 , n17071 );
xor ( n17073 , n17048 , n17072 );
xor ( n17074 , n17039 , n17073 );
xor ( n17075 , n16983 , n17074 );
and ( n17076 , n16761 , n16856 );
xor ( n17077 , n17075 , n17076 );
xor ( n17078 , n16979 , n17077 );
and ( n17079 , n16757 , n16859 );
and ( n17080 , n16860 , n16863 );
or ( n17081 , n17079 , n17080 );
xor ( n17082 , n17078 , n17081 );
buf ( n17083 , n17082 );
and ( n17084 , n16966 , n16967 );
and ( n17085 , n16874 , n16878 );
and ( n17086 , n16878 , n16964 );
and ( n17087 , n16874 , n16964 );
or ( n17088 , n17085 , n17086 , n17087 );
and ( n17089 , n16883 , n16904 );
and ( n17090 , n16904 , n16963 );
and ( n17091 , n16883 , n16963 );
or ( n17092 , n17089 , n17090 , n17091 );
and ( n17093 , n16935 , n16946 );
and ( n17094 , n16946 , n16961 );
and ( n17095 , n16935 , n16961 );
or ( n17096 , n17093 , n17094 , n17095 );
and ( n17097 , n16936 , n16940 );
and ( n17098 , n16940 , n16945 );
and ( n17099 , n16936 , n16945 );
or ( n17100 , n17097 , n17098 , n17099 );
and ( n17101 , n16951 , n16955 );
and ( n17102 , n16955 , n16960 );
and ( n17103 , n16951 , n16960 );
or ( n17104 , n17101 , n17102 , n17103 );
xor ( n17105 , n17100 , n17104 );
and ( n17106 , n12899 , n8606 );
not ( n17107 , n17106 );
xnor ( n17108 , n17107 , n8612 );
not ( n17109 , n17108 );
xor ( n17110 , n17105 , n17109 );
xor ( n17111 , n17096 , n17110 );
and ( n17112 , n16928 , n16932 );
and ( n17113 , n16932 , n16934 );
and ( n17114 , n16928 , n16934 );
or ( n17115 , n17112 , n17113 , n17114 );
and ( n17116 , n10982 , n9920 );
and ( n17117 , n11274 , n9671 );
nor ( n17118 , n17116 , n17117 );
xnor ( n17119 , n17118 , n9926 );
and ( n17120 , n9018 , n12194 );
and ( n17121 , n9240 , n11890 );
nor ( n17122 , n17120 , n17121 );
xnor ( n17123 , n17122 , n12184 );
xor ( n17124 , n17119 , n17123 );
and ( n17125 , n8643 , n12957 );
and ( n17126 , n8781 , n12511 );
nor ( n17127 , n17125 , n17126 );
xnor ( n17128 , n17127 , n12908 );
xor ( n17129 , n17124 , n17128 );
xor ( n17130 , n17115 , n17129 );
and ( n17131 , n12175 , n8992 );
and ( n17132 , n12500 , n8792 );
nor ( n17133 , n17131 , n17132 );
xnor ( n17134 , n17133 , n8998 );
and ( n17135 , n10466 , n10477 );
and ( n17136 , n10679 , n10205 );
nor ( n17137 , n17135 , n17136 );
xnor ( n17138 , n17137 , n10426 );
xor ( n17139 , n17134 , n17138 );
and ( n17140 , n8420 , n12905 );
xor ( n17141 , n17139 , n17140 );
xor ( n17142 , n17130 , n17141 );
xor ( n17143 , n17111 , n17142 );
xor ( n17144 , n17092 , n17143 );
and ( n17145 , n16887 , n16891 );
and ( n17146 , n16891 , n16903 );
and ( n17147 , n16887 , n16903 );
or ( n17148 , n17145 , n17146 , n17147 );
and ( n17149 , n16909 , n16923 );
and ( n17150 , n16923 , n16962 );
and ( n17151 , n16909 , n16962 );
or ( n17152 , n17149 , n17150 , n17151 );
xor ( n17153 , n17148 , n17152 );
and ( n17154 , n16913 , n16917 );
and ( n17155 , n16917 , n16922 );
and ( n17156 , n16913 , n16922 );
or ( n17157 , n17154 , n17155 , n17156 );
and ( n17158 , n16893 , n16897 );
and ( n17159 , n16897 , n16902 );
and ( n17160 , n16893 , n16902 );
or ( n17161 , n17158 , n17159 , n17160 );
xor ( n17162 , n17157 , n17161 );
and ( n17163 , n11539 , n9426 );
and ( n17164 , n11850 , n9251 );
nor ( n17165 , n17163 , n17164 );
xnor ( n17166 , n17165 , n9432 );
and ( n17167 , n9964 , n11052 );
and ( n17168 , n10211 , n10674 );
nor ( n17169 , n17167 , n17168 );
xnor ( n17170 , n17169 , n10952 );
xor ( n17171 , n17166 , n17170 );
and ( n17172 , n9438 , n11566 );
and ( n17173 , n9660 , n11300 );
nor ( n17174 , n17172 , n17173 );
xnor ( n17175 , n17174 , n11572 );
xor ( n17176 , n17171 , n17175 );
xor ( n17177 , n17162 , n17176 );
xor ( n17178 , n17153 , n17177 );
xor ( n17179 , n17144 , n17178 );
xor ( n17180 , n17088 , n17179 );
and ( n17181 , n16870 , n16965 );
xor ( n17182 , n17180 , n17181 );
xor ( n17183 , n17084 , n17182 );
and ( n17184 , n16866 , n16968 );
and ( n17185 , n16969 , n16972 );
or ( n17186 , n17184 , n17185 );
xor ( n17187 , n17183 , n17186 );
buf ( n17188 , n17187 );
not ( n17189 , n831 );
and ( n17190 , n17189 , n17083 );
and ( n17191 , n17188 , n831 );
or ( n17192 , n17190 , n17191 );
and ( n17193 , n16987 , n17038 );
and ( n17194 , n17038 , n17073 );
and ( n17195 , n16987 , n17073 );
or ( n17196 , n17193 , n17194 , n17195 );
and ( n17197 , n17043 , n17047 );
and ( n17198 , n17047 , n17072 );
and ( n17199 , n17043 , n17072 );
or ( n17200 , n17197 , n17198 , n17199 );
and ( n17201 , n16995 , n16999 );
and ( n17202 , n16999 , n17004 );
and ( n17203 , n16995 , n17004 );
or ( n17204 , n17201 , n17202 , n17203 );
and ( n17205 , n17010 , n17024 );
and ( n17206 , n17024 , n17036 );
and ( n17207 , n17010 , n17036 );
or ( n17208 , n17205 , n17206 , n17207 );
xor ( n17209 , n17204 , n17208 );
and ( n17210 , n17029 , n17033 );
and ( n17211 , n17033 , n17035 );
and ( n17212 , n17029 , n17035 );
or ( n17213 , n17210 , n17211 , n17212 );
and ( n17214 , n17061 , n17065 );
and ( n17215 , n17065 , n17070 );
and ( n17216 , n17061 , n17070 );
or ( n17217 , n17214 , n17215 , n17216 );
xor ( n17218 , n17213 , n17217 );
and ( n17219 , n11699 , n9311 );
and ( n17220 , n12010 , n9150 );
nor ( n17221 , n17219 , n17220 );
xnor ( n17222 , n17221 , n9317 );
and ( n17223 , n10090 , n10907 );
and ( n17224 , n10331 , n10543 );
nor ( n17225 , n17223 , n17224 );
xnor ( n17226 , n17225 , n10807 );
xor ( n17227 , n17222 , n17226 );
and ( n17228 , n8548 , n12730 );
xor ( n17229 , n17227 , n17228 );
xor ( n17230 , n17218 , n17229 );
xor ( n17231 , n17209 , n17230 );
xor ( n17232 , n17200 , n17231 );
and ( n17233 , n17052 , n17056 );
and ( n17234 , n17056 , n17071 );
and ( n17235 , n17052 , n17071 );
or ( n17236 , n17233 , n17234 , n17235 );
and ( n17237 , n16991 , n17005 );
and ( n17238 , n17005 , n17037 );
and ( n17239 , n16991 , n17037 );
or ( n17240 , n17237 , n17238 , n17239 );
xor ( n17241 , n17236 , n17240 );
and ( n17242 , n10548 , n10342 );
and ( n17243 , n10837 , n10084 );
nor ( n17244 , n17242 , n17243 );
xnor ( n17245 , n17244 , n10291 );
and ( n17246 , n9139 , n12029 );
and ( n17247 , n9323 , n11739 );
nor ( n17248 , n17246 , n17247 );
xnor ( n17249 , n17248 , n12019 );
xor ( n17250 , n17245 , n17249 );
and ( n17251 , n8690 , n12782 );
and ( n17252 , n8913 , n12350 );
nor ( n17253 , n17251 , n17252 );
xnor ( n17254 , n17253 , n12733 );
xor ( n17255 , n17250 , n17254 );
not ( n17256 , n8517 );
and ( n17257 , n12339 , n8887 );
and ( n17258 , n12724 , n8701 );
nor ( n17259 , n17257 , n17258 );
xnor ( n17260 , n17259 , n8893 );
xor ( n17261 , n17256 , n17260 );
and ( n17262 , n11133 , n9795 );
and ( n17263 , n11384 , n9560 );
nor ( n17264 , n17262 , n17263 );
xnor ( n17265 , n17264 , n9801 );
xor ( n17266 , n17261 , n17265 );
xor ( n17267 , n17255 , n17266 );
and ( n17268 , n17014 , n17018 );
and ( n17269 , n17018 , n17023 );
and ( n17270 , n17014 , n17023 );
or ( n17271 , n17268 , n17269 , n17270 );
buf ( n17272 , n17003 );
xor ( n17273 , n17271 , n17272 );
and ( n17274 , n9549 , n11411 );
and ( n17275 , n9839 , n11159 );
nor ( n17276 , n17274 , n17275 );
xnor ( n17277 , n17276 , n11417 );
xor ( n17278 , n17273 , n17277 );
xor ( n17279 , n17267 , n17278 );
xor ( n17280 , n17241 , n17279 );
xor ( n17281 , n17232 , n17280 );
xor ( n17282 , n17196 , n17281 );
and ( n17283 , n16983 , n17074 );
xor ( n17284 , n17282 , n17283 );
and ( n17285 , n17075 , n17076 );
xor ( n17286 , n17284 , n17285 );
and ( n17287 , n16979 , n17077 );
and ( n17288 , n17078 , n17081 );
or ( n17289 , n17287 , n17288 );
xor ( n17290 , n17286 , n17289 );
buf ( n17291 , n17290 );
and ( n17292 , n17092 , n17143 );
and ( n17293 , n17143 , n17178 );
and ( n17294 , n17092 , n17178 );
or ( n17295 , n17292 , n17293 , n17294 );
and ( n17296 , n17148 , n17152 );
and ( n17297 , n17152 , n17177 );
and ( n17298 , n17148 , n17177 );
or ( n17299 , n17296 , n17297 , n17298 );
and ( n17300 , n17100 , n17104 );
and ( n17301 , n17104 , n17109 );
and ( n17302 , n17100 , n17109 );
or ( n17303 , n17300 , n17301 , n17302 );
and ( n17304 , n17115 , n17129 );
and ( n17305 , n17129 , n17141 );
and ( n17306 , n17115 , n17141 );
or ( n17307 , n17304 , n17305 , n17306 );
xor ( n17308 , n17303 , n17307 );
and ( n17309 , n17134 , n17138 );
and ( n17310 , n17138 , n17140 );
and ( n17311 , n17134 , n17140 );
or ( n17312 , n17309 , n17310 , n17311 );
and ( n17313 , n17166 , n17170 );
and ( n17314 , n17170 , n17175 );
and ( n17315 , n17166 , n17175 );
or ( n17316 , n17313 , n17314 , n17315 );
xor ( n17317 , n17312 , n17316 );
and ( n17318 , n11850 , n9426 );
and ( n17319 , n12175 , n9251 );
nor ( n17320 , n17318 , n17319 );
xnor ( n17321 , n17320 , n9432 );
and ( n17322 , n10211 , n11052 );
and ( n17323 , n10466 , n10674 );
nor ( n17324 , n17322 , n17323 );
xnor ( n17325 , n17324 , n10952 );
xor ( n17326 , n17321 , n17325 );
and ( n17327 , n8643 , n12905 );
xor ( n17328 , n17326 , n17327 );
xor ( n17329 , n17317 , n17328 );
xor ( n17330 , n17308 , n17329 );
xor ( n17331 , n17299 , n17330 );
and ( n17332 , n17157 , n17161 );
and ( n17333 , n17161 , n17176 );
and ( n17334 , n17157 , n17176 );
or ( n17335 , n17332 , n17333 , n17334 );
and ( n17336 , n17096 , n17110 );
and ( n17337 , n17110 , n17142 );
and ( n17338 , n17096 , n17142 );
or ( n17339 , n17336 , n17337 , n17338 );
xor ( n17340 , n17335 , n17339 );
and ( n17341 , n10679 , n10477 );
and ( n17342 , n10982 , n10205 );
nor ( n17343 , n17341 , n17342 );
xnor ( n17344 , n17343 , n10426 );
and ( n17345 , n9240 , n12194 );
and ( n17346 , n9438 , n11890 );
nor ( n17347 , n17345 , n17346 );
xnor ( n17348 , n17347 , n12184 );
xor ( n17349 , n17344 , n17348 );
and ( n17350 , n8781 , n12957 );
and ( n17351 , n9018 , n12511 );
nor ( n17352 , n17350 , n17351 );
xnor ( n17353 , n17352 , n12908 );
xor ( n17354 , n17349 , n17353 );
not ( n17355 , n8612 );
and ( n17356 , n12500 , n8992 );
and ( n17357 , n12899 , n8792 );
nor ( n17358 , n17356 , n17357 );
xnor ( n17359 , n17358 , n8998 );
xor ( n17360 , n17355 , n17359 );
and ( n17361 , n11274 , n9920 );
and ( n17362 , n11539 , n9671 );
nor ( n17363 , n17361 , n17362 );
xnor ( n17364 , n17363 , n9926 );
xor ( n17365 , n17360 , n17364 );
xor ( n17366 , n17354 , n17365 );
and ( n17367 , n17119 , n17123 );
and ( n17368 , n17123 , n17128 );
and ( n17369 , n17119 , n17128 );
or ( n17370 , n17367 , n17368 , n17369 );
buf ( n17371 , n17108 );
xor ( n17372 , n17370 , n17371 );
and ( n17373 , n9660 , n11566 );
and ( n17374 , n9964 , n11300 );
nor ( n17375 , n17373 , n17374 );
xnor ( n17376 , n17375 , n11572 );
xor ( n17377 , n17372 , n17376 );
xor ( n17378 , n17366 , n17377 );
xor ( n17379 , n17340 , n17378 );
xor ( n17380 , n17331 , n17379 );
xor ( n17381 , n17295 , n17380 );
and ( n17382 , n17088 , n17179 );
xor ( n17383 , n17381 , n17382 );
and ( n17384 , n17180 , n17181 );
xor ( n17385 , n17383 , n17384 );
and ( n17386 , n17084 , n17182 );
and ( n17387 , n17183 , n17186 );
or ( n17388 , n17386 , n17387 );
xor ( n17389 , n17385 , n17388 );
buf ( n17390 , n17389 );
not ( n17391 , n831 );
and ( n17392 , n17391 , n17291 );
and ( n17393 , n17390 , n831 );
or ( n17394 , n17392 , n17393 );
and ( n17395 , n17282 , n17283 );
and ( n17396 , n17200 , n17231 );
and ( n17397 , n17231 , n17280 );
and ( n17398 , n17200 , n17280 );
or ( n17399 , n17396 , n17397 , n17398 );
and ( n17400 , n17236 , n17240 );
and ( n17401 , n17240 , n17279 );
and ( n17402 , n17236 , n17279 );
or ( n17403 , n17400 , n17401 , n17402 );
and ( n17404 , n17271 , n17272 );
and ( n17405 , n17272 , n17277 );
and ( n17406 , n17271 , n17277 );
or ( n17407 , n17404 , n17405 , n17406 );
and ( n17408 , n17213 , n17217 );
and ( n17409 , n17217 , n17229 );
and ( n17410 , n17213 , n17229 );
or ( n17411 , n17408 , n17409 , n17410 );
xor ( n17412 , n17407 , n17411 );
and ( n17413 , n17222 , n17226 );
and ( n17414 , n17226 , n17228 );
and ( n17415 , n17222 , n17228 );
or ( n17416 , n17413 , n17414 , n17415 );
and ( n17417 , n17245 , n17249 );
and ( n17418 , n17249 , n17254 );
and ( n17419 , n17245 , n17254 );
or ( n17420 , n17417 , n17418 , n17419 );
xor ( n17421 , n17416 , n17420 );
and ( n17422 , n17256 , n17260 );
and ( n17423 , n17260 , n17265 );
and ( n17424 , n17256 , n17265 );
or ( n17425 , n17422 , n17423 , n17424 );
xor ( n17426 , n17421 , n17425 );
xor ( n17427 , n17412 , n17426 );
xor ( n17428 , n17403 , n17427 );
and ( n17429 , n17255 , n17266 );
and ( n17430 , n17266 , n17278 );
and ( n17431 , n17255 , n17278 );
or ( n17432 , n17429 , n17430 , n17431 );
and ( n17433 , n17204 , n17208 );
and ( n17434 , n17208 , n17230 );
and ( n17435 , n17204 , n17230 );
or ( n17436 , n17433 , n17434 , n17435 );
xor ( n17437 , n17432 , n17436 );
and ( n17438 , n10837 , n10342 );
and ( n17439 , n11133 , n10084 );
nor ( n17440 , n17438 , n17439 );
xnor ( n17441 , n17440 , n10291 );
and ( n17442 , n8913 , n12782 );
and ( n17443 , n9139 , n12350 );
nor ( n17444 , n17442 , n17443 );
xnor ( n17445 , n17444 , n12733 );
xor ( n17446 , n17441 , n17445 );
and ( n17447 , n8690 , n12730 );
xor ( n17448 , n17446 , n17447 );
and ( n17449 , n12010 , n9311 );
and ( n17450 , n12339 , n9150 );
nor ( n17451 , n17449 , n17450 );
xnor ( n17452 , n17451 , n9317 );
and ( n17453 , n11384 , n9795 );
and ( n17454 , n11699 , n9560 );
nor ( n17455 , n17453 , n17454 );
xnor ( n17456 , n17455 , n9801 );
xor ( n17457 , n17452 , n17456 );
and ( n17458 , n10331 , n10907 );
and ( n17459 , n10548 , n10543 );
nor ( n17460 , n17458 , n17459 );
xnor ( n17461 , n17460 , n10807 );
xor ( n17462 , n17457 , n17461 );
xor ( n17463 , n17448 , n17462 );
and ( n17464 , n12724 , n8887 );
not ( n17465 , n17464 );
xnor ( n17466 , n17465 , n8893 );
not ( n17467 , n17466 );
and ( n17468 , n9839 , n11411 );
and ( n17469 , n10090 , n11159 );
nor ( n17470 , n17468 , n17469 );
xnor ( n17471 , n17470 , n11417 );
xor ( n17472 , n17467 , n17471 );
and ( n17473 , n9323 , n12029 );
and ( n17474 , n9549 , n11739 );
nor ( n17475 , n17473 , n17474 );
xnor ( n17476 , n17475 , n12019 );
xor ( n17477 , n17472 , n17476 );
xor ( n17478 , n17463 , n17477 );
xor ( n17479 , n17437 , n17478 );
xor ( n17480 , n17428 , n17479 );
xor ( n17481 , n17399 , n17480 );
and ( n17482 , n17196 , n17281 );
xor ( n17483 , n17481 , n17482 );
xor ( n17484 , n17395 , n17483 );
and ( n17485 , n17284 , n17285 );
and ( n17486 , n17286 , n17289 );
or ( n17487 , n17485 , n17486 );
xor ( n17488 , n17484 , n17487 );
buf ( n17489 , n17488 );
and ( n17490 , n17381 , n17382 );
and ( n17491 , n17299 , n17330 );
and ( n17492 , n17330 , n17379 );
and ( n17493 , n17299 , n17379 );
or ( n17494 , n17491 , n17492 , n17493 );
and ( n17495 , n17335 , n17339 );
and ( n17496 , n17339 , n17378 );
and ( n17497 , n17335 , n17378 );
or ( n17498 , n17495 , n17496 , n17497 );
and ( n17499 , n17370 , n17371 );
and ( n17500 , n17371 , n17376 );
and ( n17501 , n17370 , n17376 );
or ( n17502 , n17499 , n17500 , n17501 );
and ( n17503 , n17312 , n17316 );
and ( n17504 , n17316 , n17328 );
and ( n17505 , n17312 , n17328 );
or ( n17506 , n17503 , n17504 , n17505 );
xor ( n17507 , n17502 , n17506 );
and ( n17508 , n17321 , n17325 );
and ( n17509 , n17325 , n17327 );
and ( n17510 , n17321 , n17327 );
or ( n17511 , n17508 , n17509 , n17510 );
and ( n17512 , n17344 , n17348 );
and ( n17513 , n17348 , n17353 );
and ( n17514 , n17344 , n17353 );
or ( n17515 , n17512 , n17513 , n17514 );
xor ( n17516 , n17511 , n17515 );
and ( n17517 , n17355 , n17359 );
and ( n17518 , n17359 , n17364 );
and ( n17519 , n17355 , n17364 );
or ( n17520 , n17517 , n17518 , n17519 );
xor ( n17521 , n17516 , n17520 );
xor ( n17522 , n17507 , n17521 );
xor ( n17523 , n17498 , n17522 );
and ( n17524 , n17354 , n17365 );
and ( n17525 , n17365 , n17377 );
and ( n17526 , n17354 , n17377 );
or ( n17527 , n17524 , n17525 , n17526 );
and ( n17528 , n17303 , n17307 );
and ( n17529 , n17307 , n17329 );
and ( n17530 , n17303 , n17329 );
or ( n17531 , n17528 , n17529 , n17530 );
xor ( n17532 , n17527 , n17531 );
and ( n17533 , n10982 , n10477 );
and ( n17534 , n11274 , n10205 );
nor ( n17535 , n17533 , n17534 );
xnor ( n17536 , n17535 , n10426 );
and ( n17537 , n9018 , n12957 );
and ( n17538 , n9240 , n12511 );
nor ( n17539 , n17537 , n17538 );
xnor ( n17540 , n17539 , n12908 );
xor ( n17541 , n17536 , n17540 );
and ( n17542 , n8781 , n12905 );
xor ( n17543 , n17541 , n17542 );
and ( n17544 , n12175 , n9426 );
and ( n17545 , n12500 , n9251 );
nor ( n17546 , n17544 , n17545 );
xnor ( n17547 , n17546 , n9432 );
and ( n17548 , n11539 , n9920 );
and ( n17549 , n11850 , n9671 );
nor ( n17550 , n17548 , n17549 );
xnor ( n17551 , n17550 , n9926 );
xor ( n17552 , n17547 , n17551 );
and ( n17553 , n10466 , n11052 );
and ( n17554 , n10679 , n10674 );
nor ( n17555 , n17553 , n17554 );
xnor ( n17556 , n17555 , n10952 );
xor ( n17557 , n17552 , n17556 );
xor ( n17558 , n17543 , n17557 );
and ( n17559 , n12899 , n8992 );
not ( n17560 , n17559 );
xnor ( n17561 , n17560 , n8998 );
not ( n17562 , n17561 );
and ( n17563 , n9964 , n11566 );
and ( n17564 , n10211 , n11300 );
nor ( n17565 , n17563 , n17564 );
xnor ( n17566 , n17565 , n11572 );
xor ( n17567 , n17562 , n17566 );
and ( n17568 , n9438 , n12194 );
and ( n17569 , n9660 , n11890 );
nor ( n17570 , n17568 , n17569 );
xnor ( n17571 , n17570 , n12184 );
xor ( n17572 , n17567 , n17571 );
xor ( n17573 , n17558 , n17572 );
xor ( n17574 , n17532 , n17573 );
xor ( n17575 , n17523 , n17574 );
xor ( n17576 , n17494 , n17575 );
and ( n17577 , n17295 , n17380 );
xor ( n17578 , n17576 , n17577 );
xor ( n17579 , n17490 , n17578 );
and ( n17580 , n17383 , n17384 );
and ( n17581 , n17385 , n17388 );
or ( n17582 , n17580 , n17581 );
xor ( n17583 , n17579 , n17582 );
buf ( n17584 , n17583 );
not ( n17585 , n831 );
and ( n17586 , n17585 , n17489 );
and ( n17587 , n17584 , n831 );
or ( n17588 , n17586 , n17587 );
and ( n17589 , n17481 , n17482 );
and ( n17590 , n17403 , n17427 );
and ( n17591 , n17427 , n17479 );
and ( n17592 , n17403 , n17479 );
or ( n17593 , n17590 , n17591 , n17592 );
and ( n17594 , n17432 , n17436 );
and ( n17595 , n17436 , n17478 );
and ( n17596 , n17432 , n17478 );
or ( n17597 , n17594 , n17595 , n17596 );
and ( n17598 , n17416 , n17420 );
and ( n17599 , n17420 , n17425 );
and ( n17600 , n17416 , n17425 );
or ( n17601 , n17598 , n17599 , n17600 );
and ( n17602 , n17467 , n17471 );
and ( n17603 , n17471 , n17476 );
and ( n17604 , n17467 , n17476 );
or ( n17605 , n17602 , n17603 , n17604 );
xor ( n17606 , n17601 , n17605 );
and ( n17607 , n17441 , n17445 );
and ( n17608 , n17445 , n17447 );
and ( n17609 , n17441 , n17447 );
or ( n17610 , n17607 , n17608 , n17609 );
and ( n17611 , n17452 , n17456 );
and ( n17612 , n17456 , n17461 );
and ( n17613 , n17452 , n17461 );
or ( n17614 , n17611 , n17612 , n17613 );
xor ( n17615 , n17610 , n17614 );
buf ( n17616 , n17466 );
xor ( n17617 , n17615 , n17616 );
xor ( n17618 , n17606 , n17617 );
xor ( n17619 , n17597 , n17618 );
and ( n17620 , n17448 , n17462 );
and ( n17621 , n17462 , n17477 );
and ( n17622 , n17448 , n17477 );
or ( n17623 , n17620 , n17621 , n17622 );
and ( n17624 , n17407 , n17411 );
and ( n17625 , n17411 , n17426 );
and ( n17626 , n17407 , n17426 );
or ( n17627 , n17624 , n17625 , n17626 );
xor ( n17628 , n17623 , n17627 );
and ( n17629 , n10548 , n10907 );
and ( n17630 , n10837 , n10543 );
nor ( n17631 , n17629 , n17630 );
xnor ( n17632 , n17631 , n10807 );
and ( n17633 , n9139 , n12782 );
and ( n17634 , n9323 , n12350 );
nor ( n17635 , n17633 , n17634 );
xnor ( n17636 , n17635 , n12733 );
xor ( n17637 , n17632 , n17636 );
and ( n17638 , n8913 , n12730 );
xor ( n17639 , n17637 , n17638 );
and ( n17640 , n11699 , n9795 );
and ( n17641 , n12010 , n9560 );
nor ( n17642 , n17640 , n17641 );
xnor ( n17643 , n17642 , n9801 );
and ( n17644 , n10090 , n11411 );
and ( n17645 , n10331 , n11159 );
nor ( n17646 , n17644 , n17645 );
xnor ( n17647 , n17646 , n11417 );
xor ( n17648 , n17643 , n17647 );
and ( n17649 , n9549 , n12029 );
and ( n17650 , n9839 , n11739 );
nor ( n17651 , n17649 , n17650 );
xnor ( n17652 , n17651 , n12019 );
xor ( n17653 , n17648 , n17652 );
xor ( n17654 , n17639 , n17653 );
not ( n17655 , n8893 );
and ( n17656 , n12339 , n9311 );
and ( n17657 , n12724 , n9150 );
nor ( n17658 , n17656 , n17657 );
xnor ( n17659 , n17658 , n9317 );
xor ( n17660 , n17655 , n17659 );
and ( n17661 , n11133 , n10342 );
and ( n17662 , n11384 , n10084 );
nor ( n17663 , n17661 , n17662 );
xnor ( n17664 , n17663 , n10291 );
xor ( n17665 , n17660 , n17664 );
xor ( n17666 , n17654 , n17665 );
xor ( n17667 , n17628 , n17666 );
xor ( n17668 , n17619 , n17667 );
xor ( n17669 , n17593 , n17668 );
and ( n17670 , n17399 , n17480 );
xor ( n17671 , n17669 , n17670 );
xor ( n17672 , n17589 , n17671 );
and ( n17673 , n17395 , n17483 );
and ( n17674 , n17484 , n17487 );
or ( n17675 , n17673 , n17674 );
xor ( n17676 , n17672 , n17675 );
buf ( n17677 , n17676 );
and ( n17678 , n17576 , n17577 );
and ( n17679 , n17498 , n17522 );
and ( n17680 , n17522 , n17574 );
and ( n17681 , n17498 , n17574 );
or ( n17682 , n17679 , n17680 , n17681 );
and ( n17683 , n17527 , n17531 );
and ( n17684 , n17531 , n17573 );
and ( n17685 , n17527 , n17573 );
or ( n17686 , n17683 , n17684 , n17685 );
and ( n17687 , n17511 , n17515 );
and ( n17688 , n17515 , n17520 );
and ( n17689 , n17511 , n17520 );
or ( n17690 , n17687 , n17688 , n17689 );
and ( n17691 , n17562 , n17566 );
and ( n17692 , n17566 , n17571 );
and ( n17693 , n17562 , n17571 );
or ( n17694 , n17691 , n17692 , n17693 );
xor ( n17695 , n17690 , n17694 );
and ( n17696 , n17536 , n17540 );
and ( n17697 , n17540 , n17542 );
and ( n17698 , n17536 , n17542 );
or ( n17699 , n17696 , n17697 , n17698 );
and ( n17700 , n17547 , n17551 );
and ( n17701 , n17551 , n17556 );
and ( n17702 , n17547 , n17556 );
or ( n17703 , n17700 , n17701 , n17702 );
xor ( n17704 , n17699 , n17703 );
buf ( n17705 , n17561 );
xor ( n17706 , n17704 , n17705 );
xor ( n17707 , n17695 , n17706 );
xor ( n17708 , n17686 , n17707 );
and ( n17709 , n17543 , n17557 );
and ( n17710 , n17557 , n17572 );
and ( n17711 , n17543 , n17572 );
or ( n17712 , n17709 , n17710 , n17711 );
and ( n17713 , n17502 , n17506 );
and ( n17714 , n17506 , n17521 );
and ( n17715 , n17502 , n17521 );
or ( n17716 , n17713 , n17714 , n17715 );
xor ( n17717 , n17712 , n17716 );
and ( n17718 , n10679 , n11052 );
and ( n17719 , n10982 , n10674 );
nor ( n17720 , n17718 , n17719 );
xnor ( n17721 , n17720 , n10952 );
and ( n17722 , n9240 , n12957 );
and ( n17723 , n9438 , n12511 );
nor ( n17724 , n17722 , n17723 );
xnor ( n17725 , n17724 , n12908 );
xor ( n17726 , n17721 , n17725 );
and ( n17727 , n9018 , n12905 );
xor ( n17728 , n17726 , n17727 );
and ( n17729 , n11850 , n9920 );
and ( n17730 , n12175 , n9671 );
nor ( n17731 , n17729 , n17730 );
xnor ( n17732 , n17731 , n9926 );
and ( n17733 , n10211 , n11566 );
and ( n17734 , n10466 , n11300 );
nor ( n17735 , n17733 , n17734 );
xnor ( n17736 , n17735 , n11572 );
xor ( n17737 , n17732 , n17736 );
and ( n17738 , n9660 , n12194 );
and ( n17739 , n9964 , n11890 );
nor ( n17740 , n17738 , n17739 );
xnor ( n17741 , n17740 , n12184 );
xor ( n17742 , n17737 , n17741 );
xor ( n17743 , n17728 , n17742 );
not ( n17744 , n8998 );
and ( n17745 , n12500 , n9426 );
and ( n17746 , n12899 , n9251 );
nor ( n17747 , n17745 , n17746 );
xnor ( n17748 , n17747 , n9432 );
xor ( n17749 , n17744 , n17748 );
and ( n17750 , n11274 , n10477 );
and ( n17751 , n11539 , n10205 );
nor ( n17752 , n17750 , n17751 );
xnor ( n17753 , n17752 , n10426 );
xor ( n17754 , n17749 , n17753 );
xor ( n17755 , n17743 , n17754 );
xor ( n17756 , n17717 , n17755 );
xor ( n17757 , n17708 , n17756 );
xor ( n17758 , n17682 , n17757 );
and ( n17759 , n17494 , n17575 );
xor ( n17760 , n17758 , n17759 );
xor ( n17761 , n17678 , n17760 );
and ( n17762 , n17490 , n17578 );
and ( n17763 , n17579 , n17582 );
or ( n17764 , n17762 , n17763 );
xor ( n17765 , n17761 , n17764 );
buf ( n17766 , n17765 );
not ( n17767 , n831 );
and ( n17768 , n17767 , n17677 );
and ( n17769 , n17766 , n831 );
or ( n17770 , n17768 , n17769 );
and ( n17771 , n17669 , n17670 );
and ( n17772 , n17597 , n17618 );
and ( n17773 , n17618 , n17667 );
and ( n17774 , n17597 , n17667 );
or ( n17775 , n17772 , n17773 , n17774 );
and ( n17776 , n17601 , n17605 );
and ( n17777 , n17605 , n17617 );
and ( n17778 , n17601 , n17617 );
or ( n17779 , n17776 , n17777 , n17778 );
and ( n17780 , n17623 , n17627 );
and ( n17781 , n17627 , n17666 );
and ( n17782 , n17623 , n17666 );
or ( n17783 , n17780 , n17781 , n17782 );
xor ( n17784 , n17779 , n17783 );
and ( n17785 , n17639 , n17653 );
and ( n17786 , n17653 , n17665 );
and ( n17787 , n17639 , n17665 );
or ( n17788 , n17785 , n17786 , n17787 );
and ( n17789 , n17632 , n17636 );
and ( n17790 , n17636 , n17638 );
and ( n17791 , n17632 , n17638 );
or ( n17792 , n17789 , n17790 , n17791 );
and ( n17793 , n17643 , n17647 );
and ( n17794 , n17647 , n17652 );
and ( n17795 , n17643 , n17652 );
or ( n17796 , n17793 , n17794 , n17795 );
xor ( n17797 , n17792 , n17796 );
and ( n17798 , n11384 , n10342 );
and ( n17799 , n11699 , n10084 );
nor ( n17800 , n17798 , n17799 );
xnor ( n17801 , n17800 , n10291 );
and ( n17802 , n10331 , n11411 );
and ( n17803 , n10548 , n11159 );
nor ( n17804 , n17802 , n17803 );
xnor ( n17805 , n17804 , n11417 );
xor ( n17806 , n17801 , n17805 );
and ( n17807 , n9839 , n12029 );
and ( n17808 , n10090 , n11739 );
nor ( n17809 , n17807 , n17808 );
xnor ( n17810 , n17809 , n12019 );
xor ( n17811 , n17806 , n17810 );
xor ( n17812 , n17797 , n17811 );
xor ( n17813 , n17788 , n17812 );
and ( n17814 , n17610 , n17614 );
and ( n17815 , n17614 , n17616 );
and ( n17816 , n17610 , n17616 );
or ( n17817 , n17814 , n17815 , n17816 );
and ( n17818 , n12010 , n9795 );
and ( n17819 , n12339 , n9560 );
nor ( n17820 , n17818 , n17819 );
xnor ( n17821 , n17820 , n9801 );
and ( n17822 , n10837 , n10907 );
and ( n17823 , n11133 , n10543 );
nor ( n17824 , n17822 , n17823 );
xnor ( n17825 , n17824 , n10807 );
xor ( n17826 , n17821 , n17825 );
and ( n17827 , n9139 , n12730 );
xor ( n17828 , n17826 , n17827 );
xor ( n17829 , n17817 , n17828 );
and ( n17830 , n17655 , n17659 );
and ( n17831 , n17659 , n17664 );
and ( n17832 , n17655 , n17664 );
or ( n17833 , n17830 , n17831 , n17832 );
and ( n17834 , n12724 , n9311 );
not ( n17835 , n17834 );
xnor ( n17836 , n17835 , n9317 );
not ( n17837 , n17836 );
xor ( n17838 , n17833 , n17837 );
and ( n17839 , n9323 , n12782 );
and ( n17840 , n9549 , n12350 );
nor ( n17841 , n17839 , n17840 );
xnor ( n17842 , n17841 , n12733 );
xor ( n17843 , n17838 , n17842 );
xor ( n17844 , n17829 , n17843 );
xor ( n17845 , n17813 , n17844 );
xor ( n17846 , n17784 , n17845 );
xor ( n17847 , n17775 , n17846 );
and ( n17848 , n17593 , n17668 );
xor ( n17849 , n17847 , n17848 );
xor ( n17850 , n17771 , n17849 );
and ( n17851 , n17589 , n17671 );
and ( n17852 , n17672 , n17675 );
or ( n17853 , n17851 , n17852 );
xor ( n17854 , n17850 , n17853 );
buf ( n17855 , n17854 );
and ( n17856 , n17758 , n17759 );
and ( n17857 , n17686 , n17707 );
and ( n17858 , n17707 , n17756 );
and ( n17859 , n17686 , n17756 );
or ( n17860 , n17857 , n17858 , n17859 );
and ( n17861 , n17690 , n17694 );
and ( n17862 , n17694 , n17706 );
and ( n17863 , n17690 , n17706 );
or ( n17864 , n17861 , n17862 , n17863 );
and ( n17865 , n17712 , n17716 );
and ( n17866 , n17716 , n17755 );
and ( n17867 , n17712 , n17755 );
or ( n17868 , n17865 , n17866 , n17867 );
xor ( n17869 , n17864 , n17868 );
and ( n17870 , n17728 , n17742 );
and ( n17871 , n17742 , n17754 );
and ( n17872 , n17728 , n17754 );
or ( n17873 , n17870 , n17871 , n17872 );
and ( n17874 , n17721 , n17725 );
and ( n17875 , n17725 , n17727 );
and ( n17876 , n17721 , n17727 );
or ( n17877 , n17874 , n17875 , n17876 );
and ( n17878 , n17732 , n17736 );
and ( n17879 , n17736 , n17741 );
and ( n17880 , n17732 , n17741 );
or ( n17881 , n17878 , n17879 , n17880 );
xor ( n17882 , n17877 , n17881 );
and ( n17883 , n11539 , n10477 );
and ( n17884 , n11850 , n10205 );
nor ( n17885 , n17883 , n17884 );
xnor ( n17886 , n17885 , n10426 );
and ( n17887 , n10466 , n11566 );
and ( n17888 , n10679 , n11300 );
nor ( n17889 , n17887 , n17888 );
xnor ( n17890 , n17889 , n11572 );
xor ( n17891 , n17886 , n17890 );
and ( n17892 , n9964 , n12194 );
and ( n17893 , n10211 , n11890 );
nor ( n17894 , n17892 , n17893 );
xnor ( n17895 , n17894 , n12184 );
xor ( n17896 , n17891 , n17895 );
xor ( n17897 , n17882 , n17896 );
xor ( n17898 , n17873 , n17897 );
and ( n17899 , n17699 , n17703 );
and ( n17900 , n17703 , n17705 );
and ( n17901 , n17699 , n17705 );
or ( n17902 , n17899 , n17900 , n17901 );
and ( n17903 , n12175 , n9920 );
and ( n17904 , n12500 , n9671 );
nor ( n17905 , n17903 , n17904 );
xnor ( n17906 , n17905 , n9926 );
and ( n17907 , n10982 , n11052 );
and ( n17908 , n11274 , n10674 );
nor ( n17909 , n17907 , n17908 );
xnor ( n17910 , n17909 , n10952 );
xor ( n17911 , n17906 , n17910 );
and ( n17912 , n9240 , n12905 );
xor ( n17913 , n17911 , n17912 );
xor ( n17914 , n17902 , n17913 );
and ( n17915 , n17744 , n17748 );
and ( n17916 , n17748 , n17753 );
and ( n17917 , n17744 , n17753 );
or ( n17918 , n17915 , n17916 , n17917 );
and ( n17919 , n12899 , n9426 );
not ( n17920 , n17919 );
xnor ( n17921 , n17920 , n9432 );
not ( n17922 , n17921 );
xor ( n17923 , n17918 , n17922 );
and ( n17924 , n9438 , n12957 );
and ( n17925 , n9660 , n12511 );
nor ( n17926 , n17924 , n17925 );
xnor ( n17927 , n17926 , n12908 );
xor ( n17928 , n17923 , n17927 );
xor ( n17929 , n17914 , n17928 );
xor ( n17930 , n17898 , n17929 );
xor ( n17931 , n17869 , n17930 );
xor ( n17932 , n17860 , n17931 );
and ( n17933 , n17682 , n17757 );
xor ( n17934 , n17932 , n17933 );
xor ( n17935 , n17856 , n17934 );
and ( n17936 , n17678 , n17760 );
and ( n17937 , n17761 , n17764 );
or ( n17938 , n17936 , n17937 );
xor ( n17939 , n17935 , n17938 );
buf ( n17940 , n17939 );
not ( n17941 , n831 );
and ( n17942 , n17941 , n17855 );
and ( n17943 , n17940 , n831 );
or ( n17944 , n17942 , n17943 );
and ( n17945 , n17847 , n17848 );
and ( n17946 , n17779 , n17783 );
and ( n17947 , n17783 , n17845 );
and ( n17948 , n17779 , n17845 );
or ( n17949 , n17946 , n17947 , n17948 );
and ( n17950 , n17788 , n17812 );
and ( n17951 , n17812 , n17844 );
and ( n17952 , n17788 , n17844 );
or ( n17953 , n17950 , n17951 , n17952 );
and ( n17954 , n17833 , n17837 );
and ( n17955 , n17837 , n17842 );
and ( n17956 , n17833 , n17842 );
or ( n17957 , n17954 , n17955 , n17956 );
and ( n17958 , n11699 , n10342 );
and ( n17959 , n12010 , n10084 );
nor ( n17960 , n17958 , n17959 );
xnor ( n17961 , n17960 , n10291 );
and ( n17962 , n10548 , n11411 );
and ( n17963 , n10837 , n11159 );
nor ( n17964 , n17962 , n17963 );
xnor ( n17965 , n17964 , n11417 );
xor ( n17966 , n17961 , n17965 );
and ( n17967 , n9323 , n12730 );
xor ( n17968 , n17966 , n17967 );
xor ( n17969 , n17957 , n17968 );
buf ( n17970 , n17836 );
and ( n17971 , n10090 , n12029 );
and ( n17972 , n10331 , n11739 );
nor ( n17973 , n17971 , n17972 );
xnor ( n17974 , n17973 , n12019 );
xor ( n17975 , n17970 , n17974 );
and ( n17976 , n9549 , n12782 );
and ( n17977 , n9839 , n12350 );
nor ( n17978 , n17976 , n17977 );
xnor ( n17979 , n17978 , n12733 );
xor ( n17980 , n17975 , n17979 );
xor ( n17981 , n17969 , n17980 );
xor ( n17982 , n17953 , n17981 );
and ( n17983 , n17792 , n17796 );
and ( n17984 , n17796 , n17811 );
and ( n17985 , n17792 , n17811 );
or ( n17986 , n17983 , n17984 , n17985 );
and ( n17987 , n17817 , n17828 );
and ( n17988 , n17828 , n17843 );
and ( n17989 , n17817 , n17843 );
or ( n17990 , n17987 , n17988 , n17989 );
xor ( n17991 , n17986 , n17990 );
and ( n17992 , n17801 , n17805 );
and ( n17993 , n17805 , n17810 );
and ( n17994 , n17801 , n17810 );
or ( n17995 , n17992 , n17993 , n17994 );
and ( n17996 , n17821 , n17825 );
and ( n17997 , n17825 , n17827 );
and ( n17998 , n17821 , n17827 );
or ( n17999 , n17996 , n17997 , n17998 );
xor ( n18000 , n17995 , n17999 );
not ( n18001 , n9317 );
and ( n18002 , n12339 , n9795 );
and ( n18003 , n12724 , n9560 );
nor ( n18004 , n18002 , n18003 );
xnor ( n18005 , n18004 , n9801 );
xor ( n18006 , n18001 , n18005 );
and ( n18007 , n11133 , n10907 );
and ( n18008 , n11384 , n10543 );
nor ( n18009 , n18007 , n18008 );
xnor ( n18010 , n18009 , n10807 );
xor ( n18011 , n18006 , n18010 );
xor ( n18012 , n18000 , n18011 );
xor ( n18013 , n17991 , n18012 );
xor ( n18014 , n17982 , n18013 );
xor ( n18015 , n17949 , n18014 );
and ( n18016 , n17775 , n17846 );
xor ( n18017 , n18015 , n18016 );
xor ( n18018 , n17945 , n18017 );
and ( n18019 , n17771 , n17849 );
and ( n18020 , n17850 , n17853 );
or ( n18021 , n18019 , n18020 );
xor ( n18022 , n18018 , n18021 );
buf ( n18023 , n18022 );
and ( n18024 , n17932 , n17933 );
and ( n18025 , n17864 , n17868 );
and ( n18026 , n17868 , n17930 );
and ( n18027 , n17864 , n17930 );
or ( n18028 , n18025 , n18026 , n18027 );
and ( n18029 , n17873 , n17897 );
and ( n18030 , n17897 , n17929 );
and ( n18031 , n17873 , n17929 );
or ( n18032 , n18029 , n18030 , n18031 );
and ( n18033 , n17918 , n17922 );
and ( n18034 , n17922 , n17927 );
and ( n18035 , n17918 , n17927 );
or ( n18036 , n18033 , n18034 , n18035 );
and ( n18037 , n11850 , n10477 );
and ( n18038 , n12175 , n10205 );
nor ( n18039 , n18037 , n18038 );
xnor ( n18040 , n18039 , n10426 );
and ( n18041 , n10679 , n11566 );
and ( n18042 , n10982 , n11300 );
nor ( n18043 , n18041 , n18042 );
xnor ( n18044 , n18043 , n11572 );
xor ( n18045 , n18040 , n18044 );
and ( n18046 , n9438 , n12905 );
xor ( n18047 , n18045 , n18046 );
xor ( n18048 , n18036 , n18047 );
buf ( n18049 , n17921 );
and ( n18050 , n10211 , n12194 );
and ( n18051 , n10466 , n11890 );
nor ( n18052 , n18050 , n18051 );
xnor ( n18053 , n18052 , n12184 );
xor ( n18054 , n18049 , n18053 );
and ( n18055 , n9660 , n12957 );
and ( n18056 , n9964 , n12511 );
nor ( n18057 , n18055 , n18056 );
xnor ( n18058 , n18057 , n12908 );
xor ( n18059 , n18054 , n18058 );
xor ( n18060 , n18048 , n18059 );
xor ( n18061 , n18032 , n18060 );
and ( n18062 , n17877 , n17881 );
and ( n18063 , n17881 , n17896 );
and ( n18064 , n17877 , n17896 );
or ( n18065 , n18062 , n18063 , n18064 );
and ( n18066 , n17902 , n17913 );
and ( n18067 , n17913 , n17928 );
and ( n18068 , n17902 , n17928 );
or ( n18069 , n18066 , n18067 , n18068 );
xor ( n18070 , n18065 , n18069 );
and ( n18071 , n17886 , n17890 );
and ( n18072 , n17890 , n17895 );
and ( n18073 , n17886 , n17895 );
or ( n18074 , n18071 , n18072 , n18073 );
and ( n18075 , n17906 , n17910 );
and ( n18076 , n17910 , n17912 );
and ( n18077 , n17906 , n17912 );
or ( n18078 , n18075 , n18076 , n18077 );
xor ( n18079 , n18074 , n18078 );
not ( n18080 , n9432 );
and ( n18081 , n12500 , n9920 );
and ( n18082 , n12899 , n9671 );
nor ( n18083 , n18081 , n18082 );
xnor ( n18084 , n18083 , n9926 );
xor ( n18085 , n18080 , n18084 );
and ( n18086 , n11274 , n11052 );
and ( n18087 , n11539 , n10674 );
nor ( n18088 , n18086 , n18087 );
xnor ( n18089 , n18088 , n10952 );
xor ( n18090 , n18085 , n18089 );
xor ( n18091 , n18079 , n18090 );
xor ( n18092 , n18070 , n18091 );
xor ( n18093 , n18061 , n18092 );
xor ( n18094 , n18028 , n18093 );
and ( n18095 , n17860 , n17931 );
xor ( n18096 , n18094 , n18095 );
xor ( n18097 , n18024 , n18096 );
and ( n18098 , n17856 , n17934 );
and ( n18099 , n17935 , n17938 );
or ( n18100 , n18098 , n18099 );
xor ( n18101 , n18097 , n18100 );
buf ( n18102 , n18101 );
not ( n18103 , n831 );
and ( n18104 , n18103 , n18023 );
and ( n18105 , n18102 , n831 );
or ( n18106 , n18104 , n18105 );
and ( n18107 , n18015 , n18016 );
and ( n18108 , n17953 , n17981 );
and ( n18109 , n17981 , n18013 );
and ( n18110 , n17953 , n18013 );
or ( n18111 , n18108 , n18109 , n18110 );
and ( n18112 , n17957 , n17968 );
and ( n18113 , n17968 , n17980 );
and ( n18114 , n17957 , n17980 );
or ( n18115 , n18112 , n18113 , n18114 );
and ( n18116 , n17986 , n17990 );
and ( n18117 , n17990 , n18012 );
and ( n18118 , n17986 , n18012 );
or ( n18119 , n18116 , n18117 , n18118 );
xor ( n18120 , n18115 , n18119 );
and ( n18121 , n17995 , n17999 );
and ( n18122 , n17999 , n18011 );
and ( n18123 , n17995 , n18011 );
or ( n18124 , n18121 , n18122 , n18123 );
and ( n18125 , n17961 , n17965 );
and ( n18126 , n17965 , n17967 );
and ( n18127 , n17961 , n17967 );
or ( n18128 , n18125 , n18126 , n18127 );
and ( n18129 , n18001 , n18005 );
and ( n18130 , n18005 , n18010 );
and ( n18131 , n18001 , n18010 );
or ( n18132 , n18129 , n18130 , n18131 );
xor ( n18133 , n18128 , n18132 );
and ( n18134 , n12724 , n9795 );
not ( n18135 , n18134 );
xnor ( n18136 , n18135 , n9801 );
not ( n18137 , n18136 );
xor ( n18138 , n18133 , n18137 );
xor ( n18139 , n18124 , n18138 );
and ( n18140 , n17970 , n17974 );
and ( n18141 , n17974 , n17979 );
and ( n18142 , n17970 , n17979 );
or ( n18143 , n18140 , n18141 , n18142 );
and ( n18144 , n12010 , n10342 );
and ( n18145 , n12339 , n10084 );
nor ( n18146 , n18144 , n18145 );
xnor ( n18147 , n18146 , n10291 );
and ( n18148 , n10837 , n11411 );
and ( n18149 , n11133 , n11159 );
nor ( n18150 , n18148 , n18149 );
xnor ( n18151 , n18150 , n11417 );
xor ( n18152 , n18147 , n18151 );
and ( n18153 , n10331 , n12029 );
and ( n18154 , n10548 , n11739 );
nor ( n18155 , n18153 , n18154 );
xnor ( n18156 , n18155 , n12019 );
xor ( n18157 , n18152 , n18156 );
xor ( n18158 , n18143 , n18157 );
and ( n18159 , n11384 , n10907 );
and ( n18160 , n11699 , n10543 );
nor ( n18161 , n18159 , n18160 );
xnor ( n18162 , n18161 , n10807 );
and ( n18163 , n9839 , n12782 );
and ( n18164 , n10090 , n12350 );
nor ( n18165 , n18163 , n18164 );
xnor ( n18166 , n18165 , n12733 );
xor ( n18167 , n18162 , n18166 );
and ( n18168 , n9549 , n12730 );
xor ( n18169 , n18167 , n18168 );
xor ( n18170 , n18158 , n18169 );
xor ( n18171 , n18139 , n18170 );
xor ( n18172 , n18120 , n18171 );
xor ( n18173 , n18111 , n18172 );
and ( n18174 , n17949 , n18014 );
xor ( n18175 , n18173 , n18174 );
xor ( n18176 , n18107 , n18175 );
and ( n18177 , n17945 , n18017 );
and ( n18178 , n18018 , n18021 );
or ( n18179 , n18177 , n18178 );
xor ( n18180 , n18176 , n18179 );
buf ( n18181 , n18180 );
and ( n18182 , n18094 , n18095 );
and ( n18183 , n18032 , n18060 );
and ( n18184 , n18060 , n18092 );
and ( n18185 , n18032 , n18092 );
or ( n18186 , n18183 , n18184 , n18185 );
and ( n18187 , n18036 , n18047 );
and ( n18188 , n18047 , n18059 );
and ( n18189 , n18036 , n18059 );
or ( n18190 , n18187 , n18188 , n18189 );
and ( n18191 , n18065 , n18069 );
and ( n18192 , n18069 , n18091 );
and ( n18193 , n18065 , n18091 );
or ( n18194 , n18191 , n18192 , n18193 );
xor ( n18195 , n18190 , n18194 );
and ( n18196 , n18074 , n18078 );
and ( n18197 , n18078 , n18090 );
and ( n18198 , n18074 , n18090 );
or ( n18199 , n18196 , n18197 , n18198 );
and ( n18200 , n18040 , n18044 );
and ( n18201 , n18044 , n18046 );
and ( n18202 , n18040 , n18046 );
or ( n18203 , n18200 , n18201 , n18202 );
and ( n18204 , n18080 , n18084 );
and ( n18205 , n18084 , n18089 );
and ( n18206 , n18080 , n18089 );
or ( n18207 , n18204 , n18205 , n18206 );
xor ( n18208 , n18203 , n18207 );
and ( n18209 , n12899 , n9920 );
not ( n18210 , n18209 );
xnor ( n18211 , n18210 , n9926 );
not ( n18212 , n18211 );
xor ( n18213 , n18208 , n18212 );
xor ( n18214 , n18199 , n18213 );
and ( n18215 , n18049 , n18053 );
and ( n18216 , n18053 , n18058 );
and ( n18217 , n18049 , n18058 );
or ( n18218 , n18215 , n18216 , n18217 );
and ( n18219 , n12175 , n10477 );
and ( n18220 , n12500 , n10205 );
nor ( n18221 , n18219 , n18220 );
xnor ( n18222 , n18221 , n10426 );
and ( n18223 , n10982 , n11566 );
and ( n18224 , n11274 , n11300 );
nor ( n18225 , n18223 , n18224 );
xnor ( n18226 , n18225 , n11572 );
xor ( n18227 , n18222 , n18226 );
and ( n18228 , n10466 , n12194 );
and ( n18229 , n10679 , n11890 );
nor ( n18230 , n18228 , n18229 );
xnor ( n18231 , n18230 , n12184 );
xor ( n18232 , n18227 , n18231 );
xor ( n18233 , n18218 , n18232 );
and ( n18234 , n11539 , n11052 );
and ( n18235 , n11850 , n10674 );
nor ( n18236 , n18234 , n18235 );
xnor ( n18237 , n18236 , n10952 );
and ( n18238 , n9964 , n12957 );
and ( n18239 , n10211 , n12511 );
nor ( n18240 , n18238 , n18239 );
xnor ( n18241 , n18240 , n12908 );
xor ( n18242 , n18237 , n18241 );
and ( n18243 , n9660 , n12905 );
xor ( n18244 , n18242 , n18243 );
xor ( n18245 , n18233 , n18244 );
xor ( n18246 , n18214 , n18245 );
xor ( n18247 , n18195 , n18246 );
xor ( n18248 , n18186 , n18247 );
and ( n18249 , n18028 , n18093 );
xor ( n18250 , n18248 , n18249 );
xor ( n18251 , n18182 , n18250 );
and ( n18252 , n18024 , n18096 );
and ( n18253 , n18097 , n18100 );
or ( n18254 , n18252 , n18253 );
xor ( n18255 , n18251 , n18254 );
buf ( n18256 , n18255 );
not ( n18257 , n831 );
and ( n18258 , n18257 , n18181 );
and ( n18259 , n18256 , n831 );
or ( n18260 , n18258 , n18259 );
and ( n18261 , n18173 , n18174 );
and ( n18262 , n18115 , n18119 );
and ( n18263 , n18119 , n18171 );
and ( n18264 , n18115 , n18171 );
or ( n18265 , n18262 , n18263 , n18264 );
and ( n18266 , n18124 , n18138 );
and ( n18267 , n18138 , n18170 );
and ( n18268 , n18124 , n18170 );
or ( n18269 , n18266 , n18267 , n18268 );
and ( n18270 , n18162 , n18166 );
and ( n18271 , n18166 , n18168 );
and ( n18272 , n18162 , n18168 );
or ( n18273 , n18270 , n18271 , n18272 );
not ( n18274 , n9801 );
and ( n18275 , n12339 , n10342 );
and ( n18276 , n12724 , n10084 );
nor ( n18277 , n18275 , n18276 );
xnor ( n18278 , n18277 , n10291 );
xor ( n18279 , n18274 , n18278 );
and ( n18280 , n11133 , n11411 );
and ( n18281 , n11384 , n11159 );
nor ( n18282 , n18280 , n18281 );
xnor ( n18283 , n18282 , n11417 );
xor ( n18284 , n18279 , n18283 );
xor ( n18285 , n18273 , n18284 );
and ( n18286 , n11699 , n10907 );
and ( n18287 , n12010 , n10543 );
nor ( n18288 , n18286 , n18287 );
xnor ( n18289 , n18288 , n10807 );
and ( n18290 , n10548 , n12029 );
and ( n18291 , n10837 , n11739 );
nor ( n18292 , n18290 , n18291 );
xnor ( n18293 , n18292 , n12019 );
xor ( n18294 , n18289 , n18293 );
and ( n18295 , n10090 , n12782 );
and ( n18296 , n10331 , n12350 );
nor ( n18297 , n18295 , n18296 );
xnor ( n18298 , n18297 , n12733 );
xor ( n18299 , n18294 , n18298 );
xor ( n18300 , n18285 , n18299 );
xor ( n18301 , n18269 , n18300 );
and ( n18302 , n18128 , n18132 );
and ( n18303 , n18132 , n18137 );
and ( n18304 , n18128 , n18137 );
or ( n18305 , n18302 , n18303 , n18304 );
and ( n18306 , n18143 , n18157 );
and ( n18307 , n18157 , n18169 );
and ( n18308 , n18143 , n18169 );
or ( n18309 , n18306 , n18307 , n18308 );
xor ( n18310 , n18305 , n18309 );
and ( n18311 , n18147 , n18151 );
and ( n18312 , n18151 , n18156 );
and ( n18313 , n18147 , n18156 );
or ( n18314 , n18311 , n18312 , n18313 );
buf ( n18315 , n18136 );
xor ( n18316 , n18314 , n18315 );
and ( n18317 , n9839 , n12730 );
xor ( n18318 , n18316 , n18317 );
xor ( n18319 , n18310 , n18318 );
xor ( n18320 , n18301 , n18319 );
xor ( n18321 , n18265 , n18320 );
and ( n18322 , n18111 , n18172 );
xor ( n18323 , n18321 , n18322 );
xor ( n18324 , n18261 , n18323 );
and ( n18325 , n18107 , n18175 );
and ( n18326 , n18176 , n18179 );
or ( n18327 , n18325 , n18326 );
xor ( n18328 , n18324 , n18327 );
buf ( n18329 , n18328 );
and ( n18330 , n18248 , n18249 );
and ( n18331 , n18190 , n18194 );
and ( n18332 , n18194 , n18246 );
and ( n18333 , n18190 , n18246 );
or ( n18334 , n18331 , n18332 , n18333 );
and ( n18335 , n18199 , n18213 );
and ( n18336 , n18213 , n18245 );
and ( n18337 , n18199 , n18245 );
or ( n18338 , n18335 , n18336 , n18337 );
and ( n18339 , n18237 , n18241 );
and ( n18340 , n18241 , n18243 );
and ( n18341 , n18237 , n18243 );
or ( n18342 , n18339 , n18340 , n18341 );
not ( n18343 , n9926 );
and ( n18344 , n12500 , n10477 );
and ( n18345 , n12899 , n10205 );
nor ( n18346 , n18344 , n18345 );
xnor ( n18347 , n18346 , n10426 );
xor ( n18348 , n18343 , n18347 );
and ( n18349 , n11274 , n11566 );
and ( n18350 , n11539 , n11300 );
nor ( n18351 , n18349 , n18350 );
xnor ( n18352 , n18351 , n11572 );
xor ( n18353 , n18348 , n18352 );
xor ( n18354 , n18342 , n18353 );
and ( n18355 , n11850 , n11052 );
and ( n18356 , n12175 , n10674 );
nor ( n18357 , n18355 , n18356 );
xnor ( n18358 , n18357 , n10952 );
and ( n18359 , n10679 , n12194 );
and ( n18360 , n10982 , n11890 );
nor ( n18361 , n18359 , n18360 );
xnor ( n18362 , n18361 , n12184 );
xor ( n18363 , n18358 , n18362 );
and ( n18364 , n10211 , n12957 );
and ( n18365 , n10466 , n12511 );
nor ( n18366 , n18364 , n18365 );
xnor ( n18367 , n18366 , n12908 );
xor ( n18368 , n18363 , n18367 );
xor ( n18369 , n18354 , n18368 );
xor ( n18370 , n18338 , n18369 );
and ( n18371 , n18203 , n18207 );
and ( n18372 , n18207 , n18212 );
and ( n18373 , n18203 , n18212 );
or ( n18374 , n18371 , n18372 , n18373 );
and ( n18375 , n18218 , n18232 );
and ( n18376 , n18232 , n18244 );
and ( n18377 , n18218 , n18244 );
or ( n18378 , n18375 , n18376 , n18377 );
xor ( n18379 , n18374 , n18378 );
and ( n18380 , n18222 , n18226 );
and ( n18381 , n18226 , n18231 );
and ( n18382 , n18222 , n18231 );
or ( n18383 , n18380 , n18381 , n18382 );
buf ( n18384 , n18211 );
xor ( n18385 , n18383 , n18384 );
and ( n18386 , n9964 , n12905 );
xor ( n18387 , n18385 , n18386 );
xor ( n18388 , n18379 , n18387 );
xor ( n18389 , n18370 , n18388 );
xor ( n18390 , n18334 , n18389 );
and ( n18391 , n18186 , n18247 );
xor ( n18392 , n18390 , n18391 );
xor ( n18393 , n18330 , n18392 );
and ( n18394 , n18182 , n18250 );
and ( n18395 , n18251 , n18254 );
or ( n18396 , n18394 , n18395 );
xor ( n18397 , n18393 , n18396 );
buf ( n18398 , n18397 );
not ( n18399 , n831 );
and ( n18400 , n18399 , n18329 );
and ( n18401 , n18398 , n831 );
or ( n18402 , n18400 , n18401 );
and ( n18403 , n18321 , n18322 );
and ( n18404 , n18269 , n18300 );
and ( n18405 , n18300 , n18319 );
and ( n18406 , n18269 , n18319 );
or ( n18407 , n18404 , n18405 , n18406 );
and ( n18408 , n18305 , n18309 );
and ( n18409 , n18309 , n18318 );
and ( n18410 , n18305 , n18318 );
or ( n18411 , n18408 , n18409 , n18410 );
and ( n18412 , n18274 , n18278 );
and ( n18413 , n18278 , n18283 );
and ( n18414 , n18274 , n18283 );
or ( n18415 , n18412 , n18413 , n18414 );
and ( n18416 , n18289 , n18293 );
and ( n18417 , n18293 , n18298 );
and ( n18418 , n18289 , n18298 );
or ( n18419 , n18416 , n18417 , n18418 );
xor ( n18420 , n18415 , n18419 );
and ( n18421 , n12724 , n10342 );
not ( n18422 , n18421 );
xnor ( n18423 , n18422 , n10291 );
and ( n18424 , n10837 , n12029 );
and ( n18425 , n11133 , n11739 );
nor ( n18426 , n18424 , n18425 );
xnor ( n18427 , n18426 , n12019 );
xor ( n18428 , n18423 , n18427 );
and ( n18429 , n10331 , n12782 );
and ( n18430 , n10548 , n12350 );
nor ( n18431 , n18429 , n18430 );
xnor ( n18432 , n18431 , n12733 );
xor ( n18433 , n18428 , n18432 );
xor ( n18434 , n18420 , n18433 );
xor ( n18435 , n18411 , n18434 );
and ( n18436 , n18314 , n18315 );
and ( n18437 , n18315 , n18317 );
and ( n18438 , n18314 , n18317 );
or ( n18439 , n18436 , n18437 , n18438 );
and ( n18440 , n18273 , n18284 );
and ( n18441 , n18284 , n18299 );
and ( n18442 , n18273 , n18299 );
or ( n18443 , n18440 , n18441 , n18442 );
xor ( n18444 , n18439 , n18443 );
and ( n18445 , n12010 , n10907 );
and ( n18446 , n12339 , n10543 );
nor ( n18447 , n18445 , n18446 );
xnor ( n18448 , n18447 , n10807 );
not ( n18449 , n18448 );
and ( n18450 , n11384 , n11411 );
and ( n18451 , n11699 , n11159 );
nor ( n18452 , n18450 , n18451 );
xnor ( n18453 , n18452 , n11417 );
xor ( n18454 , n18449 , n18453 );
and ( n18455 , n10090 , n12730 );
xor ( n18456 , n18454 , n18455 );
xor ( n18457 , n18444 , n18456 );
xor ( n18458 , n18435 , n18457 );
xor ( n18459 , n18407 , n18458 );
and ( n18460 , n18265 , n18320 );
xor ( n18461 , n18459 , n18460 );
xor ( n18462 , n18403 , n18461 );
and ( n18463 , n18261 , n18323 );
and ( n18464 , n18324 , n18327 );
or ( n18465 , n18463 , n18464 );
xor ( n18466 , n18462 , n18465 );
buf ( n18467 , n18466 );
and ( n18468 , n18390 , n18391 );
and ( n18469 , n18338 , n18369 );
and ( n18470 , n18369 , n18388 );
and ( n18471 , n18338 , n18388 );
or ( n18472 , n18469 , n18470 , n18471 );
and ( n18473 , n18374 , n18378 );
and ( n18474 , n18378 , n18387 );
and ( n18475 , n18374 , n18387 );
or ( n18476 , n18473 , n18474 , n18475 );
and ( n18477 , n18343 , n18347 );
and ( n18478 , n18347 , n18352 );
and ( n18479 , n18343 , n18352 );
or ( n18480 , n18477 , n18478 , n18479 );
and ( n18481 , n18358 , n18362 );
and ( n18482 , n18362 , n18367 );
and ( n18483 , n18358 , n18367 );
or ( n18484 , n18481 , n18482 , n18483 );
xor ( n18485 , n18480 , n18484 );
and ( n18486 , n12899 , n10477 );
not ( n18487 , n18486 );
xnor ( n18488 , n18487 , n10426 );
and ( n18489 , n10982 , n12194 );
and ( n18490 , n11274 , n11890 );
nor ( n18491 , n18489 , n18490 );
xnor ( n18492 , n18491 , n12184 );
xor ( n18493 , n18488 , n18492 );
and ( n18494 , n10466 , n12957 );
and ( n18495 , n10679 , n12511 );
nor ( n18496 , n18494 , n18495 );
xnor ( n18497 , n18496 , n12908 );
xor ( n18498 , n18493 , n18497 );
xor ( n18499 , n18485 , n18498 );
xor ( n18500 , n18476 , n18499 );
and ( n18501 , n18383 , n18384 );
and ( n18502 , n18384 , n18386 );
and ( n18503 , n18383 , n18386 );
or ( n18504 , n18501 , n18502 , n18503 );
and ( n18505 , n18342 , n18353 );
and ( n18506 , n18353 , n18368 );
and ( n18507 , n18342 , n18368 );
or ( n18508 , n18505 , n18506 , n18507 );
xor ( n18509 , n18504 , n18508 );
and ( n18510 , n12175 , n11052 );
and ( n18511 , n12500 , n10674 );
nor ( n18512 , n18510 , n18511 );
xnor ( n18513 , n18512 , n10952 );
not ( n18514 , n18513 );
and ( n18515 , n11539 , n11566 );
and ( n18516 , n11850 , n11300 );
nor ( n18517 , n18515 , n18516 );
xnor ( n18518 , n18517 , n11572 );
xor ( n18519 , n18514 , n18518 );
and ( n18520 , n10211 , n12905 );
xor ( n18521 , n18519 , n18520 );
xor ( n18522 , n18509 , n18521 );
xor ( n18523 , n18500 , n18522 );
xor ( n18524 , n18472 , n18523 );
and ( n18525 , n18334 , n18389 );
xor ( n18526 , n18524 , n18525 );
xor ( n18527 , n18468 , n18526 );
and ( n18528 , n18330 , n18392 );
and ( n18529 , n18393 , n18396 );
or ( n18530 , n18528 , n18529 );
xor ( n18531 , n18527 , n18530 );
buf ( n18532 , n18531 );
not ( n18533 , n831 );
and ( n18534 , n18533 , n18467 );
and ( n18535 , n18532 , n831 );
or ( n18536 , n18534 , n18535 );
and ( n18537 , n18459 , n18460 );
and ( n18538 , n18411 , n18434 );
and ( n18539 , n18434 , n18457 );
and ( n18540 , n18411 , n18457 );
or ( n18541 , n18538 , n18539 , n18540 );
and ( n18542 , n18415 , n18419 );
and ( n18543 , n18419 , n18433 );
and ( n18544 , n18415 , n18433 );
or ( n18545 , n18542 , n18543 , n18544 );
and ( n18546 , n18439 , n18443 );
and ( n18547 , n18443 , n18456 );
and ( n18548 , n18439 , n18456 );
or ( n18549 , n18546 , n18547 , n18548 );
xor ( n18550 , n18545 , n18549 );
and ( n18551 , n18449 , n18453 );
and ( n18552 , n18453 , n18455 );
and ( n18553 , n18449 , n18455 );
or ( n18554 , n18551 , n18552 , n18553 );
not ( n18555 , n10291 );
and ( n18556 , n12339 , n10907 );
and ( n18557 , n12724 , n10543 );
nor ( n18558 , n18556 , n18557 );
xnor ( n18559 , n18558 , n10807 );
xor ( n18560 , n18555 , n18559 );
and ( n18561 , n11133 , n12029 );
and ( n18562 , n11384 , n11739 );
nor ( n18563 , n18561 , n18562 );
xnor ( n18564 , n18563 , n12019 );
xor ( n18565 , n18560 , n18564 );
xor ( n18566 , n18554 , n18565 );
and ( n18567 , n18423 , n18427 );
and ( n18568 , n18427 , n18432 );
and ( n18569 , n18423 , n18432 );
or ( n18570 , n18567 , n18568 , n18569 );
buf ( n18571 , n18448 );
xor ( n18572 , n18570 , n18571 );
and ( n18573 , n11699 , n11411 );
and ( n18574 , n12010 , n11159 );
nor ( n18575 , n18573 , n18574 );
xnor ( n18576 , n18575 , n11417 );
and ( n18577 , n10548 , n12782 );
and ( n18578 , n10837 , n12350 );
nor ( n18579 , n18577 , n18578 );
xnor ( n18580 , n18579 , n12733 );
xor ( n18581 , n18576 , n18580 );
and ( n18582 , n10331 , n12730 );
xor ( n18583 , n18581 , n18582 );
xor ( n18584 , n18572 , n18583 );
xor ( n18585 , n18566 , n18584 );
xor ( n18586 , n18550 , n18585 );
xor ( n18587 , n18541 , n18586 );
and ( n18588 , n18407 , n18458 );
xor ( n18589 , n18587 , n18588 );
xor ( n18590 , n18537 , n18589 );
and ( n18591 , n18403 , n18461 );
and ( n18592 , n18462 , n18465 );
or ( n18593 , n18591 , n18592 );
xor ( n18594 , n18590 , n18593 );
buf ( n18595 , n18594 );
and ( n18596 , n18524 , n18525 );
and ( n18597 , n18476 , n18499 );
and ( n18598 , n18499 , n18522 );
and ( n18599 , n18476 , n18522 );
or ( n18600 , n18597 , n18598 , n18599 );
and ( n18601 , n18480 , n18484 );
and ( n18602 , n18484 , n18498 );
and ( n18603 , n18480 , n18498 );
or ( n18604 , n18601 , n18602 , n18603 );
and ( n18605 , n18504 , n18508 );
and ( n18606 , n18508 , n18521 );
and ( n18607 , n18504 , n18521 );
or ( n18608 , n18605 , n18606 , n18607 );
xor ( n18609 , n18604 , n18608 );
and ( n18610 , n18514 , n18518 );
and ( n18611 , n18518 , n18520 );
and ( n18612 , n18514 , n18520 );
or ( n18613 , n18610 , n18611 , n18612 );
not ( n18614 , n10426 );
and ( n18615 , n12500 , n11052 );
and ( n18616 , n12899 , n10674 );
nor ( n18617 , n18615 , n18616 );
xnor ( n18618 , n18617 , n10952 );
xor ( n18619 , n18614 , n18618 );
and ( n18620 , n11274 , n12194 );
and ( n18621 , n11539 , n11890 );
nor ( n18622 , n18620 , n18621 );
xnor ( n18623 , n18622 , n12184 );
xor ( n18624 , n18619 , n18623 );
xor ( n18625 , n18613 , n18624 );
and ( n18626 , n18488 , n18492 );
and ( n18627 , n18492 , n18497 );
and ( n18628 , n18488 , n18497 );
or ( n18629 , n18626 , n18627 , n18628 );
buf ( n18630 , n18513 );
xor ( n18631 , n18629 , n18630 );
and ( n18632 , n11850 , n11566 );
and ( n18633 , n12175 , n11300 );
nor ( n18634 , n18632 , n18633 );
xnor ( n18635 , n18634 , n11572 );
and ( n18636 , n10679 , n12957 );
and ( n18637 , n10982 , n12511 );
nor ( n18638 , n18636 , n18637 );
xnor ( n18639 , n18638 , n12908 );
xor ( n18640 , n18635 , n18639 );
and ( n18641 , n10466 , n12905 );
xor ( n18642 , n18640 , n18641 );
xor ( n18643 , n18631 , n18642 );
xor ( n18644 , n18625 , n18643 );
xor ( n18645 , n18609 , n18644 );
xor ( n18646 , n18600 , n18645 );
and ( n18647 , n18472 , n18523 );
xor ( n18648 , n18646 , n18647 );
xor ( n18649 , n18596 , n18648 );
and ( n18650 , n18468 , n18526 );
and ( n18651 , n18527 , n18530 );
or ( n18652 , n18650 , n18651 );
xor ( n18653 , n18649 , n18652 );
buf ( n18654 , n18653 );
not ( n18655 , n831 );
and ( n18656 , n18655 , n18595 );
and ( n18657 , n18654 , n831 );
or ( n18658 , n18656 , n18657 );
and ( n18659 , n18587 , n18588 );
and ( n18660 , n18545 , n18549 );
and ( n18661 , n18549 , n18585 );
and ( n18662 , n18545 , n18585 );
or ( n18663 , n18660 , n18661 , n18662 );
and ( n18664 , n18570 , n18571 );
and ( n18665 , n18571 , n18583 );
and ( n18666 , n18570 , n18583 );
or ( n18667 , n18664 , n18665 , n18666 );
and ( n18668 , n18554 , n18565 );
and ( n18669 , n18565 , n18584 );
and ( n18670 , n18554 , n18584 );
or ( n18671 , n18668 , n18669 , n18670 );
xor ( n18672 , n18667 , n18671 );
and ( n18673 , n18555 , n18559 );
and ( n18674 , n18559 , n18564 );
and ( n18675 , n18555 , n18564 );
or ( n18676 , n18673 , n18674 , n18675 );
and ( n18677 , n12724 , n10907 );
not ( n18678 , n18677 );
xnor ( n18679 , n18678 , n10807 );
and ( n18680 , n10837 , n12782 );
and ( n18681 , n11133 , n12350 );
nor ( n18682 , n18680 , n18681 );
xnor ( n18683 , n18682 , n12733 );
xor ( n18684 , n18679 , n18683 );
and ( n18685 , n10548 , n12730 );
xor ( n18686 , n18684 , n18685 );
xor ( n18687 , n18676 , n18686 );
and ( n18688 , n18576 , n18580 );
and ( n18689 , n18580 , n18582 );
and ( n18690 , n18576 , n18582 );
or ( n18691 , n18688 , n18689 , n18690 );
and ( n18692 , n12010 , n11411 );
and ( n18693 , n12339 , n11159 );
nor ( n18694 , n18692 , n18693 );
xnor ( n18695 , n18694 , n11417 );
not ( n18696 , n18695 );
xor ( n18697 , n18691 , n18696 );
and ( n18698 , n11384 , n12029 );
and ( n18699 , n11699 , n11739 );
nor ( n18700 , n18698 , n18699 );
xnor ( n18701 , n18700 , n12019 );
xor ( n18702 , n18697 , n18701 );
xor ( n18703 , n18687 , n18702 );
xor ( n18704 , n18672 , n18703 );
xor ( n18705 , n18663 , n18704 );
and ( n18706 , n18541 , n18586 );
xor ( n18707 , n18705 , n18706 );
xor ( n18708 , n18659 , n18707 );
and ( n18709 , n18537 , n18589 );
and ( n18710 , n18590 , n18593 );
or ( n18711 , n18709 , n18710 );
xor ( n18712 , n18708 , n18711 );
buf ( n18713 , n18712 );
and ( n18714 , n18646 , n18647 );
and ( n18715 , n18604 , n18608 );
and ( n18716 , n18608 , n18644 );
and ( n18717 , n18604 , n18644 );
or ( n18718 , n18715 , n18716 , n18717 );
and ( n18719 , n18629 , n18630 );
and ( n18720 , n18630 , n18642 );
and ( n18721 , n18629 , n18642 );
or ( n18722 , n18719 , n18720 , n18721 );
and ( n18723 , n18613 , n18624 );
and ( n18724 , n18624 , n18643 );
and ( n18725 , n18613 , n18643 );
or ( n18726 , n18723 , n18724 , n18725 );
xor ( n18727 , n18722 , n18726 );
and ( n18728 , n18614 , n18618 );
and ( n18729 , n18618 , n18623 );
and ( n18730 , n18614 , n18623 );
or ( n18731 , n18728 , n18729 , n18730 );
and ( n18732 , n12899 , n11052 );
not ( n18733 , n18732 );
xnor ( n18734 , n18733 , n10952 );
and ( n18735 , n10982 , n12957 );
and ( n18736 , n11274 , n12511 );
nor ( n18737 , n18735 , n18736 );
xnor ( n18738 , n18737 , n12908 );
xor ( n18739 , n18734 , n18738 );
and ( n18740 , n10679 , n12905 );
xor ( n18741 , n18739 , n18740 );
xor ( n18742 , n18731 , n18741 );
and ( n18743 , n18635 , n18639 );
and ( n18744 , n18639 , n18641 );
and ( n18745 , n18635 , n18641 );
or ( n18746 , n18743 , n18744 , n18745 );
and ( n18747 , n12175 , n11566 );
and ( n18748 , n12500 , n11300 );
nor ( n18749 , n18747 , n18748 );
xnor ( n18750 , n18749 , n11572 );
not ( n18751 , n18750 );
xor ( n18752 , n18746 , n18751 );
and ( n18753 , n11539 , n12194 );
and ( n18754 , n11850 , n11890 );
nor ( n18755 , n18753 , n18754 );
xnor ( n18756 , n18755 , n12184 );
xor ( n18757 , n18752 , n18756 );
xor ( n18758 , n18742 , n18757 );
xor ( n18759 , n18727 , n18758 );
xor ( n18760 , n18718 , n18759 );
and ( n18761 , n18600 , n18645 );
xor ( n18762 , n18760 , n18761 );
xor ( n18763 , n18714 , n18762 );
and ( n18764 , n18596 , n18648 );
and ( n18765 , n18649 , n18652 );
or ( n18766 , n18764 , n18765 );
xor ( n18767 , n18763 , n18766 );
buf ( n18768 , n18767 );
not ( n18769 , n831 );
and ( n18770 , n18769 , n18713 );
and ( n18771 , n18768 , n831 );
or ( n18772 , n18770 , n18771 );
and ( n18773 , n18667 , n18671 );
and ( n18774 , n18671 , n18703 );
and ( n18775 , n18667 , n18703 );
or ( n18776 , n18773 , n18774 , n18775 );
and ( n18777 , n18691 , n18696 );
and ( n18778 , n18696 , n18701 );
and ( n18779 , n18691 , n18701 );
or ( n18780 , n18777 , n18778 , n18779 );
and ( n18781 , n18676 , n18686 );
and ( n18782 , n18686 , n18702 );
and ( n18783 , n18676 , n18702 );
or ( n18784 , n18781 , n18782 , n18783 );
xor ( n18785 , n18780 , n18784 );
and ( n18786 , n18679 , n18683 );
and ( n18787 , n18683 , n18685 );
and ( n18788 , n18679 , n18685 );
or ( n18789 , n18786 , n18787 , n18788 );
not ( n18790 , n10807 );
and ( n18791 , n12339 , n11411 );
and ( n18792 , n12724 , n11159 );
nor ( n18793 , n18791 , n18792 );
xnor ( n18794 , n18793 , n11417 );
xor ( n18795 , n18790 , n18794 );
and ( n18796 , n11133 , n12782 );
and ( n18797 , n11384 , n12350 );
nor ( n18798 , n18796 , n18797 );
xnor ( n18799 , n18798 , n12733 );
xor ( n18800 , n18795 , n18799 );
xor ( n18801 , n18789 , n18800 );
buf ( n18802 , n18695 );
and ( n18803 , n11699 , n12029 );
and ( n18804 , n12010 , n11739 );
nor ( n18805 , n18803 , n18804 );
xnor ( n18806 , n18805 , n12019 );
xor ( n18807 , n18802 , n18806 );
and ( n18808 , n10837 , n12730 );
xor ( n18809 , n18807 , n18808 );
xor ( n18810 , n18801 , n18809 );
xor ( n18811 , n18785 , n18810 );
xor ( n18812 , n18776 , n18811 );
and ( n18813 , n18663 , n18704 );
xor ( n18814 , n18812 , n18813 );
and ( n18815 , n18705 , n18706 );
xor ( n18816 , n18814 , n18815 );
and ( n18817 , n18659 , n18707 );
and ( n18818 , n18708 , n18711 );
or ( n18819 , n18817 , n18818 );
xor ( n18820 , n18816 , n18819 );
buf ( n18821 , n18820 );
and ( n18822 , n18722 , n18726 );
and ( n18823 , n18726 , n18758 );
and ( n18824 , n18722 , n18758 );
or ( n18825 , n18822 , n18823 , n18824 );
and ( n18826 , n18746 , n18751 );
and ( n18827 , n18751 , n18756 );
and ( n18828 , n18746 , n18756 );
or ( n18829 , n18826 , n18827 , n18828 );
and ( n18830 , n18731 , n18741 );
and ( n18831 , n18741 , n18757 );
and ( n18832 , n18731 , n18757 );
or ( n18833 , n18830 , n18831 , n18832 );
xor ( n18834 , n18829 , n18833 );
and ( n18835 , n18734 , n18738 );
and ( n18836 , n18738 , n18740 );
and ( n18837 , n18734 , n18740 );
or ( n18838 , n18835 , n18836 , n18837 );
not ( n18839 , n10952 );
and ( n18840 , n12500 , n11566 );
and ( n18841 , n12899 , n11300 );
nor ( n18842 , n18840 , n18841 );
xnor ( n18843 , n18842 , n11572 );
xor ( n18844 , n18839 , n18843 );
and ( n18845 , n11274 , n12957 );
and ( n18846 , n11539 , n12511 );
nor ( n18847 , n18845 , n18846 );
xnor ( n18848 , n18847 , n12908 );
xor ( n18849 , n18844 , n18848 );
xor ( n18850 , n18838 , n18849 );
buf ( n18851 , n18750 );
and ( n18852 , n11850 , n12194 );
and ( n18853 , n12175 , n11890 );
nor ( n18854 , n18852 , n18853 );
xnor ( n18855 , n18854 , n12184 );
xor ( n18856 , n18851 , n18855 );
and ( n18857 , n10982 , n12905 );
xor ( n18858 , n18856 , n18857 );
xor ( n18859 , n18850 , n18858 );
xor ( n18860 , n18834 , n18859 );
xor ( n18861 , n18825 , n18860 );
and ( n18862 , n18718 , n18759 );
xor ( n18863 , n18861 , n18862 );
and ( n18864 , n18760 , n18761 );
xor ( n18865 , n18863 , n18864 );
and ( n18866 , n18714 , n18762 );
and ( n18867 , n18763 , n18766 );
or ( n18868 , n18866 , n18867 );
xor ( n18869 , n18865 , n18868 );
buf ( n18870 , n18869 );
not ( n18871 , n831 );
and ( n18872 , n18871 , n18821 );
and ( n18873 , n18870 , n831 );
or ( n18874 , n18872 , n18873 );
and ( n18875 , n18812 , n18813 );
and ( n18876 , n18780 , n18784 );
and ( n18877 , n18784 , n18810 );
and ( n18878 , n18780 , n18810 );
or ( n18879 , n18876 , n18877 , n18878 );
and ( n18880 , n18802 , n18806 );
and ( n18881 , n18806 , n18808 );
and ( n18882 , n18802 , n18808 );
or ( n18883 , n18880 , n18881 , n18882 );
and ( n18884 , n18789 , n18800 );
and ( n18885 , n18800 , n18809 );
and ( n18886 , n18789 , n18809 );
or ( n18887 , n18884 , n18885 , n18886 );
xor ( n18888 , n18883 , n18887 );
and ( n18889 , n18790 , n18794 );
and ( n18890 , n18794 , n18799 );
and ( n18891 , n18790 , n18799 );
or ( n18892 , n18889 , n18890 , n18891 );
and ( n18893 , n12724 , n11411 );
not ( n18894 , n18893 );
xnor ( n18895 , n18894 , n11417 );
not ( n18896 , n18895 );
xor ( n18897 , n18892 , n18896 );
and ( n18898 , n12010 , n12029 );
and ( n18899 , n12339 , n11739 );
nor ( n18900 , n18898 , n18899 );
xnor ( n18901 , n18900 , n12019 );
and ( n18902 , n11384 , n12782 );
and ( n18903 , n11699 , n12350 );
nor ( n18904 , n18902 , n18903 );
xnor ( n18905 , n18904 , n12733 );
xor ( n18906 , n18901 , n18905 );
and ( n18907 , n11133 , n12730 );
xor ( n18908 , n18906 , n18907 );
xor ( n18909 , n18897 , n18908 );
xor ( n18910 , n18888 , n18909 );
xor ( n18911 , n18879 , n18910 );
and ( n18912 , n18776 , n18811 );
xor ( n18913 , n18911 , n18912 );
xor ( n18914 , n18875 , n18913 );
and ( n18915 , n18814 , n18815 );
and ( n18916 , n18816 , n18819 );
or ( n18917 , n18915 , n18916 );
xor ( n18918 , n18914 , n18917 );
buf ( n18919 , n18918 );
and ( n18920 , n18861 , n18862 );
and ( n18921 , n18829 , n18833 );
and ( n18922 , n18833 , n18859 );
and ( n18923 , n18829 , n18859 );
or ( n18924 , n18921 , n18922 , n18923 );
and ( n18925 , n18851 , n18855 );
and ( n18926 , n18855 , n18857 );
and ( n18927 , n18851 , n18857 );
or ( n18928 , n18925 , n18926 , n18927 );
and ( n18929 , n18838 , n18849 );
and ( n18930 , n18849 , n18858 );
and ( n18931 , n18838 , n18858 );
or ( n18932 , n18929 , n18930 , n18931 );
xor ( n18933 , n18928 , n18932 );
and ( n18934 , n18839 , n18843 );
and ( n18935 , n18843 , n18848 );
and ( n18936 , n18839 , n18848 );
or ( n18937 , n18934 , n18935 , n18936 );
and ( n18938 , n12899 , n11566 );
not ( n18939 , n18938 );
xnor ( n18940 , n18939 , n11572 );
not ( n18941 , n18940 );
xor ( n18942 , n18937 , n18941 );
and ( n18943 , n12175 , n12194 );
and ( n18944 , n12500 , n11890 );
nor ( n18945 , n18943 , n18944 );
xnor ( n18946 , n18945 , n12184 );
and ( n18947 , n11539 , n12957 );
and ( n18948 , n11850 , n12511 );
nor ( n18949 , n18947 , n18948 );
xnor ( n18950 , n18949 , n12908 );
xor ( n18951 , n18946 , n18950 );
and ( n18952 , n11274 , n12905 );
xor ( n18953 , n18951 , n18952 );
xor ( n18954 , n18942 , n18953 );
xor ( n18955 , n18933 , n18954 );
xor ( n18956 , n18924 , n18955 );
and ( n18957 , n18825 , n18860 );
xor ( n18958 , n18956 , n18957 );
xor ( n18959 , n18920 , n18958 );
and ( n18960 , n18863 , n18864 );
and ( n18961 , n18865 , n18868 );
or ( n18962 , n18960 , n18961 );
xor ( n18963 , n18959 , n18962 );
buf ( n18964 , n18963 );
not ( n18965 , n831 );
and ( n18966 , n18965 , n18919 );
and ( n18967 , n18964 , n831 );
or ( n18968 , n18966 , n18967 );
and ( n18969 , n18911 , n18912 );
and ( n18970 , n18883 , n18887 );
and ( n18971 , n18887 , n18909 );
and ( n18972 , n18883 , n18909 );
or ( n18973 , n18970 , n18971 , n18972 );
and ( n18974 , n18892 , n18896 );
and ( n18975 , n18896 , n18908 );
and ( n18976 , n18892 , n18908 );
or ( n18977 , n18974 , n18975 , n18976 );
not ( n18978 , n11417 );
and ( n18979 , n12339 , n12029 );
and ( n18980 , n12724 , n11739 );
nor ( n18981 , n18979 , n18980 );
xnor ( n18982 , n18981 , n12019 );
xor ( n18983 , n18978 , n18982 );
and ( n18984 , n11384 , n12730 );
xor ( n18985 , n18983 , n18984 );
xor ( n18986 , n18977 , n18985 );
and ( n18987 , n18901 , n18905 );
and ( n18988 , n18905 , n18907 );
and ( n18989 , n18901 , n18907 );
or ( n18990 , n18987 , n18988 , n18989 );
buf ( n18991 , n18895 );
xor ( n18992 , n18990 , n18991 );
and ( n18993 , n11699 , n12782 );
and ( n18994 , n12010 , n12350 );
nor ( n18995 , n18993 , n18994 );
xnor ( n18996 , n18995 , n12733 );
xor ( n18997 , n18992 , n18996 );
xor ( n18998 , n18986 , n18997 );
xor ( n18999 , n18973 , n18998 );
and ( n19000 , n18879 , n18910 );
xor ( n19001 , n18999 , n19000 );
xor ( n19002 , n18969 , n19001 );
and ( n19003 , n18875 , n18913 );
and ( n19004 , n18914 , n18917 );
or ( n19005 , n19003 , n19004 );
xor ( n19006 , n19002 , n19005 );
buf ( n19007 , n19006 );
and ( n19008 , n18956 , n18957 );
and ( n19009 , n18928 , n18932 );
and ( n19010 , n18932 , n18954 );
and ( n19011 , n18928 , n18954 );
or ( n19012 , n19009 , n19010 , n19011 );
and ( n19013 , n18937 , n18941 );
and ( n19014 , n18941 , n18953 );
and ( n19015 , n18937 , n18953 );
or ( n19016 , n19013 , n19014 , n19015 );
not ( n19017 , n11572 );
and ( n19018 , n12500 , n12194 );
and ( n19019 , n12899 , n11890 );
nor ( n19020 , n19018 , n19019 );
xnor ( n19021 , n19020 , n12184 );
xor ( n19022 , n19017 , n19021 );
and ( n19023 , n11539 , n12905 );
xor ( n19024 , n19022 , n19023 );
xor ( n19025 , n19016 , n19024 );
and ( n19026 , n18946 , n18950 );
and ( n19027 , n18950 , n18952 );
and ( n19028 , n18946 , n18952 );
or ( n19029 , n19026 , n19027 , n19028 );
buf ( n19030 , n18940 );
xor ( n19031 , n19029 , n19030 );
and ( n19032 , n11850 , n12957 );
and ( n19033 , n12175 , n12511 );
nor ( n19034 , n19032 , n19033 );
xnor ( n19035 , n19034 , n12908 );
xor ( n19036 , n19031 , n19035 );
xor ( n19037 , n19025 , n19036 );
xor ( n19038 , n19012 , n19037 );
and ( n19039 , n18924 , n18955 );
xor ( n19040 , n19038 , n19039 );
xor ( n19041 , n19008 , n19040 );
and ( n19042 , n18920 , n18958 );
and ( n19043 , n18959 , n18962 );
or ( n19044 , n19042 , n19043 );
xor ( n19045 , n19041 , n19044 );
buf ( n19046 , n19045 );
not ( n19047 , n831 );
and ( n19048 , n19047 , n19007 );
and ( n19049 , n19046 , n831 );
or ( n19050 , n19048 , n19049 );
and ( n19051 , n18999 , n19000 );
and ( n19052 , n18977 , n18985 );
and ( n19053 , n18985 , n18997 );
and ( n19054 , n18977 , n18997 );
or ( n19055 , n19052 , n19053 , n19054 );
and ( n19056 , n18978 , n18982 );
and ( n19057 , n18982 , n18984 );
and ( n19058 , n18978 , n18984 );
or ( n19059 , n19056 , n19057 , n19058 );
and ( n19060 , n18990 , n18991 );
and ( n19061 , n18991 , n18996 );
and ( n19062 , n18990 , n18996 );
or ( n19063 , n19060 , n19061 , n19062 );
xor ( n19064 , n19059 , n19063 );
and ( n19065 , n12724 , n12029 );
not ( n19066 , n19065 );
xnor ( n19067 , n19066 , n12019 );
not ( n19068 , n19067 );
and ( n19069 , n12010 , n12782 );
and ( n19070 , n12339 , n12350 );
nor ( n19071 , n19069 , n19070 );
xnor ( n19072 , n19071 , n12733 );
xor ( n19073 , n19068 , n19072 );
and ( n19074 , n11699 , n12730 );
xor ( n19075 , n19073 , n19074 );
xor ( n19076 , n19064 , n19075 );
xor ( n19077 , n19055 , n19076 );
and ( n19078 , n18973 , n18998 );
xor ( n19079 , n19077 , n19078 );
xor ( n19080 , n19051 , n19079 );
and ( n19081 , n18969 , n19001 );
and ( n19082 , n19002 , n19005 );
or ( n19083 , n19081 , n19082 );
xor ( n19084 , n19080 , n19083 );
buf ( n19085 , n19084 );
and ( n19086 , n19038 , n19039 );
and ( n19087 , n19016 , n19024 );
and ( n19088 , n19024 , n19036 );
and ( n19089 , n19016 , n19036 );
or ( n19090 , n19087 , n19088 , n19089 );
and ( n19091 , n19017 , n19021 );
and ( n19092 , n19021 , n19023 );
and ( n19093 , n19017 , n19023 );
or ( n19094 , n19091 , n19092 , n19093 );
and ( n19095 , n19029 , n19030 );
and ( n19096 , n19030 , n19035 );
and ( n19097 , n19029 , n19035 );
or ( n19098 , n19095 , n19096 , n19097 );
xor ( n19099 , n19094 , n19098 );
and ( n19100 , n12899 , n12194 );
not ( n19101 , n19100 );
xnor ( n19102 , n19101 , n12184 );
not ( n19103 , n19102 );
and ( n19104 , n12175 , n12957 );
and ( n19105 , n12500 , n12511 );
nor ( n19106 , n19104 , n19105 );
xnor ( n19107 , n19106 , n12908 );
xor ( n19108 , n19103 , n19107 );
and ( n19109 , n11850 , n12905 );
xor ( n19110 , n19108 , n19109 );
xor ( n19111 , n19099 , n19110 );
xor ( n19112 , n19090 , n19111 );
and ( n19113 , n19012 , n19037 );
xor ( n19114 , n19112 , n19113 );
xor ( n19115 , n19086 , n19114 );
and ( n19116 , n19008 , n19040 );
and ( n19117 , n19041 , n19044 );
or ( n19118 , n19116 , n19117 );
xor ( n19119 , n19115 , n19118 );
buf ( n19120 , n19119 );
not ( n19121 , n831 );
and ( n19122 , n19121 , n19085 );
and ( n19123 , n19120 , n831 );
or ( n19124 , n19122 , n19123 );
and ( n19125 , n19059 , n19063 );
and ( n19126 , n19063 , n19075 );
and ( n19127 , n19059 , n19075 );
or ( n19128 , n19125 , n19126 , n19127 );
and ( n19129 , n19068 , n19072 );
and ( n19130 , n19072 , n19074 );
and ( n19131 , n19068 , n19074 );
or ( n19132 , n19129 , n19130 , n19131 );
buf ( n19133 , n19067 );
xor ( n19134 , n19132 , n19133 );
not ( n19135 , n12019 );
and ( n19136 , n12339 , n12782 );
and ( n19137 , n12724 , n12350 );
nor ( n19138 , n19136 , n19137 );
xnor ( n19139 , n19138 , n12733 );
xor ( n19140 , n19135 , n19139 );
and ( n19141 , n12010 , n12730 );
xor ( n19142 , n19140 , n19141 );
xor ( n19143 , n19134 , n19142 );
xor ( n19144 , n19128 , n19143 );
and ( n19145 , n19055 , n19076 );
xor ( n19146 , n19144 , n19145 );
and ( n19147 , n19077 , n19078 );
xor ( n19148 , n19146 , n19147 );
and ( n19149 , n19051 , n19079 );
and ( n19150 , n19080 , n19083 );
or ( n19151 , n19149 , n19150 );
xor ( n19152 , n19148 , n19151 );
buf ( n19153 , n19152 );
and ( n19154 , n19094 , n19098 );
and ( n19155 , n19098 , n19110 );
and ( n19156 , n19094 , n19110 );
or ( n19157 , n19154 , n19155 , n19156 );
and ( n19158 , n19103 , n19107 );
and ( n19159 , n19107 , n19109 );
and ( n19160 , n19103 , n19109 );
or ( n19161 , n19158 , n19159 , n19160 );
buf ( n19162 , n19102 );
xor ( n19163 , n19161 , n19162 );
not ( n19164 , n12184 );
and ( n19165 , n12500 , n12957 );
and ( n19166 , n12899 , n12511 );
nor ( n19167 , n19165 , n19166 );
xnor ( n19168 , n19167 , n12908 );
xor ( n19169 , n19164 , n19168 );
and ( n19170 , n12175 , n12905 );
xor ( n19171 , n19169 , n19170 );
xor ( n19172 , n19163 , n19171 );
xor ( n19173 , n19157 , n19172 );
and ( n19174 , n19090 , n19111 );
xor ( n19175 , n19173 , n19174 );
and ( n19176 , n19112 , n19113 );
xor ( n19177 , n19175 , n19176 );
and ( n19178 , n19086 , n19114 );
and ( n19179 , n19115 , n19118 );
or ( n19180 , n19178 , n19179 );
xor ( n19181 , n19177 , n19180 );
buf ( n19182 , n19181 );
not ( n19183 , n831 );
and ( n19184 , n19183 , n19153 );
and ( n19185 , n19182 , n831 );
or ( n19186 , n19184 , n19185 );
and ( n19187 , n19144 , n19145 );
and ( n19188 , n19132 , n19133 );
and ( n19189 , n19133 , n19142 );
and ( n19190 , n19132 , n19142 );
or ( n19191 , n19188 , n19189 , n19190 );
and ( n19192 , n19135 , n19139 );
and ( n19193 , n19139 , n19141 );
and ( n19194 , n19135 , n19141 );
or ( n19195 , n19192 , n19193 , n19194 );
and ( n19196 , n12724 , n12782 );
not ( n19197 , n19196 );
xnor ( n19198 , n19197 , n12733 );
xor ( n19199 , n19195 , n19198 );
and ( n19200 , n12339 , n12730 );
not ( n19201 , n19200 );
xor ( n19202 , n19199 , n19201 );
xor ( n19203 , n19191 , n19202 );
and ( n19204 , n19128 , n19143 );
xor ( n19205 , n19203 , n19204 );
xor ( n19206 , n19187 , n19205 );
and ( n19207 , n19146 , n19147 );
and ( n19208 , n19148 , n19151 );
or ( n19209 , n19207 , n19208 );
xor ( n19210 , n19206 , n19209 );
buf ( n19211 , n19210 );
and ( n19212 , n19173 , n19174 );
and ( n19213 , n19161 , n19162 );
and ( n19214 , n19162 , n19171 );
and ( n19215 , n19161 , n19171 );
or ( n19216 , n19213 , n19214 , n19215 );
and ( n19217 , n19164 , n19168 );
and ( n19218 , n19168 , n19170 );
and ( n19219 , n19164 , n19170 );
or ( n19220 , n19217 , n19218 , n19219 );
and ( n19221 , n12899 , n12957 );
not ( n19222 , n19221 );
xnor ( n19223 , n19222 , n12908 );
xor ( n19224 , n19220 , n19223 );
and ( n19225 , n12500 , n12905 );
not ( n19226 , n19225 );
xor ( n19227 , n19224 , n19226 );
xor ( n19228 , n19216 , n19227 );
and ( n19229 , n19157 , n19172 );
xor ( n19230 , n19228 , n19229 );
xor ( n19231 , n19212 , n19230 );
and ( n19232 , n19175 , n19176 );
and ( n19233 , n19177 , n19180 );
or ( n19234 , n19232 , n19233 );
xor ( n19235 , n19231 , n19234 );
buf ( n19236 , n19235 );
not ( n19237 , n831 );
and ( n19238 , n19237 , n19211 );
and ( n19239 , n19236 , n831 );
or ( n19240 , n19238 , n19239 );
and ( n19241 , n19195 , n19198 );
and ( n19242 , n19198 , n19201 );
and ( n19243 , n19195 , n19201 );
or ( n19244 , n19241 , n19242 , n19243 );
and ( n19245 , n19191 , n19202 );
xor ( n19246 , n19244 , n19245 );
buf ( n19247 , n19200 );
not ( n19248 , n12733 );
xor ( n19249 , n19247 , n19248 );
and ( n19250 , n12724 , n12730 );
xor ( n19251 , n19249 , n19250 );
xor ( n19252 , n19246 , n19251 );
and ( n19253 , n19203 , n19204 );
xor ( n19254 , n19252 , n19253 );
and ( n19255 , n19187 , n19205 );
and ( n19256 , n19206 , n19209 );
or ( n19257 , n19255 , n19256 );
xor ( n19258 , n19254 , n19257 );
buf ( n19259 , n19258 );
and ( n19260 , n19220 , n19223 );
and ( n19261 , n19223 , n19226 );
and ( n19262 , n19220 , n19226 );
or ( n19263 , n19260 , n19261 , n19262 );
and ( n19264 , n19216 , n19227 );
xor ( n19265 , n19263 , n19264 );
buf ( n19266 , n19225 );
not ( n19267 , n12908 );
xor ( n19268 , n19266 , n19267 );
and ( n19269 , n12899 , n12905 );
xor ( n19270 , n19268 , n19269 );
xor ( n19271 , n19265 , n19270 );
and ( n19272 , n19228 , n19229 );
xor ( n19273 , n19271 , n19272 );
and ( n19274 , n19212 , n19230 );
and ( n19275 , n19231 , n19234 );
or ( n19276 , n19274 , n19275 );
xor ( n19277 , n19273 , n19276 );
buf ( n19278 , n19277 );
not ( n19279 , n831 );
and ( n19280 , n19279 , n19259 );
and ( n19281 , n19278 , n831 );
or ( n19282 , n19280 , n19281 );
buf ( n19283 , n19282 );
buf ( n19284 , n19240 );
buf ( n19285 , n19186 );
buf ( n19286 , n19124 );
buf ( n19287 , n19050 );
buf ( n19288 , n18968 );
buf ( n19289 , n18874 );
buf ( n19290 , n18772 );
buf ( n19291 , n18658 );
buf ( n19292 , n18536 );
buf ( n19293 , n18402 );
buf ( n19294 , n18260 );
buf ( n19295 , n18106 );
buf ( n19296 , n17944 );
buf ( n19297 , n17770 );
buf ( n19298 , n17588 );
buf ( n19299 , n17394 );
buf ( n19300 , n17192 );
buf ( n19301 , n16978 );
buf ( n19302 , n16756 );
buf ( n19303 , n16522 );
buf ( n19304 , n16280 );
buf ( n19305 , n16026 );
buf ( n19306 , n15764 );
buf ( n19307 , n15490 );
buf ( n19308 , n15208 );
buf ( n19309 , n14914 );
buf ( n19310 , n14612 );
buf ( n19311 , n14298 );
buf ( n19312 , n13976 );
buf ( n19313 , n13646 );
buf ( n19314 , n13324 );
buf ( n19315 , n12996 );
buf ( n19316 , n12642 );
buf ( n19317 , n12316 );
buf ( n19318 , n11982 );
buf ( n19319 , n11676 );
buf ( n19320 , n11362 );
buf ( n19321 , n11076 );
buf ( n19322 , n10782 );
buf ( n19323 , n10516 );
buf ( n19324 , n10242 );
buf ( n19325 , n9996 );
buf ( n19326 , n9742 );
buf ( n19327 , n9516 );
buf ( n19328 , n9282 );
buf ( n19329 , n9076 );
buf ( n19330 , n8862 );
buf ( n19331 , n8676 );
buf ( n19332 , n8482 );
buf ( n19333 , n8316 );
buf ( n19334 , n8142 );
buf ( n19335 , n7996 );
buf ( n19336 , n7842 );
buf ( n19337 , n7716 );
buf ( n19338 , n7582 );
buf ( n19339 , n7476 );
buf ( n19340 , n7362 );
buf ( n19341 , n7276 );
buf ( n19342 , n7182 );
buf ( n19343 , n7116 );
buf ( n19344 , n7042 );
buf ( n19345 , n6996 );
buf ( n19346 , n6952 );
buf ( n19347 , n6804 );
buf ( n19348 , n6806 );
buf ( n19349 , n6808 );
buf ( n19350 , n6810 );
buf ( n19351 , n6812 );
buf ( n19352 , n6814 );
buf ( n19353 , n6816 );
buf ( n19354 , n6818 );
buf ( n19355 , n6820 );
buf ( n19356 , n6822 );
buf ( n19357 , n6824 );
buf ( n19358 , n6826 );
buf ( n19359 , n6828 );
buf ( n19360 , n6830 );
buf ( n19361 , n6832 );
buf ( n19362 , n6834 );
buf ( n19363 , n6836 );
buf ( n19364 , n6838 );
buf ( n19365 , n6840 );
buf ( n19366 , n6842 );
buf ( n19367 , n6844 );
buf ( n19368 , n6846 );
buf ( n19369 , n6848 );
buf ( n19370 , n6850 );
buf ( n19371 , n6852 );
buf ( n19372 , n6854 );
buf ( n19373 , n6856 );
buf ( n19374 , n6858 );
buf ( n19375 , n6860 );
buf ( n19376 , n6862 );
buf ( n19377 , n6864 );
buf ( n19378 , n6866 );
buf ( n19379 , n6868 );
buf ( n19380 , n6870 );
buf ( n19381 , n6872 );
buf ( n19382 , n6874 );
buf ( n19383 , n6876 );
buf ( n19384 , n6878 );
buf ( n19385 , n6880 );
buf ( n19386 , n6882 );
buf ( n19387 , n6884 );
buf ( n19388 , n6886 );
buf ( n19389 , n6888 );
buf ( n19390 , n6890 );
buf ( n19391 , n6892 );
buf ( n19392 , n6894 );
buf ( n19393 , n6896 );
buf ( n19394 , n6898 );
buf ( n19395 , n6900 );
buf ( n19396 , n6902 );
buf ( n19397 , n6904 );
buf ( n19398 , n6906 );
buf ( n19399 , n6908 );
buf ( n19400 , n6910 );
buf ( n19401 , n6912 );
buf ( n19402 , n6914 );
buf ( n19403 , n6916 );
buf ( n19404 , n6918 );
buf ( n19405 , n6920 );
buf ( n19406 , n6922 );
buf ( n19407 , n6924 );
buf ( n19408 , n6926 );
buf ( n19409 , n6928 );
buf ( n19410 , n6930 );
buf ( n19411 , n19349 );
buf ( n19412 , n19350 );
buf ( n19413 , n19351 );
and ( n19414 , n19412 , n19413 );
not ( n19415 , n19414 );
and ( n19416 , n19411 , n19415 );
not ( n19417 , n19416 );
buf ( n19418 , n19284 );
buf ( n19419 , n19347 );
buf ( n19420 , n19348 );
xor ( n19421 , n19419 , n19420 );
xor ( n19422 , n19420 , n19411 );
not ( n19423 , n19422 );
and ( n19424 , n19421 , n19423 );
and ( n19425 , n19418 , n19424 );
buf ( n19426 , n19283 );
and ( n19427 , n19426 , n19422 );
nor ( n19428 , n19425 , n19427 );
and ( n19429 , n19420 , n19411 );
not ( n19430 , n19429 );
and ( n19431 , n19419 , n19430 );
xnor ( n19432 , n19428 , n19431 );
and ( n19433 , n19417 , n19432 );
buf ( n19434 , n19285 );
and ( n19435 , n19434 , n19419 );
and ( n19436 , n19432 , n19435 );
and ( n19437 , n19417 , n19435 );
or ( n19438 , n19433 , n19436 , n19437 );
and ( n19439 , n19426 , n19424 );
not ( n19440 , n19439 );
xnor ( n19441 , n19440 , n19431 );
and ( n19442 , n19438 , n19441 );
and ( n19443 , n19418 , n19419 );
not ( n19444 , n19443 );
and ( n19445 , n19441 , n19444 );
and ( n19446 , n19438 , n19444 );
or ( n19447 , n19442 , n19445 , n19446 );
buf ( n19448 , n19443 );
not ( n19449 , n19431 );
xor ( n19450 , n19448 , n19449 );
and ( n19451 , n19426 , n19419 );
xor ( n19452 , n19450 , n19451 );
xor ( n19453 , n19447 , n19452 );
xor ( n19454 , n19438 , n19441 );
xor ( n19455 , n19454 , n19444 );
xor ( n19456 , n19411 , n19412 );
xor ( n19457 , n19412 , n19413 );
not ( n19458 , n19457 );
and ( n19459 , n19456 , n19458 );
and ( n19460 , n19426 , n19459 );
not ( n19461 , n19460 );
xnor ( n19462 , n19461 , n19416 );
not ( n19463 , n19462 );
and ( n19464 , n19434 , n19424 );
and ( n19465 , n19418 , n19422 );
nor ( n19466 , n19464 , n19465 );
xnor ( n19467 , n19466 , n19431 );
and ( n19468 , n19463 , n19467 );
buf ( n19469 , n19286 );
and ( n19470 , n19469 , n19419 );
and ( n19471 , n19467 , n19470 );
and ( n19472 , n19463 , n19470 );
or ( n19473 , n19468 , n19471 , n19472 );
buf ( n19474 , n19462 );
and ( n19475 , n19473 , n19474 );
xor ( n19476 , n19417 , n19432 );
xor ( n19477 , n19476 , n19435 );
and ( n19478 , n19474 , n19477 );
and ( n19479 , n19473 , n19477 );
or ( n19480 , n19475 , n19478 , n19479 );
and ( n19481 , n19455 , n19480 );
xor ( n19482 , n19455 , n19480 );
xor ( n19483 , n19473 , n19474 );
xor ( n19484 , n19483 , n19477 );
buf ( n19485 , n19352 );
buf ( n19486 , n19353 );
and ( n19487 , n19485 , n19486 );
not ( n19488 , n19487 );
and ( n19489 , n19413 , n19488 );
not ( n19490 , n19489 );
and ( n19491 , n19418 , n19459 );
and ( n19492 , n19426 , n19457 );
nor ( n19493 , n19491 , n19492 );
xnor ( n19494 , n19493 , n19416 );
and ( n19495 , n19490 , n19494 );
buf ( n19496 , n19287 );
and ( n19497 , n19496 , n19419 );
and ( n19498 , n19494 , n19497 );
and ( n19499 , n19490 , n19497 );
or ( n19500 , n19495 , n19498 , n19499 );
and ( n19501 , n19434 , n19459 );
and ( n19502 , n19418 , n19457 );
nor ( n19503 , n19501 , n19502 );
xnor ( n19504 , n19503 , n19416 );
and ( n19505 , n19496 , n19424 );
and ( n19506 , n19469 , n19422 );
nor ( n19507 , n19505 , n19506 );
xnor ( n19508 , n19507 , n19431 );
and ( n19509 , n19504 , n19508 );
buf ( n19510 , n19288 );
and ( n19511 , n19510 , n19419 );
and ( n19512 , n19508 , n19511 );
and ( n19513 , n19504 , n19511 );
or ( n19514 , n19509 , n19512 , n19513 );
xor ( n19515 , n19413 , n19485 );
xor ( n19516 , n19485 , n19486 );
not ( n19517 , n19516 );
and ( n19518 , n19515 , n19517 );
and ( n19519 , n19426 , n19518 );
not ( n19520 , n19519 );
xnor ( n19521 , n19520 , n19489 );
buf ( n19522 , n19521 );
and ( n19523 , n19514 , n19522 );
and ( n19524 , n19469 , n19424 );
and ( n19525 , n19434 , n19422 );
nor ( n19526 , n19524 , n19525 );
xnor ( n19527 , n19526 , n19431 );
and ( n19528 , n19522 , n19527 );
and ( n19529 , n19514 , n19527 );
or ( n19530 , n19523 , n19528 , n19529 );
and ( n19531 , n19500 , n19530 );
xor ( n19532 , n19463 , n19467 );
xor ( n19533 , n19532 , n19470 );
and ( n19534 , n19530 , n19533 );
and ( n19535 , n19500 , n19533 );
or ( n19536 , n19531 , n19534 , n19535 );
and ( n19537 , n19484 , n19536 );
xor ( n19538 , n19484 , n19536 );
xor ( n19539 , n19500 , n19530 );
xor ( n19540 , n19539 , n19533 );
buf ( n19541 , n19354 );
buf ( n19542 , n19355 );
and ( n19543 , n19541 , n19542 );
not ( n19544 , n19543 );
and ( n19545 , n19486 , n19544 );
not ( n19546 , n19545 );
and ( n19547 , n19418 , n19518 );
and ( n19548 , n19426 , n19516 );
nor ( n19549 , n19547 , n19548 );
xnor ( n19550 , n19549 , n19489 );
and ( n19551 , n19546 , n19550 );
and ( n19552 , n19510 , n19424 );
and ( n19553 , n19496 , n19422 );
nor ( n19554 , n19552 , n19553 );
xnor ( n19555 , n19554 , n19431 );
and ( n19556 , n19550 , n19555 );
and ( n19557 , n19546 , n19555 );
or ( n19558 , n19551 , n19556 , n19557 );
not ( n19559 , n19521 );
and ( n19560 , n19558 , n19559 );
xor ( n19561 , n19504 , n19508 );
xor ( n19562 , n19561 , n19511 );
and ( n19563 , n19559 , n19562 );
and ( n19564 , n19558 , n19562 );
or ( n19565 , n19560 , n19563 , n19564 );
xor ( n19566 , n19490 , n19494 );
xor ( n19567 , n19566 , n19497 );
and ( n19568 , n19565 , n19567 );
xor ( n19569 , n19514 , n19522 );
xor ( n19570 , n19569 , n19527 );
and ( n19571 , n19567 , n19570 );
and ( n19572 , n19565 , n19570 );
or ( n19573 , n19568 , n19571 , n19572 );
and ( n19574 , n19540 , n19573 );
xor ( n19575 , n19540 , n19573 );
xor ( n19576 , n19565 , n19567 );
xor ( n19577 , n19576 , n19570 );
and ( n19578 , n19434 , n19518 );
and ( n19579 , n19418 , n19516 );
nor ( n19580 , n19578 , n19579 );
xnor ( n19581 , n19580 , n19489 );
buf ( n19582 , n19581 );
and ( n19583 , n19469 , n19459 );
and ( n19584 , n19434 , n19457 );
nor ( n19585 , n19583 , n19584 );
xnor ( n19586 , n19585 , n19416 );
and ( n19587 , n19582 , n19586 );
buf ( n19588 , n19289 );
and ( n19589 , n19588 , n19419 );
and ( n19590 , n19586 , n19589 );
and ( n19591 , n19582 , n19589 );
or ( n19592 , n19587 , n19590 , n19591 );
xor ( n19593 , n19486 , n19541 );
xor ( n19594 , n19541 , n19542 );
not ( n19595 , n19594 );
and ( n19596 , n19593 , n19595 );
and ( n19597 , n19426 , n19596 );
not ( n19598 , n19597 );
xnor ( n19599 , n19598 , n19545 );
and ( n19600 , n19588 , n19424 );
and ( n19601 , n19510 , n19422 );
nor ( n19602 , n19600 , n19601 );
xnor ( n19603 , n19602 , n19431 );
and ( n19604 , n19599 , n19603 );
buf ( n19605 , n19290 );
and ( n19606 , n19605 , n19419 );
and ( n19607 , n19603 , n19606 );
and ( n19608 , n19599 , n19606 );
or ( n19609 , n19604 , n19607 , n19608 );
xor ( n19610 , n19546 , n19550 );
xor ( n19611 , n19610 , n19555 );
and ( n19612 , n19609 , n19611 );
xor ( n19613 , n19582 , n19586 );
xor ( n19614 , n19613 , n19589 );
and ( n19615 , n19611 , n19614 );
and ( n19616 , n19609 , n19614 );
or ( n19617 , n19612 , n19615 , n19616 );
and ( n19618 , n19592 , n19617 );
xor ( n19619 , n19558 , n19559 );
xor ( n19620 , n19619 , n19562 );
and ( n19621 , n19617 , n19620 );
and ( n19622 , n19592 , n19620 );
or ( n19623 , n19618 , n19621 , n19622 );
and ( n19624 , n19577 , n19623 );
xor ( n19625 , n19577 , n19623 );
xor ( n19626 , n19592 , n19617 );
xor ( n19627 , n19626 , n19620 );
and ( n19628 , n19469 , n19518 );
and ( n19629 , n19434 , n19516 );
nor ( n19630 , n19628 , n19629 );
xnor ( n19631 , n19630 , n19489 );
and ( n19632 , n19605 , n19424 );
and ( n19633 , n19588 , n19422 );
nor ( n19634 , n19632 , n19633 );
xnor ( n19635 , n19634 , n19431 );
and ( n19636 , n19631 , n19635 );
buf ( n19637 , n19291 );
and ( n19638 , n19637 , n19419 );
and ( n19639 , n19635 , n19638 );
and ( n19640 , n19631 , n19638 );
or ( n19641 , n19636 , n19639 , n19640 );
not ( n19642 , n19581 );
and ( n19643 , n19641 , n19642 );
and ( n19644 , n19496 , n19459 );
and ( n19645 , n19469 , n19457 );
nor ( n19646 , n19644 , n19645 );
xnor ( n19647 , n19646 , n19416 );
and ( n19648 , n19642 , n19647 );
and ( n19649 , n19641 , n19647 );
or ( n19650 , n19643 , n19648 , n19649 );
buf ( n19651 , n19356 );
buf ( n19652 , n19357 );
and ( n19653 , n19651 , n19652 );
not ( n19654 , n19653 );
and ( n19655 , n19542 , n19654 );
not ( n19656 , n19655 );
and ( n19657 , n19418 , n19596 );
and ( n19658 , n19426 , n19594 );
nor ( n19659 , n19657 , n19658 );
xnor ( n19660 , n19659 , n19545 );
and ( n19661 , n19656 , n19660 );
and ( n19662 , n19510 , n19459 );
and ( n19663 , n19496 , n19457 );
nor ( n19664 , n19662 , n19663 );
xnor ( n19665 , n19664 , n19416 );
and ( n19666 , n19660 , n19665 );
and ( n19667 , n19656 , n19665 );
or ( n19668 , n19661 , n19666 , n19667 );
xor ( n19669 , n19599 , n19603 );
xor ( n19670 , n19669 , n19606 );
and ( n19671 , n19668 , n19670 );
xor ( n19672 , n19641 , n19642 );
xor ( n19673 , n19672 , n19647 );
and ( n19674 , n19670 , n19673 );
and ( n19675 , n19668 , n19673 );
or ( n19676 , n19671 , n19674 , n19675 );
and ( n19677 , n19650 , n19676 );
xor ( n19678 , n19609 , n19611 );
xor ( n19679 , n19678 , n19614 );
and ( n19680 , n19676 , n19679 );
and ( n19681 , n19650 , n19679 );
or ( n19682 , n19677 , n19680 , n19681 );
and ( n19683 , n19627 , n19682 );
xor ( n19684 , n19627 , n19682 );
xor ( n19685 , n19542 , n19651 );
xor ( n19686 , n19651 , n19652 );
not ( n19687 , n19686 );
and ( n19688 , n19685 , n19687 );
and ( n19689 , n19426 , n19688 );
not ( n19690 , n19689 );
xnor ( n19691 , n19690 , n19655 );
and ( n19692 , n19588 , n19459 );
and ( n19693 , n19510 , n19457 );
nor ( n19694 , n19692 , n19693 );
xnor ( n19695 , n19694 , n19416 );
and ( n19696 , n19691 , n19695 );
and ( n19697 , n19637 , n19424 );
and ( n19698 , n19605 , n19422 );
nor ( n19699 , n19697 , n19698 );
xnor ( n19700 , n19699 , n19431 );
and ( n19701 , n19695 , n19700 );
and ( n19702 , n19691 , n19700 );
or ( n19703 , n19696 , n19701 , n19702 );
and ( n19704 , n19434 , n19596 );
and ( n19705 , n19418 , n19594 );
nor ( n19706 , n19704 , n19705 );
xnor ( n19707 , n19706 , n19545 );
buf ( n19708 , n19707 );
and ( n19709 , n19703 , n19708 );
xor ( n19710 , n19631 , n19635 );
xor ( n19711 , n19710 , n19638 );
and ( n19712 , n19708 , n19711 );
and ( n19713 , n19703 , n19711 );
or ( n19714 , n19709 , n19712 , n19713 );
not ( n19715 , n19707 );
and ( n19716 , n19496 , n19518 );
and ( n19717 , n19469 , n19516 );
nor ( n19718 , n19716 , n19717 );
xnor ( n19719 , n19718 , n19489 );
and ( n19720 , n19715 , n19719 );
buf ( n19721 , n19292 );
and ( n19722 , n19721 , n19419 );
and ( n19723 , n19719 , n19722 );
and ( n19724 , n19715 , n19722 );
or ( n19725 , n19720 , n19723 , n19724 );
xor ( n19726 , n19656 , n19660 );
xor ( n19727 , n19726 , n19665 );
and ( n19728 , n19725 , n19727 );
xor ( n19729 , n19703 , n19708 );
xor ( n19730 , n19729 , n19711 );
and ( n19731 , n19727 , n19730 );
and ( n19732 , n19725 , n19730 );
or ( n19733 , n19728 , n19731 , n19732 );
and ( n19734 , n19714 , n19733 );
xor ( n19735 , n19668 , n19670 );
xor ( n19736 , n19735 , n19673 );
and ( n19737 , n19733 , n19736 );
and ( n19738 , n19714 , n19736 );
or ( n19739 , n19734 , n19737 , n19738 );
xor ( n19740 , n19650 , n19676 );
xor ( n19741 , n19740 , n19679 );
and ( n19742 , n19739 , n19741 );
xor ( n19743 , n19739 , n19741 );
xor ( n19744 , n19714 , n19733 );
xor ( n19745 , n19744 , n19736 );
buf ( n19746 , n19358 );
buf ( n19747 , n19359 );
and ( n19748 , n19746 , n19747 );
not ( n19749 , n19748 );
and ( n19750 , n19652 , n19749 );
not ( n19751 , n19750 );
and ( n19752 , n19418 , n19688 );
and ( n19753 , n19426 , n19686 );
nor ( n19754 , n19752 , n19753 );
xnor ( n19755 , n19754 , n19655 );
and ( n19756 , n19751 , n19755 );
and ( n19757 , n19510 , n19518 );
and ( n19758 , n19496 , n19516 );
nor ( n19759 , n19757 , n19758 );
xnor ( n19760 , n19759 , n19489 );
and ( n19761 , n19755 , n19760 );
and ( n19762 , n19751 , n19760 );
or ( n19763 , n19756 , n19761 , n19762 );
and ( n19764 , n19469 , n19596 );
and ( n19765 , n19434 , n19594 );
nor ( n19766 , n19764 , n19765 );
xnor ( n19767 , n19766 , n19545 );
and ( n19768 , n19605 , n19459 );
and ( n19769 , n19588 , n19457 );
nor ( n19770 , n19768 , n19769 );
xnor ( n19771 , n19770 , n19416 );
and ( n19772 , n19767 , n19771 );
and ( n19773 , n19721 , n19424 );
and ( n19774 , n19637 , n19422 );
nor ( n19775 , n19773 , n19774 );
xnor ( n19776 , n19775 , n19431 );
and ( n19777 , n19771 , n19776 );
and ( n19778 , n19767 , n19776 );
or ( n19779 , n19772 , n19777 , n19778 );
and ( n19780 , n19763 , n19779 );
xor ( n19781 , n19691 , n19695 );
xor ( n19782 , n19781 , n19700 );
and ( n19783 , n19779 , n19782 );
and ( n19784 , n19763 , n19782 );
or ( n19785 , n19780 , n19783 , n19784 );
and ( n19786 , n19434 , n19688 );
and ( n19787 , n19418 , n19686 );
nor ( n19788 , n19786 , n19787 );
xnor ( n19789 , n19788 , n19655 );
and ( n19790 , n19588 , n19518 );
and ( n19791 , n19510 , n19516 );
nor ( n19792 , n19790 , n19791 );
xnor ( n19793 , n19792 , n19489 );
and ( n19794 , n19789 , n19793 );
and ( n19795 , n19637 , n19459 );
and ( n19796 , n19605 , n19457 );
nor ( n19797 , n19795 , n19796 );
xnor ( n19798 , n19797 , n19416 );
and ( n19799 , n19793 , n19798 );
and ( n19800 , n19789 , n19798 );
or ( n19801 , n19794 , n19799 , n19800 );
xor ( n19802 , n19652 , n19746 );
xor ( n19803 , n19746 , n19747 );
not ( n19804 , n19803 );
and ( n19805 , n19802 , n19804 );
and ( n19806 , n19426 , n19805 );
not ( n19807 , n19806 );
xnor ( n19808 , n19807 , n19750 );
buf ( n19809 , n19808 );
and ( n19810 , n19801 , n19809 );
buf ( n19811 , n19293 );
and ( n19812 , n19811 , n19419 );
and ( n19813 , n19809 , n19812 );
and ( n19814 , n19801 , n19812 );
or ( n19815 , n19810 , n19813 , n19814 );
and ( n19816 , n19496 , n19596 );
and ( n19817 , n19469 , n19594 );
nor ( n19818 , n19816 , n19817 );
xnor ( n19819 , n19818 , n19545 );
and ( n19820 , n19811 , n19424 );
and ( n19821 , n19721 , n19422 );
nor ( n19822 , n19820 , n19821 );
xnor ( n19823 , n19822 , n19431 );
and ( n19824 , n19819 , n19823 );
buf ( n19825 , n19294 );
and ( n19826 , n19825 , n19419 );
and ( n19827 , n19823 , n19826 );
and ( n19828 , n19819 , n19826 );
or ( n19829 , n19824 , n19827 , n19828 );
xor ( n19830 , n19751 , n19755 );
xor ( n19831 , n19830 , n19760 );
and ( n19832 , n19829 , n19831 );
xor ( n19833 , n19767 , n19771 );
xor ( n19834 , n19833 , n19776 );
and ( n19835 , n19831 , n19834 );
and ( n19836 , n19829 , n19834 );
or ( n19837 , n19832 , n19835 , n19836 );
and ( n19838 , n19815 , n19837 );
xor ( n19839 , n19715 , n19719 );
xor ( n19840 , n19839 , n19722 );
and ( n19841 , n19837 , n19840 );
and ( n19842 , n19815 , n19840 );
or ( n19843 , n19838 , n19841 , n19842 );
and ( n19844 , n19785 , n19843 );
xor ( n19845 , n19725 , n19727 );
xor ( n19846 , n19845 , n19730 );
and ( n19847 , n19843 , n19846 );
and ( n19848 , n19785 , n19846 );
or ( n19849 , n19844 , n19847 , n19848 );
and ( n19850 , n19745 , n19849 );
xor ( n19851 , n19745 , n19849 );
xor ( n19852 , n19785 , n19843 );
xor ( n19853 , n19852 , n19846 );
buf ( n19854 , n19360 );
buf ( n19855 , n19361 );
and ( n19856 , n19854 , n19855 );
not ( n19857 , n19856 );
and ( n19858 , n19747 , n19857 );
not ( n19859 , n19858 );
and ( n19860 , n19418 , n19805 );
and ( n19861 , n19426 , n19803 );
nor ( n19862 , n19860 , n19861 );
xnor ( n19863 , n19862 , n19750 );
and ( n19864 , n19859 , n19863 );
and ( n19865 , n19510 , n19596 );
and ( n19866 , n19496 , n19594 );
nor ( n19867 , n19865 , n19866 );
xnor ( n19868 , n19867 , n19545 );
and ( n19869 , n19863 , n19868 );
and ( n19870 , n19859 , n19868 );
or ( n19871 , n19864 , n19869 , n19870 );
and ( n19872 , n19469 , n19688 );
and ( n19873 , n19434 , n19686 );
nor ( n19874 , n19872 , n19873 );
xnor ( n19875 , n19874 , n19655 );
and ( n19876 , n19605 , n19518 );
and ( n19877 , n19588 , n19516 );
nor ( n19878 , n19876 , n19877 );
xnor ( n19879 , n19878 , n19489 );
and ( n19880 , n19875 , n19879 );
buf ( n19881 , n19295 );
and ( n19882 , n19881 , n19419 );
and ( n19883 , n19879 , n19882 );
and ( n19884 , n19875 , n19882 );
or ( n19885 , n19880 , n19883 , n19884 );
and ( n19886 , n19871 , n19885 );
not ( n19887 , n19808 );
and ( n19888 , n19885 , n19887 );
and ( n19889 , n19871 , n19887 );
or ( n19890 , n19886 , n19888 , n19889 );
xor ( n19891 , n19747 , n19854 );
xor ( n19892 , n19854 , n19855 );
not ( n19893 , n19892 );
and ( n19894 , n19891 , n19893 );
and ( n19895 , n19426 , n19894 );
not ( n19896 , n19895 );
xnor ( n19897 , n19896 , n19858 );
buf ( n19898 , n19897 );
and ( n19899 , n19721 , n19459 );
and ( n19900 , n19637 , n19457 );
nor ( n19901 , n19899 , n19900 );
xnor ( n19902 , n19901 , n19416 );
and ( n19903 , n19898 , n19902 );
and ( n19904 , n19825 , n19424 );
and ( n19905 , n19811 , n19422 );
nor ( n19906 , n19904 , n19905 );
xnor ( n19907 , n19906 , n19431 );
and ( n19908 , n19902 , n19907 );
and ( n19909 , n19898 , n19907 );
or ( n19910 , n19903 , n19908 , n19909 );
xor ( n19911 , n19789 , n19793 );
xor ( n19912 , n19911 , n19798 );
and ( n19913 , n19910 , n19912 );
xor ( n19914 , n19819 , n19823 );
xor ( n19915 , n19914 , n19826 );
and ( n19916 , n19912 , n19915 );
and ( n19917 , n19910 , n19915 );
or ( n19918 , n19913 , n19916 , n19917 );
and ( n19919 , n19890 , n19918 );
xor ( n19920 , n19801 , n19809 );
xor ( n19921 , n19920 , n19812 );
and ( n19922 , n19918 , n19921 );
and ( n19923 , n19890 , n19921 );
or ( n19924 , n19919 , n19922 , n19923 );
xor ( n19925 , n19763 , n19779 );
xor ( n19926 , n19925 , n19782 );
and ( n19927 , n19924 , n19926 );
xor ( n19928 , n19815 , n19837 );
xor ( n19929 , n19928 , n19840 );
and ( n19930 , n19926 , n19929 );
and ( n19931 , n19924 , n19929 );
or ( n19932 , n19927 , n19930 , n19931 );
and ( n19933 , n19853 , n19932 );
xor ( n19934 , n19853 , n19932 );
xor ( n19935 , n19924 , n19926 );
xor ( n19936 , n19935 , n19929 );
and ( n19937 , n19434 , n19805 );
and ( n19938 , n19418 , n19803 );
nor ( n19939 , n19937 , n19938 );
xnor ( n19940 , n19939 , n19750 );
and ( n19941 , n19588 , n19596 );
and ( n19942 , n19510 , n19594 );
nor ( n19943 , n19941 , n19942 );
xnor ( n19944 , n19943 , n19545 );
and ( n19945 , n19940 , n19944 );
buf ( n19946 , n19296 );
and ( n19947 , n19946 , n19419 );
and ( n19948 , n19944 , n19947 );
and ( n19949 , n19940 , n19947 );
or ( n19950 , n19945 , n19948 , n19949 );
and ( n19951 , n19496 , n19688 );
and ( n19952 , n19469 , n19686 );
nor ( n19953 , n19951 , n19952 );
xnor ( n19954 , n19953 , n19655 );
and ( n19955 , n19637 , n19518 );
and ( n19956 , n19605 , n19516 );
nor ( n19957 , n19955 , n19956 );
xnor ( n19958 , n19957 , n19489 );
and ( n19959 , n19954 , n19958 );
and ( n19960 , n19811 , n19459 );
and ( n19961 , n19721 , n19457 );
nor ( n19962 , n19960 , n19961 );
xnor ( n19963 , n19962 , n19416 );
and ( n19964 , n19958 , n19963 );
and ( n19965 , n19954 , n19963 );
or ( n19966 , n19959 , n19964 , n19965 );
and ( n19967 , n19950 , n19966 );
xor ( n19968 , n19859 , n19863 );
xor ( n19969 , n19968 , n19868 );
and ( n19970 , n19966 , n19969 );
and ( n19971 , n19950 , n19969 );
or ( n19972 , n19967 , n19970 , n19971 );
xor ( n19973 , n19871 , n19885 );
xor ( n19974 , n19973 , n19887 );
and ( n19975 , n19972 , n19974 );
xor ( n19976 , n19910 , n19912 );
xor ( n19977 , n19976 , n19915 );
and ( n19978 , n19974 , n19977 );
and ( n19979 , n19972 , n19977 );
or ( n19980 , n19975 , n19978 , n19979 );
xor ( n19981 , n19829 , n19831 );
xor ( n19982 , n19981 , n19834 );
and ( n19983 , n19980 , n19982 );
xor ( n19984 , n19890 , n19918 );
xor ( n19985 , n19984 , n19921 );
and ( n19986 , n19982 , n19985 );
and ( n19987 , n19980 , n19985 );
or ( n19988 , n19983 , n19986 , n19987 );
and ( n19989 , n19936 , n19988 );
xor ( n19990 , n19936 , n19988 );
xor ( n19991 , n19980 , n19982 );
xor ( n19992 , n19991 , n19985 );
buf ( n19993 , n19362 );
buf ( n19994 , n19363 );
and ( n19995 , n19993 , n19994 );
not ( n19996 , n19995 );
and ( n19997 , n19855 , n19996 );
not ( n19998 , n19997 );
and ( n19999 , n19418 , n19894 );
and ( n20000 , n19426 , n19892 );
nor ( n20001 , n19999 , n20000 );
xnor ( n20002 , n20001 , n19858 );
and ( n20003 , n19998 , n20002 );
buf ( n20004 , n19297 );
and ( n20005 , n20004 , n19419 );
and ( n20006 , n20002 , n20005 );
and ( n20007 , n19998 , n20005 );
or ( n20008 , n20003 , n20006 , n20007 );
not ( n20009 , n19897 );
and ( n20010 , n20008 , n20009 );
and ( n20011 , n19881 , n19424 );
and ( n20012 , n19825 , n19422 );
nor ( n20013 , n20011 , n20012 );
xnor ( n20014 , n20013 , n19431 );
and ( n20015 , n20009 , n20014 );
and ( n20016 , n20008 , n20014 );
or ( n20017 , n20010 , n20015 , n20016 );
xor ( n20018 , n19875 , n19879 );
xor ( n20019 , n20018 , n19882 );
and ( n20020 , n20017 , n20019 );
xor ( n20021 , n19898 , n19902 );
xor ( n20022 , n20021 , n19907 );
and ( n20023 , n20019 , n20022 );
and ( n20024 , n20017 , n20022 );
or ( n20025 , n20020 , n20023 , n20024 );
and ( n20026 , n19510 , n19688 );
and ( n20027 , n19496 , n19686 );
nor ( n20028 , n20026 , n20027 );
xnor ( n20029 , n20028 , n19655 );
and ( n20030 , n19605 , n19596 );
and ( n20031 , n19588 , n19594 );
nor ( n20032 , n20030 , n20031 );
xnor ( n20033 , n20032 , n19545 );
and ( n20034 , n20029 , n20033 );
and ( n20035 , n19946 , n19424 );
and ( n20036 , n19881 , n19422 );
nor ( n20037 , n20035 , n20036 );
xnor ( n20038 , n20037 , n19431 );
and ( n20039 , n20033 , n20038 );
and ( n20040 , n20029 , n20038 );
or ( n20041 , n20034 , n20039 , n20040 );
and ( n20042 , n19469 , n19805 );
and ( n20043 , n19434 , n19803 );
nor ( n20044 , n20042 , n20043 );
xnor ( n20045 , n20044 , n19750 );
and ( n20046 , n19721 , n19518 );
and ( n20047 , n19637 , n19516 );
nor ( n20048 , n20046 , n20047 );
xnor ( n20049 , n20048 , n19489 );
and ( n20050 , n20045 , n20049 );
and ( n20051 , n19825 , n19459 );
and ( n20052 , n19811 , n19457 );
nor ( n20053 , n20051 , n20052 );
xnor ( n20054 , n20053 , n19416 );
and ( n20055 , n20049 , n20054 );
and ( n20056 , n20045 , n20054 );
or ( n20057 , n20050 , n20055 , n20056 );
and ( n20058 , n20041 , n20057 );
xor ( n20059 , n19954 , n19958 );
xor ( n20060 , n20059 , n19963 );
and ( n20061 , n20057 , n20060 );
and ( n20062 , n20041 , n20060 );
or ( n20063 , n20058 , n20061 , n20062 );
and ( n20064 , n19434 , n19894 );
and ( n20065 , n19418 , n19892 );
nor ( n20066 , n20064 , n20065 );
xnor ( n20067 , n20066 , n19858 );
and ( n20068 , n19588 , n19688 );
and ( n20069 , n19510 , n19686 );
nor ( n20070 , n20068 , n20069 );
xnor ( n20071 , n20070 , n19655 );
and ( n20072 , n20067 , n20071 );
and ( n20073 , n20004 , n19424 );
and ( n20074 , n19946 , n19422 );
nor ( n20075 , n20073 , n20074 );
xnor ( n20076 , n20075 , n19431 );
and ( n20077 , n20071 , n20076 );
and ( n20078 , n20067 , n20076 );
or ( n20079 , n20072 , n20077 , n20078 );
buf ( n20080 , n19298 );
and ( n20081 , n20080 , n19419 );
buf ( n20082 , n20081 );
and ( n20083 , n20079 , n20082 );
xor ( n20084 , n19998 , n20002 );
xor ( n20085 , n20084 , n20005 );
and ( n20086 , n20082 , n20085 );
and ( n20087 , n20079 , n20085 );
or ( n20088 , n20083 , n20086 , n20087 );
xor ( n20089 , n19940 , n19944 );
xor ( n20090 , n20089 , n19947 );
and ( n20091 , n20088 , n20090 );
xor ( n20092 , n20008 , n20009 );
xor ( n20093 , n20092 , n20014 );
and ( n20094 , n20090 , n20093 );
and ( n20095 , n20088 , n20093 );
or ( n20096 , n20091 , n20094 , n20095 );
and ( n20097 , n20063 , n20096 );
xor ( n20098 , n19950 , n19966 );
xor ( n20099 , n20098 , n19969 );
and ( n20100 , n20096 , n20099 );
and ( n20101 , n20063 , n20099 );
or ( n20102 , n20097 , n20100 , n20101 );
and ( n20103 , n20025 , n20102 );
xor ( n20104 , n19972 , n19974 );
xor ( n20105 , n20104 , n19977 );
and ( n20106 , n20102 , n20105 );
and ( n20107 , n20025 , n20105 );
or ( n20108 , n20103 , n20106 , n20107 );
and ( n20109 , n19992 , n20108 );
xor ( n20110 , n19992 , n20108 );
xor ( n20111 , n19855 , n19993 );
xor ( n20112 , n19993 , n19994 );
not ( n20113 , n20112 );
and ( n20114 , n20111 , n20113 );
and ( n20115 , n19426 , n20114 );
not ( n20116 , n20115 );
xnor ( n20117 , n20116 , n19997 );
and ( n20118 , n19496 , n19805 );
and ( n20119 , n19469 , n19803 );
nor ( n20120 , n20118 , n20119 );
xnor ( n20121 , n20120 , n19750 );
and ( n20122 , n20117 , n20121 );
and ( n20123 , n19637 , n19596 );
and ( n20124 , n19605 , n19594 );
nor ( n20125 , n20123 , n20124 );
xnor ( n20126 , n20125 , n19545 );
and ( n20127 , n20121 , n20126 );
and ( n20128 , n20117 , n20126 );
or ( n20129 , n20122 , n20127 , n20128 );
and ( n20130 , n19811 , n19518 );
and ( n20131 , n19721 , n19516 );
nor ( n20132 , n20130 , n20131 );
xnor ( n20133 , n20132 , n19489 );
and ( n20134 , n19881 , n19459 );
and ( n20135 , n19825 , n19457 );
nor ( n20136 , n20134 , n20135 );
xnor ( n20137 , n20136 , n19416 );
and ( n20138 , n20133 , n20137 );
not ( n20139 , n20081 );
and ( n20140 , n20137 , n20139 );
and ( n20141 , n20133 , n20139 );
or ( n20142 , n20138 , n20140 , n20141 );
and ( n20143 , n20129 , n20142 );
xor ( n20144 , n20045 , n20049 );
xor ( n20145 , n20144 , n20054 );
and ( n20146 , n20142 , n20145 );
and ( n20147 , n20129 , n20145 );
or ( n20148 , n20143 , n20146 , n20147 );
xor ( n20149 , n20041 , n20057 );
xor ( n20150 , n20149 , n20060 );
and ( n20151 , n20148 , n20150 );
xor ( n20152 , n20088 , n20090 );
xor ( n20153 , n20152 , n20093 );
and ( n20154 , n20150 , n20153 );
and ( n20155 , n20148 , n20153 );
or ( n20156 , n20151 , n20154 , n20155 );
xor ( n20157 , n20017 , n20019 );
xor ( n20158 , n20157 , n20022 );
and ( n20159 , n20156 , n20158 );
xor ( n20160 , n20063 , n20096 );
xor ( n20161 , n20160 , n20099 );
and ( n20162 , n20158 , n20161 );
and ( n20163 , n20156 , n20161 );
or ( n20164 , n20159 , n20162 , n20163 );
xor ( n20165 , n20025 , n20102 );
xor ( n20166 , n20165 , n20105 );
and ( n20167 , n20164 , n20166 );
xor ( n20168 , n20164 , n20166 );
xor ( n20169 , n20156 , n20158 );
xor ( n20170 , n20169 , n20161 );
buf ( n20171 , n19364 );
buf ( n20172 , n19365 );
and ( n20173 , n20171 , n20172 );
not ( n20174 , n20173 );
and ( n20175 , n19994 , n20174 );
not ( n20176 , n20175 );
and ( n20177 , n20080 , n19424 );
and ( n20178 , n20004 , n19422 );
nor ( n20179 , n20177 , n20178 );
xnor ( n20180 , n20179 , n19431 );
and ( n20181 , n20176 , n20180 );
buf ( n20182 , n19299 );
and ( n20183 , n20182 , n19419 );
and ( n20184 , n20180 , n20183 );
and ( n20185 , n20176 , n20183 );
or ( n20186 , n20181 , n20184 , n20185 );
and ( n20187 , n19418 , n20114 );
and ( n20188 , n19426 , n20112 );
nor ( n20189 , n20187 , n20188 );
xnor ( n20190 , n20189 , n19997 );
and ( n20191 , n19510 , n19805 );
and ( n20192 , n19496 , n19803 );
nor ( n20193 , n20191 , n20192 );
xnor ( n20194 , n20193 , n19750 );
and ( n20195 , n20190 , n20194 );
and ( n20196 , n19946 , n19459 );
and ( n20197 , n19881 , n19457 );
nor ( n20198 , n20196 , n20197 );
xnor ( n20199 , n20198 , n19416 );
and ( n20200 , n20194 , n20199 );
and ( n20201 , n20190 , n20199 );
or ( n20202 , n20195 , n20200 , n20201 );
and ( n20203 , n20186 , n20202 );
and ( n20204 , n19469 , n19894 );
and ( n20205 , n19434 , n19892 );
nor ( n20206 , n20204 , n20205 );
xnor ( n20207 , n20206 , n19858 );
and ( n20208 , n19605 , n19688 );
and ( n20209 , n19588 , n19686 );
nor ( n20210 , n20208 , n20209 );
xnor ( n20211 , n20210 , n19655 );
and ( n20212 , n20207 , n20211 );
and ( n20213 , n19721 , n19596 );
and ( n20214 , n19637 , n19594 );
nor ( n20215 , n20213 , n20214 );
xnor ( n20216 , n20215 , n19545 );
and ( n20217 , n20211 , n20216 );
and ( n20218 , n20207 , n20216 );
or ( n20219 , n20212 , n20217 , n20218 );
and ( n20220 , n20202 , n20219 );
and ( n20221 , n20186 , n20219 );
or ( n20222 , n20203 , n20220 , n20221 );
xor ( n20223 , n20029 , n20033 );
xor ( n20224 , n20223 , n20038 );
and ( n20225 , n20222 , n20224 );
xor ( n20226 , n20079 , n20082 );
xor ( n20227 , n20226 , n20085 );
and ( n20228 , n20224 , n20227 );
and ( n20229 , n20222 , n20227 );
or ( n20230 , n20225 , n20228 , n20229 );
xor ( n20231 , n20067 , n20071 );
xor ( n20232 , n20231 , n20076 );
xor ( n20233 , n20117 , n20121 );
xor ( n20234 , n20233 , n20126 );
and ( n20235 , n20232 , n20234 );
xor ( n20236 , n20133 , n20137 );
xor ( n20237 , n20236 , n20139 );
and ( n20238 , n20234 , n20237 );
and ( n20239 , n20232 , n20237 );
or ( n20240 , n20235 , n20238 , n20239 );
xor ( n20241 , n20129 , n20142 );
xor ( n20242 , n20241 , n20145 );
and ( n20243 , n20240 , n20242 );
xor ( n20244 , n20222 , n20224 );
xor ( n20245 , n20244 , n20227 );
and ( n20246 , n20242 , n20245 );
and ( n20247 , n20240 , n20245 );
or ( n20248 , n20243 , n20246 , n20247 );
and ( n20249 , n20230 , n20248 );
xor ( n20250 , n20148 , n20150 );
xor ( n20251 , n20250 , n20153 );
and ( n20252 , n20248 , n20251 );
and ( n20253 , n20230 , n20251 );
or ( n20254 , n20249 , n20252 , n20253 );
and ( n20255 , n20170 , n20254 );
xor ( n20256 , n20170 , n20254 );
xor ( n20257 , n20230 , n20248 );
xor ( n20258 , n20257 , n20251 );
and ( n20259 , n19434 , n20114 );
and ( n20260 , n19418 , n20112 );
nor ( n20261 , n20259 , n20260 );
xnor ( n20262 , n20261 , n19997 );
and ( n20263 , n20004 , n19459 );
and ( n20264 , n19946 , n19457 );
nor ( n20265 , n20263 , n20264 );
xnor ( n20266 , n20265 , n19416 );
and ( n20267 , n20262 , n20266 );
buf ( n20268 , n19300 );
and ( n20269 , n20268 , n19419 );
and ( n20270 , n20266 , n20269 );
and ( n20271 , n20262 , n20269 );
or ( n20272 , n20267 , n20270 , n20271 );
xor ( n20273 , n19994 , n20171 );
xor ( n20274 , n20171 , n20172 );
not ( n20275 , n20274 );
and ( n20276 , n20273 , n20275 );
and ( n20277 , n19426 , n20276 );
not ( n20278 , n20277 );
xnor ( n20279 , n20278 , n20175 );
and ( n20280 , n19588 , n19805 );
and ( n20281 , n19510 , n19803 );
nor ( n20282 , n20280 , n20281 );
xnor ( n20283 , n20282 , n19750 );
and ( n20284 , n20279 , n20283 );
and ( n20285 , n19637 , n19688 );
and ( n20286 , n19605 , n19686 );
nor ( n20287 , n20285 , n20286 );
xnor ( n20288 , n20287 , n19655 );
and ( n20289 , n20283 , n20288 );
and ( n20290 , n20279 , n20288 );
or ( n20291 , n20284 , n20289 , n20290 );
and ( n20292 , n20272 , n20291 );
and ( n20293 , n19496 , n19894 );
and ( n20294 , n19469 , n19892 );
nor ( n20295 , n20293 , n20294 );
xnor ( n20296 , n20295 , n19858 );
and ( n20297 , n19811 , n19596 );
and ( n20298 , n19721 , n19594 );
nor ( n20299 , n20297 , n20298 );
xnor ( n20300 , n20299 , n19545 );
and ( n20301 , n20296 , n20300 );
and ( n20302 , n19881 , n19518 );
and ( n20303 , n19825 , n19516 );
nor ( n20304 , n20302 , n20303 );
xnor ( n20305 , n20304 , n19489 );
and ( n20306 , n20300 , n20305 );
and ( n20307 , n20296 , n20305 );
or ( n20308 , n20301 , n20306 , n20307 );
and ( n20309 , n20291 , n20308 );
and ( n20310 , n20272 , n20308 );
or ( n20311 , n20292 , n20309 , n20310 );
and ( n20312 , n20182 , n19424 );
and ( n20313 , n20080 , n19422 );
nor ( n20314 , n20312 , n20313 );
xnor ( n20315 , n20314 , n19431 );
buf ( n20316 , n20315 );
and ( n20317 , n19825 , n19518 );
and ( n20318 , n19811 , n19516 );
nor ( n20319 , n20317 , n20318 );
xnor ( n20320 , n20319 , n19489 );
and ( n20321 , n20316 , n20320 );
xor ( n20322 , n20176 , n20180 );
xor ( n20323 , n20322 , n20183 );
and ( n20324 , n20320 , n20323 );
and ( n20325 , n20316 , n20323 );
or ( n20326 , n20321 , n20324 , n20325 );
and ( n20327 , n20311 , n20326 );
xor ( n20328 , n20186 , n20202 );
xor ( n20329 , n20328 , n20219 );
and ( n20330 , n20326 , n20329 );
and ( n20331 , n20311 , n20329 );
or ( n20332 , n20327 , n20330 , n20331 );
buf ( n20333 , n19366 );
buf ( n20334 , n19367 );
and ( n20335 , n20333 , n20334 );
not ( n20336 , n20335 );
and ( n20337 , n20172 , n20336 );
not ( n20338 , n20337 );
and ( n20339 , n20080 , n19459 );
and ( n20340 , n20004 , n19457 );
nor ( n20341 , n20339 , n20340 );
xnor ( n20342 , n20341 , n19416 );
and ( n20343 , n20338 , n20342 );
and ( n20344 , n20268 , n19424 );
and ( n20345 , n20182 , n19422 );
nor ( n20346 , n20344 , n20345 );
xnor ( n20347 , n20346 , n19431 );
and ( n20348 , n20342 , n20347 );
and ( n20349 , n20338 , n20347 );
or ( n20350 , n20343 , n20348 , n20349 );
and ( n20351 , n19418 , n20276 );
and ( n20352 , n19426 , n20274 );
nor ( n20353 , n20351 , n20352 );
xnor ( n20354 , n20353 , n20175 );
and ( n20355 , n19946 , n19518 );
and ( n20356 , n19881 , n19516 );
nor ( n20357 , n20355 , n20356 );
xnor ( n20358 , n20357 , n19489 );
and ( n20359 , n20354 , n20358 );
buf ( n20360 , n19301 );
and ( n20361 , n20360 , n19419 );
and ( n20362 , n20358 , n20361 );
and ( n20363 , n20354 , n20361 );
or ( n20364 , n20359 , n20362 , n20363 );
and ( n20365 , n20350 , n20364 );
not ( n20366 , n20315 );
and ( n20367 , n20364 , n20366 );
and ( n20368 , n20350 , n20366 );
or ( n20369 , n20365 , n20367 , n20368 );
xor ( n20370 , n20190 , n20194 );
xor ( n20371 , n20370 , n20199 );
and ( n20372 , n20369 , n20371 );
xor ( n20373 , n20207 , n20211 );
xor ( n20374 , n20373 , n20216 );
and ( n20375 , n20371 , n20374 );
and ( n20376 , n20369 , n20374 );
or ( n20377 , n20372 , n20375 , n20376 );
and ( n20378 , n19469 , n20114 );
and ( n20379 , n19434 , n20112 );
nor ( n20380 , n20378 , n20379 );
xnor ( n20381 , n20380 , n19997 );
and ( n20382 , n19510 , n19894 );
and ( n20383 , n19496 , n19892 );
nor ( n20384 , n20382 , n20383 );
xnor ( n20385 , n20384 , n19858 );
and ( n20386 , n20381 , n20385 );
and ( n20387 , n19605 , n19805 );
and ( n20388 , n19588 , n19803 );
nor ( n20389 , n20387 , n20388 );
xnor ( n20390 , n20389 , n19750 );
and ( n20391 , n20385 , n20390 );
and ( n20392 , n20381 , n20390 );
or ( n20393 , n20386 , n20391 , n20392 );
xor ( n20394 , n20262 , n20266 );
xor ( n20395 , n20394 , n20269 );
and ( n20396 , n20393 , n20395 );
xor ( n20397 , n20279 , n20283 );
xor ( n20398 , n20397 , n20288 );
and ( n20399 , n20395 , n20398 );
and ( n20400 , n20393 , n20398 );
or ( n20401 , n20396 , n20399 , n20400 );
xor ( n20402 , n20272 , n20291 );
xor ( n20403 , n20402 , n20308 );
and ( n20404 , n20401 , n20403 );
xor ( n20405 , n20316 , n20320 );
xor ( n20406 , n20405 , n20323 );
and ( n20407 , n20403 , n20406 );
and ( n20408 , n20401 , n20406 );
or ( n20409 , n20404 , n20407 , n20408 );
and ( n20410 , n20377 , n20409 );
xor ( n20411 , n20232 , n20234 );
xor ( n20412 , n20411 , n20237 );
and ( n20413 , n20409 , n20412 );
and ( n20414 , n20377 , n20412 );
or ( n20415 , n20410 , n20413 , n20414 );
and ( n20416 , n20332 , n20415 );
xor ( n20417 , n20240 , n20242 );
xor ( n20418 , n20417 , n20245 );
and ( n20419 , n20415 , n20418 );
and ( n20420 , n20332 , n20418 );
or ( n20421 , n20416 , n20419 , n20420 );
and ( n20422 , n20258 , n20421 );
xor ( n20423 , n20258 , n20421 );
xor ( n20424 , n20332 , n20415 );
xor ( n20425 , n20424 , n20418 );
and ( n20426 , n20360 , n19424 );
and ( n20427 , n20268 , n19422 );
nor ( n20428 , n20426 , n20427 );
xnor ( n20429 , n20428 , n19431 );
buf ( n20430 , n20429 );
and ( n20431 , n19721 , n19688 );
and ( n20432 , n19637 , n19686 );
nor ( n20433 , n20431 , n20432 );
xnor ( n20434 , n20433 , n19655 );
and ( n20435 , n20430 , n20434 );
and ( n20436 , n19825 , n19596 );
and ( n20437 , n19811 , n19594 );
nor ( n20438 , n20436 , n20437 );
xnor ( n20439 , n20438 , n19545 );
and ( n20440 , n20434 , n20439 );
and ( n20441 , n20430 , n20439 );
or ( n20442 , n20435 , n20440 , n20441 );
and ( n20443 , n19434 , n20276 );
and ( n20444 , n19418 , n20274 );
nor ( n20445 , n20443 , n20444 );
xnor ( n20446 , n20445 , n20175 );
and ( n20447 , n20182 , n19459 );
and ( n20448 , n20080 , n19457 );
nor ( n20449 , n20447 , n20448 );
xnor ( n20450 , n20449 , n19416 );
and ( n20451 , n20446 , n20450 );
buf ( n20452 , n19302 );
and ( n20453 , n20452 , n19419 );
and ( n20454 , n20450 , n20453 );
and ( n20455 , n20446 , n20453 );
or ( n20456 , n20451 , n20454 , n20455 );
xor ( n20457 , n20172 , n20333 );
xor ( n20458 , n20333 , n20334 );
not ( n20459 , n20458 );
and ( n20460 , n20457 , n20459 );
and ( n20461 , n19426 , n20460 );
not ( n20462 , n20461 );
xnor ( n20463 , n20462 , n20337 );
and ( n20464 , n19496 , n20114 );
and ( n20465 , n19469 , n20112 );
nor ( n20466 , n20464 , n20465 );
xnor ( n20467 , n20466 , n19997 );
and ( n20468 , n20463 , n20467 );
and ( n20469 , n19811 , n19688 );
and ( n20470 , n19721 , n19686 );
nor ( n20471 , n20469 , n20470 );
xnor ( n20472 , n20471 , n19655 );
and ( n20473 , n20467 , n20472 );
and ( n20474 , n20463 , n20472 );
or ( n20475 , n20468 , n20473 , n20474 );
and ( n20476 , n20456 , n20475 );
xor ( n20477 , n20338 , n20342 );
xor ( n20478 , n20477 , n20347 );
and ( n20479 , n20475 , n20478 );
and ( n20480 , n20456 , n20478 );
or ( n20481 , n20476 , n20479 , n20480 );
and ( n20482 , n20442 , n20481 );
xor ( n20483 , n20296 , n20300 );
xor ( n20484 , n20483 , n20305 );
and ( n20485 , n20481 , n20484 );
and ( n20486 , n20442 , n20484 );
or ( n20487 , n20482 , n20485 , n20486 );
and ( n20488 , n19588 , n19894 );
and ( n20489 , n19510 , n19892 );
nor ( n20490 , n20488 , n20489 );
xnor ( n20491 , n20490 , n19858 );
and ( n20492 , n19637 , n19805 );
and ( n20493 , n19605 , n19803 );
nor ( n20494 , n20492 , n20493 );
xnor ( n20495 , n20494 , n19750 );
and ( n20496 , n20491 , n20495 );
and ( n20497 , n20004 , n19518 );
and ( n20498 , n19946 , n19516 );
nor ( n20499 , n20497 , n20498 );
xnor ( n20500 , n20499 , n19489 );
and ( n20501 , n20495 , n20500 );
and ( n20502 , n20491 , n20500 );
or ( n20503 , n20496 , n20501 , n20502 );
xor ( n20504 , n20354 , n20358 );
xor ( n20505 , n20504 , n20361 );
and ( n20506 , n20503 , n20505 );
xor ( n20507 , n20381 , n20385 );
xor ( n20508 , n20507 , n20390 );
and ( n20509 , n20505 , n20508 );
and ( n20510 , n20503 , n20508 );
or ( n20511 , n20506 , n20509 , n20510 );
xor ( n20512 , n20350 , n20364 );
xor ( n20513 , n20512 , n20366 );
and ( n20514 , n20511 , n20513 );
xor ( n20515 , n20393 , n20395 );
xor ( n20516 , n20515 , n20398 );
and ( n20517 , n20513 , n20516 );
and ( n20518 , n20511 , n20516 );
or ( n20519 , n20514 , n20517 , n20518 );
and ( n20520 , n20487 , n20519 );
xor ( n20521 , n20369 , n20371 );
xor ( n20522 , n20521 , n20374 );
and ( n20523 , n20519 , n20522 );
and ( n20524 , n20487 , n20522 );
or ( n20525 , n20520 , n20523 , n20524 );
xor ( n20526 , n20311 , n20326 );
xor ( n20527 , n20526 , n20329 );
and ( n20528 , n20525 , n20527 );
xor ( n20529 , n20377 , n20409 );
xor ( n20530 , n20529 , n20412 );
and ( n20531 , n20527 , n20530 );
and ( n20532 , n20525 , n20530 );
or ( n20533 , n20528 , n20531 , n20532 );
and ( n20534 , n20425 , n20533 );
xor ( n20535 , n20425 , n20533 );
xor ( n20536 , n20525 , n20527 );
xor ( n20537 , n20536 , n20530 );
buf ( n20538 , n19368 );
buf ( n20539 , n19369 );
and ( n20540 , n20538 , n20539 );
not ( n20541 , n20540 );
and ( n20542 , n20334 , n20541 );
not ( n20543 , n20542 );
and ( n20544 , n20080 , n19518 );
and ( n20545 , n20004 , n19516 );
nor ( n20546 , n20544 , n20545 );
xnor ( n20547 , n20546 , n19489 );
and ( n20548 , n20543 , n20547 );
and ( n20549 , n20268 , n19459 );
and ( n20550 , n20182 , n19457 );
nor ( n20551 , n20549 , n20550 );
xnor ( n20552 , n20551 , n19416 );
and ( n20553 , n20547 , n20552 );
and ( n20554 , n20543 , n20552 );
or ( n20555 , n20548 , n20553 , n20554 );
and ( n20556 , n19881 , n19596 );
and ( n20557 , n19825 , n19594 );
nor ( n20558 , n20556 , n20557 );
xnor ( n20559 , n20558 , n19545 );
and ( n20560 , n20555 , n20559 );
not ( n20561 , n20429 );
and ( n20562 , n20559 , n20561 );
and ( n20563 , n20555 , n20561 );
or ( n20564 , n20560 , n20562 , n20563 );
and ( n20565 , n19469 , n20276 );
and ( n20566 , n19434 , n20274 );
nor ( n20567 , n20565 , n20566 );
xnor ( n20568 , n20567 , n20175 );
and ( n20569 , n19721 , n19805 );
and ( n20570 , n19637 , n19803 );
nor ( n20571 , n20569 , n20570 );
xnor ( n20572 , n20571 , n19750 );
and ( n20573 , n20568 , n20572 );
and ( n20574 , n19825 , n19688 );
and ( n20575 , n19811 , n19686 );
nor ( n20576 , n20574 , n20575 );
xnor ( n20577 , n20576 , n19655 );
and ( n20578 , n20572 , n20577 );
and ( n20579 , n20568 , n20577 );
or ( n20580 , n20573 , n20578 , n20579 );
and ( n20581 , n19510 , n20114 );
and ( n20582 , n19496 , n20112 );
nor ( n20583 , n20581 , n20582 );
xnor ( n20584 , n20583 , n19997 );
and ( n20585 , n19605 , n19894 );
and ( n20586 , n19588 , n19892 );
nor ( n20587 , n20585 , n20586 );
xnor ( n20588 , n20587 , n19858 );
and ( n20589 , n20584 , n20588 );
and ( n20590 , n19946 , n19596 );
and ( n20591 , n19881 , n19594 );
nor ( n20592 , n20590 , n20591 );
xnor ( n20593 , n20592 , n19545 );
and ( n20594 , n20588 , n20593 );
and ( n20595 , n20584 , n20593 );
or ( n20596 , n20589 , n20594 , n20595 );
and ( n20597 , n20580 , n20596 );
xor ( n20598 , n20446 , n20450 );
xor ( n20599 , n20598 , n20453 );
and ( n20600 , n20596 , n20599 );
and ( n20601 , n20580 , n20599 );
or ( n20602 , n20597 , n20600 , n20601 );
and ( n20603 , n20564 , n20602 );
xor ( n20604 , n20430 , n20434 );
xor ( n20605 , n20604 , n20439 );
and ( n20606 , n20602 , n20605 );
and ( n20607 , n20564 , n20605 );
or ( n20608 , n20603 , n20606 , n20607 );
and ( n20609 , n19418 , n20460 );
and ( n20610 , n19426 , n20458 );
nor ( n20611 , n20609 , n20610 );
xnor ( n20612 , n20611 , n20337 );
and ( n20613 , n20452 , n19424 );
and ( n20614 , n20360 , n19422 );
nor ( n20615 , n20613 , n20614 );
xnor ( n20616 , n20615 , n19431 );
and ( n20617 , n20612 , n20616 );
buf ( n20618 , n19303 );
and ( n20619 , n20618 , n19419 );
and ( n20620 , n20616 , n20619 );
and ( n20621 , n20612 , n20619 );
or ( n20622 , n20617 , n20620 , n20621 );
xor ( n20623 , n20491 , n20495 );
xor ( n20624 , n20623 , n20500 );
and ( n20625 , n20622 , n20624 );
xor ( n20626 , n20463 , n20467 );
xor ( n20627 , n20626 , n20472 );
and ( n20628 , n20624 , n20627 );
and ( n20629 , n20622 , n20627 );
or ( n20630 , n20625 , n20628 , n20629 );
xor ( n20631 , n20456 , n20475 );
xor ( n20632 , n20631 , n20478 );
and ( n20633 , n20630 , n20632 );
xor ( n20634 , n20503 , n20505 );
xor ( n20635 , n20634 , n20508 );
and ( n20636 , n20632 , n20635 );
and ( n20637 , n20630 , n20635 );
or ( n20638 , n20633 , n20636 , n20637 );
and ( n20639 , n20608 , n20638 );
xor ( n20640 , n20442 , n20481 );
xor ( n20641 , n20640 , n20484 );
and ( n20642 , n20638 , n20641 );
and ( n20643 , n20608 , n20641 );
or ( n20644 , n20639 , n20642 , n20643 );
xor ( n20645 , n20401 , n20403 );
xor ( n20646 , n20645 , n20406 );
and ( n20647 , n20644 , n20646 );
xor ( n20648 , n20487 , n20519 );
xor ( n20649 , n20648 , n20522 );
and ( n20650 , n20646 , n20649 );
and ( n20651 , n20644 , n20649 );
or ( n20652 , n20647 , n20650 , n20651 );
and ( n20653 , n20537 , n20652 );
xor ( n20654 , n20537 , n20652 );
xor ( n20655 , n20644 , n20646 );
xor ( n20656 , n20655 , n20649 );
and ( n20657 , n20182 , n19518 );
and ( n20658 , n20080 , n19516 );
nor ( n20659 , n20657 , n20658 );
xnor ( n20660 , n20659 , n19489 );
and ( n20661 , n20618 , n19424 );
and ( n20662 , n20452 , n19422 );
nor ( n20663 , n20661 , n20662 );
xnor ( n20664 , n20663 , n19431 );
and ( n20665 , n20660 , n20664 );
buf ( n20666 , n19304 );
and ( n20667 , n20666 , n19419 );
and ( n20668 , n20664 , n20667 );
and ( n20669 , n20660 , n20667 );
or ( n20670 , n20665 , n20668 , n20669 );
xor ( n20671 , n20334 , n20538 );
xor ( n20672 , n20538 , n20539 );
not ( n20673 , n20672 );
and ( n20674 , n20671 , n20673 );
and ( n20675 , n19426 , n20674 );
not ( n20676 , n20675 );
xnor ( n20677 , n20676 , n20542 );
and ( n20678 , n19637 , n19894 );
and ( n20679 , n19605 , n19892 );
nor ( n20680 , n20678 , n20679 );
xnor ( n20681 , n20680 , n19858 );
and ( n20682 , n20677 , n20681 );
and ( n20683 , n19811 , n19805 );
and ( n20684 , n19721 , n19803 );
nor ( n20685 , n20683 , n20684 );
xnor ( n20686 , n20685 , n19750 );
and ( n20687 , n20681 , n20686 );
and ( n20688 , n20677 , n20686 );
or ( n20689 , n20682 , n20687 , n20688 );
and ( n20690 , n20670 , n20689 );
and ( n20691 , n20360 , n19459 );
and ( n20692 , n20268 , n19457 );
nor ( n20693 , n20691 , n20692 );
xnor ( n20694 , n20693 , n19416 );
buf ( n20695 , n20694 );
and ( n20696 , n20689 , n20695 );
and ( n20697 , n20670 , n20695 );
or ( n20698 , n20690 , n20696 , n20697 );
and ( n20699 , n19434 , n20460 );
and ( n20700 , n19418 , n20458 );
nor ( n20701 , n20699 , n20700 );
xnor ( n20702 , n20701 , n20337 );
and ( n20703 , n19588 , n20114 );
and ( n20704 , n19510 , n20112 );
nor ( n20705 , n20703 , n20704 );
xnor ( n20706 , n20705 , n19997 );
and ( n20707 , n20702 , n20706 );
and ( n20708 , n20004 , n19596 );
and ( n20709 , n19946 , n19594 );
nor ( n20710 , n20708 , n20709 );
xnor ( n20711 , n20710 , n19545 );
and ( n20712 , n20706 , n20711 );
and ( n20713 , n20702 , n20711 );
or ( n20714 , n20707 , n20712 , n20713 );
xor ( n20715 , n20543 , n20547 );
xor ( n20716 , n20715 , n20552 );
and ( n20717 , n20714 , n20716 );
xor ( n20718 , n20612 , n20616 );
xor ( n20719 , n20718 , n20619 );
and ( n20720 , n20716 , n20719 );
and ( n20721 , n20714 , n20719 );
or ( n20722 , n20717 , n20720 , n20721 );
and ( n20723 , n20698 , n20722 );
xor ( n20724 , n20555 , n20559 );
xor ( n20725 , n20724 , n20561 );
and ( n20726 , n20722 , n20725 );
and ( n20727 , n20698 , n20725 );
or ( n20728 , n20723 , n20726 , n20727 );
and ( n20729 , n19496 , n20276 );
and ( n20730 , n19469 , n20274 );
nor ( n20731 , n20729 , n20730 );
xnor ( n20732 , n20731 , n20175 );
and ( n20733 , n19881 , n19688 );
and ( n20734 , n19825 , n19686 );
nor ( n20735 , n20733 , n20734 );
xnor ( n20736 , n20735 , n19655 );
and ( n20737 , n20732 , n20736 );
not ( n20738 , n20694 );
and ( n20739 , n20736 , n20738 );
and ( n20740 , n20732 , n20738 );
or ( n20741 , n20737 , n20739 , n20740 );
xor ( n20742 , n20568 , n20572 );
xor ( n20743 , n20742 , n20577 );
and ( n20744 , n20741 , n20743 );
xor ( n20745 , n20584 , n20588 );
xor ( n20746 , n20745 , n20593 );
and ( n20747 , n20743 , n20746 );
and ( n20748 , n20741 , n20746 );
or ( n20749 , n20744 , n20747 , n20748 );
xor ( n20750 , n20580 , n20596 );
xor ( n20751 , n20750 , n20599 );
and ( n20752 , n20749 , n20751 );
xor ( n20753 , n20622 , n20624 );
xor ( n20754 , n20753 , n20627 );
and ( n20755 , n20751 , n20754 );
and ( n20756 , n20749 , n20754 );
or ( n20757 , n20752 , n20755 , n20756 );
and ( n20758 , n20728 , n20757 );
xor ( n20759 , n20564 , n20602 );
xor ( n20760 , n20759 , n20605 );
and ( n20761 , n20757 , n20760 );
and ( n20762 , n20728 , n20760 );
or ( n20763 , n20758 , n20761 , n20762 );
xor ( n20764 , n20511 , n20513 );
xor ( n20765 , n20764 , n20516 );
and ( n20766 , n20763 , n20765 );
xor ( n20767 , n20608 , n20638 );
xor ( n20768 , n20767 , n20641 );
and ( n20769 , n20765 , n20768 );
and ( n20770 , n20763 , n20768 );
or ( n20771 , n20766 , n20769 , n20770 );
and ( n20772 , n20656 , n20771 );
xor ( n20773 , n20656 , n20771 );
xor ( n20774 , n20763 , n20765 );
xor ( n20775 , n20774 , n20768 );
buf ( n20776 , n19370 );
buf ( n20777 , n19371 );
and ( n20778 , n20776 , n20777 );
not ( n20779 , n20778 );
and ( n20780 , n20539 , n20779 );
not ( n20781 , n20780 );
and ( n20782 , n20080 , n19596 );
and ( n20783 , n20004 , n19594 );
nor ( n20784 , n20782 , n20783 );
xnor ( n20785 , n20784 , n19545 );
and ( n20786 , n20781 , n20785 );
and ( n20787 , n20268 , n19518 );
and ( n20788 , n20182 , n19516 );
nor ( n20789 , n20787 , n20788 );
xnor ( n20790 , n20789 , n19489 );
and ( n20791 , n20785 , n20790 );
and ( n20792 , n20781 , n20790 );
or ( n20793 , n20786 , n20791 , n20792 );
and ( n20794 , n20452 , n19459 );
and ( n20795 , n20360 , n19457 );
nor ( n20796 , n20794 , n20795 );
xnor ( n20797 , n20796 , n19416 );
and ( n20798 , n20666 , n19424 );
and ( n20799 , n20618 , n19422 );
nor ( n20800 , n20798 , n20799 );
xnor ( n20801 , n20800 , n19431 );
and ( n20802 , n20797 , n20801 );
buf ( n20803 , n19305 );
and ( n20804 , n20803 , n19419 );
and ( n20805 , n20801 , n20804 );
and ( n20806 , n20797 , n20804 );
or ( n20807 , n20802 , n20805 , n20806 );
and ( n20808 , n20793 , n20807 );
xor ( n20809 , n20660 , n20664 );
xor ( n20810 , n20809 , n20667 );
and ( n20811 , n20807 , n20810 );
and ( n20812 , n20793 , n20810 );
or ( n20813 , n20808 , n20811 , n20812 );
and ( n20814 , n19418 , n20674 );
and ( n20815 , n19426 , n20672 );
nor ( n20816 , n20814 , n20815 );
xnor ( n20817 , n20816 , n20542 );
and ( n20818 , n19510 , n20276 );
and ( n20819 , n19496 , n20274 );
nor ( n20820 , n20818 , n20819 );
xnor ( n20821 , n20820 , n20175 );
and ( n20822 , n20817 , n20821 );
and ( n20823 , n19946 , n19688 );
and ( n20824 , n19881 , n19686 );
nor ( n20825 , n20823 , n20824 );
xnor ( n20826 , n20825 , n19655 );
and ( n20827 , n20821 , n20826 );
and ( n20828 , n20817 , n20826 );
or ( n20829 , n20822 , n20827 , n20828 );
and ( n20830 , n19469 , n20460 );
and ( n20831 , n19434 , n20458 );
nor ( n20832 , n20830 , n20831 );
xnor ( n20833 , n20832 , n20337 );
and ( n20834 , n19605 , n20114 );
and ( n20835 , n19588 , n20112 );
nor ( n20836 , n20834 , n20835 );
xnor ( n20837 , n20836 , n19997 );
and ( n20838 , n20833 , n20837 );
and ( n20839 , n19721 , n19894 );
and ( n20840 , n19637 , n19892 );
nor ( n20841 , n20839 , n20840 );
xnor ( n20842 , n20841 , n19858 );
and ( n20843 , n20837 , n20842 );
and ( n20844 , n20833 , n20842 );
or ( n20845 , n20838 , n20843 , n20844 );
and ( n20846 , n20829 , n20845 );
xor ( n20847 , n20677 , n20681 );
xor ( n20848 , n20847 , n20686 );
and ( n20849 , n20845 , n20848 );
and ( n20850 , n20829 , n20848 );
or ( n20851 , n20846 , n20849 , n20850 );
and ( n20852 , n20813 , n20851 );
xor ( n20853 , n20670 , n20689 );
xor ( n20854 , n20853 , n20695 );
and ( n20855 , n20851 , n20854 );
and ( n20856 , n20813 , n20854 );
or ( n20857 , n20852 , n20855 , n20856 );
and ( n20858 , n20182 , n19596 );
and ( n20859 , n20080 , n19594 );
nor ( n20860 , n20858 , n20859 );
xnor ( n20861 , n20860 , n19545 );
and ( n20862 , n20618 , n19459 );
and ( n20863 , n20452 , n19457 );
nor ( n20864 , n20862 , n20863 );
xnor ( n20865 , n20864 , n19416 );
and ( n20866 , n20861 , n20865 );
buf ( n20867 , n19306 );
and ( n20868 , n20867 , n19419 );
and ( n20869 , n20865 , n20868 );
and ( n20870 , n20861 , n20868 );
or ( n20871 , n20866 , n20869 , n20870 );
and ( n20872 , n20360 , n19518 );
and ( n20873 , n20268 , n19516 );
nor ( n20874 , n20872 , n20873 );
xnor ( n20875 , n20874 , n19489 );
buf ( n20876 , n20875 );
and ( n20877 , n20871 , n20876 );
and ( n20878 , n19825 , n19805 );
and ( n20879 , n19811 , n19803 );
nor ( n20880 , n20878 , n20879 );
xnor ( n20881 , n20880 , n19750 );
and ( n20882 , n20876 , n20881 );
and ( n20883 , n20871 , n20881 );
or ( n20884 , n20877 , n20882 , n20883 );
xor ( n20885 , n20702 , n20706 );
xor ( n20886 , n20885 , n20711 );
and ( n20887 , n20884 , n20886 );
xor ( n20888 , n20732 , n20736 );
xor ( n20889 , n20888 , n20738 );
and ( n20890 , n20886 , n20889 );
and ( n20891 , n20884 , n20889 );
or ( n20892 , n20887 , n20890 , n20891 );
xor ( n20893 , n20714 , n20716 );
xor ( n20894 , n20893 , n20719 );
and ( n20895 , n20892 , n20894 );
xor ( n20896 , n20741 , n20743 );
xor ( n20897 , n20896 , n20746 );
and ( n20898 , n20894 , n20897 );
and ( n20899 , n20892 , n20897 );
or ( n20900 , n20895 , n20898 , n20899 );
and ( n20901 , n20857 , n20900 );
xor ( n20902 , n20698 , n20722 );
xor ( n20903 , n20902 , n20725 );
and ( n20904 , n20900 , n20903 );
and ( n20905 , n20857 , n20903 );
or ( n20906 , n20901 , n20904 , n20905 );
xor ( n20907 , n20630 , n20632 );
xor ( n20908 , n20907 , n20635 );
and ( n20909 , n20906 , n20908 );
xor ( n20910 , n20728 , n20757 );
xor ( n20911 , n20910 , n20760 );
and ( n20912 , n20908 , n20911 );
and ( n20913 , n20906 , n20911 );
or ( n20914 , n20909 , n20912 , n20913 );
and ( n20915 , n20775 , n20914 );
xor ( n20916 , n20775 , n20914 );
xor ( n20917 , n20906 , n20908 );
xor ( n20918 , n20917 , n20911 );
and ( n20919 , n19434 , n20674 );
and ( n20920 , n19418 , n20672 );
nor ( n20921 , n20919 , n20920 );
xnor ( n20922 , n20921 , n20542 );
and ( n20923 , n20004 , n19688 );
and ( n20924 , n19946 , n19686 );
nor ( n20925 , n20923 , n20924 );
xnor ( n20926 , n20925 , n19655 );
and ( n20927 , n20922 , n20926 );
and ( n20928 , n20803 , n19424 );
and ( n20929 , n20666 , n19422 );
nor ( n20930 , n20928 , n20929 );
xnor ( n20931 , n20930 , n19431 );
and ( n20932 , n20926 , n20931 );
and ( n20933 , n20922 , n20931 );
or ( n20934 , n20927 , n20932 , n20933 );
and ( n20935 , n19496 , n20460 );
and ( n20936 , n19469 , n20458 );
nor ( n20937 , n20935 , n20936 );
xnor ( n20938 , n20937 , n20337 );
and ( n20939 , n19811 , n19894 );
and ( n20940 , n19721 , n19892 );
nor ( n20941 , n20939 , n20940 );
xnor ( n20942 , n20941 , n19858 );
and ( n20943 , n20938 , n20942 );
and ( n20944 , n19881 , n19805 );
and ( n20945 , n19825 , n19803 );
nor ( n20946 , n20944 , n20945 );
xnor ( n20947 , n20946 , n19750 );
and ( n20948 , n20942 , n20947 );
and ( n20949 , n20938 , n20947 );
or ( n20950 , n20943 , n20948 , n20949 );
and ( n20951 , n20934 , n20950 );
xor ( n20952 , n20539 , n20776 );
xor ( n20953 , n20776 , n20777 );
not ( n20954 , n20953 );
and ( n20955 , n20952 , n20954 );
and ( n20956 , n19426 , n20955 );
not ( n20957 , n20956 );
xnor ( n20958 , n20957 , n20780 );
and ( n20959 , n19588 , n20276 );
and ( n20960 , n19510 , n20274 );
nor ( n20961 , n20959 , n20960 );
xnor ( n20962 , n20961 , n20175 );
and ( n20963 , n20958 , n20962 );
and ( n20964 , n19637 , n20114 );
and ( n20965 , n19605 , n20112 );
nor ( n20966 , n20964 , n20965 );
xnor ( n20967 , n20966 , n19997 );
and ( n20968 , n20962 , n20967 );
and ( n20969 , n20958 , n20967 );
or ( n20970 , n20963 , n20968 , n20969 );
and ( n20971 , n20950 , n20970 );
and ( n20972 , n20934 , n20970 );
or ( n20973 , n20951 , n20971 , n20972 );
xor ( n20974 , n20781 , n20785 );
xor ( n20975 , n20974 , n20790 );
xor ( n20976 , n20797 , n20801 );
xor ( n20977 , n20976 , n20804 );
and ( n20978 , n20975 , n20977 );
xor ( n20979 , n20817 , n20821 );
xor ( n20980 , n20979 , n20826 );
and ( n20981 , n20977 , n20980 );
and ( n20982 , n20975 , n20980 );
or ( n20983 , n20978 , n20981 , n20982 );
and ( n20984 , n20973 , n20983 );
xor ( n20985 , n20793 , n20807 );
xor ( n20986 , n20985 , n20810 );
and ( n20987 , n20983 , n20986 );
and ( n20988 , n20973 , n20986 );
or ( n20989 , n20984 , n20987 , n20988 );
buf ( n20990 , n19372 );
buf ( n20991 , n19373 );
and ( n20992 , n20990 , n20991 );
not ( n20993 , n20992 );
and ( n20994 , n20777 , n20993 );
not ( n20995 , n20994 );
and ( n20996 , n20080 , n19688 );
and ( n20997 , n20004 , n19686 );
nor ( n20998 , n20996 , n20997 );
xnor ( n20999 , n20998 , n19655 );
and ( n21000 , n20995 , n20999 );
and ( n21001 , n20268 , n19596 );
and ( n21002 , n20182 , n19594 );
nor ( n21003 , n21001 , n21002 );
xnor ( n21004 , n21003 , n19545 );
and ( n21005 , n20999 , n21004 );
and ( n21006 , n20995 , n21004 );
or ( n21007 , n21000 , n21005 , n21006 );
and ( n21008 , n20452 , n19518 );
and ( n21009 , n20360 , n19516 );
nor ( n21010 , n21008 , n21009 );
xnor ( n21011 , n21010 , n19489 );
and ( n21012 , n20666 , n19459 );
and ( n21013 , n20618 , n19457 );
nor ( n21014 , n21012 , n21013 );
xnor ( n21015 , n21014 , n19416 );
and ( n21016 , n21011 , n21015 );
and ( n21017 , n20867 , n19424 );
and ( n21018 , n20803 , n19422 );
nor ( n21019 , n21017 , n21018 );
xnor ( n21020 , n21019 , n19431 );
and ( n21021 , n21015 , n21020 );
and ( n21022 , n21011 , n21020 );
or ( n21023 , n21016 , n21021 , n21022 );
and ( n21024 , n21007 , n21023 );
not ( n21025 , n20875 );
and ( n21026 , n21023 , n21025 );
and ( n21027 , n21007 , n21025 );
or ( n21028 , n21024 , n21026 , n21027 );
xor ( n21029 , n20833 , n20837 );
xor ( n21030 , n21029 , n20842 );
and ( n21031 , n21028 , n21030 );
xor ( n21032 , n20871 , n20876 );
xor ( n21033 , n21032 , n20881 );
and ( n21034 , n21030 , n21033 );
and ( n21035 , n21028 , n21033 );
or ( n21036 , n21031 , n21034 , n21035 );
xor ( n21037 , n20829 , n20845 );
xor ( n21038 , n21037 , n20848 );
and ( n21039 , n21036 , n21038 );
xor ( n21040 , n20884 , n20886 );
xor ( n21041 , n21040 , n20889 );
and ( n21042 , n21038 , n21041 );
and ( n21043 , n21036 , n21041 );
or ( n21044 , n21039 , n21042 , n21043 );
and ( n21045 , n20989 , n21044 );
xor ( n21046 , n20813 , n20851 );
xor ( n21047 , n21046 , n20854 );
and ( n21048 , n21044 , n21047 );
and ( n21049 , n20989 , n21047 );
or ( n21050 , n21045 , n21048 , n21049 );
xor ( n21051 , n20749 , n20751 );
xor ( n21052 , n21051 , n20754 );
and ( n21053 , n21050 , n21052 );
xor ( n21054 , n20857 , n20900 );
xor ( n21055 , n21054 , n20903 );
and ( n21056 , n21052 , n21055 );
and ( n21057 , n21050 , n21055 );
or ( n21058 , n21053 , n21056 , n21057 );
and ( n21059 , n20918 , n21058 );
xor ( n21060 , n20918 , n21058 );
xor ( n21061 , n21050 , n21052 );
xor ( n21062 , n21061 , n21055 );
and ( n21063 , n19418 , n20955 );
and ( n21064 , n19426 , n20953 );
nor ( n21065 , n21063 , n21064 );
xnor ( n21066 , n21065 , n20780 );
and ( n21067 , n19946 , n19805 );
and ( n21068 , n19881 , n19803 );
nor ( n21069 , n21067 , n21068 );
xnor ( n21070 , n21069 , n19750 );
and ( n21071 , n21066 , n21070 );
buf ( n21072 , n19307 );
and ( n21073 , n21072 , n19419 );
and ( n21074 , n21070 , n21073 );
and ( n21075 , n21066 , n21073 );
or ( n21076 , n21071 , n21074 , n21075 );
and ( n21077 , n19510 , n20460 );
and ( n21078 , n19496 , n20458 );
nor ( n21079 , n21077 , n21078 );
xnor ( n21080 , n21079 , n20337 );
and ( n21081 , n19605 , n20276 );
and ( n21082 , n19588 , n20274 );
nor ( n21083 , n21081 , n21082 );
xnor ( n21084 , n21083 , n20175 );
and ( n21085 , n21080 , n21084 );
and ( n21086 , n19721 , n20114 );
and ( n21087 , n19637 , n20112 );
nor ( n21088 , n21086 , n21087 );
xnor ( n21089 , n21088 , n19997 );
and ( n21090 , n21084 , n21089 );
and ( n21091 , n21080 , n21089 );
or ( n21092 , n21085 , n21090 , n21091 );
and ( n21093 , n21076 , n21092 );
xor ( n21094 , n20861 , n20865 );
xor ( n21095 , n21094 , n20868 );
and ( n21096 , n21092 , n21095 );
and ( n21097 , n21076 , n21095 );
or ( n21098 , n21093 , n21096 , n21097 );
xor ( n21099 , n20922 , n20926 );
xor ( n21100 , n21099 , n20931 );
xor ( n21101 , n20938 , n20942 );
xor ( n21102 , n21101 , n20947 );
and ( n21103 , n21100 , n21102 );
xor ( n21104 , n20958 , n20962 );
xor ( n21105 , n21104 , n20967 );
and ( n21106 , n21102 , n21105 );
and ( n21107 , n21100 , n21105 );
or ( n21108 , n21103 , n21106 , n21107 );
and ( n21109 , n21098 , n21108 );
xor ( n21110 , n20975 , n20977 );
xor ( n21111 , n21110 , n20980 );
and ( n21112 , n21108 , n21111 );
and ( n21113 , n21098 , n21111 );
or ( n21114 , n21109 , n21112 , n21113 );
xor ( n21115 , n20973 , n20983 );
xor ( n21116 , n21115 , n20986 );
and ( n21117 , n21114 , n21116 );
xor ( n21118 , n21036 , n21038 );
xor ( n21119 , n21118 , n21041 );
and ( n21120 , n21116 , n21119 );
and ( n21121 , n21114 , n21119 );
or ( n21122 , n21117 , n21120 , n21121 );
xor ( n21123 , n20892 , n20894 );
xor ( n21124 , n21123 , n20897 );
and ( n21125 , n21122 , n21124 );
xor ( n21126 , n20989 , n21044 );
xor ( n21127 , n21126 , n21047 );
and ( n21128 , n21124 , n21127 );
and ( n21129 , n21122 , n21127 );
or ( n21130 , n21125 , n21128 , n21129 );
and ( n21131 , n21062 , n21130 );
xor ( n21132 , n21062 , n21130 );
xor ( n21133 , n21122 , n21124 );
xor ( n21134 , n21133 , n21127 );
and ( n21135 , n20360 , n19596 );
and ( n21136 , n20268 , n19594 );
nor ( n21137 , n21135 , n21136 );
xnor ( n21138 , n21137 , n19545 );
buf ( n21139 , n21138 );
and ( n21140 , n19469 , n20674 );
and ( n21141 , n19434 , n20672 );
nor ( n21142 , n21140 , n21141 );
xnor ( n21143 , n21142 , n20542 );
and ( n21144 , n21139 , n21143 );
and ( n21145 , n19825 , n19894 );
and ( n21146 , n19811 , n19892 );
nor ( n21147 , n21145 , n21146 );
xnor ( n21148 , n21147 , n19858 );
and ( n21149 , n21143 , n21148 );
and ( n21150 , n21139 , n21148 );
or ( n21151 , n21144 , n21149 , n21150 );
xor ( n21152 , n20777 , n20990 );
xor ( n21153 , n20990 , n20991 );
not ( n21154 , n21153 );
and ( n21155 , n21152 , n21154 );
and ( n21156 , n19426 , n21155 );
not ( n21157 , n21156 );
xnor ( n21158 , n21157 , n20994 );
and ( n21159 , n19496 , n20674 );
and ( n21160 , n19469 , n20672 );
nor ( n21161 , n21159 , n21160 );
xnor ( n21162 , n21161 , n20542 );
and ( n21163 , n21158 , n21162 );
and ( n21164 , n19811 , n20114 );
and ( n21165 , n19721 , n20112 );
nor ( n21166 , n21164 , n21165 );
xnor ( n21167 , n21166 , n19997 );
and ( n21168 , n21162 , n21167 );
and ( n21169 , n21158 , n21167 );
or ( n21170 , n21163 , n21168 , n21169 );
xor ( n21171 , n20995 , n20999 );
xor ( n21172 , n21171 , n21004 );
and ( n21173 , n21170 , n21172 );
xor ( n21174 , n21011 , n21015 );
xor ( n21175 , n21174 , n21020 );
and ( n21176 , n21172 , n21175 );
and ( n21177 , n21170 , n21175 );
or ( n21178 , n21173 , n21176 , n21177 );
and ( n21179 , n21151 , n21178 );
xor ( n21180 , n21007 , n21023 );
xor ( n21181 , n21180 , n21025 );
and ( n21182 , n21178 , n21181 );
and ( n21183 , n21151 , n21181 );
or ( n21184 , n21179 , n21182 , n21183 );
xor ( n21185 , n20934 , n20950 );
xor ( n21186 , n21185 , n20970 );
and ( n21187 , n21184 , n21186 );
xor ( n21188 , n21028 , n21030 );
xor ( n21189 , n21188 , n21033 );
and ( n21190 , n21186 , n21189 );
and ( n21191 , n21184 , n21189 );
or ( n21192 , n21187 , n21190 , n21191 );
and ( n21193 , n20182 , n19688 );
and ( n21194 , n20080 , n19686 );
nor ( n21195 , n21193 , n21194 );
xnor ( n21196 , n21195 , n19655 );
and ( n21197 , n20618 , n19518 );
and ( n21198 , n20452 , n19516 );
nor ( n21199 , n21197 , n21198 );
xnor ( n21200 , n21199 , n19489 );
and ( n21201 , n21196 , n21200 );
and ( n21202 , n21072 , n19424 );
and ( n21203 , n20867 , n19422 );
nor ( n21204 , n21202 , n21203 );
xnor ( n21205 , n21204 , n19431 );
and ( n21206 , n21200 , n21205 );
and ( n21207 , n21196 , n21205 );
or ( n21208 , n21201 , n21206 , n21207 );
and ( n21209 , n19434 , n20955 );
and ( n21210 , n19418 , n20953 );
nor ( n21211 , n21209 , n21210 );
xnor ( n21212 , n21211 , n20780 );
and ( n21213 , n20803 , n19459 );
and ( n21214 , n20666 , n19457 );
nor ( n21215 , n21213 , n21214 );
xnor ( n21216 , n21215 , n19416 );
and ( n21217 , n21212 , n21216 );
buf ( n21218 , n19308 );
and ( n21219 , n21218 , n19419 );
and ( n21220 , n21216 , n21219 );
and ( n21221 , n21212 , n21219 );
or ( n21222 , n21217 , n21220 , n21221 );
and ( n21223 , n21208 , n21222 );
and ( n21224 , n19588 , n20460 );
and ( n21225 , n19510 , n20458 );
nor ( n21226 , n21224 , n21225 );
xnor ( n21227 , n21226 , n20337 );
and ( n21228 , n19637 , n20276 );
and ( n21229 , n19605 , n20274 );
nor ( n21230 , n21228 , n21229 );
xnor ( n21231 , n21230 , n20175 );
and ( n21232 , n21227 , n21231 );
and ( n21233 , n20004 , n19805 );
and ( n21234 , n19946 , n19803 );
nor ( n21235 , n21233 , n21234 );
xnor ( n21236 , n21235 , n19750 );
and ( n21237 , n21231 , n21236 );
and ( n21238 , n21227 , n21236 );
or ( n21239 , n21232 , n21237 , n21238 );
and ( n21240 , n21222 , n21239 );
and ( n21241 , n21208 , n21239 );
or ( n21242 , n21223 , n21240 , n21241 );
xor ( n21243 , n21066 , n21070 );
xor ( n21244 , n21243 , n21073 );
xor ( n21245 , n21080 , n21084 );
xor ( n21246 , n21245 , n21089 );
and ( n21247 , n21244 , n21246 );
xor ( n21248 , n21139 , n21143 );
xor ( n21249 , n21248 , n21148 );
and ( n21250 , n21246 , n21249 );
and ( n21251 , n21244 , n21249 );
or ( n21252 , n21247 , n21250 , n21251 );
and ( n21253 , n21242 , n21252 );
xor ( n21254 , n21076 , n21092 );
xor ( n21255 , n21254 , n21095 );
and ( n21256 , n21252 , n21255 );
and ( n21257 , n21242 , n21255 );
or ( n21258 , n21253 , n21256 , n21257 );
xor ( n21259 , n21098 , n21108 );
xor ( n21260 , n21259 , n21111 );
and ( n21261 , n21258 , n21260 );
xor ( n21262 , n21184 , n21186 );
xor ( n21263 , n21262 , n21189 );
and ( n21264 , n21260 , n21263 );
and ( n21265 , n21258 , n21263 );
or ( n21266 , n21261 , n21264 , n21265 );
and ( n21267 , n21192 , n21266 );
xor ( n21268 , n21114 , n21116 );
xor ( n21269 , n21268 , n21119 );
and ( n21270 , n21266 , n21269 );
and ( n21271 , n21192 , n21269 );
or ( n21272 , n21267 , n21270 , n21271 );
and ( n21273 , n21134 , n21272 );
xor ( n21274 , n21134 , n21272 );
xor ( n21275 , n21192 , n21266 );
xor ( n21276 , n21275 , n21269 );
and ( n21277 , n20452 , n19596 );
and ( n21278 , n20360 , n19594 );
nor ( n21279 , n21277 , n21278 );
xnor ( n21280 , n21279 , n19545 );
and ( n21281 , n20666 , n19518 );
and ( n21282 , n20618 , n19516 );
nor ( n21283 , n21281 , n21282 );
xnor ( n21284 , n21283 , n19489 );
and ( n21285 , n21280 , n21284 );
and ( n21286 , n20867 , n19459 );
and ( n21287 , n20803 , n19457 );
nor ( n21288 , n21286 , n21287 );
xnor ( n21289 , n21288 , n19416 );
and ( n21290 , n21284 , n21289 );
and ( n21291 , n21280 , n21289 );
or ( n21292 , n21285 , n21290 , n21291 );
and ( n21293 , n19418 , n21155 );
and ( n21294 , n19426 , n21153 );
nor ( n21295 , n21293 , n21294 );
xnor ( n21296 , n21295 , n20994 );
and ( n21297 , n21218 , n19424 );
and ( n21298 , n21072 , n19422 );
nor ( n21299 , n21297 , n21298 );
xnor ( n21300 , n21299 , n19431 );
and ( n21301 , n21296 , n21300 );
buf ( n21302 , n19309 );
and ( n21303 , n21302 , n19419 );
and ( n21304 , n21300 , n21303 );
and ( n21305 , n21296 , n21303 );
or ( n21306 , n21301 , n21304 , n21305 );
and ( n21307 , n21292 , n21306 );
and ( n21308 , n19510 , n20674 );
and ( n21309 , n19496 , n20672 );
nor ( n21310 , n21308 , n21309 );
xnor ( n21311 , n21310 , n20542 );
and ( n21312 , n19605 , n20460 );
and ( n21313 , n19588 , n20458 );
nor ( n21314 , n21312 , n21313 );
xnor ( n21315 , n21314 , n20337 );
and ( n21316 , n21311 , n21315 );
and ( n21317 , n19946 , n19894 );
and ( n21318 , n19881 , n19892 );
nor ( n21319 , n21317 , n21318 );
xnor ( n21320 , n21319 , n19858 );
and ( n21321 , n21315 , n21320 );
and ( n21322 , n21311 , n21320 );
or ( n21323 , n21316 , n21321 , n21322 );
and ( n21324 , n21306 , n21323 );
and ( n21325 , n21292 , n21323 );
or ( n21326 , n21307 , n21324 , n21325 );
buf ( n21327 , n19374 );
buf ( n21328 , n19375 );
and ( n21329 , n21327 , n21328 );
not ( n21330 , n21329 );
and ( n21331 , n20991 , n21330 );
not ( n21332 , n21331 );
and ( n21333 , n20080 , n19805 );
and ( n21334 , n20004 , n19803 );
nor ( n21335 , n21333 , n21334 );
xnor ( n21336 , n21335 , n19750 );
and ( n21337 , n21332 , n21336 );
and ( n21338 , n20268 , n19688 );
and ( n21339 , n20182 , n19686 );
nor ( n21340 , n21338 , n21339 );
xnor ( n21341 , n21340 , n19655 );
and ( n21342 , n21336 , n21341 );
and ( n21343 , n21332 , n21341 );
or ( n21344 , n21337 , n21342 , n21343 );
and ( n21345 , n19881 , n19894 );
and ( n21346 , n19825 , n19892 );
nor ( n21347 , n21345 , n21346 );
xnor ( n21348 , n21347 , n19858 );
and ( n21349 , n21344 , n21348 );
not ( n21350 , n21138 );
and ( n21351 , n21348 , n21350 );
and ( n21352 , n21344 , n21350 );
or ( n21353 , n21349 , n21351 , n21352 );
and ( n21354 , n21326 , n21353 );
and ( n21355 , n19469 , n20955 );
and ( n21356 , n19434 , n20953 );
nor ( n21357 , n21355 , n21356 );
xnor ( n21358 , n21357 , n20780 );
and ( n21359 , n19721 , n20276 );
and ( n21360 , n19637 , n20274 );
nor ( n21361 , n21359 , n21360 );
xnor ( n21362 , n21361 , n20175 );
and ( n21363 , n21358 , n21362 );
and ( n21364 , n19825 , n20114 );
and ( n21365 , n19811 , n20112 );
nor ( n21366 , n21364 , n21365 );
xnor ( n21367 , n21366 , n19997 );
and ( n21368 , n21362 , n21367 );
and ( n21369 , n21358 , n21367 );
or ( n21370 , n21363 , n21368 , n21369 );
xor ( n21371 , n21196 , n21200 );
xor ( n21372 , n21371 , n21205 );
and ( n21373 , n21370 , n21372 );
xor ( n21374 , n21212 , n21216 );
xor ( n21375 , n21374 , n21219 );
and ( n21376 , n21372 , n21375 );
and ( n21377 , n21370 , n21375 );
or ( n21378 , n21373 , n21376 , n21377 );
and ( n21379 , n21353 , n21378 );
and ( n21380 , n21326 , n21378 );
or ( n21381 , n21354 , n21379 , n21380 );
xor ( n21382 , n21100 , n21102 );
xor ( n21383 , n21382 , n21105 );
and ( n21384 , n21381 , n21383 );
xor ( n21385 , n21151 , n21178 );
xor ( n21386 , n21385 , n21181 );
and ( n21387 , n21383 , n21386 );
and ( n21388 , n21381 , n21386 );
or ( n21389 , n21384 , n21387 , n21388 );
xor ( n21390 , n21158 , n21162 );
xor ( n21391 , n21390 , n21167 );
xor ( n21392 , n21227 , n21231 );
xor ( n21393 , n21392 , n21236 );
and ( n21394 , n21391 , n21393 );
xor ( n21395 , n21344 , n21348 );
xor ( n21396 , n21395 , n21350 );
and ( n21397 , n21393 , n21396 );
and ( n21398 , n21391 , n21396 );
or ( n21399 , n21394 , n21397 , n21398 );
xor ( n21400 , n21208 , n21222 );
xor ( n21401 , n21400 , n21239 );
and ( n21402 , n21399 , n21401 );
xor ( n21403 , n21170 , n21172 );
xor ( n21404 , n21403 , n21175 );
and ( n21405 , n21401 , n21404 );
and ( n21406 , n21399 , n21404 );
or ( n21407 , n21402 , n21405 , n21406 );
xor ( n21408 , n21242 , n21252 );
xor ( n21409 , n21408 , n21255 );
and ( n21410 , n21407 , n21409 );
xor ( n21411 , n21381 , n21383 );
xor ( n21412 , n21411 , n21386 );
and ( n21413 , n21409 , n21412 );
and ( n21414 , n21407 , n21412 );
or ( n21415 , n21410 , n21413 , n21414 );
and ( n21416 , n21389 , n21415 );
xor ( n21417 , n21258 , n21260 );
xor ( n21418 , n21417 , n21263 );
and ( n21419 , n21415 , n21418 );
and ( n21420 , n21389 , n21418 );
or ( n21421 , n21416 , n21419 , n21420 );
and ( n21422 , n21276 , n21421 );
xor ( n21423 , n21276 , n21421 );
xor ( n21424 , n21389 , n21415 );
xor ( n21425 , n21424 , n21418 );
and ( n21426 , n20360 , n19688 );
and ( n21427 , n20268 , n19686 );
nor ( n21428 , n21426 , n21427 );
xnor ( n21429 , n21428 , n19655 );
and ( n21430 , n20618 , n19596 );
and ( n21431 , n20452 , n19594 );
nor ( n21432 , n21430 , n21431 );
xnor ( n21433 , n21432 , n19545 );
and ( n21434 , n21429 , n21433 );
and ( n21435 , n20803 , n19518 );
and ( n21436 , n20666 , n19516 );
nor ( n21437 , n21435 , n21436 );
xnor ( n21438 , n21437 , n19489 );
and ( n21439 , n21433 , n21438 );
and ( n21440 , n21429 , n21438 );
or ( n21441 , n21434 , n21439 , n21440 );
and ( n21442 , n21072 , n19459 );
and ( n21443 , n20867 , n19457 );
nor ( n21444 , n21442 , n21443 );
xnor ( n21445 , n21444 , n19416 );
and ( n21446 , n21302 , n19424 );
and ( n21447 , n21218 , n19422 );
nor ( n21448 , n21446 , n21447 );
xnor ( n21449 , n21448 , n19431 );
and ( n21450 , n21445 , n21449 );
buf ( n21451 , n19310 );
and ( n21452 , n21451 , n19419 );
and ( n21453 , n21449 , n21452 );
and ( n21454 , n21445 , n21452 );
or ( n21455 , n21450 , n21453 , n21454 );
and ( n21456 , n21441 , n21455 );
and ( n21457 , n20182 , n19805 );
and ( n21458 , n20080 , n19803 );
nor ( n21459 , n21457 , n21458 );
xnor ( n21460 , n21459 , n19750 );
buf ( n21461 , n21460 );
and ( n21462 , n21455 , n21461 );
and ( n21463 , n21441 , n21461 );
or ( n21464 , n21456 , n21462 , n21463 );
xor ( n21465 , n20991 , n21327 );
xor ( n21466 , n21327 , n21328 );
not ( n21467 , n21466 );
and ( n21468 , n21465 , n21467 );
and ( n21469 , n19426 , n21468 );
not ( n21470 , n21469 );
xnor ( n21471 , n21470 , n21331 );
and ( n21472 , n19637 , n20460 );
and ( n21473 , n19605 , n20458 );
nor ( n21474 , n21472 , n21473 );
xnor ( n21475 , n21474 , n20337 );
and ( n21476 , n21471 , n21475 );
and ( n21477 , n19811 , n20276 );
and ( n21478 , n19721 , n20274 );
nor ( n21479 , n21477 , n21478 );
xnor ( n21480 , n21479 , n20175 );
and ( n21481 , n21475 , n21480 );
and ( n21482 , n21471 , n21480 );
or ( n21483 , n21476 , n21481 , n21482 );
and ( n21484 , n19434 , n21155 );
and ( n21485 , n19418 , n21153 );
nor ( n21486 , n21484 , n21485 );
xnor ( n21487 , n21486 , n20994 );
and ( n21488 , n19588 , n20674 );
and ( n21489 , n19510 , n20672 );
nor ( n21490 , n21488 , n21489 );
xnor ( n21491 , n21490 , n20542 );
and ( n21492 , n21487 , n21491 );
and ( n21493 , n20004 , n19894 );
and ( n21494 , n19946 , n19892 );
nor ( n21495 , n21493 , n21494 );
xnor ( n21496 , n21495 , n19858 );
and ( n21497 , n21491 , n21496 );
and ( n21498 , n21487 , n21496 );
or ( n21499 , n21492 , n21497 , n21498 );
and ( n21500 , n21483 , n21499 );
xor ( n21501 , n21296 , n21300 );
xor ( n21502 , n21501 , n21303 );
and ( n21503 , n21499 , n21502 );
and ( n21504 , n21483 , n21502 );
or ( n21505 , n21500 , n21503 , n21504 );
and ( n21506 , n21464 , n21505 );
xor ( n21507 , n21292 , n21306 );
xor ( n21508 , n21507 , n21323 );
and ( n21509 , n21505 , n21508 );
and ( n21510 , n21464 , n21508 );
or ( n21511 , n21506 , n21509 , n21510 );
xor ( n21512 , n21326 , n21353 );
xor ( n21513 , n21512 , n21378 );
and ( n21514 , n21511 , n21513 );
xor ( n21515 , n21244 , n21246 );
xor ( n21516 , n21515 , n21249 );
and ( n21517 , n21513 , n21516 );
and ( n21518 , n21511 , n21516 );
or ( n21519 , n21514 , n21517 , n21518 );
xor ( n21520 , n21429 , n21433 );
xor ( n21521 , n21520 , n21438 );
xor ( n21522 , n21471 , n21475 );
xor ( n21523 , n21522 , n21480 );
and ( n21524 , n21521 , n21523 );
and ( n21525 , n19496 , n20955 );
and ( n21526 , n19469 , n20953 );
nor ( n21527 , n21525 , n21526 );
xnor ( n21528 , n21527 , n20780 );
and ( n21529 , n19881 , n20114 );
and ( n21530 , n19825 , n20112 );
nor ( n21531 , n21529 , n21530 );
xnor ( n21532 , n21531 , n19997 );
xor ( n21533 , n21528 , n21532 );
not ( n21534 , n21460 );
xor ( n21535 , n21533 , n21534 );
and ( n21536 , n21523 , n21535 );
and ( n21537 , n21521 , n21535 );
or ( n21538 , n21524 , n21536 , n21537 );
and ( n21539 , n19469 , n21155 );
and ( n21540 , n19434 , n21153 );
nor ( n21541 , n21539 , n21540 );
xnor ( n21542 , n21541 , n20994 );
and ( n21543 , n19605 , n20674 );
and ( n21544 , n19588 , n20672 );
nor ( n21545 , n21543 , n21544 );
xnor ( n21546 , n21545 , n20542 );
and ( n21547 , n21542 , n21546 );
and ( n21548 , n19721 , n20460 );
and ( n21549 , n19637 , n20458 );
nor ( n21550 , n21548 , n21549 );
xnor ( n21551 , n21550 , n20337 );
and ( n21552 , n21546 , n21551 );
and ( n21553 , n21542 , n21551 );
or ( n21554 , n21547 , n21552 , n21553 );
and ( n21555 , n19418 , n21468 );
and ( n21556 , n19426 , n21466 );
nor ( n21557 , n21555 , n21556 );
xnor ( n21558 , n21557 , n21331 );
and ( n21559 , n19510 , n20955 );
and ( n21560 , n19496 , n20953 );
nor ( n21561 , n21559 , n21560 );
xnor ( n21562 , n21561 , n20780 );
and ( n21563 , n21558 , n21562 );
and ( n21564 , n19946 , n20114 );
and ( n21565 , n19881 , n20112 );
nor ( n21566 , n21564 , n21565 );
xnor ( n21567 , n21566 , n19997 );
and ( n21568 , n21562 , n21567 );
and ( n21569 , n21558 , n21567 );
or ( n21570 , n21563 , n21568 , n21569 );
and ( n21571 , n21554 , n21570 );
xor ( n21572 , n21445 , n21449 );
xor ( n21573 , n21572 , n21452 );
and ( n21574 , n21570 , n21573 );
and ( n21575 , n21554 , n21573 );
or ( n21576 , n21571 , n21574 , n21575 );
and ( n21577 , n21538 , n21576 );
xor ( n21578 , n21441 , n21455 );
xor ( n21579 , n21578 , n21461 );
and ( n21580 , n21576 , n21579 );
and ( n21581 , n21538 , n21579 );
or ( n21582 , n21577 , n21580 , n21581 );
xor ( n21583 , n21391 , n21393 );
xor ( n21584 , n21583 , n21396 );
and ( n21585 , n21582 , n21584 );
xor ( n21586 , n21464 , n21505 );
xor ( n21587 , n21586 , n21508 );
and ( n21588 , n21584 , n21587 );
and ( n21589 , n21582 , n21587 );
or ( n21590 , n21585 , n21588 , n21589 );
xor ( n21591 , n21332 , n21336 );
xor ( n21592 , n21591 , n21341 );
xor ( n21593 , n21280 , n21284 );
xor ( n21594 , n21593 , n21289 );
and ( n21595 , n21592 , n21594 );
xor ( n21596 , n21358 , n21362 );
xor ( n21597 , n21596 , n21367 );
and ( n21598 , n21594 , n21597 );
and ( n21599 , n21592 , n21597 );
or ( n21600 , n21595 , n21598 , n21599 );
buf ( n21601 , n19376 );
buf ( n21602 , n19377 );
and ( n21603 , n21601 , n21602 );
not ( n21604 , n21603 );
and ( n21605 , n21328 , n21604 );
not ( n21606 , n21605 );
and ( n21607 , n20080 , n19894 );
and ( n21608 , n20004 , n19892 );
nor ( n21609 , n21607 , n21608 );
xnor ( n21610 , n21609 , n19858 );
and ( n21611 , n21606 , n21610 );
buf ( n21612 , n19311 );
and ( n21613 , n21612 , n19419 );
and ( n21614 , n21610 , n21613 );
and ( n21615 , n21606 , n21613 );
or ( n21616 , n21611 , n21614 , n21615 );
and ( n21617 , n20268 , n19805 );
and ( n21618 , n20182 , n19803 );
nor ( n21619 , n21617 , n21618 );
xnor ( n21620 , n21619 , n19750 );
and ( n21621 , n20452 , n19688 );
and ( n21622 , n20360 , n19686 );
nor ( n21623 , n21621 , n21622 );
xnor ( n21624 , n21623 , n19655 );
and ( n21625 , n21620 , n21624 );
and ( n21626 , n20666 , n19596 );
and ( n21627 , n20618 , n19594 );
nor ( n21628 , n21626 , n21627 );
xnor ( n21629 , n21628 , n19545 );
and ( n21630 , n21624 , n21629 );
and ( n21631 , n21620 , n21629 );
or ( n21632 , n21625 , n21630 , n21631 );
and ( n21633 , n21616 , n21632 );
and ( n21634 , n20867 , n19518 );
and ( n21635 , n20803 , n19516 );
nor ( n21636 , n21634 , n21635 );
xnor ( n21637 , n21636 , n19489 );
and ( n21638 , n21218 , n19459 );
and ( n21639 , n21072 , n19457 );
nor ( n21640 , n21638 , n21639 );
xnor ( n21641 , n21640 , n19416 );
and ( n21642 , n21637 , n21641 );
and ( n21643 , n21451 , n19424 );
and ( n21644 , n21302 , n19422 );
nor ( n21645 , n21643 , n21644 );
xnor ( n21646 , n21645 , n19431 );
and ( n21647 , n21641 , n21646 );
and ( n21648 , n21637 , n21646 );
or ( n21649 , n21642 , n21647 , n21648 );
and ( n21650 , n21632 , n21649 );
and ( n21651 , n21616 , n21649 );
or ( n21652 , n21633 , n21650 , n21651 );
and ( n21653 , n21528 , n21532 );
and ( n21654 , n21532 , n21534 );
and ( n21655 , n21528 , n21534 );
or ( n21656 , n21653 , n21654 , n21655 );
and ( n21657 , n21652 , n21656 );
xor ( n21658 , n21311 , n21315 );
xor ( n21659 , n21658 , n21320 );
and ( n21660 , n21656 , n21659 );
and ( n21661 , n21652 , n21659 );
or ( n21662 , n21657 , n21660 , n21661 );
and ( n21663 , n21600 , n21662 );
xor ( n21664 , n21370 , n21372 );
xor ( n21665 , n21664 , n21375 );
and ( n21666 , n21662 , n21665 );
and ( n21667 , n21600 , n21665 );
or ( n21668 , n21663 , n21666 , n21667 );
and ( n21669 , n21590 , n21668 );
xor ( n21670 , n21399 , n21401 );
xor ( n21671 , n21670 , n21404 );
and ( n21672 , n21668 , n21671 );
and ( n21673 , n21590 , n21671 );
or ( n21674 , n21669 , n21672 , n21673 );
and ( n21675 , n21519 , n21674 );
xor ( n21676 , n21407 , n21409 );
xor ( n21677 , n21676 , n21412 );
and ( n21678 , n21674 , n21677 );
and ( n21679 , n21519 , n21677 );
or ( n21680 , n21675 , n21678 , n21679 );
and ( n21681 , n21425 , n21680 );
xor ( n21682 , n21425 , n21680 );
xor ( n21683 , n21519 , n21674 );
xor ( n21684 , n21683 , n21677 );
xor ( n21685 , n21483 , n21499 );
xor ( n21686 , n21685 , n21502 );
xor ( n21687 , n21592 , n21594 );
xor ( n21688 , n21687 , n21597 );
and ( n21689 , n21686 , n21688 );
xor ( n21690 , n21652 , n21656 );
xor ( n21691 , n21690 , n21659 );
and ( n21692 , n21688 , n21691 );
and ( n21693 , n21686 , n21691 );
or ( n21694 , n21689 , n21692 , n21693 );
and ( n21695 , n20360 , n19805 );
and ( n21696 , n20268 , n19803 );
nor ( n21697 , n21695 , n21696 );
xnor ( n21698 , n21697 , n19750 );
and ( n21699 , n20618 , n19688 );
and ( n21700 , n20452 , n19686 );
nor ( n21701 , n21699 , n21700 );
xnor ( n21702 , n21701 , n19655 );
and ( n21703 , n21698 , n21702 );
buf ( n21704 , n19312 );
and ( n21705 , n21704 , n19419 );
and ( n21706 , n21702 , n21705 );
and ( n21707 , n21698 , n21705 );
or ( n21708 , n21703 , n21706 , n21707 );
and ( n21709 , n20182 , n19894 );
and ( n21710 , n20080 , n19892 );
nor ( n21711 , n21709 , n21710 );
xnor ( n21712 , n21711 , n19858 );
buf ( n21713 , n21712 );
and ( n21714 , n21708 , n21713 );
and ( n21715 , n19825 , n20276 );
and ( n21716 , n19811 , n20274 );
nor ( n21717 , n21715 , n21716 );
xnor ( n21718 , n21717 , n20175 );
and ( n21719 , n21713 , n21718 );
and ( n21720 , n21708 , n21718 );
or ( n21721 , n21714 , n21719 , n21720 );
and ( n21722 , n19496 , n21155 );
and ( n21723 , n19469 , n21153 );
nor ( n21724 , n21722 , n21723 );
xnor ( n21725 , n21724 , n20994 );
and ( n21726 , n19811 , n20460 );
and ( n21727 , n19721 , n20458 );
nor ( n21728 , n21726 , n21727 );
xnor ( n21729 , n21728 , n20337 );
and ( n21730 , n21725 , n21729 );
and ( n21731 , n19881 , n20276 );
and ( n21732 , n19825 , n20274 );
nor ( n21733 , n21731 , n21732 );
xnor ( n21734 , n21733 , n20175 );
and ( n21735 , n21729 , n21734 );
and ( n21736 , n21725 , n21734 );
or ( n21737 , n21730 , n21735 , n21736 );
xor ( n21738 , n21328 , n21601 );
xor ( n21739 , n21601 , n21602 );
not ( n21740 , n21739 );
and ( n21741 , n21738 , n21740 );
and ( n21742 , n19426 , n21741 );
not ( n21743 , n21742 );
xnor ( n21744 , n21743 , n21605 );
and ( n21745 , n19588 , n20955 );
and ( n21746 , n19510 , n20953 );
nor ( n21747 , n21745 , n21746 );
xnor ( n21748 , n21747 , n20780 );
and ( n21749 , n21744 , n21748 );
and ( n21750 , n19637 , n20674 );
and ( n21751 , n19605 , n20672 );
nor ( n21752 , n21750 , n21751 );
xnor ( n21753 , n21752 , n20542 );
and ( n21754 , n21748 , n21753 );
and ( n21755 , n21744 , n21753 );
or ( n21756 , n21749 , n21754 , n21755 );
and ( n21757 , n21737 , n21756 );
xor ( n21758 , n21637 , n21641 );
xor ( n21759 , n21758 , n21646 );
and ( n21760 , n21756 , n21759 );
and ( n21761 , n21737 , n21759 );
or ( n21762 , n21757 , n21760 , n21761 );
and ( n21763 , n21721 , n21762 );
xor ( n21764 , n21487 , n21491 );
xor ( n21765 , n21764 , n21496 );
and ( n21766 , n21762 , n21765 );
and ( n21767 , n21721 , n21765 );
or ( n21768 , n21763 , n21766 , n21767 );
and ( n21769 , n20803 , n19596 );
and ( n21770 , n20666 , n19594 );
nor ( n21771 , n21769 , n21770 );
xnor ( n21772 , n21771 , n19545 );
and ( n21773 , n21072 , n19518 );
and ( n21774 , n20867 , n19516 );
nor ( n21775 , n21773 , n21774 );
xnor ( n21776 , n21775 , n19489 );
and ( n21777 , n21772 , n21776 );
and ( n21778 , n21302 , n19459 );
and ( n21779 , n21218 , n19457 );
nor ( n21780 , n21778 , n21779 );
xnor ( n21781 , n21780 , n19416 );
and ( n21782 , n21776 , n21781 );
and ( n21783 , n21772 , n21781 );
or ( n21784 , n21777 , n21782 , n21783 );
and ( n21785 , n19434 , n21468 );
and ( n21786 , n19418 , n21466 );
nor ( n21787 , n21785 , n21786 );
xnor ( n21788 , n21787 , n21331 );
and ( n21789 , n20004 , n20114 );
and ( n21790 , n19946 , n20112 );
nor ( n21791 , n21789 , n21790 );
xnor ( n21792 , n21791 , n19997 );
and ( n21793 , n21788 , n21792 );
and ( n21794 , n21612 , n19424 );
and ( n21795 , n21451 , n19422 );
nor ( n21796 , n21794 , n21795 );
xnor ( n21797 , n21796 , n19431 );
and ( n21798 , n21792 , n21797 );
and ( n21799 , n21788 , n21797 );
or ( n21800 , n21793 , n21798 , n21799 );
and ( n21801 , n21784 , n21800 );
xor ( n21802 , n21606 , n21610 );
xor ( n21803 , n21802 , n21613 );
and ( n21804 , n21800 , n21803 );
and ( n21805 , n21784 , n21803 );
or ( n21806 , n21801 , n21804 , n21805 );
xor ( n21807 , n21616 , n21632 );
xor ( n21808 , n21807 , n21649 );
and ( n21809 , n21806 , n21808 );
xor ( n21810 , n21554 , n21570 );
xor ( n21811 , n21810 , n21573 );
and ( n21812 , n21808 , n21811 );
and ( n21813 , n21806 , n21811 );
or ( n21814 , n21809 , n21812 , n21813 );
and ( n21815 , n21768 , n21814 );
xor ( n21816 , n21538 , n21576 );
xor ( n21817 , n21816 , n21579 );
and ( n21818 , n21814 , n21817 );
and ( n21819 , n21768 , n21817 );
or ( n21820 , n21815 , n21818 , n21819 );
and ( n21821 , n21694 , n21820 );
xor ( n21822 , n21600 , n21662 );
xor ( n21823 , n21822 , n21665 );
and ( n21824 , n21820 , n21823 );
and ( n21825 , n21694 , n21823 );
or ( n21826 , n21821 , n21824 , n21825 );
xor ( n21827 , n21511 , n21513 );
xor ( n21828 , n21827 , n21516 );
and ( n21829 , n21826 , n21828 );
xor ( n21830 , n21590 , n21668 );
xor ( n21831 , n21830 , n21671 );
and ( n21832 , n21828 , n21831 );
and ( n21833 , n21826 , n21831 );
or ( n21834 , n21829 , n21832 , n21833 );
and ( n21835 , n21684 , n21834 );
xor ( n21836 , n21684 , n21834 );
xor ( n21837 , n21826 , n21828 );
xor ( n21838 , n21837 , n21831 );
xor ( n21839 , n21620 , n21624 );
xor ( n21840 , n21839 , n21629 );
xor ( n21841 , n21542 , n21546 );
xor ( n21842 , n21841 , n21551 );
and ( n21843 , n21840 , n21842 );
xor ( n21844 , n21558 , n21562 );
xor ( n21845 , n21844 , n21567 );
and ( n21846 , n21842 , n21845 );
and ( n21847 , n21840 , n21845 );
or ( n21848 , n21843 , n21846 , n21847 );
buf ( n21849 , n19378 );
buf ( n21850 , n19379 );
and ( n21851 , n21849 , n21850 );
not ( n21852 , n21851 );
and ( n21853 , n21602 , n21852 );
not ( n21854 , n21853 );
and ( n21855 , n20080 , n20114 );
and ( n21856 , n20004 , n20112 );
nor ( n21857 , n21855 , n21856 );
xnor ( n21858 , n21857 , n19997 );
and ( n21859 , n21854 , n21858 );
and ( n21860 , n21704 , n19424 );
and ( n21861 , n21612 , n19422 );
nor ( n21862 , n21860 , n21861 );
xnor ( n21863 , n21862 , n19431 );
and ( n21864 , n21858 , n21863 );
and ( n21865 , n21854 , n21863 );
or ( n21866 , n21859 , n21864 , n21865 );
and ( n21867 , n20268 , n19894 );
and ( n21868 , n20182 , n19892 );
nor ( n21869 , n21867 , n21868 );
xnor ( n21870 , n21869 , n19858 );
and ( n21871 , n20452 , n19805 );
and ( n21872 , n20360 , n19803 );
nor ( n21873 , n21871 , n21872 );
xnor ( n21874 , n21873 , n19750 );
and ( n21875 , n21870 , n21874 );
buf ( n21876 , n19313 );
and ( n21877 , n21876 , n19419 );
and ( n21878 , n21874 , n21877 );
and ( n21879 , n21870 , n21877 );
or ( n21880 , n21875 , n21878 , n21879 );
and ( n21881 , n21866 , n21880 );
not ( n21882 , n21712 );
and ( n21883 , n21880 , n21882 );
and ( n21884 , n21866 , n21882 );
or ( n21885 , n21881 , n21883 , n21884 );
and ( n21886 , n19469 , n21468 );
and ( n21887 , n19434 , n21466 );
nor ( n21888 , n21886 , n21887 );
xnor ( n21889 , n21888 , n21331 );
and ( n21890 , n19721 , n20674 );
and ( n21891 , n19637 , n20672 );
nor ( n21892 , n21890 , n21891 );
xnor ( n21893 , n21892 , n20542 );
and ( n21894 , n21889 , n21893 );
and ( n21895 , n19825 , n20460 );
and ( n21896 , n19811 , n20458 );
nor ( n21897 , n21895 , n21896 );
xnor ( n21898 , n21897 , n20337 );
and ( n21899 , n21893 , n21898 );
and ( n21900 , n21889 , n21898 );
or ( n21901 , n21894 , n21899 , n21900 );
xor ( n21902 , n21698 , n21702 );
xor ( n21903 , n21902 , n21705 );
and ( n21904 , n21901 , n21903 );
xor ( n21905 , n21772 , n21776 );
xor ( n21906 , n21905 , n21781 );
and ( n21907 , n21903 , n21906 );
and ( n21908 , n21901 , n21906 );
or ( n21909 , n21904 , n21907 , n21908 );
and ( n21910 , n21885 , n21909 );
xor ( n21911 , n21708 , n21713 );
xor ( n21912 , n21911 , n21718 );
and ( n21913 , n21909 , n21912 );
and ( n21914 , n21885 , n21912 );
or ( n21915 , n21910 , n21913 , n21914 );
and ( n21916 , n21848 , n21915 );
xor ( n21917 , n21521 , n21523 );
xor ( n21918 , n21917 , n21535 );
and ( n21919 , n21915 , n21918 );
and ( n21920 , n21848 , n21918 );
or ( n21921 , n21916 , n21919 , n21920 );
and ( n21922 , n20666 , n19688 );
and ( n21923 , n20618 , n19686 );
nor ( n21924 , n21922 , n21923 );
xnor ( n21925 , n21924 , n19655 );
and ( n21926 , n20867 , n19596 );
and ( n21927 , n20803 , n19594 );
nor ( n21928 , n21926 , n21927 );
xnor ( n21929 , n21928 , n19545 );
and ( n21930 , n21925 , n21929 );
and ( n21931 , n21218 , n19518 );
and ( n21932 , n21072 , n19516 );
nor ( n21933 , n21931 , n21932 );
xnor ( n21934 , n21933 , n19489 );
and ( n21935 , n21929 , n21934 );
and ( n21936 , n21925 , n21934 );
or ( n21937 , n21930 , n21935 , n21936 );
and ( n21938 , n19418 , n21741 );
and ( n21939 , n19426 , n21739 );
nor ( n21940 , n21938 , n21939 );
xnor ( n21941 , n21940 , n21605 );
and ( n21942 , n19946 , n20276 );
and ( n21943 , n19881 , n20274 );
nor ( n21944 , n21942 , n21943 );
xnor ( n21945 , n21944 , n20175 );
and ( n21946 , n21941 , n21945 );
and ( n21947 , n21451 , n19459 );
and ( n21948 , n21302 , n19457 );
nor ( n21949 , n21947 , n21948 );
xnor ( n21950 , n21949 , n19416 );
and ( n21951 , n21945 , n21950 );
and ( n21952 , n21941 , n21950 );
or ( n21953 , n21946 , n21951 , n21952 );
and ( n21954 , n21937 , n21953 );
buf ( n21955 , n19314 );
and ( n21956 , n21955 , n19419 );
buf ( n21957 , n21956 );
and ( n21958 , n19510 , n21155 );
and ( n21959 , n19496 , n21153 );
nor ( n21960 , n21958 , n21959 );
xnor ( n21961 , n21960 , n20994 );
and ( n21962 , n21957 , n21961 );
and ( n21963 , n19605 , n20955 );
and ( n21964 , n19588 , n20953 );
nor ( n21965 , n21963 , n21964 );
xnor ( n21966 , n21965 , n20780 );
and ( n21967 , n21961 , n21966 );
and ( n21968 , n21957 , n21966 );
or ( n21969 , n21962 , n21967 , n21968 );
and ( n21970 , n21953 , n21969 );
and ( n21971 , n21937 , n21969 );
or ( n21972 , n21954 , n21970 , n21971 );
xor ( n21973 , n21725 , n21729 );
xor ( n21974 , n21973 , n21734 );
xor ( n21975 , n21788 , n21792 );
xor ( n21976 , n21975 , n21797 );
and ( n21977 , n21974 , n21976 );
xor ( n21978 , n21744 , n21748 );
xor ( n21979 , n21978 , n21753 );
and ( n21980 , n21976 , n21979 );
and ( n21981 , n21974 , n21979 );
or ( n21982 , n21977 , n21980 , n21981 );
and ( n21983 , n21972 , n21982 );
xor ( n21984 , n21784 , n21800 );
xor ( n21985 , n21984 , n21803 );
and ( n21986 , n21982 , n21985 );
and ( n21987 , n21972 , n21985 );
or ( n21988 , n21983 , n21986 , n21987 );
xor ( n21989 , n21721 , n21762 );
xor ( n21990 , n21989 , n21765 );
and ( n21991 , n21988 , n21990 );
xor ( n21992 , n21806 , n21808 );
xor ( n21993 , n21992 , n21811 );
and ( n21994 , n21990 , n21993 );
and ( n21995 , n21988 , n21993 );
or ( n21996 , n21991 , n21994 , n21995 );
and ( n21997 , n21921 , n21996 );
xor ( n21998 , n21686 , n21688 );
xor ( n21999 , n21998 , n21691 );
and ( n22000 , n21996 , n21999 );
and ( n22001 , n21921 , n21999 );
or ( n22002 , n21997 , n22000 , n22001 );
xor ( n22003 , n21582 , n21584 );
xor ( n22004 , n22003 , n21587 );
and ( n22005 , n22002 , n22004 );
xor ( n22006 , n21694 , n21820 );
xor ( n22007 , n22006 , n21823 );
and ( n22008 , n22004 , n22007 );
and ( n22009 , n22002 , n22007 );
or ( n22010 , n22005 , n22008 , n22009 );
and ( n22011 , n21838 , n22010 );
xor ( n22012 , n21838 , n22010 );
xor ( n22013 , n22002 , n22004 );
xor ( n22014 , n22013 , n22007 );
xor ( n22015 , n21737 , n21756 );
xor ( n22016 , n22015 , n21759 );
xor ( n22017 , n21840 , n21842 );
xor ( n22018 , n22017 , n21845 );
and ( n22019 , n22016 , n22018 );
xor ( n22020 , n21885 , n21909 );
xor ( n22021 , n22020 , n21912 );
and ( n22022 , n22018 , n22021 );
and ( n22023 , n22016 , n22021 );
or ( n22024 , n22019 , n22022 , n22023 );
xor ( n22025 , n21848 , n21915 );
xor ( n22026 , n22025 , n21918 );
and ( n22027 , n22024 , n22026 );
xor ( n22028 , n21988 , n21990 );
xor ( n22029 , n22028 , n21993 );
and ( n22030 , n22026 , n22029 );
and ( n22031 , n22024 , n22029 );
or ( n22032 , n22027 , n22030 , n22031 );
xor ( n22033 , n21768 , n21814 );
xor ( n22034 , n22033 , n21817 );
and ( n22035 , n22032 , n22034 );
xor ( n22036 , n21921 , n21996 );
xor ( n22037 , n22036 , n21999 );
and ( n22038 , n22034 , n22037 );
and ( n22039 , n22032 , n22037 );
or ( n22040 , n22035 , n22038 , n22039 );
and ( n22041 , n22014 , n22040 );
xor ( n22042 , n22014 , n22040 );
xor ( n22043 , n22032 , n22034 );
xor ( n22044 , n22043 , n22037 );
xor ( n22045 , n21602 , n21849 );
xor ( n22046 , n21849 , n21850 );
not ( n22047 , n22046 );
and ( n22048 , n22045 , n22047 );
and ( n22049 , n19426 , n22048 );
not ( n22050 , n22049 );
xnor ( n22051 , n22050 , n21853 );
and ( n22052 , n19637 , n20955 );
and ( n22053 , n19605 , n20953 );
nor ( n22054 , n22052 , n22053 );
xnor ( n22055 , n22054 , n20780 );
and ( n22056 , n22051 , n22055 );
and ( n22057 , n19811 , n20674 );
and ( n22058 , n19721 , n20672 );
nor ( n22059 , n22057 , n22058 );
xnor ( n22060 , n22059 , n20542 );
and ( n22061 , n22055 , n22060 );
and ( n22062 , n22051 , n22060 );
or ( n22063 , n22056 , n22061 , n22062 );
and ( n22064 , n19434 , n21741 );
and ( n22065 , n19418 , n21739 );
nor ( n22066 , n22064 , n22065 );
xnor ( n22067 , n22066 , n21605 );
and ( n22068 , n19588 , n21155 );
and ( n22069 , n19510 , n21153 );
nor ( n22070 , n22068 , n22069 );
xnor ( n22071 , n22070 , n20994 );
and ( n22072 , n22067 , n22071 );
and ( n22073 , n20004 , n20276 );
and ( n22074 , n19946 , n20274 );
nor ( n22075 , n22073 , n22074 );
xnor ( n22076 , n22075 , n20175 );
and ( n22077 , n22071 , n22076 );
and ( n22078 , n22067 , n22076 );
or ( n22079 , n22072 , n22077 , n22078 );
and ( n22080 , n22063 , n22079 );
and ( n22081 , n21302 , n19518 );
and ( n22082 , n21218 , n19516 );
nor ( n22083 , n22081 , n22082 );
xnor ( n22084 , n22083 , n19489 );
and ( n22085 , n21612 , n19459 );
and ( n22086 , n21451 , n19457 );
nor ( n22087 , n22085 , n22086 );
xnor ( n22088 , n22087 , n19416 );
and ( n22089 , n22084 , n22088 );
not ( n22090 , n21956 );
and ( n22091 , n22088 , n22090 );
and ( n22092 , n22084 , n22090 );
or ( n22093 , n22089 , n22091 , n22092 );
and ( n22094 , n22079 , n22093 );
and ( n22095 , n22063 , n22093 );
or ( n22096 , n22080 , n22094 , n22095 );
and ( n22097 , n20182 , n20114 );
and ( n22098 , n20080 , n20112 );
nor ( n22099 , n22097 , n22098 );
xnor ( n22100 , n22099 , n19997 );
and ( n22101 , n20360 , n19894 );
and ( n22102 , n20268 , n19892 );
nor ( n22103 , n22101 , n22102 );
xnor ( n22104 , n22103 , n19858 );
and ( n22105 , n22100 , n22104 );
and ( n22106 , n21876 , n19424 );
and ( n22107 , n21704 , n19422 );
nor ( n22108 , n22106 , n22107 );
xnor ( n22109 , n22108 , n19431 );
and ( n22110 , n22104 , n22109 );
and ( n22111 , n22100 , n22109 );
or ( n22112 , n22105 , n22110 , n22111 );
and ( n22113 , n20618 , n19805 );
and ( n22114 , n20452 , n19803 );
nor ( n22115 , n22113 , n22114 );
xnor ( n22116 , n22115 , n19750 );
and ( n22117 , n20803 , n19688 );
and ( n22118 , n20666 , n19686 );
nor ( n22119 , n22117 , n22118 );
xnor ( n22120 , n22119 , n19655 );
and ( n22121 , n22116 , n22120 );
and ( n22122 , n21072 , n19596 );
and ( n22123 , n20867 , n19594 );
nor ( n22124 , n22122 , n22123 );
xnor ( n22125 , n22124 , n19545 );
and ( n22126 , n22120 , n22125 );
and ( n22127 , n22116 , n22125 );
or ( n22128 , n22121 , n22126 , n22127 );
and ( n22129 , n22112 , n22128 );
xor ( n22130 , n21854 , n21858 );
xor ( n22131 , n22130 , n21863 );
and ( n22132 , n22128 , n22131 );
and ( n22133 , n22112 , n22131 );
or ( n22134 , n22129 , n22132 , n22133 );
and ( n22135 , n22096 , n22134 );
xor ( n22136 , n21866 , n21880 );
xor ( n22137 , n22136 , n21882 );
and ( n22138 , n22134 , n22137 );
and ( n22139 , n22096 , n22137 );
or ( n22140 , n22135 , n22138 , n22139 );
xor ( n22141 , n21870 , n21874 );
xor ( n22142 , n22141 , n21877 );
xor ( n22143 , n21925 , n21929 );
xor ( n22144 , n22143 , n21934 );
and ( n22145 , n22142 , n22144 );
xor ( n22146 , n21889 , n21893 );
xor ( n22147 , n22146 , n21898 );
and ( n22148 , n22144 , n22147 );
and ( n22149 , n22142 , n22147 );
or ( n22150 , n22145 , n22148 , n22149 );
xor ( n22151 , n21937 , n21953 );
xor ( n22152 , n22151 , n21969 );
and ( n22153 , n22150 , n22152 );
xor ( n22154 , n21901 , n21903 );
xor ( n22155 , n22154 , n21906 );
and ( n22156 , n22152 , n22155 );
and ( n22157 , n22150 , n22155 );
or ( n22158 , n22153 , n22156 , n22157 );
and ( n22159 , n22140 , n22158 );
xor ( n22160 , n21972 , n21982 );
xor ( n22161 , n22160 , n21985 );
and ( n22162 , n22158 , n22161 );
and ( n22163 , n22140 , n22161 );
or ( n22164 , n22159 , n22162 , n22163 );
and ( n22165 , n20867 , n19688 );
and ( n22166 , n20803 , n19686 );
nor ( n22167 , n22165 , n22166 );
xnor ( n22168 , n22167 , n19655 );
and ( n22169 , n21218 , n19596 );
and ( n22170 , n21072 , n19594 );
nor ( n22171 , n22169 , n22170 );
xnor ( n22172 , n22171 , n19545 );
and ( n22173 , n22168 , n22172 );
and ( n22174 , n21451 , n19518 );
and ( n22175 , n21302 , n19516 );
nor ( n22176 , n22174 , n22175 );
xnor ( n22177 , n22176 , n19489 );
and ( n22178 , n22172 , n22177 );
and ( n22179 , n22168 , n22177 );
or ( n22180 , n22173 , n22178 , n22179 );
and ( n22181 , n20268 , n20114 );
and ( n22182 , n20182 , n20112 );
nor ( n22183 , n22181 , n22182 );
xnor ( n22184 , n22183 , n19997 );
and ( n22185 , n20452 , n19894 );
and ( n22186 , n20360 , n19892 );
nor ( n22187 , n22185 , n22186 );
xnor ( n22188 , n22187 , n19858 );
and ( n22189 , n22184 , n22188 );
and ( n22190 , n20666 , n19805 );
and ( n22191 , n20618 , n19803 );
nor ( n22192 , n22190 , n22191 );
xnor ( n22193 , n22192 , n19750 );
and ( n22194 , n22188 , n22193 );
and ( n22195 , n22184 , n22193 );
or ( n22196 , n22189 , n22194 , n22195 );
and ( n22197 , n22180 , n22196 );
buf ( n22198 , n19316 );
and ( n22199 , n22198 , n19419 );
buf ( n22200 , n22199 );
and ( n22201 , n21704 , n19459 );
and ( n22202 , n21612 , n19457 );
nor ( n22203 , n22201 , n22202 );
xnor ( n22204 , n22203 , n19416 );
and ( n22205 , n22200 , n22204 );
and ( n22206 , n21955 , n19424 );
and ( n22207 , n21876 , n19422 );
nor ( n22208 , n22206 , n22207 );
xnor ( n22209 , n22208 , n19431 );
and ( n22210 , n22204 , n22209 );
and ( n22211 , n22200 , n22209 );
or ( n22212 , n22205 , n22210 , n22211 );
and ( n22213 , n22196 , n22212 );
and ( n22214 , n22180 , n22212 );
or ( n22215 , n22197 , n22213 , n22214 );
xor ( n22216 , n21941 , n21945 );
xor ( n22217 , n22216 , n21950 );
and ( n22218 , n22215 , n22217 );
xor ( n22219 , n21957 , n21961 );
xor ( n22220 , n22219 , n21966 );
and ( n22221 , n22217 , n22220 );
and ( n22222 , n22215 , n22220 );
or ( n22223 , n22218 , n22221 , n22222 );
buf ( n22224 , n19380 );
buf ( n22225 , n19381 );
and ( n22226 , n22224 , n22225 );
not ( n22227 , n22226 );
and ( n22228 , n21850 , n22227 );
not ( n22229 , n22228 );
and ( n22230 , n20080 , n20276 );
and ( n22231 , n20004 , n20274 );
nor ( n22232 , n22230 , n22231 );
xnor ( n22233 , n22232 , n20175 );
and ( n22234 , n22229 , n22233 );
buf ( n22235 , n19315 );
and ( n22236 , n22235 , n19419 );
and ( n22237 , n22233 , n22236 );
and ( n22238 , n22229 , n22236 );
or ( n22239 , n22234 , n22237 , n22238 );
and ( n22240 , n19496 , n21468 );
and ( n22241 , n19469 , n21466 );
nor ( n22242 , n22240 , n22241 );
xnor ( n22243 , n22242 , n21331 );
and ( n22244 , n22239 , n22243 );
and ( n22245 , n19881 , n20460 );
and ( n22246 , n19825 , n20458 );
nor ( n22247 , n22245 , n22246 );
xnor ( n22248 , n22247 , n20337 );
and ( n22249 , n22243 , n22248 );
and ( n22250 , n22239 , n22248 );
or ( n22251 , n22244 , n22249 , n22250 );
and ( n22252 , n19418 , n22048 );
and ( n22253 , n19426 , n22046 );
nor ( n22254 , n22252 , n22253 );
xnor ( n22255 , n22254 , n21853 );
and ( n22256 , n19510 , n21468 );
and ( n22257 , n19496 , n21466 );
nor ( n22258 , n22256 , n22257 );
xnor ( n22259 , n22258 , n21331 );
and ( n22260 , n22255 , n22259 );
and ( n22261 , n19946 , n20460 );
and ( n22262 , n19881 , n20458 );
nor ( n22263 , n22261 , n22262 );
xnor ( n22264 , n22263 , n20337 );
and ( n22265 , n22259 , n22264 );
and ( n22266 , n22255 , n22264 );
or ( n22267 , n22260 , n22265 , n22266 );
and ( n22268 , n19469 , n21741 );
and ( n22269 , n19434 , n21739 );
nor ( n22270 , n22268 , n22269 );
xnor ( n22271 , n22270 , n21605 );
and ( n22272 , n19605 , n21155 );
and ( n22273 , n19588 , n21153 );
nor ( n22274 , n22272 , n22273 );
xnor ( n22275 , n22274 , n20994 );
and ( n22276 , n22271 , n22275 );
and ( n22277 , n19721 , n20955 );
and ( n22278 , n19637 , n20953 );
nor ( n22279 , n22277 , n22278 );
xnor ( n22280 , n22279 , n20780 );
and ( n22281 , n22275 , n22280 );
and ( n22282 , n22271 , n22280 );
or ( n22283 , n22276 , n22281 , n22282 );
and ( n22284 , n22267 , n22283 );
xor ( n22285 , n22100 , n22104 );
xor ( n22286 , n22285 , n22109 );
and ( n22287 , n22283 , n22286 );
and ( n22288 , n22267 , n22286 );
or ( n22289 , n22284 , n22287 , n22288 );
and ( n22290 , n22251 , n22289 );
xor ( n22291 , n22112 , n22128 );
xor ( n22292 , n22291 , n22131 );
and ( n22293 , n22289 , n22292 );
and ( n22294 , n22251 , n22292 );
or ( n22295 , n22290 , n22293 , n22294 );
and ( n22296 , n22223 , n22295 );
xor ( n22297 , n21974 , n21976 );
xor ( n22298 , n22297 , n21979 );
and ( n22299 , n22295 , n22298 );
and ( n22300 , n22223 , n22298 );
or ( n22301 , n22296 , n22299 , n22300 );
xor ( n22302 , n22116 , n22120 );
xor ( n22303 , n22302 , n22125 );
xor ( n22304 , n22051 , n22055 );
xor ( n22305 , n22304 , n22060 );
and ( n22306 , n22303 , n22305 );
xor ( n22307 , n22084 , n22088 );
xor ( n22308 , n22307 , n22090 );
and ( n22309 , n22305 , n22308 );
and ( n22310 , n22303 , n22308 );
or ( n22311 , n22306 , n22309 , n22310 );
xor ( n22312 , n22063 , n22079 );
xor ( n22313 , n22312 , n22093 );
and ( n22314 , n22311 , n22313 );
xor ( n22315 , n22142 , n22144 );
xor ( n22316 , n22315 , n22147 );
and ( n22317 , n22313 , n22316 );
and ( n22318 , n22311 , n22316 );
or ( n22319 , n22314 , n22317 , n22318 );
xor ( n22320 , n22096 , n22134 );
xor ( n22321 , n22320 , n22137 );
and ( n22322 , n22319 , n22321 );
xor ( n22323 , n22150 , n22152 );
xor ( n22324 , n22323 , n22155 );
and ( n22325 , n22321 , n22324 );
and ( n22326 , n22319 , n22324 );
or ( n22327 , n22322 , n22325 , n22326 );
and ( n22328 , n22301 , n22327 );
xor ( n22329 , n22016 , n22018 );
xor ( n22330 , n22329 , n22021 );
and ( n22331 , n22327 , n22330 );
and ( n22332 , n22301 , n22330 );
or ( n22333 , n22328 , n22331 , n22332 );
and ( n22334 , n22164 , n22333 );
xor ( n22335 , n22024 , n22026 );
xor ( n22336 , n22335 , n22029 );
and ( n22337 , n22333 , n22336 );
and ( n22338 , n22164 , n22336 );
or ( n22339 , n22334 , n22337 , n22338 );
and ( n22340 , n22044 , n22339 );
xor ( n22341 , n22044 , n22339 );
xor ( n22342 , n22164 , n22333 );
xor ( n22343 , n22342 , n22336 );
and ( n22344 , n20182 , n20276 );
and ( n22345 , n20080 , n20274 );
nor ( n22346 , n22344 , n22345 );
xnor ( n22347 , n22346 , n20175 );
and ( n22348 , n21876 , n19459 );
and ( n22349 , n21704 , n19457 );
nor ( n22350 , n22348 , n22349 );
xnor ( n22351 , n22350 , n19416 );
and ( n22352 , n22347 , n22351 );
and ( n22353 , n22235 , n19424 );
and ( n22354 , n21955 , n19422 );
nor ( n22355 , n22353 , n22354 );
xnor ( n22356 , n22355 , n19431 );
and ( n22357 , n22351 , n22356 );
and ( n22358 , n22347 , n22356 );
or ( n22359 , n22352 , n22357 , n22358 );
and ( n22360 , n19825 , n20674 );
and ( n22361 , n19811 , n20672 );
nor ( n22362 , n22360 , n22361 );
xnor ( n22363 , n22362 , n20542 );
and ( n22364 , n22359 , n22363 );
xor ( n22365 , n22229 , n22233 );
xor ( n22366 , n22365 , n22236 );
and ( n22367 , n22363 , n22366 );
and ( n22368 , n22359 , n22366 );
or ( n22369 , n22364 , n22367 , n22368 );
xor ( n22370 , n22067 , n22071 );
xor ( n22371 , n22370 , n22076 );
and ( n22372 , n22369 , n22371 );
xor ( n22373 , n22239 , n22243 );
xor ( n22374 , n22373 , n22248 );
and ( n22375 , n22371 , n22374 );
and ( n22376 , n22369 , n22374 );
or ( n22377 , n22372 , n22375 , n22376 );
xor ( n22378 , n21850 , n22224 );
xor ( n22379 , n22224 , n22225 );
not ( n22380 , n22379 );
and ( n22381 , n22378 , n22380 );
and ( n22382 , n19426 , n22381 );
not ( n22383 , n22382 );
xnor ( n22384 , n22383 , n22228 );
and ( n22385 , n19496 , n21741 );
and ( n22386 , n19469 , n21739 );
nor ( n22387 , n22385 , n22386 );
xnor ( n22388 , n22387 , n21605 );
and ( n22389 , n22384 , n22388 );
and ( n22390 , n19811 , n20955 );
and ( n22391 , n19721 , n20953 );
nor ( n22392 , n22390 , n22391 );
xnor ( n22393 , n22392 , n20780 );
and ( n22394 , n22388 , n22393 );
and ( n22395 , n22384 , n22393 );
or ( n22396 , n22389 , n22394 , n22395 );
and ( n22397 , n19434 , n22048 );
and ( n22398 , n19418 , n22046 );
nor ( n22399 , n22397 , n22398 );
xnor ( n22400 , n22399 , n21853 );
and ( n22401 , n20004 , n20460 );
and ( n22402 , n19946 , n20458 );
nor ( n22403 , n22401 , n22402 );
xnor ( n22404 , n22403 , n20337 );
and ( n22405 , n22400 , n22404 );
and ( n22406 , n21612 , n19518 );
and ( n22407 , n21451 , n19516 );
nor ( n22408 , n22406 , n22407 );
xnor ( n22409 , n22408 , n19489 );
and ( n22410 , n22404 , n22409 );
and ( n22411 , n22400 , n22409 );
or ( n22412 , n22405 , n22410 , n22411 );
and ( n22413 , n22396 , n22412 );
buf ( n22414 , n19382 );
buf ( n22415 , n19383 );
and ( n22416 , n22414 , n22415 );
not ( n22417 , n22416 );
and ( n22418 , n22225 , n22417 );
not ( n22419 , n22418 );
and ( n22420 , n22198 , n19424 );
and ( n22421 , n22235 , n19422 );
nor ( n22422 , n22420 , n22421 );
xnor ( n22423 , n22422 , n19431 );
and ( n22424 , n22419 , n22423 );
buf ( n22425 , n19317 );
and ( n22426 , n22425 , n19419 );
and ( n22427 , n22423 , n22426 );
and ( n22428 , n22419 , n22426 );
or ( n22429 , n22424 , n22427 , n22428 );
and ( n22430 , n19588 , n21468 );
and ( n22431 , n19510 , n21466 );
nor ( n22432 , n22430 , n22431 );
xnor ( n22433 , n22432 , n21331 );
and ( n22434 , n22429 , n22433 );
and ( n22435 , n19637 , n21155 );
and ( n22436 , n19605 , n21153 );
nor ( n22437 , n22435 , n22436 );
xnor ( n22438 , n22437 , n20994 );
and ( n22439 , n22433 , n22438 );
and ( n22440 , n22429 , n22438 );
or ( n22441 , n22434 , n22439 , n22440 );
and ( n22442 , n22412 , n22441 );
and ( n22443 , n22396 , n22441 );
or ( n22444 , n22413 , n22442 , n22443 );
and ( n22445 , n20803 , n19805 );
and ( n22446 , n20666 , n19803 );
nor ( n22447 , n22445 , n22446 );
xnor ( n22448 , n22447 , n19750 );
and ( n22449 , n21072 , n19688 );
and ( n22450 , n20867 , n19686 );
nor ( n22451 , n22449 , n22450 );
xnor ( n22452 , n22451 , n19655 );
and ( n22453 , n22448 , n22452 );
and ( n22454 , n21302 , n19596 );
and ( n22455 , n21218 , n19594 );
nor ( n22456 , n22454 , n22455 );
xnor ( n22457 , n22456 , n19545 );
and ( n22458 , n22452 , n22457 );
and ( n22459 , n22448 , n22457 );
or ( n22460 , n22453 , n22458 , n22459 );
and ( n22461 , n20360 , n20114 );
and ( n22462 , n20268 , n20112 );
nor ( n22463 , n22461 , n22462 );
xnor ( n22464 , n22463 , n19997 );
and ( n22465 , n20618 , n19894 );
and ( n22466 , n20452 , n19892 );
nor ( n22467 , n22465 , n22466 );
xnor ( n22468 , n22467 , n19858 );
and ( n22469 , n22464 , n22468 );
not ( n22470 , n22199 );
and ( n22471 , n22468 , n22470 );
and ( n22472 , n22464 , n22470 );
or ( n22473 , n22469 , n22471 , n22472 );
and ( n22474 , n22460 , n22473 );
xor ( n22475 , n22200 , n22204 );
xor ( n22476 , n22475 , n22209 );
and ( n22477 , n22473 , n22476 );
and ( n22478 , n22460 , n22476 );
or ( n22479 , n22474 , n22477 , n22478 );
and ( n22480 , n22444 , n22479 );
xor ( n22481 , n22180 , n22196 );
xor ( n22482 , n22481 , n22212 );
and ( n22483 , n22479 , n22482 );
and ( n22484 , n22444 , n22482 );
or ( n22485 , n22480 , n22483 , n22484 );
and ( n22486 , n22377 , n22485 );
xor ( n22487 , n22215 , n22217 );
xor ( n22488 , n22487 , n22220 );
and ( n22489 , n22485 , n22488 );
and ( n22490 , n22377 , n22488 );
or ( n22491 , n22486 , n22489 , n22490 );
xor ( n22492 , n22168 , n22172 );
xor ( n22493 , n22492 , n22177 );
xor ( n22494 , n22184 , n22188 );
xor ( n22495 , n22494 , n22193 );
and ( n22496 , n22493 , n22495 );
xor ( n22497 , n22271 , n22275 );
xor ( n22498 , n22497 , n22280 );
and ( n22499 , n22495 , n22498 );
and ( n22500 , n22493 , n22498 );
or ( n22501 , n22496 , n22499 , n22500 );
xor ( n22502 , n22303 , n22305 );
xor ( n22503 , n22502 , n22308 );
and ( n22504 , n22501 , n22503 );
xor ( n22505 , n22267 , n22283 );
xor ( n22506 , n22505 , n22286 );
and ( n22507 , n22503 , n22506 );
and ( n22508 , n22501 , n22506 );
or ( n22509 , n22504 , n22507 , n22508 );
xor ( n22510 , n22251 , n22289 );
xor ( n22511 , n22510 , n22292 );
and ( n22512 , n22509 , n22511 );
xor ( n22513 , n22311 , n22313 );
xor ( n22514 , n22513 , n22316 );
and ( n22515 , n22511 , n22514 );
and ( n22516 , n22509 , n22514 );
or ( n22517 , n22512 , n22515 , n22516 );
and ( n22518 , n22491 , n22517 );
xor ( n22519 , n22223 , n22295 );
xor ( n22520 , n22519 , n22298 );
and ( n22521 , n22517 , n22520 );
and ( n22522 , n22491 , n22520 );
or ( n22523 , n22518 , n22521 , n22522 );
xor ( n22524 , n22140 , n22158 );
xor ( n22525 , n22524 , n22161 );
and ( n22526 , n22523 , n22525 );
xor ( n22527 , n22301 , n22327 );
xor ( n22528 , n22527 , n22330 );
and ( n22529 , n22525 , n22528 );
and ( n22530 , n22523 , n22528 );
or ( n22531 , n22526 , n22529 , n22530 );
and ( n22532 , n22343 , n22531 );
xor ( n22533 , n22343 , n22531 );
xor ( n22534 , n22523 , n22525 );
xor ( n22535 , n22534 , n22528 );
and ( n22536 , n20080 , n20460 );
and ( n22537 , n20004 , n20458 );
nor ( n22538 , n22536 , n22537 );
xnor ( n22539 , n22538 , n20337 );
and ( n22540 , n21704 , n19518 );
and ( n22541 , n21612 , n19516 );
nor ( n22542 , n22540 , n22541 );
xnor ( n22543 , n22542 , n19489 );
and ( n22544 , n22539 , n22543 );
and ( n22545 , n21955 , n19459 );
and ( n22546 , n21876 , n19457 );
nor ( n22547 , n22545 , n22546 );
xnor ( n22548 , n22547 , n19416 );
and ( n22549 , n22543 , n22548 );
and ( n22550 , n22539 , n22548 );
or ( n22551 , n22544 , n22549 , n22550 );
and ( n22552 , n22425 , n19424 );
and ( n22553 , n22198 , n19422 );
nor ( n22554 , n22552 , n22553 );
xnor ( n22555 , n22554 , n19431 );
buf ( n22556 , n22555 );
and ( n22557 , n20268 , n20276 );
and ( n22558 , n20182 , n20274 );
nor ( n22559 , n22557 , n22558 );
xnor ( n22560 , n22559 , n20175 );
and ( n22561 , n22556 , n22560 );
and ( n22562 , n20452 , n20114 );
and ( n22563 , n20360 , n20112 );
nor ( n22564 , n22562 , n22563 );
xnor ( n22565 , n22564 , n19997 );
and ( n22566 , n22560 , n22565 );
and ( n22567 , n22556 , n22565 );
or ( n22568 , n22561 , n22566 , n22567 );
and ( n22569 , n22551 , n22568 );
and ( n22570 , n19881 , n20674 );
and ( n22571 , n19825 , n20672 );
nor ( n22572 , n22570 , n22571 );
xnor ( n22573 , n22572 , n20542 );
and ( n22574 , n22568 , n22573 );
and ( n22575 , n22551 , n22573 );
or ( n22576 , n22569 , n22574 , n22575 );
and ( n22577 , n19510 , n21741 );
and ( n22578 , n19496 , n21739 );
nor ( n22579 , n22577 , n22578 );
xnor ( n22580 , n22579 , n21605 );
and ( n22581 , n19605 , n21468 );
and ( n22582 , n19588 , n21466 );
nor ( n22583 , n22581 , n22582 );
xnor ( n22584 , n22583 , n21331 );
and ( n22585 , n22580 , n22584 );
and ( n22586 , n19721 , n21155 );
and ( n22587 , n19637 , n21153 );
nor ( n22588 , n22586 , n22587 );
xnor ( n22589 , n22588 , n20994 );
and ( n22590 , n22584 , n22589 );
and ( n22591 , n22580 , n22589 );
or ( n22592 , n22585 , n22590 , n22591 );
and ( n22593 , n19418 , n22381 );
and ( n22594 , n19426 , n22379 );
nor ( n22595 , n22593 , n22594 );
xnor ( n22596 , n22595 , n22228 );
and ( n22597 , n19946 , n20674 );
and ( n22598 , n19881 , n20672 );
nor ( n22599 , n22597 , n22598 );
xnor ( n22600 , n22599 , n20542 );
and ( n22601 , n22596 , n22600 );
and ( n22602 , n21451 , n19596 );
and ( n22603 , n21302 , n19594 );
nor ( n22604 , n22602 , n22603 );
xnor ( n22605 , n22604 , n19545 );
and ( n22606 , n22600 , n22605 );
and ( n22607 , n22596 , n22605 );
or ( n22608 , n22601 , n22606 , n22607 );
and ( n22609 , n22592 , n22608 );
xor ( n22610 , n22448 , n22452 );
xor ( n22611 , n22610 , n22457 );
and ( n22612 , n22608 , n22611 );
and ( n22613 , n22592 , n22611 );
or ( n22614 , n22609 , n22612 , n22613 );
and ( n22615 , n22576 , n22614 );
xor ( n22616 , n22255 , n22259 );
xor ( n22617 , n22616 , n22264 );
and ( n22618 , n22614 , n22617 );
and ( n22619 , n22576 , n22617 );
or ( n22620 , n22615 , n22618 , n22619 );
and ( n22621 , n20666 , n19894 );
and ( n22622 , n20618 , n19892 );
nor ( n22623 , n22621 , n22622 );
xnor ( n22624 , n22623 , n19858 );
and ( n22625 , n20867 , n19805 );
and ( n22626 , n20803 , n19803 );
nor ( n22627 , n22625 , n22626 );
xnor ( n22628 , n22627 , n19750 );
and ( n22629 , n22624 , n22628 );
and ( n22630 , n21218 , n19688 );
and ( n22631 , n21072 , n19686 );
nor ( n22632 , n22630 , n22631 );
xnor ( n22633 , n22632 , n19655 );
and ( n22634 , n22628 , n22633 );
and ( n22635 , n22624 , n22633 );
or ( n22636 , n22629 , n22634 , n22635 );
xor ( n22637 , n22347 , n22351 );
xor ( n22638 , n22637 , n22356 );
and ( n22639 , n22636 , n22638 );
xor ( n22640 , n22464 , n22468 );
xor ( n22641 , n22640 , n22470 );
and ( n22642 , n22638 , n22641 );
and ( n22643 , n22636 , n22641 );
or ( n22644 , n22639 , n22642 , n22643 );
xor ( n22645 , n22359 , n22363 );
xor ( n22646 , n22645 , n22366 );
and ( n22647 , n22644 , n22646 );
xor ( n22648 , n22460 , n22473 );
xor ( n22649 , n22648 , n22476 );
and ( n22650 , n22646 , n22649 );
and ( n22651 , n22644 , n22649 );
or ( n22652 , n22647 , n22650 , n22651 );
and ( n22653 , n22620 , n22652 );
xor ( n22654 , n22369 , n22371 );
xor ( n22655 , n22654 , n22374 );
and ( n22656 , n22652 , n22655 );
and ( n22657 , n22620 , n22655 );
or ( n22658 , n22653 , n22656 , n22657 );
xor ( n22659 , n22377 , n22485 );
xor ( n22660 , n22659 , n22488 );
and ( n22661 , n22658 , n22660 );
xor ( n22662 , n22509 , n22511 );
xor ( n22663 , n22662 , n22514 );
and ( n22664 , n22660 , n22663 );
and ( n22665 , n22658 , n22663 );
or ( n22666 , n22661 , n22664 , n22665 );
xor ( n22667 , n22319 , n22321 );
xor ( n22668 , n22667 , n22324 );
and ( n22669 , n22666 , n22668 );
xor ( n22670 , n22491 , n22517 );
xor ( n22671 , n22670 , n22520 );
and ( n22672 , n22668 , n22671 );
and ( n22673 , n22666 , n22671 );
or ( n22674 , n22669 , n22672 , n22673 );
and ( n22675 , n22535 , n22674 );
xor ( n22676 , n22535 , n22674 );
xor ( n22677 , n22666 , n22668 );
xor ( n22678 , n22677 , n22671 );
and ( n22679 , n19469 , n22048 );
and ( n22680 , n19434 , n22046 );
nor ( n22681 , n22679 , n22680 );
xnor ( n22682 , n22681 , n21853 );
and ( n22683 , n19825 , n20955 );
and ( n22684 , n19811 , n20953 );
nor ( n22685 , n22683 , n22684 );
xnor ( n22686 , n22685 , n20780 );
and ( n22687 , n22682 , n22686 );
xor ( n22688 , n22419 , n22423 );
xor ( n22689 , n22688 , n22426 );
and ( n22690 , n22686 , n22689 );
and ( n22691 , n22682 , n22689 );
or ( n22692 , n22687 , n22690 , n22691 );
xor ( n22693 , n22384 , n22388 );
xor ( n22694 , n22693 , n22393 );
and ( n22695 , n22692 , n22694 );
xor ( n22696 , n22400 , n22404 );
xor ( n22697 , n22696 , n22409 );
and ( n22698 , n22694 , n22697 );
and ( n22699 , n22692 , n22697 );
or ( n22700 , n22695 , n22698 , n22699 );
xor ( n22701 , n22396 , n22412 );
xor ( n22702 , n22701 , n22441 );
and ( n22703 , n22700 , n22702 );
xor ( n22704 , n22493 , n22495 );
xor ( n22705 , n22704 , n22498 );
and ( n22706 , n22702 , n22705 );
and ( n22707 , n22700 , n22705 );
or ( n22708 , n22703 , n22706 , n22707 );
xor ( n22709 , n22444 , n22479 );
xor ( n22710 , n22709 , n22482 );
and ( n22711 , n22708 , n22710 );
xor ( n22712 , n22501 , n22503 );
xor ( n22713 , n22712 , n22506 );
and ( n22714 , n22710 , n22713 );
and ( n22715 , n22708 , n22713 );
or ( n22716 , n22711 , n22714 , n22715 );
and ( n22717 , n20182 , n20460 );
and ( n22718 , n20080 , n20458 );
nor ( n22719 , n22717 , n22718 );
xnor ( n22720 , n22719 , n20337 );
and ( n22721 , n20360 , n20276 );
and ( n22722 , n20268 , n20274 );
nor ( n22723 , n22721 , n22722 );
xnor ( n22724 , n22723 , n20175 );
and ( n22725 , n22720 , n22724 );
and ( n22726 , n21876 , n19518 );
and ( n22727 , n21704 , n19516 );
nor ( n22728 , n22726 , n22727 );
xnor ( n22729 , n22728 , n19489 );
and ( n22730 , n22724 , n22729 );
and ( n22731 , n22720 , n22729 );
or ( n22732 , n22725 , n22730 , n22731 );
and ( n22733 , n20618 , n20114 );
and ( n22734 , n20452 , n20112 );
nor ( n22735 , n22733 , n22734 );
xnor ( n22736 , n22735 , n19997 );
and ( n22737 , n20803 , n19894 );
and ( n22738 , n20666 , n19892 );
nor ( n22739 , n22737 , n22738 );
xnor ( n22740 , n22739 , n19858 );
and ( n22741 , n22736 , n22740 );
and ( n22742 , n21072 , n19805 );
and ( n22743 , n20867 , n19803 );
nor ( n22744 , n22742 , n22743 );
xnor ( n22745 , n22744 , n19750 );
and ( n22746 , n22740 , n22745 );
and ( n22747 , n22736 , n22745 );
or ( n22748 , n22741 , n22746 , n22747 );
and ( n22749 , n22732 , n22748 );
and ( n22750 , n22235 , n19459 );
and ( n22751 , n21955 , n19457 );
nor ( n22752 , n22750 , n22751 );
xnor ( n22753 , n22752 , n19416 );
not ( n22754 , n22555 );
and ( n22755 , n22753 , n22754 );
buf ( n22756 , n19318 );
and ( n22757 , n22756 , n19419 );
and ( n22758 , n22754 , n22757 );
and ( n22759 , n22753 , n22757 );
or ( n22760 , n22755 , n22758 , n22759 );
and ( n22761 , n22748 , n22760 );
and ( n22762 , n22732 , n22760 );
or ( n22763 , n22749 , n22761 , n22762 );
xor ( n22764 , n22429 , n22433 );
xor ( n22765 , n22764 , n22438 );
and ( n22766 , n22763 , n22765 );
xor ( n22767 , n22551 , n22568 );
xor ( n22768 , n22767 , n22573 );
and ( n22769 , n22765 , n22768 );
and ( n22770 , n22763 , n22768 );
or ( n22771 , n22766 , n22769 , n22770 );
xor ( n22772 , n22576 , n22614 );
xor ( n22773 , n22772 , n22617 );
and ( n22774 , n22771 , n22773 );
xor ( n22775 , n22644 , n22646 );
xor ( n22776 , n22775 , n22649 );
and ( n22777 , n22773 , n22776 );
and ( n22778 , n22771 , n22776 );
or ( n22779 , n22774 , n22777 , n22778 );
xor ( n22780 , n22620 , n22652 );
xor ( n22781 , n22780 , n22655 );
and ( n22782 , n22779 , n22781 );
xor ( n22783 , n22708 , n22710 );
xor ( n22784 , n22783 , n22713 );
and ( n22785 , n22781 , n22784 );
and ( n22786 , n22779 , n22784 );
or ( n22787 , n22782 , n22785 , n22786 );
and ( n22788 , n22716 , n22787 );
xor ( n22789 , n22658 , n22660 );
xor ( n22790 , n22789 , n22663 );
and ( n22791 , n22787 , n22790 );
and ( n22792 , n22716 , n22790 );
or ( n22793 , n22788 , n22791 , n22792 );
and ( n22794 , n22678 , n22793 );
xor ( n22795 , n22678 , n22793 );
xor ( n22796 , n22716 , n22787 );
xor ( n22797 , n22796 , n22790 );
and ( n22798 , n20004 , n20674 );
and ( n22799 , n19946 , n20672 );
nor ( n22800 , n22798 , n22799 );
xnor ( n22801 , n22800 , n20542 );
and ( n22802 , n21302 , n19688 );
and ( n22803 , n21218 , n19686 );
nor ( n22804 , n22802 , n22803 );
xnor ( n22805 , n22804 , n19655 );
and ( n22806 , n22801 , n22805 );
and ( n22807 , n21612 , n19596 );
and ( n22808 , n21451 , n19594 );
nor ( n22809 , n22807 , n22808 );
xnor ( n22810 , n22809 , n19545 );
and ( n22811 , n22805 , n22810 );
and ( n22812 , n22801 , n22810 );
or ( n22813 , n22806 , n22811 , n22812 );
xor ( n22814 , n22539 , n22543 );
xor ( n22815 , n22814 , n22548 );
and ( n22816 , n22813 , n22815 );
xor ( n22817 , n22556 , n22560 );
xor ( n22818 , n22817 , n22565 );
and ( n22819 , n22815 , n22818 );
and ( n22820 , n22813 , n22818 );
or ( n22821 , n22816 , n22819 , n22820 );
and ( n22822 , n19434 , n22381 );
and ( n22823 , n19418 , n22379 );
nor ( n22824 , n22822 , n22823 );
xnor ( n22825 , n22824 , n22228 );
and ( n22826 , n19588 , n21741 );
and ( n22827 , n19510 , n21739 );
nor ( n22828 , n22826 , n22827 );
xnor ( n22829 , n22828 , n21605 );
and ( n22830 , n22825 , n22829 );
and ( n22831 , n19637 , n21468 );
and ( n22832 , n19605 , n21466 );
nor ( n22833 , n22831 , n22832 );
xnor ( n22834 , n22833 , n21331 );
and ( n22835 , n22829 , n22834 );
and ( n22836 , n22825 , n22834 );
or ( n22837 , n22830 , n22835 , n22836 );
buf ( n22838 , n19384 );
buf ( n22839 , n19385 );
and ( n22840 , n22838 , n22839 );
not ( n22841 , n22840 );
and ( n22842 , n22415 , n22841 );
not ( n22843 , n22842 );
and ( n22844 , n22198 , n19459 );
and ( n22845 , n22235 , n19457 );
nor ( n22846 , n22844 , n22845 );
xnor ( n22847 , n22846 , n19416 );
and ( n22848 , n22843 , n22847 );
and ( n22849 , n22756 , n19424 );
and ( n22850 , n22425 , n19422 );
nor ( n22851 , n22849 , n22850 );
xnor ( n22852 , n22851 , n19431 );
and ( n22853 , n22847 , n22852 );
and ( n22854 , n22843 , n22852 );
or ( n22855 , n22848 , n22853 , n22854 );
xor ( n22856 , n22225 , n22414 );
xor ( n22857 , n22414 , n22415 );
not ( n22858 , n22857 );
and ( n22859 , n22856 , n22858 );
and ( n22860 , n19426 , n22859 );
not ( n22861 , n22860 );
xnor ( n22862 , n22861 , n22418 );
and ( n22863 , n22855 , n22862 );
and ( n22864 , n19811 , n21155 );
and ( n22865 , n19721 , n21153 );
nor ( n22866 , n22864 , n22865 );
xnor ( n22867 , n22866 , n20994 );
and ( n22868 , n22862 , n22867 );
and ( n22869 , n22855 , n22867 );
or ( n22870 , n22863 , n22868 , n22869 );
and ( n22871 , n22837 , n22870 );
xor ( n22872 , n22624 , n22628 );
xor ( n22873 , n22872 , n22633 );
and ( n22874 , n22870 , n22873 );
and ( n22875 , n22837 , n22873 );
or ( n22876 , n22871 , n22874 , n22875 );
and ( n22877 , n22821 , n22876 );
xor ( n22878 , n22580 , n22584 );
xor ( n22879 , n22878 , n22589 );
xor ( n22880 , n22596 , n22600 );
xor ( n22881 , n22880 , n22605 );
and ( n22882 , n22879 , n22881 );
xor ( n22883 , n22682 , n22686 );
xor ( n22884 , n22883 , n22689 );
and ( n22885 , n22881 , n22884 );
and ( n22886 , n22879 , n22884 );
or ( n22887 , n22882 , n22885 , n22886 );
and ( n22888 , n22876 , n22887 );
and ( n22889 , n22821 , n22887 );
or ( n22890 , n22877 , n22888 , n22889 );
xor ( n22891 , n22636 , n22638 );
xor ( n22892 , n22891 , n22641 );
xor ( n22893 , n22592 , n22608 );
xor ( n22894 , n22893 , n22611 );
and ( n22895 , n22892 , n22894 );
xor ( n22896 , n22692 , n22694 );
xor ( n22897 , n22896 , n22697 );
and ( n22898 , n22894 , n22897 );
and ( n22899 , n22892 , n22897 );
or ( n22900 , n22895 , n22898 , n22899 );
and ( n22901 , n22890 , n22900 );
xor ( n22902 , n22700 , n22702 );
xor ( n22903 , n22902 , n22705 );
and ( n22904 , n22900 , n22903 );
and ( n22905 , n22890 , n22903 );
or ( n22906 , n22901 , n22904 , n22905 );
and ( n22907 , n20080 , n20674 );
and ( n22908 , n20004 , n20672 );
nor ( n22909 , n22907 , n22908 );
xnor ( n22910 , n22909 , n20542 );
and ( n22911 , n21955 , n19518 );
and ( n22912 , n21876 , n19516 );
nor ( n22913 , n22911 , n22912 );
xnor ( n22914 , n22913 , n19489 );
and ( n22915 , n22910 , n22914 );
buf ( n22916 , n19319 );
and ( n22917 , n22916 , n19419 );
and ( n22918 , n22914 , n22917 );
and ( n22919 , n22910 , n22917 );
or ( n22920 , n22915 , n22918 , n22919 );
and ( n22921 , n20452 , n20276 );
and ( n22922 , n20360 , n20274 );
nor ( n22923 , n22921 , n22922 );
xnor ( n22924 , n22923 , n20175 );
and ( n22925 , n20666 , n20114 );
and ( n22926 , n20618 , n20112 );
nor ( n22927 , n22925 , n22926 );
xnor ( n22928 , n22927 , n19997 );
and ( n22929 , n22924 , n22928 );
and ( n22930 , n20867 , n19894 );
and ( n22931 , n20803 , n19892 );
nor ( n22932 , n22930 , n22931 );
xnor ( n22933 , n22932 , n19858 );
and ( n22934 , n22928 , n22933 );
and ( n22935 , n22924 , n22933 );
or ( n22936 , n22929 , n22934 , n22935 );
and ( n22937 , n22920 , n22936 );
and ( n22938 , n22425 , n19459 );
and ( n22939 , n22198 , n19457 );
nor ( n22940 , n22938 , n22939 );
xnor ( n22941 , n22940 , n19416 );
buf ( n22942 , n22941 );
and ( n22943 , n20268 , n20460 );
and ( n22944 , n20182 , n20458 );
nor ( n22945 , n22943 , n22944 );
xnor ( n22946 , n22945 , n20337 );
and ( n22947 , n22942 , n22946 );
and ( n22948 , n21704 , n19596 );
and ( n22949 , n21612 , n19594 );
nor ( n22950 , n22948 , n22949 );
xnor ( n22951 , n22950 , n19545 );
and ( n22952 , n22946 , n22951 );
and ( n22953 , n22942 , n22951 );
or ( n22954 , n22947 , n22952 , n22953 );
and ( n22955 , n22936 , n22954 );
and ( n22956 , n22920 , n22954 );
or ( n22957 , n22937 , n22955 , n22956 );
and ( n22958 , n19496 , n22048 );
and ( n22959 , n19469 , n22046 );
nor ( n22960 , n22958 , n22959 );
xnor ( n22961 , n22960 , n21853 );
and ( n22962 , n19881 , n20955 );
and ( n22963 , n19825 , n20953 );
nor ( n22964 , n22962 , n22963 );
xnor ( n22965 , n22964 , n20780 );
and ( n22966 , n22961 , n22965 );
xor ( n22967 , n22753 , n22754 );
xor ( n22968 , n22967 , n22757 );
and ( n22969 , n22965 , n22968 );
and ( n22970 , n22961 , n22968 );
or ( n22971 , n22966 , n22969 , n22970 );
and ( n22972 , n22957 , n22971 );
and ( n22973 , n19946 , n20955 );
and ( n22974 , n19881 , n20953 );
nor ( n22975 , n22973 , n22974 );
xnor ( n22976 , n22975 , n20780 );
and ( n22977 , n21218 , n19805 );
and ( n22978 , n21072 , n19803 );
nor ( n22979 , n22977 , n22978 );
xnor ( n22980 , n22979 , n19750 );
and ( n22981 , n22976 , n22980 );
and ( n22982 , n21451 , n19688 );
and ( n22983 , n21302 , n19686 );
nor ( n22984 , n22982 , n22983 );
xnor ( n22985 , n22984 , n19655 );
and ( n22986 , n22980 , n22985 );
and ( n22987 , n22976 , n22985 );
or ( n22988 , n22981 , n22986 , n22987 );
and ( n22989 , n19418 , n22859 );
and ( n22990 , n19426 , n22857 );
nor ( n22991 , n22989 , n22990 );
xnor ( n22992 , n22991 , n22418 );
and ( n22993 , n19510 , n22048 );
and ( n22994 , n19496 , n22046 );
nor ( n22995 , n22993 , n22994 );
xnor ( n22996 , n22995 , n21853 );
and ( n22997 , n22992 , n22996 );
and ( n22998 , n19605 , n21741 );
and ( n22999 , n19588 , n21739 );
nor ( n23000 , n22998 , n22999 );
xnor ( n23001 , n23000 , n21605 );
and ( n23002 , n22996 , n23001 );
and ( n23003 , n22992 , n23001 );
or ( n23004 , n22997 , n23002 , n23003 );
and ( n23005 , n22988 , n23004 );
xor ( n23006 , n22801 , n22805 );
xor ( n23007 , n23006 , n22810 );
and ( n23008 , n23004 , n23007 );
and ( n23009 , n22988 , n23007 );
or ( n23010 , n23005 , n23008 , n23009 );
and ( n23011 , n22971 , n23010 );
and ( n23012 , n22957 , n23010 );
or ( n23013 , n22972 , n23011 , n23012 );
and ( n23014 , n19469 , n22381 );
and ( n23015 , n19434 , n22379 );
nor ( n23016 , n23014 , n23015 );
xnor ( n23017 , n23016 , n22228 );
and ( n23018 , n19721 , n21468 );
and ( n23019 , n19637 , n21466 );
nor ( n23020 , n23018 , n23019 );
xnor ( n23021 , n23020 , n21331 );
and ( n23022 , n23017 , n23021 );
and ( n23023 , n19825 , n21155 );
and ( n23024 , n19811 , n21153 );
nor ( n23025 , n23023 , n23024 );
xnor ( n23026 , n23025 , n20994 );
and ( n23027 , n23021 , n23026 );
and ( n23028 , n23017 , n23026 );
or ( n23029 , n23022 , n23027 , n23028 );
xor ( n23030 , n22720 , n22724 );
xor ( n23031 , n23030 , n22729 );
and ( n23032 , n23029 , n23031 );
xor ( n23033 , n22736 , n22740 );
xor ( n23034 , n23033 , n22745 );
and ( n23035 , n23031 , n23034 );
and ( n23036 , n23029 , n23034 );
or ( n23037 , n23032 , n23035 , n23036 );
xor ( n23038 , n22732 , n22748 );
xor ( n23039 , n23038 , n22760 );
and ( n23040 , n23037 , n23039 );
xor ( n23041 , n22813 , n22815 );
xor ( n23042 , n23041 , n22818 );
and ( n23043 , n23039 , n23042 );
and ( n23044 , n23037 , n23042 );
or ( n23045 , n23040 , n23043 , n23044 );
and ( n23046 , n23013 , n23045 );
xor ( n23047 , n22763 , n22765 );
xor ( n23048 , n23047 , n22768 );
and ( n23049 , n23045 , n23048 );
and ( n23050 , n23013 , n23048 );
or ( n23051 , n23046 , n23049 , n23050 );
xor ( n23052 , n22825 , n22829 );
xor ( n23053 , n23052 , n22834 );
xor ( n23054 , n22855 , n22862 );
xor ( n23055 , n23054 , n22867 );
and ( n23056 , n23053 , n23055 );
xor ( n23057 , n22961 , n22965 );
xor ( n23058 , n23057 , n22968 );
and ( n23059 , n23055 , n23058 );
and ( n23060 , n23053 , n23058 );
or ( n23061 , n23056 , n23059 , n23060 );
xor ( n23062 , n22837 , n22870 );
xor ( n23063 , n23062 , n22873 );
and ( n23064 , n23061 , n23063 );
xor ( n23065 , n22879 , n22881 );
xor ( n23066 , n23065 , n22884 );
and ( n23067 , n23063 , n23066 );
and ( n23068 , n23061 , n23066 );
or ( n23069 , n23064 , n23067 , n23068 );
xor ( n23070 , n22821 , n22876 );
xor ( n23071 , n23070 , n22887 );
and ( n23072 , n23069 , n23071 );
xor ( n23073 , n22892 , n22894 );
xor ( n23074 , n23073 , n22897 );
and ( n23075 , n23071 , n23074 );
and ( n23076 , n23069 , n23074 );
or ( n23077 , n23072 , n23075 , n23076 );
and ( n23078 , n23051 , n23077 );
xor ( n23079 , n22771 , n22773 );
xor ( n23080 , n23079 , n22776 );
and ( n23081 , n23077 , n23080 );
and ( n23082 , n23051 , n23080 );
or ( n23083 , n23078 , n23081 , n23082 );
and ( n23084 , n22906 , n23083 );
xor ( n23085 , n22779 , n22781 );
xor ( n23086 , n23085 , n22784 );
and ( n23087 , n23083 , n23086 );
and ( n23088 , n22906 , n23086 );
or ( n23089 , n23084 , n23087 , n23088 );
and ( n23090 , n22797 , n23089 );
xor ( n23091 , n22797 , n23089 );
xor ( n23092 , n22906 , n23083 );
xor ( n23093 , n23092 , n23086 );
and ( n23094 , n19496 , n22381 );
and ( n23095 , n19469 , n22379 );
nor ( n23096 , n23094 , n23095 );
xnor ( n23097 , n23096 , n22228 );
and ( n23098 , n19811 , n21468 );
and ( n23099 , n19721 , n21466 );
nor ( n23100 , n23098 , n23099 );
xnor ( n23101 , n23100 , n21331 );
and ( n23102 , n23097 , n23101 );
and ( n23103 , n19881 , n21155 );
and ( n23104 , n19825 , n21153 );
nor ( n23105 , n23103 , n23104 );
xnor ( n23106 , n23105 , n20994 );
and ( n23107 , n23101 , n23106 );
and ( n23108 , n23097 , n23106 );
or ( n23109 , n23102 , n23107 , n23108 );
and ( n23110 , n19434 , n22859 );
and ( n23111 , n19418 , n22857 );
nor ( n23112 , n23110 , n23111 );
xnor ( n23113 , n23112 , n22418 );
and ( n23114 , n19588 , n22048 );
and ( n23115 , n19510 , n22046 );
nor ( n23116 , n23114 , n23115 );
xnor ( n23117 , n23116 , n21853 );
and ( n23118 , n23113 , n23117 );
and ( n23119 , n20004 , n20955 );
and ( n23120 , n19946 , n20953 );
nor ( n23121 , n23119 , n23120 );
xnor ( n23122 , n23121 , n20780 );
and ( n23123 , n23117 , n23122 );
and ( n23124 , n23113 , n23122 );
or ( n23125 , n23118 , n23123 , n23124 );
and ( n23126 , n23109 , n23125 );
xor ( n23127 , n22976 , n22980 );
xor ( n23128 , n23127 , n22985 );
and ( n23129 , n23125 , n23128 );
and ( n23130 , n23109 , n23128 );
or ( n23131 , n23126 , n23129 , n23130 );
and ( n23132 , n22235 , n19518 );
and ( n23133 , n21955 , n19516 );
nor ( n23134 , n23132 , n23133 );
xnor ( n23135 , n23134 , n19489 );
and ( n23136 , n22916 , n19424 );
and ( n23137 , n22756 , n19422 );
nor ( n23138 , n23136 , n23137 );
xnor ( n23139 , n23138 , n19431 );
and ( n23140 , n23135 , n23139 );
buf ( n23141 , n19320 );
and ( n23142 , n23141 , n19419 );
and ( n23143 , n23139 , n23142 );
and ( n23144 , n23135 , n23142 );
or ( n23145 , n23140 , n23143 , n23144 );
and ( n23146 , n20182 , n20674 );
and ( n23147 , n20080 , n20672 );
nor ( n23148 , n23146 , n23147 );
xnor ( n23149 , n23148 , n20542 );
and ( n23150 , n20360 , n20460 );
and ( n23151 , n20268 , n20458 );
nor ( n23152 , n23150 , n23151 );
xnor ( n23153 , n23152 , n20337 );
and ( n23154 , n23149 , n23153 );
and ( n23155 , n21876 , n19596 );
and ( n23156 , n21704 , n19594 );
nor ( n23157 , n23155 , n23156 );
xnor ( n23158 , n23157 , n19545 );
and ( n23159 , n23153 , n23158 );
and ( n23160 , n23149 , n23158 );
or ( n23161 , n23154 , n23159 , n23160 );
and ( n23162 , n23145 , n23161 );
xor ( n23163 , n22843 , n22847 );
xor ( n23164 , n23163 , n22852 );
and ( n23165 , n23161 , n23164 );
and ( n23166 , n23145 , n23164 );
or ( n23167 , n23162 , n23165 , n23166 );
and ( n23168 , n23131 , n23167 );
xor ( n23169 , n22920 , n22936 );
xor ( n23170 , n23169 , n22954 );
and ( n23171 , n23167 , n23170 );
and ( n23172 , n23131 , n23170 );
or ( n23173 , n23168 , n23171 , n23172 );
and ( n23174 , n21072 , n19894 );
and ( n23175 , n20867 , n19892 );
nor ( n23176 , n23174 , n23175 );
xnor ( n23177 , n23176 , n19858 );
and ( n23178 , n21302 , n19805 );
and ( n23179 , n21218 , n19803 );
nor ( n23180 , n23178 , n23179 );
xnor ( n23181 , n23180 , n19750 );
and ( n23182 , n23177 , n23181 );
and ( n23183 , n21612 , n19688 );
and ( n23184 , n21451 , n19686 );
nor ( n23185 , n23183 , n23184 );
xnor ( n23186 , n23185 , n19655 );
and ( n23187 , n23181 , n23186 );
and ( n23188 , n23177 , n23186 );
or ( n23189 , n23182 , n23187 , n23188 );
and ( n23190 , n20618 , n20276 );
and ( n23191 , n20452 , n20274 );
nor ( n23192 , n23190 , n23191 );
xnor ( n23193 , n23192 , n20175 );
and ( n23194 , n20803 , n20114 );
and ( n23195 , n20666 , n20112 );
nor ( n23196 , n23194 , n23195 );
xnor ( n23197 , n23196 , n19997 );
and ( n23198 , n23193 , n23197 );
not ( n23199 , n22941 );
and ( n23200 , n23197 , n23199 );
and ( n23201 , n23193 , n23199 );
or ( n23202 , n23198 , n23200 , n23201 );
and ( n23203 , n23189 , n23202 );
xor ( n23204 , n22942 , n22946 );
xor ( n23205 , n23204 , n22951 );
and ( n23206 , n23202 , n23205 );
and ( n23207 , n23189 , n23205 );
or ( n23208 , n23203 , n23206 , n23207 );
buf ( n23209 , n19386 );
buf ( n23210 , n19387 );
and ( n23211 , n23209 , n23210 );
not ( n23212 , n23211 );
and ( n23213 , n22839 , n23212 );
not ( n23214 , n23213 );
and ( n23215 , n22198 , n19518 );
and ( n23216 , n22235 , n19516 );
nor ( n23217 , n23215 , n23216 );
xnor ( n23218 , n23217 , n19489 );
and ( n23219 , n23214 , n23218 );
and ( n23220 , n22756 , n19459 );
and ( n23221 , n22425 , n19457 );
nor ( n23222 , n23220 , n23221 );
xnor ( n23223 , n23222 , n19416 );
and ( n23224 , n23218 , n23223 );
and ( n23225 , n23214 , n23223 );
or ( n23226 , n23219 , n23224 , n23225 );
xor ( n23227 , n22415 , n22838 );
xor ( n23228 , n22838 , n22839 );
not ( n23229 , n23228 );
and ( n23230 , n23227 , n23229 );
and ( n23231 , n19426 , n23230 );
not ( n23232 , n23231 );
xnor ( n23233 , n23232 , n22842 );
and ( n23234 , n23226 , n23233 );
and ( n23235 , n19637 , n21741 );
and ( n23236 , n19605 , n21739 );
nor ( n23237 , n23235 , n23236 );
xnor ( n23238 , n23237 , n21605 );
and ( n23239 , n23233 , n23238 );
and ( n23240 , n23226 , n23238 );
or ( n23241 , n23234 , n23239 , n23240 );
xor ( n23242 , n22910 , n22914 );
xor ( n23243 , n23242 , n22917 );
and ( n23244 , n23241 , n23243 );
xor ( n23245 , n22924 , n22928 );
xor ( n23246 , n23245 , n22933 );
and ( n23247 , n23243 , n23246 );
and ( n23248 , n23241 , n23246 );
or ( n23249 , n23244 , n23247 , n23248 );
and ( n23250 , n23208 , n23249 );
xor ( n23251 , n22988 , n23004 );
xor ( n23252 , n23251 , n23007 );
and ( n23253 , n23249 , n23252 );
and ( n23254 , n23208 , n23252 );
or ( n23255 , n23250 , n23253 , n23254 );
and ( n23256 , n23173 , n23255 );
xor ( n23257 , n22957 , n22971 );
xor ( n23258 , n23257 , n23010 );
and ( n23259 , n23255 , n23258 );
and ( n23260 , n23173 , n23258 );
or ( n23261 , n23256 , n23259 , n23260 );
and ( n23262 , n21955 , n19596 );
and ( n23263 , n21876 , n19594 );
nor ( n23264 , n23262 , n23263 );
xnor ( n23265 , n23264 , n19545 );
and ( n23266 , n23141 , n19424 );
and ( n23267 , n22916 , n19422 );
nor ( n23268 , n23266 , n23267 );
xnor ( n23269 , n23268 , n19431 );
and ( n23270 , n23265 , n23269 );
buf ( n23271 , n19321 );
and ( n23272 , n23271 , n19419 );
and ( n23273 , n23269 , n23272 );
and ( n23274 , n23265 , n23272 );
or ( n23275 , n23270 , n23273 , n23274 );
and ( n23276 , n20080 , n20955 );
and ( n23277 , n20004 , n20953 );
nor ( n23278 , n23276 , n23277 );
xnor ( n23279 , n23278 , n20780 );
and ( n23280 , n20268 , n20674 );
and ( n23281 , n20182 , n20672 );
nor ( n23282 , n23280 , n23281 );
xnor ( n23283 , n23282 , n20542 );
and ( n23284 , n23279 , n23283 );
and ( n23285 , n21704 , n19688 );
and ( n23286 , n21612 , n19686 );
nor ( n23287 , n23285 , n23286 );
xnor ( n23288 , n23287 , n19655 );
and ( n23289 , n23283 , n23288 );
and ( n23290 , n23279 , n23288 );
or ( n23291 , n23284 , n23289 , n23290 );
and ( n23292 , n23275 , n23291 );
xor ( n23293 , n23135 , n23139 );
xor ( n23294 , n23293 , n23142 );
and ( n23295 , n23291 , n23294 );
and ( n23296 , n23275 , n23294 );
or ( n23297 , n23292 , n23295 , n23296 );
xor ( n23298 , n23017 , n23021 );
xor ( n23299 , n23298 , n23026 );
and ( n23300 , n23297 , n23299 );
xor ( n23301 , n22992 , n22996 );
xor ( n23302 , n23301 , n23001 );
and ( n23303 , n23299 , n23302 );
and ( n23304 , n23297 , n23302 );
or ( n23305 , n23300 , n23303 , n23304 );
xor ( n23306 , n23029 , n23031 );
xor ( n23307 , n23306 , n23034 );
and ( n23308 , n23305 , n23307 );
xor ( n23309 , n23053 , n23055 );
xor ( n23310 , n23309 , n23058 );
and ( n23311 , n23307 , n23310 );
and ( n23312 , n23305 , n23310 );
or ( n23313 , n23308 , n23311 , n23312 );
xor ( n23314 , n23037 , n23039 );
xor ( n23315 , n23314 , n23042 );
and ( n23316 , n23313 , n23315 );
xor ( n23317 , n23061 , n23063 );
xor ( n23318 , n23317 , n23066 );
and ( n23319 , n23315 , n23318 );
and ( n23320 , n23313 , n23318 );
or ( n23321 , n23316 , n23319 , n23320 );
and ( n23322 , n23261 , n23321 );
xor ( n23323 , n23013 , n23045 );
xor ( n23324 , n23323 , n23048 );
and ( n23325 , n23321 , n23324 );
and ( n23326 , n23261 , n23324 );
or ( n23327 , n23322 , n23325 , n23326 );
xor ( n23328 , n22890 , n22900 );
xor ( n23329 , n23328 , n22903 );
and ( n23330 , n23327 , n23329 );
xor ( n23331 , n23051 , n23077 );
xor ( n23332 , n23331 , n23080 );
and ( n23333 , n23329 , n23332 );
and ( n23334 , n23327 , n23332 );
or ( n23335 , n23330 , n23333 , n23334 );
and ( n23336 , n23093 , n23335 );
xor ( n23337 , n23093 , n23335 );
xor ( n23338 , n23327 , n23329 );
xor ( n23339 , n23338 , n23332 );
and ( n23340 , n19418 , n23230 );
and ( n23341 , n19426 , n23228 );
nor ( n23342 , n23340 , n23341 );
xnor ( n23343 , n23342 , n22842 );
and ( n23344 , n19510 , n22381 );
and ( n23345 , n19496 , n22379 );
nor ( n23346 , n23344 , n23345 );
xnor ( n23347 , n23346 , n22228 );
and ( n23348 , n23343 , n23347 );
and ( n23349 , n19946 , n21155 );
and ( n23350 , n19881 , n21153 );
nor ( n23351 , n23349 , n23350 );
xnor ( n23352 , n23351 , n20994 );
and ( n23353 , n23347 , n23352 );
and ( n23354 , n23343 , n23352 );
or ( n23355 , n23348 , n23353 , n23354 );
xor ( n23356 , n23149 , n23153 );
xor ( n23357 , n23356 , n23158 );
and ( n23358 , n23355 , n23357 );
xor ( n23359 , n23177 , n23181 );
xor ( n23360 , n23359 , n23186 );
and ( n23361 , n23357 , n23360 );
and ( n23362 , n23355 , n23360 );
or ( n23363 , n23358 , n23361 , n23362 );
xor ( n23364 , n23145 , n23161 );
xor ( n23365 , n23364 , n23164 );
and ( n23366 , n23363 , n23365 );
xor ( n23367 , n23189 , n23202 );
xor ( n23368 , n23367 , n23205 );
and ( n23369 , n23365 , n23368 );
and ( n23370 , n23363 , n23368 );
or ( n23371 , n23366 , n23369 , n23370 );
and ( n23372 , n22916 , n19459 );
and ( n23373 , n22756 , n19457 );
nor ( n23374 , n23372 , n23373 );
xnor ( n23375 , n23374 , n19416 );
and ( n23376 , n23271 , n19424 );
and ( n23377 , n23141 , n19422 );
nor ( n23378 , n23376 , n23377 );
xnor ( n23379 , n23378 , n19431 );
and ( n23380 , n23375 , n23379 );
buf ( n23381 , n19322 );
and ( n23382 , n23381 , n19419 );
and ( n23383 , n23379 , n23382 );
and ( n23384 , n23375 , n23382 );
or ( n23385 , n23380 , n23383 , n23384 );
and ( n23386 , n19605 , n22048 );
and ( n23387 , n19588 , n22046 );
nor ( n23388 , n23386 , n23387 );
xnor ( n23389 , n23388 , n21853 );
and ( n23390 , n23385 , n23389 );
and ( n23391 , n19721 , n21741 );
and ( n23392 , n19637 , n21739 );
nor ( n23393 , n23391 , n23392 );
xnor ( n23394 , n23393 , n21605 );
and ( n23395 , n23389 , n23394 );
and ( n23396 , n23385 , n23394 );
or ( n23397 , n23390 , n23395 , n23396 );
and ( n23398 , n19469 , n22859 );
and ( n23399 , n19434 , n22857 );
nor ( n23400 , n23398 , n23399 );
xnor ( n23401 , n23400 , n22418 );
and ( n23402 , n19825 , n21468 );
and ( n23403 , n19811 , n21466 );
nor ( n23404 , n23402 , n23403 );
xnor ( n23405 , n23404 , n21331 );
and ( n23406 , n23401 , n23405 );
xor ( n23407 , n23214 , n23218 );
xor ( n23408 , n23407 , n23223 );
and ( n23409 , n23405 , n23408 );
and ( n23410 , n23401 , n23408 );
or ( n23411 , n23406 , n23409 , n23410 );
and ( n23412 , n23397 , n23411 );
xor ( n23413 , n23097 , n23101 );
xor ( n23414 , n23413 , n23106 );
and ( n23415 , n23411 , n23414 );
and ( n23416 , n23397 , n23414 );
or ( n23417 , n23412 , n23415 , n23416 );
and ( n23418 , n20867 , n20114 );
and ( n23419 , n20803 , n20112 );
nor ( n23420 , n23418 , n23419 );
xnor ( n23421 , n23420 , n19997 );
and ( n23422 , n21218 , n19894 );
and ( n23423 , n21072 , n19892 );
nor ( n23424 , n23422 , n23423 );
xnor ( n23425 , n23424 , n19858 );
and ( n23426 , n23421 , n23425 );
and ( n23427 , n21451 , n19805 );
and ( n23428 , n21302 , n19803 );
nor ( n23429 , n23427 , n23428 );
xnor ( n23430 , n23429 , n19750 );
and ( n23431 , n23425 , n23430 );
and ( n23432 , n23421 , n23430 );
or ( n23433 , n23426 , n23431 , n23432 );
and ( n23434 , n22425 , n19518 );
and ( n23435 , n22198 , n19516 );
nor ( n23436 , n23434 , n23435 );
xnor ( n23437 , n23436 , n19489 );
buf ( n23438 , n23437 );
and ( n23439 , n20452 , n20460 );
and ( n23440 , n20360 , n20458 );
nor ( n23441 , n23439 , n23440 );
xnor ( n23442 , n23441 , n20337 );
and ( n23443 , n23438 , n23442 );
and ( n23444 , n20666 , n20276 );
and ( n23445 , n20618 , n20274 );
nor ( n23446 , n23444 , n23445 );
xnor ( n23447 , n23446 , n20175 );
and ( n23448 , n23442 , n23447 );
and ( n23449 , n23438 , n23447 );
or ( n23450 , n23443 , n23448 , n23449 );
and ( n23451 , n23433 , n23450 );
xor ( n23452 , n23193 , n23197 );
xor ( n23453 , n23452 , n23199 );
and ( n23454 , n23450 , n23453 );
and ( n23455 , n23433 , n23453 );
or ( n23456 , n23451 , n23454 , n23455 );
and ( n23457 , n23417 , n23456 );
xor ( n23458 , n23109 , n23125 );
xor ( n23459 , n23458 , n23128 );
and ( n23460 , n23456 , n23459 );
and ( n23461 , n23417 , n23459 );
or ( n23462 , n23457 , n23460 , n23461 );
and ( n23463 , n23371 , n23462 );
xor ( n23464 , n23131 , n23167 );
xor ( n23465 , n23464 , n23170 );
and ( n23466 , n23462 , n23465 );
and ( n23467 , n23371 , n23465 );
or ( n23468 , n23463 , n23466 , n23467 );
and ( n23469 , n20182 , n20955 );
and ( n23470 , n20080 , n20953 );
nor ( n23471 , n23469 , n23470 );
xnor ( n23472 , n23471 , n20780 );
and ( n23473 , n21876 , n19688 );
and ( n23474 , n21704 , n19686 );
nor ( n23475 , n23473 , n23474 );
xnor ( n23476 , n23475 , n19655 );
and ( n23477 , n23472 , n23476 );
and ( n23478 , n22235 , n19596 );
and ( n23479 , n21955 , n19594 );
nor ( n23480 , n23478 , n23479 );
xnor ( n23481 , n23480 , n19545 );
and ( n23482 , n23476 , n23481 );
and ( n23483 , n23472 , n23481 );
or ( n23484 , n23477 , n23482 , n23483 );
and ( n23485 , n20360 , n20674 );
and ( n23486 , n20268 , n20672 );
nor ( n23487 , n23485 , n23486 );
xnor ( n23488 , n23487 , n20542 );
and ( n23489 , n20618 , n20460 );
and ( n23490 , n20452 , n20458 );
nor ( n23491 , n23489 , n23490 );
xnor ( n23492 , n23491 , n20337 );
and ( n23493 , n23488 , n23492 );
not ( n23494 , n23437 );
and ( n23495 , n23492 , n23494 );
and ( n23496 , n23488 , n23494 );
or ( n23497 , n23493 , n23495 , n23496 );
and ( n23498 , n23484 , n23497 );
xor ( n23499 , n23265 , n23269 );
xor ( n23500 , n23499 , n23272 );
and ( n23501 , n23497 , n23500 );
and ( n23502 , n23484 , n23500 );
or ( n23503 , n23498 , n23501 , n23502 );
xor ( n23504 , n23113 , n23117 );
xor ( n23505 , n23504 , n23122 );
and ( n23506 , n23503 , n23505 );
xor ( n23507 , n23226 , n23233 );
xor ( n23508 , n23507 , n23238 );
and ( n23509 , n23505 , n23508 );
and ( n23510 , n23503 , n23508 );
or ( n23511 , n23506 , n23509 , n23510 );
xor ( n23512 , n23297 , n23299 );
xor ( n23513 , n23512 , n23302 );
and ( n23514 , n23511 , n23513 );
xor ( n23515 , n23241 , n23243 );
xor ( n23516 , n23515 , n23246 );
and ( n23517 , n23513 , n23516 );
and ( n23518 , n23511 , n23516 );
or ( n23519 , n23514 , n23517 , n23518 );
xor ( n23520 , n23208 , n23249 );
xor ( n23521 , n23520 , n23252 );
and ( n23522 , n23519 , n23521 );
xor ( n23523 , n23305 , n23307 );
xor ( n23524 , n23523 , n23310 );
and ( n23525 , n23521 , n23524 );
and ( n23526 , n23519 , n23524 );
or ( n23527 , n23522 , n23525 , n23526 );
and ( n23528 , n23468 , n23527 );
xor ( n23529 , n23173 , n23255 );
xor ( n23530 , n23529 , n23258 );
and ( n23531 , n23527 , n23530 );
and ( n23532 , n23468 , n23530 );
or ( n23533 , n23528 , n23531 , n23532 );
xor ( n23534 , n23069 , n23071 );
xor ( n23535 , n23534 , n23074 );
and ( n23536 , n23533 , n23535 );
xor ( n23537 , n23261 , n23321 );
xor ( n23538 , n23537 , n23324 );
and ( n23539 , n23535 , n23538 );
and ( n23540 , n23533 , n23538 );
or ( n23541 , n23536 , n23539 , n23540 );
and ( n23542 , n23339 , n23541 );
xor ( n23543 , n23339 , n23541 );
xor ( n23544 , n23533 , n23535 );
xor ( n23545 , n23544 , n23538 );
buf ( n23546 , n19388 );
buf ( n23547 , n19389 );
and ( n23548 , n23546 , n23547 );
not ( n23549 , n23548 );
and ( n23550 , n23210 , n23549 );
not ( n23551 , n23550 );
and ( n23552 , n22198 , n19596 );
and ( n23553 , n22235 , n19594 );
nor ( n23554 , n23552 , n23553 );
xnor ( n23555 , n23554 , n19545 );
and ( n23556 , n23551 , n23555 );
and ( n23557 , n22756 , n19518 );
and ( n23558 , n22425 , n19516 );
nor ( n23559 , n23557 , n23558 );
xnor ( n23560 , n23559 , n19489 );
and ( n23561 , n23555 , n23560 );
and ( n23562 , n23551 , n23560 );
or ( n23563 , n23556 , n23561 , n23562 );
and ( n23564 , n23141 , n19459 );
and ( n23565 , n22916 , n19457 );
nor ( n23566 , n23564 , n23565 );
xnor ( n23567 , n23566 , n19416 );
and ( n23568 , n23381 , n19424 );
and ( n23569 , n23271 , n19422 );
nor ( n23570 , n23568 , n23569 );
xnor ( n23571 , n23570 , n19431 );
and ( n23572 , n23567 , n23571 );
buf ( n23573 , n19323 );
and ( n23574 , n23573 , n19419 );
and ( n23575 , n23571 , n23574 );
and ( n23576 , n23567 , n23574 );
or ( n23577 , n23572 , n23575 , n23576 );
and ( n23578 , n23563 , n23577 );
and ( n23579 , n19811 , n21741 );
and ( n23580 , n19721 , n21739 );
nor ( n23581 , n23579 , n23580 );
xnor ( n23582 , n23581 , n21605 );
and ( n23583 , n23577 , n23582 );
and ( n23584 , n23563 , n23582 );
or ( n23585 , n23578 , n23583 , n23584 );
xor ( n23586 , n23421 , n23425 );
xor ( n23587 , n23586 , n23430 );
and ( n23588 , n23585 , n23587 );
xor ( n23589 , n23279 , n23283 );
xor ( n23590 , n23589 , n23288 );
and ( n23591 , n23587 , n23590 );
and ( n23592 , n23585 , n23590 );
or ( n23593 , n23588 , n23591 , n23592 );
and ( n23594 , n19434 , n23230 );
and ( n23595 , n19418 , n23228 );
nor ( n23596 , n23594 , n23595 );
xnor ( n23597 , n23596 , n22842 );
and ( n23598 , n20004 , n21155 );
and ( n23599 , n19946 , n21153 );
nor ( n23600 , n23598 , n23599 );
xnor ( n23601 , n23600 , n20994 );
and ( n23602 , n23597 , n23601 );
and ( n23603 , n21612 , n19805 );
and ( n23604 , n21451 , n19803 );
nor ( n23605 , n23603 , n23604 );
xnor ( n23606 , n23605 , n19750 );
and ( n23607 , n23601 , n23606 );
and ( n23608 , n23597 , n23606 );
or ( n23609 , n23602 , n23607 , n23608 );
and ( n23610 , n20803 , n20276 );
and ( n23611 , n20666 , n20274 );
nor ( n23612 , n23610 , n23611 );
xnor ( n23613 , n23612 , n20175 );
and ( n23614 , n21072 , n20114 );
and ( n23615 , n20867 , n20112 );
nor ( n23616 , n23614 , n23615 );
xnor ( n23617 , n23616 , n19997 );
and ( n23618 , n23613 , n23617 );
and ( n23619 , n21302 , n19894 );
and ( n23620 , n21218 , n19892 );
nor ( n23621 , n23619 , n23620 );
xnor ( n23622 , n23621 , n19858 );
and ( n23623 , n23617 , n23622 );
and ( n23624 , n23613 , n23622 );
or ( n23625 , n23618 , n23623 , n23624 );
and ( n23626 , n23609 , n23625 );
xor ( n23627 , n23438 , n23442 );
xor ( n23628 , n23627 , n23447 );
and ( n23629 , n23625 , n23628 );
and ( n23630 , n23609 , n23628 );
or ( n23631 , n23626 , n23629 , n23630 );
and ( n23632 , n23593 , n23631 );
xor ( n23633 , n23433 , n23450 );
xor ( n23634 , n23633 , n23453 );
and ( n23635 , n23631 , n23634 );
and ( n23636 , n23593 , n23634 );
or ( n23637 , n23632 , n23635 , n23636 );
xor ( n23638 , n22839 , n23209 );
xor ( n23639 , n23209 , n23210 );
not ( n23640 , n23639 );
and ( n23641 , n23638 , n23640 );
and ( n23642 , n19426 , n23641 );
not ( n23643 , n23642 );
xnor ( n23644 , n23643 , n23213 );
and ( n23645 , n19588 , n22381 );
and ( n23646 , n19510 , n22379 );
nor ( n23647 , n23645 , n23646 );
xnor ( n23648 , n23647 , n22228 );
and ( n23649 , n23644 , n23648 );
and ( n23650 , n19637 , n22048 );
and ( n23651 , n19605 , n22046 );
nor ( n23652 , n23650 , n23651 );
xnor ( n23653 , n23652 , n21853 );
and ( n23654 , n23648 , n23653 );
and ( n23655 , n23644 , n23653 );
or ( n23656 , n23649 , n23654 , n23655 );
xor ( n23657 , n23343 , n23347 );
xor ( n23658 , n23657 , n23352 );
and ( n23659 , n23656 , n23658 );
xor ( n23660 , n23401 , n23405 );
xor ( n23661 , n23660 , n23408 );
and ( n23662 , n23658 , n23661 );
and ( n23663 , n23656 , n23661 );
or ( n23664 , n23659 , n23662 , n23663 );
xor ( n23665 , n23275 , n23291 );
xor ( n23666 , n23665 , n23294 );
and ( n23667 , n23664 , n23666 );
xor ( n23668 , n23355 , n23357 );
xor ( n23669 , n23668 , n23360 );
and ( n23670 , n23666 , n23669 );
and ( n23671 , n23664 , n23669 );
or ( n23672 , n23667 , n23670 , n23671 );
and ( n23673 , n23637 , n23672 );
xor ( n23674 , n23363 , n23365 );
xor ( n23675 , n23674 , n23368 );
and ( n23676 , n23672 , n23675 );
and ( n23677 , n23637 , n23675 );
or ( n23678 , n23673 , n23676 , n23677 );
and ( n23679 , n20080 , n21155 );
and ( n23680 , n20004 , n21153 );
nor ( n23681 , n23679 , n23680 );
xnor ( n23682 , n23681 , n20994 );
and ( n23683 , n21704 , n19805 );
and ( n23684 , n21612 , n19803 );
nor ( n23685 , n23683 , n23684 );
xnor ( n23686 , n23685 , n19750 );
and ( n23687 , n23682 , n23686 );
and ( n23688 , n21955 , n19688 );
and ( n23689 , n21876 , n19686 );
nor ( n23690 , n23688 , n23689 );
xnor ( n23691 , n23690 , n19655 );
and ( n23692 , n23686 , n23691 );
and ( n23693 , n23682 , n23691 );
or ( n23694 , n23687 , n23692 , n23693 );
and ( n23695 , n20666 , n20460 );
and ( n23696 , n20618 , n20458 );
nor ( n23697 , n23695 , n23696 );
xnor ( n23698 , n23697 , n20337 );
and ( n23699 , n20867 , n20276 );
and ( n23700 , n20803 , n20274 );
nor ( n23701 , n23699 , n23700 );
xnor ( n23702 , n23701 , n20175 );
and ( n23703 , n23698 , n23702 );
and ( n23704 , n21218 , n20114 );
and ( n23705 , n21072 , n20112 );
nor ( n23706 , n23704 , n23705 );
xnor ( n23707 , n23706 , n19997 );
and ( n23708 , n23702 , n23707 );
and ( n23709 , n23698 , n23707 );
or ( n23710 , n23703 , n23708 , n23709 );
and ( n23711 , n23694 , n23710 );
and ( n23712 , n22425 , n19596 );
and ( n23713 , n22198 , n19594 );
nor ( n23714 , n23712 , n23713 );
xnor ( n23715 , n23714 , n19545 );
buf ( n23716 , n23715 );
and ( n23717 , n20268 , n20955 );
and ( n23718 , n20182 , n20953 );
nor ( n23719 , n23717 , n23718 );
xnor ( n23720 , n23719 , n20780 );
and ( n23721 , n23716 , n23720 );
and ( n23722 , n20452 , n20674 );
and ( n23723 , n20360 , n20672 );
nor ( n23724 , n23722 , n23723 );
xnor ( n23725 , n23724 , n20542 );
and ( n23726 , n23720 , n23725 );
and ( n23727 , n23716 , n23725 );
or ( n23728 , n23721 , n23726 , n23727 );
and ( n23729 , n23710 , n23728 );
and ( n23730 , n23694 , n23728 );
or ( n23731 , n23711 , n23729 , n23730 );
and ( n23732 , n19496 , n22859 );
and ( n23733 , n19469 , n22857 );
nor ( n23734 , n23732 , n23733 );
xnor ( n23735 , n23734 , n22418 );
and ( n23736 , n19881 , n21468 );
and ( n23737 , n19825 , n21466 );
nor ( n23738 , n23736 , n23737 );
xnor ( n23739 , n23738 , n21331 );
and ( n23740 , n23735 , n23739 );
xor ( n23741 , n23375 , n23379 );
xor ( n23742 , n23741 , n23382 );
and ( n23743 , n23739 , n23742 );
and ( n23744 , n23735 , n23742 );
or ( n23745 , n23740 , n23743 , n23744 );
and ( n23746 , n23731 , n23745 );
xor ( n23747 , n23385 , n23389 );
xor ( n23748 , n23747 , n23394 );
and ( n23749 , n23745 , n23748 );
and ( n23750 , n23731 , n23748 );
or ( n23751 , n23746 , n23749 , n23750 );
xor ( n23752 , n23397 , n23411 );
xor ( n23753 , n23752 , n23414 );
and ( n23754 , n23751 , n23753 );
xor ( n23755 , n23503 , n23505 );
xor ( n23756 , n23755 , n23508 );
and ( n23757 , n23753 , n23756 );
and ( n23758 , n23751 , n23756 );
or ( n23759 , n23754 , n23757 , n23758 );
xor ( n23760 , n23417 , n23456 );
xor ( n23761 , n23760 , n23459 );
and ( n23762 , n23759 , n23761 );
xor ( n23763 , n23511 , n23513 );
xor ( n23764 , n23763 , n23516 );
and ( n23765 , n23761 , n23764 );
and ( n23766 , n23759 , n23764 );
or ( n23767 , n23762 , n23765 , n23766 );
and ( n23768 , n23678 , n23767 );
xor ( n23769 , n23371 , n23462 );
xor ( n23770 , n23769 , n23465 );
and ( n23771 , n23767 , n23770 );
and ( n23772 , n23678 , n23770 );
or ( n23773 , n23768 , n23771 , n23772 );
xor ( n23774 , n23468 , n23527 );
xor ( n23775 , n23774 , n23530 );
and ( n23776 , n23773 , n23775 );
xor ( n23777 , n23313 , n23315 );
xor ( n23778 , n23777 , n23318 );
and ( n23779 , n23775 , n23778 );
and ( n23780 , n23773 , n23778 );
or ( n23781 , n23776 , n23779 , n23780 );
and ( n23782 , n23545 , n23781 );
xor ( n23783 , n23545 , n23781 );
xor ( n23784 , n23773 , n23775 );
xor ( n23785 , n23784 , n23778 );
and ( n23786 , n19418 , n23641 );
and ( n23787 , n19426 , n23639 );
nor ( n23788 , n23786 , n23787 );
xnor ( n23789 , n23788 , n23213 );
and ( n23790 , n19946 , n21468 );
and ( n23791 , n19881 , n21466 );
nor ( n23792 , n23790 , n23791 );
xnor ( n23793 , n23792 , n21331 );
and ( n23794 , n23789 , n23793 );
and ( n23795 , n21451 , n19894 );
and ( n23796 , n21302 , n19892 );
nor ( n23797 , n23795 , n23796 );
xnor ( n23798 , n23797 , n19858 );
and ( n23799 , n23793 , n23798 );
and ( n23800 , n23789 , n23798 );
or ( n23801 , n23794 , n23799 , n23800 );
and ( n23802 , n19510 , n22859 );
and ( n23803 , n19496 , n22857 );
nor ( n23804 , n23802 , n23803 );
xnor ( n23805 , n23804 , n22418 );
and ( n23806 , n19605 , n22381 );
and ( n23807 , n19588 , n22379 );
nor ( n23808 , n23806 , n23807 );
xnor ( n23809 , n23808 , n22228 );
and ( n23810 , n23805 , n23809 );
and ( n23811 , n19721 , n22048 );
and ( n23812 , n19637 , n22046 );
nor ( n23813 , n23811 , n23812 );
xnor ( n23814 , n23813 , n21853 );
and ( n23815 , n23809 , n23814 );
and ( n23816 , n23805 , n23814 );
or ( n23817 , n23810 , n23815 , n23816 );
and ( n23818 , n23801 , n23817 );
xor ( n23819 , n23488 , n23492 );
xor ( n23820 , n23819 , n23494 );
and ( n23821 , n23817 , n23820 );
and ( n23822 , n23801 , n23820 );
or ( n23823 , n23818 , n23821 , n23822 );
and ( n23824 , n22916 , n19518 );
and ( n23825 , n22756 , n19516 );
nor ( n23826 , n23824 , n23825 );
xnor ( n23827 , n23826 , n19489 );
and ( n23828 , n23271 , n19459 );
and ( n23829 , n23141 , n19457 );
nor ( n23830 , n23828 , n23829 );
xnor ( n23831 , n23830 , n19416 );
and ( n23832 , n23827 , n23831 );
and ( n23833 , n23573 , n19424 );
and ( n23834 , n23381 , n19422 );
nor ( n23835 , n23833 , n23834 );
xnor ( n23836 , n23835 , n19431 );
and ( n23837 , n23831 , n23836 );
and ( n23838 , n23827 , n23836 );
or ( n23839 , n23832 , n23837 , n23838 );
and ( n23840 , n19469 , n23230 );
and ( n23841 , n19434 , n23228 );
nor ( n23842 , n23840 , n23841 );
xnor ( n23843 , n23842 , n22842 );
and ( n23844 , n23839 , n23843 );
and ( n23845 , n19825 , n21741 );
and ( n23846 , n19811 , n21739 );
nor ( n23847 , n23845 , n23846 );
xnor ( n23848 , n23847 , n21605 );
and ( n23849 , n23843 , n23848 );
and ( n23850 , n23839 , n23848 );
or ( n23851 , n23844 , n23849 , n23850 );
xor ( n23852 , n23472 , n23476 );
xor ( n23853 , n23852 , n23481 );
and ( n23854 , n23851 , n23853 );
xor ( n23855 , n23613 , n23617 );
xor ( n23856 , n23855 , n23622 );
and ( n23857 , n23853 , n23856 );
and ( n23858 , n23851 , n23856 );
or ( n23859 , n23854 , n23857 , n23858 );
and ( n23860 , n23823 , n23859 );
xor ( n23861 , n23484 , n23497 );
xor ( n23862 , n23861 , n23500 );
and ( n23863 , n23859 , n23862 );
and ( n23864 , n23823 , n23862 );
or ( n23865 , n23860 , n23863 , n23864 );
xor ( n23866 , n23597 , n23601 );
xor ( n23867 , n23866 , n23606 );
xor ( n23868 , n23644 , n23648 );
xor ( n23869 , n23868 , n23653 );
and ( n23870 , n23867 , n23869 );
xor ( n23871 , n23735 , n23739 );
xor ( n23872 , n23871 , n23742 );
and ( n23873 , n23869 , n23872 );
and ( n23874 , n23867 , n23872 );
or ( n23875 , n23870 , n23873 , n23874 );
xor ( n23876 , n23585 , n23587 );
xor ( n23877 , n23876 , n23590 );
and ( n23878 , n23875 , n23877 );
xor ( n23879 , n23609 , n23625 );
xor ( n23880 , n23879 , n23628 );
and ( n23881 , n23877 , n23880 );
and ( n23882 , n23875 , n23880 );
or ( n23883 , n23878 , n23881 , n23882 );
and ( n23884 , n23865 , n23883 );
xor ( n23885 , n23593 , n23631 );
xor ( n23886 , n23885 , n23634 );
and ( n23887 , n23883 , n23886 );
and ( n23888 , n23865 , n23886 );
or ( n23889 , n23884 , n23887 , n23888 );
and ( n23890 , n20004 , n21468 );
and ( n23891 , n19946 , n21466 );
nor ( n23892 , n23890 , n23891 );
xnor ( n23893 , n23892 , n21331 );
and ( n23894 , n21302 , n20114 );
and ( n23895 , n21218 , n20112 );
nor ( n23896 , n23894 , n23895 );
xnor ( n23897 , n23896 , n19997 );
and ( n23898 , n23893 , n23897 );
and ( n23899 , n21612 , n19894 );
and ( n23900 , n21451 , n19892 );
nor ( n23901 , n23899 , n23900 );
xnor ( n23902 , n23901 , n19858 );
and ( n23903 , n23897 , n23902 );
and ( n23904 , n23893 , n23902 );
or ( n23905 , n23898 , n23903 , n23904 );
and ( n23906 , n19434 , n23641 );
and ( n23907 , n19418 , n23639 );
nor ( n23908 , n23906 , n23907 );
xnor ( n23909 , n23908 , n23213 );
and ( n23910 , n19588 , n22859 );
and ( n23911 , n19510 , n22857 );
nor ( n23912 , n23910 , n23911 );
xnor ( n23913 , n23912 , n22418 );
and ( n23914 , n23909 , n23913 );
and ( n23915 , n19637 , n22381 );
and ( n23916 , n19605 , n22379 );
nor ( n23917 , n23915 , n23916 );
xnor ( n23918 , n23917 , n22228 );
and ( n23919 , n23913 , n23918 );
and ( n23920 , n23909 , n23918 );
or ( n23921 , n23914 , n23919 , n23920 );
and ( n23922 , n23905 , n23921 );
buf ( n23923 , n19390 );
buf ( n23924 , n19391 );
and ( n23925 , n23923 , n23924 );
not ( n23926 , n23925 );
and ( n23927 , n23547 , n23926 );
not ( n23928 , n23927 );
and ( n23929 , n22198 , n19688 );
and ( n23930 , n22235 , n19686 );
nor ( n23931 , n23929 , n23930 );
xnor ( n23932 , n23931 , n19655 );
and ( n23933 , n23928 , n23932 );
and ( n23934 , n22756 , n19596 );
and ( n23935 , n22425 , n19594 );
nor ( n23936 , n23934 , n23935 );
xnor ( n23937 , n23936 , n19545 );
and ( n23938 , n23932 , n23937 );
and ( n23939 , n23928 , n23937 );
or ( n23940 , n23933 , n23938 , n23939 );
xor ( n23941 , n23210 , n23546 );
xor ( n23942 , n23546 , n23547 );
not ( n23943 , n23942 );
and ( n23944 , n23941 , n23943 );
and ( n23945 , n19426 , n23944 );
not ( n23946 , n23945 );
xnor ( n23947 , n23946 , n23550 );
and ( n23948 , n23940 , n23947 );
and ( n23949 , n19811 , n22048 );
and ( n23950 , n19721 , n22046 );
nor ( n23951 , n23949 , n23950 );
xnor ( n23952 , n23951 , n21853 );
and ( n23953 , n23947 , n23952 );
and ( n23954 , n23940 , n23952 );
or ( n23955 , n23948 , n23953 , n23954 );
and ( n23956 , n23921 , n23955 );
and ( n23957 , n23905 , n23955 );
or ( n23958 , n23922 , n23956 , n23957 );
and ( n23959 , n23141 , n19518 );
and ( n23960 , n22916 , n19516 );
nor ( n23961 , n23959 , n23960 );
xnor ( n23962 , n23961 , n19489 );
and ( n23963 , n23381 , n19459 );
and ( n23964 , n23271 , n19457 );
nor ( n23965 , n23963 , n23964 );
xnor ( n23966 , n23965 , n19416 );
and ( n23967 , n23962 , n23966 );
buf ( n23968 , n19324 );
and ( n23969 , n23968 , n19424 );
and ( n23970 , n23573 , n19422 );
nor ( n23971 , n23969 , n23970 );
xnor ( n23972 , n23971 , n19431 );
and ( n23973 , n23966 , n23972 );
and ( n23974 , n23962 , n23972 );
or ( n23975 , n23967 , n23973 , n23974 );
and ( n23976 , n19496 , n23230 );
and ( n23977 , n19469 , n23228 );
nor ( n23978 , n23976 , n23977 );
xnor ( n23979 , n23978 , n22842 );
and ( n23980 , n23975 , n23979 );
and ( n23981 , n19881 , n21741 );
and ( n23982 , n19825 , n21739 );
nor ( n23983 , n23981 , n23982 );
xnor ( n23984 , n23983 , n21605 );
and ( n23985 , n23979 , n23984 );
and ( n23986 , n23975 , n23984 );
or ( n23987 , n23980 , n23985 , n23986 );
xor ( n23988 , n23682 , n23686 );
xor ( n23989 , n23988 , n23691 );
and ( n23990 , n23987 , n23989 );
xor ( n23991 , n23716 , n23720 );
xor ( n23992 , n23991 , n23725 );
and ( n23993 , n23989 , n23992 );
and ( n23994 , n23987 , n23992 );
or ( n23995 , n23990 , n23993 , n23994 );
and ( n23996 , n23958 , n23995 );
xor ( n23997 , n23694 , n23710 );
xor ( n23998 , n23997 , n23728 );
and ( n23999 , n23995 , n23998 );
and ( n24000 , n23958 , n23998 );
or ( n24001 , n23996 , n23999 , n24000 );
xor ( n24002 , n23731 , n23745 );
xor ( n24003 , n24002 , n23748 );
and ( n24004 , n24001 , n24003 );
xor ( n24005 , n23656 , n23658 );
xor ( n24006 , n24005 , n23661 );
and ( n24007 , n24003 , n24006 );
and ( n24008 , n24001 , n24006 );
or ( n24009 , n24004 , n24007 , n24008 );
xor ( n24010 , n23664 , n23666 );
xor ( n24011 , n24010 , n23669 );
and ( n24012 , n24009 , n24011 );
xor ( n24013 , n23751 , n23753 );
xor ( n24014 , n24013 , n23756 );
and ( n24015 , n24011 , n24014 );
and ( n24016 , n24009 , n24014 );
or ( n24017 , n24012 , n24015 , n24016 );
and ( n24018 , n23889 , n24017 );
xor ( n24019 , n23637 , n23672 );
xor ( n24020 , n24019 , n23675 );
and ( n24021 , n24017 , n24020 );
and ( n24022 , n23889 , n24020 );
or ( n24023 , n24018 , n24021 , n24022 );
xor ( n24024 , n23678 , n23767 );
xor ( n24025 , n24024 , n23770 );
and ( n24026 , n24023 , n24025 );
xor ( n24027 , n23519 , n23521 );
xor ( n24028 , n24027 , n23524 );
and ( n24029 , n24025 , n24028 );
and ( n24030 , n24023 , n24028 );
or ( n24031 , n24026 , n24029 , n24030 );
and ( n24032 , n23785 , n24031 );
xor ( n24033 , n23785 , n24031 );
xor ( n24034 , n24023 , n24025 );
xor ( n24035 , n24034 , n24028 );
and ( n24036 , n21876 , n19805 );
and ( n24037 , n21704 , n19803 );
nor ( n24038 , n24036 , n24037 );
xnor ( n24039 , n24038 , n19750 );
and ( n24040 , n22235 , n19688 );
and ( n24041 , n21955 , n19686 );
nor ( n24042 , n24040 , n24041 );
xnor ( n24043 , n24042 , n19655 );
and ( n24044 , n24039 , n24043 );
and ( n24045 , n23968 , n19419 );
and ( n24046 , n24043 , n24045 );
and ( n24047 , n24039 , n24045 );
or ( n24048 , n24044 , n24046 , n24047 );
xor ( n24049 , n23551 , n23555 );
xor ( n24050 , n24049 , n23560 );
and ( n24051 , n24048 , n24050 );
xor ( n24052 , n23567 , n23571 );
xor ( n24053 , n24052 , n23574 );
and ( n24054 , n24050 , n24053 );
and ( n24055 , n24048 , n24053 );
or ( n24056 , n24051 , n24054 , n24055 );
and ( n24057 , n20182 , n21155 );
and ( n24058 , n20080 , n21153 );
nor ( n24059 , n24057 , n24058 );
xnor ( n24060 , n24059 , n20994 );
and ( n24061 , n20360 , n20955 );
and ( n24062 , n20268 , n20953 );
nor ( n24063 , n24061 , n24062 );
xnor ( n24064 , n24063 , n20780 );
and ( n24065 , n24060 , n24064 );
and ( n24066 , n20618 , n20674 );
and ( n24067 , n20452 , n20672 );
nor ( n24068 , n24066 , n24067 );
xnor ( n24069 , n24068 , n20542 );
and ( n24070 , n24064 , n24069 );
and ( n24071 , n24060 , n24069 );
or ( n24072 , n24065 , n24070 , n24071 );
and ( n24073 , n20803 , n20460 );
and ( n24074 , n20666 , n20458 );
nor ( n24075 , n24073 , n24074 );
xnor ( n24076 , n24075 , n20337 );
and ( n24077 , n21072 , n20276 );
and ( n24078 , n20867 , n20274 );
nor ( n24079 , n24077 , n24078 );
xnor ( n24080 , n24079 , n20175 );
and ( n24081 , n24076 , n24080 );
not ( n24082 , n23715 );
and ( n24083 , n24080 , n24082 );
and ( n24084 , n24076 , n24082 );
or ( n24085 , n24081 , n24083 , n24084 );
and ( n24086 , n24072 , n24085 );
xor ( n24087 , n23698 , n23702 );
xor ( n24088 , n24087 , n23707 );
and ( n24089 , n24085 , n24088 );
and ( n24090 , n24072 , n24088 );
or ( n24091 , n24086 , n24089 , n24090 );
and ( n24092 , n24056 , n24091 );
xor ( n24093 , n23563 , n23577 );
xor ( n24094 , n24093 , n23582 );
and ( n24095 , n24091 , n24094 );
and ( n24096 , n24056 , n24094 );
or ( n24097 , n24092 , n24095 , n24096 );
xor ( n24098 , n23789 , n23793 );
xor ( n24099 , n24098 , n23798 );
xor ( n24100 , n23805 , n23809 );
xor ( n24101 , n24100 , n23814 );
and ( n24102 , n24099 , n24101 );
xor ( n24103 , n23839 , n23843 );
xor ( n24104 , n24103 , n23848 );
and ( n24105 , n24101 , n24104 );
and ( n24106 , n24099 , n24104 );
or ( n24107 , n24102 , n24105 , n24106 );
xor ( n24108 , n23801 , n23817 );
xor ( n24109 , n24108 , n23820 );
and ( n24110 , n24107 , n24109 );
xor ( n24111 , n23851 , n23853 );
xor ( n24112 , n24111 , n23856 );
and ( n24113 , n24109 , n24112 );
and ( n24114 , n24107 , n24112 );
or ( n24115 , n24110 , n24113 , n24114 );
and ( n24116 , n24097 , n24115 );
xor ( n24117 , n23823 , n23859 );
xor ( n24118 , n24117 , n23862 );
and ( n24119 , n24115 , n24118 );
and ( n24120 , n24097 , n24118 );
or ( n24121 , n24116 , n24119 , n24120 );
and ( n24122 , n20080 , n21468 );
and ( n24123 , n20004 , n21466 );
nor ( n24124 , n24122 , n24123 );
xnor ( n24125 , n24124 , n21331 );
and ( n24126 , n21955 , n19805 );
and ( n24127 , n21876 , n19803 );
nor ( n24128 , n24126 , n24127 );
xnor ( n24129 , n24128 , n19750 );
and ( n24130 , n24125 , n24129 );
buf ( n24131 , n19325 );
and ( n24132 , n24131 , n19419 );
and ( n24133 , n24129 , n24132 );
and ( n24134 , n24125 , n24132 );
or ( n24135 , n24130 , n24133 , n24134 );
xor ( n24136 , n23827 , n23831 );
xor ( n24137 , n24136 , n23836 );
and ( n24138 , n24135 , n24137 );
xor ( n24139 , n24039 , n24043 );
xor ( n24140 , n24139 , n24045 );
and ( n24141 , n24137 , n24140 );
and ( n24142 , n24135 , n24140 );
or ( n24143 , n24138 , n24141 , n24142 );
and ( n24144 , n23271 , n19518 );
and ( n24145 , n23141 , n19516 );
nor ( n24146 , n24144 , n24145 );
xnor ( n24147 , n24146 , n19489 );
and ( n24148 , n23573 , n19459 );
and ( n24149 , n23381 , n19457 );
nor ( n24150 , n24148 , n24149 );
xnor ( n24151 , n24150 , n19416 );
and ( n24152 , n24147 , n24151 );
and ( n24153 , n24131 , n19424 );
and ( n24154 , n23968 , n19422 );
nor ( n24155 , n24153 , n24154 );
xnor ( n24156 , n24155 , n19431 );
and ( n24157 , n24151 , n24156 );
and ( n24158 , n24147 , n24156 );
or ( n24159 , n24152 , n24157 , n24158 );
and ( n24160 , n19469 , n23641 );
and ( n24161 , n19434 , n23639 );
nor ( n24162 , n24160 , n24161 );
xnor ( n24163 , n24162 , n23213 );
and ( n24164 , n24159 , n24163 );
and ( n24165 , n19721 , n22381 );
and ( n24166 , n19637 , n22379 );
nor ( n24167 , n24165 , n24166 );
xnor ( n24168 , n24167 , n22228 );
and ( n24169 , n24163 , n24168 );
and ( n24170 , n24159 , n24168 );
or ( n24171 , n24164 , n24169 , n24170 );
xor ( n24172 , n23893 , n23897 );
xor ( n24173 , n24172 , n23902 );
and ( n24174 , n24171 , n24173 );
xor ( n24175 , n24060 , n24064 );
xor ( n24176 , n24175 , n24069 );
and ( n24177 , n24173 , n24176 );
and ( n24178 , n24171 , n24176 );
or ( n24179 , n24174 , n24177 , n24178 );
and ( n24180 , n24143 , n24179 );
xor ( n24181 , n24048 , n24050 );
xor ( n24182 , n24181 , n24053 );
and ( n24183 , n24179 , n24182 );
and ( n24184 , n24143 , n24182 );
or ( n24185 , n24180 , n24183 , n24184 );
xor ( n24186 , n24056 , n24091 );
xor ( n24187 , n24186 , n24094 );
and ( n24188 , n24185 , n24187 );
xor ( n24189 , n23867 , n23869 );
xor ( n24190 , n24189 , n23872 );
and ( n24191 , n24187 , n24190 );
and ( n24192 , n24185 , n24190 );
or ( n24193 , n24188 , n24191 , n24192 );
xor ( n24194 , n23875 , n23877 );
xor ( n24195 , n24194 , n23880 );
and ( n24196 , n24193 , n24195 );
xor ( n24197 , n24001 , n24003 );
xor ( n24198 , n24197 , n24006 );
and ( n24199 , n24195 , n24198 );
and ( n24200 , n24193 , n24198 );
or ( n24201 , n24196 , n24199 , n24200 );
and ( n24202 , n24121 , n24201 );
xor ( n24203 , n23865 , n23883 );
xor ( n24204 , n24203 , n23886 );
and ( n24205 , n24201 , n24204 );
and ( n24206 , n24121 , n24204 );
or ( n24207 , n24202 , n24205 , n24206 );
xor ( n24208 , n23759 , n23761 );
xor ( n24209 , n24208 , n23764 );
and ( n24210 , n24207 , n24209 );
xor ( n24211 , n23889 , n24017 );
xor ( n24212 , n24211 , n24020 );
and ( n24213 , n24209 , n24212 );
and ( n24214 , n24207 , n24212 );
or ( n24215 , n24210 , n24213 , n24214 );
and ( n24216 , n24035 , n24215 );
xor ( n24217 , n24035 , n24215 );
xor ( n24218 , n24207 , n24209 );
xor ( n24219 , n24218 , n24212 );
and ( n24220 , n19825 , n22048 );
and ( n24221 , n19811 , n22046 );
nor ( n24222 , n24220 , n24221 );
xnor ( n24223 , n24222 , n21853 );
xor ( n24224 , n23928 , n23932 );
xor ( n24225 , n24224 , n23937 );
and ( n24226 , n24223 , n24225 );
xor ( n24227 , n23962 , n23966 );
xor ( n24228 , n24227 , n23972 );
and ( n24229 , n24225 , n24228 );
and ( n24230 , n24223 , n24228 );
or ( n24231 , n24226 , n24229 , n24230 );
xor ( n24232 , n23909 , n23913 );
xor ( n24233 , n24232 , n23918 );
and ( n24234 , n24231 , n24233 );
xor ( n24235 , n23940 , n23947 );
xor ( n24236 , n24235 , n23952 );
and ( n24237 , n24233 , n24236 );
and ( n24238 , n24231 , n24236 );
or ( n24239 , n24234 , n24237 , n24238 );
and ( n24240 , n20268 , n21155 );
and ( n24241 , n20182 , n21153 );
nor ( n24242 , n24240 , n24241 );
xnor ( n24243 , n24242 , n20994 );
and ( n24244 , n20452 , n20955 );
and ( n24245 , n20360 , n20953 );
nor ( n24246 , n24244 , n24245 );
xnor ( n24247 , n24246 , n20780 );
and ( n24248 , n24243 , n24247 );
and ( n24249 , n21704 , n19894 );
and ( n24250 , n21612 , n19892 );
nor ( n24251 , n24249 , n24250 );
xnor ( n24252 , n24251 , n19858 );
and ( n24253 , n24247 , n24252 );
and ( n24254 , n24243 , n24252 );
or ( n24255 , n24248 , n24253 , n24254 );
and ( n24256 , n22916 , n19596 );
and ( n24257 , n22756 , n19594 );
nor ( n24258 , n24256 , n24257 );
xnor ( n24259 , n24258 , n19545 );
buf ( n24260 , n24259 );
and ( n24261 , n20666 , n20674 );
and ( n24262 , n20618 , n20672 );
nor ( n24263 , n24261 , n24262 );
xnor ( n24264 , n24263 , n20542 );
and ( n24265 , n24260 , n24264 );
and ( n24266 , n20867 , n20460 );
and ( n24267 , n20803 , n20458 );
nor ( n24268 , n24266 , n24267 );
xnor ( n24269 , n24268 , n20337 );
and ( n24270 , n24264 , n24269 );
and ( n24271 , n24260 , n24269 );
or ( n24272 , n24265 , n24270 , n24271 );
and ( n24273 , n24255 , n24272 );
xor ( n24274 , n24076 , n24080 );
xor ( n24275 , n24274 , n24082 );
and ( n24276 , n24272 , n24275 );
and ( n24277 , n24255 , n24275 );
or ( n24278 , n24273 , n24276 , n24277 );
and ( n24279 , n24239 , n24278 );
xor ( n24280 , n24072 , n24085 );
xor ( n24281 , n24280 , n24088 );
and ( n24282 , n24278 , n24281 );
and ( n24283 , n24239 , n24281 );
or ( n24284 , n24279 , n24282 , n24283 );
and ( n24285 , n19946 , n21741 );
and ( n24286 , n19881 , n21739 );
nor ( n24287 , n24285 , n24286 );
xnor ( n24288 , n24287 , n21605 );
and ( n24289 , n21218 , n20276 );
and ( n24290 , n21072 , n20274 );
nor ( n24291 , n24289 , n24290 );
xnor ( n24292 , n24291 , n20175 );
and ( n24293 , n24288 , n24292 );
and ( n24294 , n21451 , n20114 );
and ( n24295 , n21302 , n20112 );
nor ( n24296 , n24294 , n24295 );
xnor ( n24297 , n24296 , n19997 );
and ( n24298 , n24292 , n24297 );
and ( n24299 , n24288 , n24297 );
or ( n24300 , n24293 , n24298 , n24299 );
and ( n24301 , n19418 , n23944 );
and ( n24302 , n19426 , n23942 );
nor ( n24303 , n24301 , n24302 );
xnor ( n24304 , n24303 , n23550 );
and ( n24305 , n19510 , n23230 );
and ( n24306 , n19496 , n23228 );
nor ( n24307 , n24305 , n24306 );
xnor ( n24308 , n24307 , n22842 );
and ( n24309 , n24304 , n24308 );
and ( n24310 , n19605 , n22859 );
and ( n24311 , n19588 , n22857 );
nor ( n24312 , n24310 , n24311 );
xnor ( n24313 , n24312 , n22418 );
and ( n24314 , n24308 , n24313 );
and ( n24315 , n24304 , n24313 );
or ( n24316 , n24309 , n24314 , n24315 );
and ( n24317 , n24300 , n24316 );
xor ( n24318 , n23975 , n23979 );
xor ( n24319 , n24318 , n23984 );
and ( n24320 , n24316 , n24319 );
and ( n24321 , n24300 , n24319 );
or ( n24322 , n24317 , n24320 , n24321 );
xor ( n24323 , n23905 , n23921 );
xor ( n24324 , n24323 , n23955 );
and ( n24325 , n24322 , n24324 );
xor ( n24326 , n23987 , n23989 );
xor ( n24327 , n24326 , n23992 );
and ( n24328 , n24324 , n24327 );
and ( n24329 , n24322 , n24327 );
or ( n24330 , n24325 , n24328 , n24329 );
and ( n24331 , n24284 , n24330 );
xor ( n24332 , n23958 , n23995 );
xor ( n24333 , n24332 , n23998 );
and ( n24334 , n24330 , n24333 );
and ( n24335 , n24284 , n24333 );
or ( n24336 , n24331 , n24334 , n24335 );
xor ( n24337 , n24097 , n24115 );
xor ( n24338 , n24337 , n24118 );
and ( n24339 , n24336 , n24338 );
xor ( n24340 , n24193 , n24195 );
xor ( n24341 , n24340 , n24198 );
and ( n24342 , n24338 , n24341 );
and ( n24343 , n24336 , n24341 );
or ( n24344 , n24339 , n24342 , n24343 );
xor ( n24345 , n24009 , n24011 );
xor ( n24346 , n24345 , n24014 );
and ( n24347 , n24344 , n24346 );
xor ( n24348 , n24121 , n24201 );
xor ( n24349 , n24348 , n24204 );
and ( n24350 , n24346 , n24349 );
and ( n24351 , n24344 , n24349 );
or ( n24352 , n24347 , n24350 , n24351 );
and ( n24353 , n24219 , n24352 );
xor ( n24354 , n24219 , n24352 );
xor ( n24355 , n24344 , n24346 );
xor ( n24356 , n24355 , n24349 );
and ( n24357 , n21072 , n20460 );
and ( n24358 , n20867 , n20458 );
nor ( n24359 , n24357 , n24358 );
xnor ( n24360 , n24359 , n20337 );
and ( n24361 , n21302 , n20276 );
and ( n24362 , n21218 , n20274 );
nor ( n24363 , n24361 , n24362 );
xnor ( n24364 , n24363 , n20175 );
and ( n24365 , n24360 , n24364 );
and ( n24366 , n21612 , n20114 );
and ( n24367 , n21451 , n20112 );
nor ( n24368 , n24366 , n24367 );
xnor ( n24369 , n24368 , n19997 );
and ( n24370 , n24364 , n24369 );
and ( n24371 , n24360 , n24369 );
or ( n24372 , n24365 , n24370 , n24371 );
xor ( n24373 , n23547 , n23923 );
xor ( n24374 , n23923 , n23924 );
not ( n24375 , n24374 );
and ( n24376 , n24373 , n24375 );
and ( n24377 , n19426 , n24376 );
not ( n24378 , n24377 );
xnor ( n24379 , n24378 , n23927 );
and ( n24380 , n19637 , n22859 );
and ( n24381 , n19605 , n22857 );
nor ( n24382 , n24380 , n24381 );
xnor ( n24383 , n24382 , n22418 );
and ( n24384 , n24379 , n24383 );
and ( n24385 , n19811 , n22381 );
and ( n24386 , n19721 , n22379 );
nor ( n24387 , n24385 , n24386 );
xnor ( n24388 , n24387 , n22228 );
and ( n24389 , n24383 , n24388 );
and ( n24390 , n24379 , n24388 );
or ( n24391 , n24384 , n24389 , n24390 );
and ( n24392 , n24372 , n24391 );
buf ( n24393 , n19392 );
buf ( n24394 , n19393 );
and ( n24395 , n24393 , n24394 );
not ( n24396 , n24395 );
and ( n24397 , n23924 , n24396 );
not ( n24398 , n24397 );
and ( n24399 , n22198 , n19805 );
and ( n24400 , n22235 , n19803 );
nor ( n24401 , n24399 , n24400 );
xnor ( n24402 , n24401 , n19750 );
and ( n24403 , n24398 , n24402 );
and ( n24404 , n22756 , n19688 );
and ( n24405 , n22425 , n19686 );
nor ( n24406 , n24404 , n24405 );
xnor ( n24407 , n24406 , n19655 );
and ( n24408 , n24402 , n24407 );
and ( n24409 , n24398 , n24407 );
or ( n24410 , n24403 , n24408 , n24409 );
and ( n24411 , n23141 , n19596 );
and ( n24412 , n22916 , n19594 );
nor ( n24413 , n24411 , n24412 );
xnor ( n24414 , n24413 , n19545 );
and ( n24415 , n23381 , n19518 );
and ( n24416 , n23271 , n19516 );
nor ( n24417 , n24415 , n24416 );
xnor ( n24418 , n24417 , n19489 );
and ( n24419 , n24414 , n24418 );
and ( n24420 , n23968 , n19459 );
and ( n24421 , n23573 , n19457 );
nor ( n24422 , n24420 , n24421 );
xnor ( n24423 , n24422 , n19416 );
and ( n24424 , n24418 , n24423 );
and ( n24425 , n24414 , n24423 );
or ( n24426 , n24419 , n24424 , n24425 );
and ( n24427 , n24410 , n24426 );
and ( n24428 , n19496 , n23641 );
and ( n24429 , n19469 , n23639 );
nor ( n24430 , n24428 , n24429 );
xnor ( n24431 , n24430 , n23213 );
and ( n24432 , n24426 , n24431 );
and ( n24433 , n24410 , n24431 );
or ( n24434 , n24427 , n24432 , n24433 );
and ( n24435 , n24391 , n24434 );
and ( n24436 , n24372 , n24434 );
or ( n24437 , n24392 , n24435 , n24436 );
and ( n24438 , n19434 , n23944 );
and ( n24439 , n19418 , n23942 );
nor ( n24440 , n24438 , n24439 );
xnor ( n24441 , n24440 , n23550 );
and ( n24442 , n19588 , n23230 );
and ( n24443 , n19510 , n23228 );
nor ( n24444 , n24442 , n24443 );
xnor ( n24445 , n24444 , n22842 );
and ( n24446 , n24441 , n24445 );
and ( n24447 , n20004 , n21741 );
and ( n24448 , n19946 , n21739 );
nor ( n24449 , n24447 , n24448 );
xnor ( n24450 , n24449 , n21605 );
and ( n24451 , n24445 , n24450 );
and ( n24452 , n24441 , n24450 );
or ( n24453 , n24446 , n24451 , n24452 );
xor ( n24454 , n24125 , n24129 );
xor ( n24455 , n24454 , n24132 );
and ( n24456 , n24453 , n24455 );
xor ( n24457 , n24304 , n24308 );
xor ( n24458 , n24457 , n24313 );
and ( n24459 , n24455 , n24458 );
and ( n24460 , n24453 , n24458 );
or ( n24461 , n24456 , n24459 , n24460 );
and ( n24462 , n24437 , n24461 );
xor ( n24463 , n24135 , n24137 );
xor ( n24464 , n24463 , n24140 );
and ( n24465 , n24461 , n24464 );
and ( n24466 , n24437 , n24464 );
or ( n24467 , n24462 , n24465 , n24466 );
xor ( n24468 , n24171 , n24173 );
xor ( n24469 , n24468 , n24176 );
xor ( n24470 , n24300 , n24316 );
xor ( n24471 , n24470 , n24319 );
and ( n24472 , n24469 , n24471 );
xor ( n24473 , n24231 , n24233 );
xor ( n24474 , n24473 , n24236 );
and ( n24475 , n24471 , n24474 );
and ( n24476 , n24469 , n24474 );
or ( n24477 , n24472 , n24475 , n24476 );
and ( n24478 , n24467 , n24477 );
xor ( n24479 , n24239 , n24278 );
xor ( n24480 , n24479 , n24281 );
and ( n24481 , n24477 , n24480 );
and ( n24482 , n24467 , n24480 );
or ( n24483 , n24478 , n24481 , n24482 );
and ( n24484 , n20452 , n21155 );
and ( n24485 , n20360 , n21153 );
nor ( n24486 , n24484 , n24485 );
xnor ( n24487 , n24486 , n20994 );
and ( n24488 , n20666 , n20955 );
and ( n24489 , n20618 , n20953 );
nor ( n24490 , n24488 , n24489 );
xnor ( n24491 , n24490 , n20780 );
and ( n24492 , n24487 , n24491 );
and ( n24493 , n20867 , n20674 );
and ( n24494 , n20803 , n20672 );
nor ( n24495 , n24493 , n24494 );
xnor ( n24496 , n24495 , n20542 );
and ( n24497 , n24491 , n24496 );
and ( n24498 , n24487 , n24496 );
or ( n24499 , n24492 , n24497 , n24498 );
and ( n24500 , n20080 , n21741 );
and ( n24501 , n20004 , n21739 );
nor ( n24502 , n24500 , n24501 );
xnor ( n24503 , n24502 , n21605 );
and ( n24504 , n20268 , n21468 );
and ( n24505 , n20182 , n21466 );
nor ( n24506 , n24504 , n24505 );
xnor ( n24507 , n24506 , n21331 );
and ( n24508 , n24503 , n24507 );
and ( n24509 , n21704 , n20114 );
and ( n24510 , n21612 , n20112 );
nor ( n24511 , n24509 , n24510 );
xnor ( n24512 , n24511 , n19997 );
and ( n24513 , n24507 , n24512 );
and ( n24514 , n24503 , n24512 );
or ( n24515 , n24508 , n24513 , n24514 );
and ( n24516 , n24499 , n24515 );
and ( n24517 , n21955 , n19894 );
and ( n24518 , n21876 , n19892 );
nor ( n24519 , n24517 , n24518 );
xnor ( n24520 , n24519 , n19858 );
buf ( n24521 , n19326 );
and ( n24522 , n24521 , n19424 );
and ( n24523 , n24131 , n19422 );
nor ( n24524 , n24522 , n24523 );
xnor ( n24525 , n24524 , n19431 );
and ( n24526 , n24520 , n24525 );
buf ( n24527 , n19327 );
and ( n24528 , n24527 , n19419 );
and ( n24529 , n24525 , n24528 );
and ( n24530 , n24520 , n24528 );
or ( n24531 , n24526 , n24529 , n24530 );
and ( n24532 , n24515 , n24531 );
and ( n24533 , n24499 , n24531 );
or ( n24534 , n24516 , n24532 , n24533 );
and ( n24535 , n19881 , n22048 );
and ( n24536 , n19825 , n22046 );
nor ( n24537 , n24535 , n24536 );
xnor ( n24538 , n24537 , n21853 );
xor ( n24539 , n24147 , n24151 );
xor ( n24540 , n24539 , n24156 );
and ( n24541 , n24538 , n24540 );
and ( n24542 , n22235 , n19805 );
and ( n24543 , n21955 , n19803 );
nor ( n24544 , n24542 , n24543 );
xnor ( n24545 , n24544 , n19750 );
and ( n24546 , n22425 , n19688 );
and ( n24547 , n22198 , n19686 );
nor ( n24548 , n24546 , n24547 );
xnor ( n24549 , n24548 , n19655 );
xor ( n24550 , n24545 , n24549 );
and ( n24551 , n24521 , n19419 );
xor ( n24552 , n24550 , n24551 );
and ( n24553 , n24540 , n24552 );
and ( n24554 , n24538 , n24552 );
or ( n24555 , n24541 , n24553 , n24554 );
and ( n24556 , n24534 , n24555 );
xor ( n24557 , n24159 , n24163 );
xor ( n24558 , n24557 , n24168 );
and ( n24559 , n24555 , n24558 );
and ( n24560 , n24534 , n24558 );
or ( n24561 , n24556 , n24559 , n24560 );
and ( n24562 , n19469 , n23944 );
and ( n24563 , n19434 , n23942 );
nor ( n24564 , n24562 , n24563 );
xnor ( n24565 , n24564 , n23550 );
and ( n24566 , n19605 , n23230 );
and ( n24567 , n19588 , n23228 );
nor ( n24568 , n24566 , n24567 );
xnor ( n24569 , n24568 , n22842 );
and ( n24570 , n24565 , n24569 );
and ( n24571 , n19721 , n22859 );
and ( n24572 , n19637 , n22857 );
nor ( n24573 , n24571 , n24572 );
xnor ( n24574 , n24573 , n22418 );
and ( n24575 , n24569 , n24574 );
and ( n24576 , n24565 , n24574 );
or ( n24577 , n24570 , n24575 , n24576 );
and ( n24578 , n22916 , n19688 );
and ( n24579 , n22756 , n19686 );
nor ( n24580 , n24578 , n24579 );
xnor ( n24581 , n24580 , n19655 );
buf ( n24582 , n24581 );
and ( n24583 , n21218 , n20460 );
and ( n24584 , n21072 , n20458 );
nor ( n24585 , n24583 , n24584 );
xnor ( n24586 , n24585 , n20337 );
and ( n24587 , n24582 , n24586 );
and ( n24588 , n21451 , n20276 );
and ( n24589 , n21302 , n20274 );
nor ( n24590 , n24588 , n24589 );
xnor ( n24591 , n24590 , n20175 );
and ( n24592 , n24586 , n24591 );
and ( n24593 , n24582 , n24591 );
or ( n24594 , n24587 , n24592 , n24593 );
and ( n24595 , n24577 , n24594 );
and ( n24596 , n23271 , n19596 );
and ( n24597 , n23141 , n19594 );
nor ( n24598 , n24596 , n24597 );
xnor ( n24599 , n24598 , n19545 );
and ( n24600 , n23573 , n19518 );
and ( n24601 , n23381 , n19516 );
nor ( n24602 , n24600 , n24601 );
xnor ( n24603 , n24602 , n19489 );
and ( n24604 , n24599 , n24603 );
and ( n24605 , n24131 , n19459 );
and ( n24606 , n23968 , n19457 );
nor ( n24607 , n24605 , n24606 );
xnor ( n24608 , n24607 , n19416 );
and ( n24609 , n24603 , n24608 );
and ( n24610 , n24599 , n24608 );
or ( n24611 , n24604 , n24609 , n24610 );
and ( n24612 , n22425 , n19805 );
and ( n24613 , n22198 , n19803 );
nor ( n24614 , n24612 , n24613 );
xnor ( n24615 , n24614 , n19750 );
and ( n24616 , n24527 , n19424 );
and ( n24617 , n24521 , n19422 );
nor ( n24618 , n24616 , n24617 );
xnor ( n24619 , n24618 , n19431 );
and ( n24620 , n24615 , n24619 );
buf ( n24621 , n19328 );
and ( n24622 , n24621 , n19419 );
and ( n24623 , n24619 , n24622 );
and ( n24624 , n24615 , n24622 );
or ( n24625 , n24620 , n24623 , n24624 );
and ( n24626 , n24611 , n24625 );
and ( n24627 , n19825 , n22381 );
and ( n24628 , n19811 , n22379 );
nor ( n24629 , n24627 , n24628 );
xnor ( n24630 , n24629 , n22228 );
and ( n24631 , n24625 , n24630 );
and ( n24632 , n24611 , n24630 );
or ( n24633 , n24626 , n24631 , n24632 );
and ( n24634 , n24594 , n24633 );
and ( n24635 , n24577 , n24633 );
or ( n24636 , n24595 , n24634 , n24635 );
xor ( n24637 , n24360 , n24364 );
xor ( n24638 , n24637 , n24369 );
and ( n24639 , n20182 , n21468 );
and ( n24640 , n20080 , n21466 );
nor ( n24641 , n24639 , n24640 );
xnor ( n24642 , n24641 , n21331 );
and ( n24643 , n20360 , n21155 );
and ( n24644 , n20268 , n21153 );
nor ( n24645 , n24643 , n24644 );
xnor ( n24646 , n24645 , n20994 );
xor ( n24647 , n24642 , n24646 );
and ( n24648 , n21876 , n19894 );
and ( n24649 , n21704 , n19892 );
nor ( n24650 , n24648 , n24649 );
xnor ( n24651 , n24650 , n19858 );
xor ( n24652 , n24647 , n24651 );
and ( n24653 , n24638 , n24652 );
and ( n24654 , n20618 , n20955 );
and ( n24655 , n20452 , n20953 );
nor ( n24656 , n24654 , n24655 );
xnor ( n24657 , n24656 , n20780 );
and ( n24658 , n20803 , n20674 );
and ( n24659 , n20666 , n20672 );
nor ( n24660 , n24658 , n24659 );
xnor ( n24661 , n24660 , n20542 );
xor ( n24662 , n24657 , n24661 );
not ( n24663 , n24259 );
xor ( n24664 , n24662 , n24663 );
and ( n24665 , n24652 , n24664 );
and ( n24666 , n24638 , n24664 );
or ( n24667 , n24653 , n24665 , n24666 );
and ( n24668 , n24636 , n24667 );
xor ( n24669 , n24223 , n24225 );
xor ( n24670 , n24669 , n24228 );
and ( n24671 , n24667 , n24670 );
and ( n24672 , n24636 , n24670 );
or ( n24673 , n24668 , n24671 , n24672 );
and ( n24674 , n24561 , n24673 );
xor ( n24675 , n24437 , n24461 );
xor ( n24676 , n24675 , n24464 );
and ( n24677 , n24673 , n24676 );
and ( n24678 , n24561 , n24676 );
or ( n24679 , n24674 , n24677 , n24678 );
xor ( n24680 , n24322 , n24324 );
xor ( n24681 , n24680 , n24327 );
and ( n24682 , n24679 , n24681 );
and ( n24683 , n24545 , n24549 );
and ( n24684 , n24549 , n24551 );
and ( n24685 , n24545 , n24551 );
or ( n24686 , n24683 , n24684 , n24685 );
and ( n24687 , n24642 , n24646 );
and ( n24688 , n24646 , n24651 );
and ( n24689 , n24642 , n24651 );
or ( n24690 , n24687 , n24688 , n24689 );
and ( n24691 , n24686 , n24690 );
and ( n24692 , n24657 , n24661 );
and ( n24693 , n24661 , n24663 );
and ( n24694 , n24657 , n24663 );
or ( n24695 , n24692 , n24693 , n24694 );
and ( n24696 , n24690 , n24695 );
and ( n24697 , n24686 , n24695 );
or ( n24698 , n24691 , n24696 , n24697 );
xor ( n24699 , n24288 , n24292 );
xor ( n24700 , n24699 , n24297 );
xor ( n24701 , n24243 , n24247 );
xor ( n24702 , n24701 , n24252 );
and ( n24703 , n24700 , n24702 );
xor ( n24704 , n24260 , n24264 );
xor ( n24705 , n24704 , n24269 );
and ( n24706 , n24702 , n24705 );
and ( n24707 , n24700 , n24705 );
or ( n24708 , n24703 , n24706 , n24707 );
and ( n24709 , n24698 , n24708 );
xor ( n24710 , n24255 , n24272 );
xor ( n24711 , n24710 , n24275 );
and ( n24712 , n24708 , n24711 );
and ( n24713 , n24698 , n24711 );
or ( n24714 , n24709 , n24712 , n24713 );
xor ( n24715 , n24099 , n24101 );
xor ( n24716 , n24715 , n24104 );
xor ( n24717 , n24714 , n24716 );
xor ( n24718 , n24143 , n24179 );
xor ( n24719 , n24718 , n24182 );
xor ( n24720 , n24717 , n24719 );
and ( n24721 , n24681 , n24720 );
and ( n24722 , n24679 , n24720 );
or ( n24723 , n24682 , n24721 , n24722 );
and ( n24724 , n24483 , n24723 );
xor ( n24725 , n24284 , n24330 );
xor ( n24726 , n24725 , n24333 );
and ( n24727 , n24723 , n24726 );
and ( n24728 , n24483 , n24726 );
or ( n24729 , n24724 , n24727 , n24728 );
and ( n24730 , n24714 , n24716 );
and ( n24731 , n24716 , n24719 );
and ( n24732 , n24714 , n24719 );
or ( n24733 , n24730 , n24731 , n24732 );
xor ( n24734 , n24107 , n24109 );
xor ( n24735 , n24734 , n24112 );
and ( n24736 , n24733 , n24735 );
xor ( n24737 , n24185 , n24187 );
xor ( n24738 , n24737 , n24190 );
and ( n24739 , n24735 , n24738 );
and ( n24740 , n24733 , n24738 );
or ( n24741 , n24736 , n24739 , n24740 );
and ( n24742 , n24729 , n24741 );
xor ( n24743 , n24336 , n24338 );
xor ( n24744 , n24743 , n24341 );
and ( n24745 , n24741 , n24744 );
and ( n24746 , n24729 , n24744 );
or ( n24747 , n24742 , n24745 , n24746 );
and ( n24748 , n24356 , n24747 );
xor ( n24749 , n24356 , n24747 );
xor ( n24750 , n24729 , n24741 );
xor ( n24751 , n24750 , n24744 );
and ( n24752 , n19418 , n24376 );
and ( n24753 , n19426 , n24374 );
nor ( n24754 , n24752 , n24753 );
xnor ( n24755 , n24754 , n23927 );
and ( n24756 , n19510 , n23641 );
and ( n24757 , n19496 , n23639 );
nor ( n24758 , n24756 , n24757 );
xnor ( n24759 , n24758 , n23213 );
and ( n24760 , n24755 , n24759 );
and ( n24761 , n19946 , n22048 );
and ( n24762 , n19881 , n22046 );
nor ( n24763 , n24761 , n24762 );
xnor ( n24764 , n24763 , n21853 );
and ( n24765 , n24759 , n24764 );
and ( n24766 , n24755 , n24764 );
or ( n24767 , n24760 , n24765 , n24766 );
xor ( n24768 , n24379 , n24383 );
xor ( n24769 , n24768 , n24388 );
and ( n24770 , n24767 , n24769 );
xor ( n24771 , n24410 , n24426 );
xor ( n24772 , n24771 , n24431 );
and ( n24773 , n24769 , n24772 );
and ( n24774 , n24767 , n24772 );
or ( n24775 , n24770 , n24773 , n24774 );
xor ( n24776 , n24686 , n24690 );
xor ( n24777 , n24776 , n24695 );
and ( n24778 , n24775 , n24777 );
xor ( n24779 , n24453 , n24455 );
xor ( n24780 , n24779 , n24458 );
and ( n24781 , n24777 , n24780 );
and ( n24782 , n24775 , n24780 );
or ( n24783 , n24778 , n24781 , n24782 );
xor ( n24784 , n24698 , n24708 );
xor ( n24785 , n24784 , n24711 );
and ( n24786 , n24783 , n24785 );
xor ( n24787 , n24469 , n24471 );
xor ( n24788 , n24787 , n24474 );
and ( n24789 , n24785 , n24788 );
and ( n24790 , n24783 , n24788 );
or ( n24791 , n24786 , n24789 , n24790 );
and ( n24792 , n20182 , n21741 );
and ( n24793 , n20080 , n21739 );
nor ( n24794 , n24792 , n24793 );
xnor ( n24795 , n24794 , n21605 );
and ( n24796 , n21876 , n20114 );
and ( n24797 , n21704 , n20112 );
nor ( n24798 , n24796 , n24797 );
xnor ( n24799 , n24798 , n19997 );
and ( n24800 , n24795 , n24799 );
and ( n24801 , n22235 , n19894 );
and ( n24802 , n21955 , n19892 );
nor ( n24803 , n24801 , n24802 );
xnor ( n24804 , n24803 , n19858 );
and ( n24805 , n24799 , n24804 );
and ( n24806 , n24795 , n24804 );
or ( n24807 , n24800 , n24805 , n24806 );
and ( n24808 , n20360 , n21468 );
and ( n24809 , n20268 , n21466 );
nor ( n24810 , n24808 , n24809 );
xnor ( n24811 , n24810 , n21331 );
and ( n24812 , n20618 , n21155 );
and ( n24813 , n20452 , n21153 );
nor ( n24814 , n24812 , n24813 );
xnor ( n24815 , n24814 , n20994 );
and ( n24816 , n24811 , n24815 );
and ( n24817 , n20803 , n20955 );
and ( n24818 , n20666 , n20953 );
nor ( n24819 , n24817 , n24818 );
xnor ( n24820 , n24819 , n20780 );
and ( n24821 , n24815 , n24820 );
and ( n24822 , n24811 , n24820 );
or ( n24823 , n24816 , n24821 , n24822 );
and ( n24824 , n24807 , n24823 );
and ( n24825 , n21072 , n20674 );
and ( n24826 , n20867 , n20672 );
nor ( n24827 , n24825 , n24826 );
xnor ( n24828 , n24827 , n20542 );
and ( n24829 , n21302 , n20460 );
and ( n24830 , n21218 , n20458 );
nor ( n24831 , n24829 , n24830 );
xnor ( n24832 , n24831 , n20337 );
and ( n24833 , n24828 , n24832 );
not ( n24834 , n24581 );
and ( n24835 , n24832 , n24834 );
and ( n24836 , n24828 , n24834 );
or ( n24837 , n24833 , n24835 , n24836 );
and ( n24838 , n24823 , n24837 );
and ( n24839 , n24807 , n24837 );
or ( n24840 , n24824 , n24838 , n24839 );
xor ( n24841 , n24398 , n24402 );
xor ( n24842 , n24841 , n24407 );
xor ( n24843 , n24414 , n24418 );
xor ( n24844 , n24843 , n24423 );
and ( n24845 , n24842 , n24844 );
xor ( n24846 , n24520 , n24525 );
xor ( n24847 , n24846 , n24528 );
and ( n24848 , n24844 , n24847 );
and ( n24849 , n24842 , n24847 );
or ( n24850 , n24845 , n24848 , n24849 );
and ( n24851 , n24840 , n24850 );
xor ( n24852 , n24441 , n24445 );
xor ( n24853 , n24852 , n24450 );
and ( n24854 , n24850 , n24853 );
and ( n24855 , n24840 , n24853 );
or ( n24856 , n24851 , n24854 , n24855 );
xor ( n24857 , n24372 , n24391 );
xor ( n24858 , n24857 , n24434 );
and ( n24859 , n24856 , n24858 );
xor ( n24860 , n24700 , n24702 );
xor ( n24861 , n24860 , n24705 );
and ( n24862 , n24858 , n24861 );
and ( n24863 , n24856 , n24861 );
or ( n24864 , n24859 , n24862 , n24863 );
and ( n24865 , n19588 , n23641 );
and ( n24866 , n19510 , n23639 );
nor ( n24867 , n24865 , n24866 );
xnor ( n24868 , n24867 , n23213 );
and ( n24869 , n19637 , n23230 );
and ( n24870 , n19605 , n23228 );
nor ( n24871 , n24869 , n24870 );
xnor ( n24872 , n24871 , n22842 );
and ( n24873 , n24868 , n24872 );
and ( n24874 , n19811 , n22859 );
and ( n24875 , n19721 , n22857 );
nor ( n24876 , n24874 , n24875 );
xnor ( n24877 , n24876 , n22418 );
and ( n24878 , n24872 , n24877 );
and ( n24879 , n24868 , n24877 );
or ( n24880 , n24873 , n24878 , n24879 );
buf ( n24881 , n19394 );
buf ( n24882 , n19395 );
and ( n24883 , n24881 , n24882 );
not ( n24884 , n24883 );
and ( n24885 , n24394 , n24884 );
not ( n24886 , n24885 );
and ( n24887 , n22198 , n19894 );
and ( n24888 , n22235 , n19892 );
nor ( n24889 , n24887 , n24888 );
xnor ( n24890 , n24889 , n19858 );
and ( n24891 , n24886 , n24890 );
and ( n24892 , n22756 , n19805 );
and ( n24893 , n22425 , n19803 );
nor ( n24894 , n24892 , n24893 );
xnor ( n24895 , n24894 , n19750 );
and ( n24896 , n24890 , n24895 );
and ( n24897 , n24886 , n24895 );
or ( n24898 , n24891 , n24896 , n24897 );
xor ( n24899 , n23924 , n24393 );
xor ( n24900 , n24393 , n24394 );
not ( n24901 , n24900 );
and ( n24902 , n24899 , n24901 );
and ( n24903 , n19426 , n24902 );
not ( n24904 , n24903 );
xnor ( n24905 , n24904 , n24397 );
and ( n24906 , n24898 , n24905 );
and ( n24907 , n19496 , n23944 );
and ( n24908 , n19469 , n23942 );
nor ( n24909 , n24907 , n24908 );
xnor ( n24910 , n24909 , n23550 );
and ( n24911 , n24905 , n24910 );
and ( n24912 , n24898 , n24910 );
or ( n24913 , n24906 , n24911 , n24912 );
and ( n24914 , n24880 , n24913 );
and ( n24915 , n23141 , n19688 );
and ( n24916 , n22916 , n19686 );
nor ( n24917 , n24915 , n24916 );
xnor ( n24918 , n24917 , n19655 );
and ( n24919 , n23381 , n19596 );
and ( n24920 , n23271 , n19594 );
nor ( n24921 , n24919 , n24920 );
xnor ( n24922 , n24921 , n19545 );
and ( n24923 , n24918 , n24922 );
and ( n24924 , n23968 , n19518 );
and ( n24925 , n23573 , n19516 );
nor ( n24926 , n24924 , n24925 );
xnor ( n24927 , n24926 , n19489 );
and ( n24928 , n24922 , n24927 );
and ( n24929 , n24918 , n24927 );
or ( n24930 , n24923 , n24928 , n24929 );
and ( n24931 , n24521 , n19459 );
and ( n24932 , n24131 , n19457 );
nor ( n24933 , n24931 , n24932 );
xnor ( n24934 , n24933 , n19416 );
and ( n24935 , n24621 , n19424 );
and ( n24936 , n24527 , n19422 );
nor ( n24937 , n24935 , n24936 );
xnor ( n24938 , n24937 , n19431 );
and ( n24939 , n24934 , n24938 );
buf ( n24940 , n19329 );
and ( n24941 , n24940 , n19419 );
and ( n24942 , n24938 , n24941 );
and ( n24943 , n24934 , n24941 );
or ( n24944 , n24939 , n24942 , n24943 );
and ( n24945 , n24930 , n24944 );
and ( n24946 , n19881 , n22381 );
and ( n24947 , n19825 , n22379 );
nor ( n24948 , n24946 , n24947 );
xnor ( n24949 , n24948 , n22228 );
and ( n24950 , n24944 , n24949 );
and ( n24951 , n24930 , n24949 );
or ( n24952 , n24945 , n24950 , n24951 );
and ( n24953 , n24913 , n24952 );
and ( n24954 , n24880 , n24952 );
or ( n24955 , n24914 , n24953 , n24954 );
xor ( n24956 , n24487 , n24491 );
xor ( n24957 , n24956 , n24496 );
xor ( n24958 , n24503 , n24507 );
xor ( n24959 , n24958 , n24512 );
and ( n24960 , n24957 , n24959 );
xor ( n24961 , n24582 , n24586 );
xor ( n24962 , n24961 , n24591 );
and ( n24963 , n24959 , n24962 );
and ( n24964 , n24957 , n24962 );
or ( n24965 , n24960 , n24963 , n24964 );
and ( n24966 , n24955 , n24965 );
xor ( n24967 , n24538 , n24540 );
xor ( n24968 , n24967 , n24552 );
and ( n24969 , n24965 , n24968 );
and ( n24970 , n24955 , n24968 );
or ( n24971 , n24966 , n24969 , n24970 );
xor ( n24972 , n24499 , n24515 );
xor ( n24973 , n24972 , n24531 );
xor ( n24974 , n24577 , n24594 );
xor ( n24975 , n24974 , n24633 );
and ( n24976 , n24973 , n24975 );
xor ( n24977 , n24638 , n24652 );
xor ( n24978 , n24977 , n24664 );
and ( n24979 , n24975 , n24978 );
and ( n24980 , n24973 , n24978 );
or ( n24981 , n24976 , n24979 , n24980 );
and ( n24982 , n24971 , n24981 );
xor ( n24983 , n24534 , n24555 );
xor ( n24984 , n24983 , n24558 );
and ( n24985 , n24981 , n24984 );
and ( n24986 , n24971 , n24984 );
or ( n24987 , n24982 , n24985 , n24986 );
and ( n24988 , n24864 , n24987 );
xor ( n24989 , n24561 , n24673 );
xor ( n24990 , n24989 , n24676 );
and ( n24991 , n24987 , n24990 );
and ( n24992 , n24864 , n24990 );
or ( n24993 , n24988 , n24991 , n24992 );
and ( n24994 , n24791 , n24993 );
xor ( n24995 , n24467 , n24477 );
xor ( n24996 , n24995 , n24480 );
and ( n24997 , n24993 , n24996 );
and ( n24998 , n24791 , n24996 );
or ( n24999 , n24994 , n24997 , n24998 );
xor ( n25000 , n24483 , n24723 );
xor ( n25001 , n25000 , n24726 );
and ( n25002 , n24999 , n25001 );
xor ( n25003 , n24733 , n24735 );
xor ( n25004 , n25003 , n24738 );
and ( n25005 , n25001 , n25004 );
and ( n25006 , n24999 , n25004 );
or ( n25007 , n25002 , n25005 , n25006 );
and ( n25008 , n24751 , n25007 );
xor ( n25009 , n24751 , n25007 );
xor ( n25010 , n24999 , n25001 );
xor ( n25011 , n25010 , n25004 );
and ( n25012 , n19434 , n24376 );
and ( n25013 , n19418 , n24374 );
nor ( n25014 , n25012 , n25013 );
xnor ( n25015 , n25014 , n23927 );
and ( n25016 , n20004 , n22048 );
and ( n25017 , n19946 , n22046 );
nor ( n25018 , n25016 , n25017 );
xnor ( n25019 , n25018 , n21853 );
and ( n25020 , n25015 , n25019 );
and ( n25021 , n21612 , n20276 );
and ( n25022 , n21451 , n20274 );
nor ( n25023 , n25021 , n25022 );
xnor ( n25024 , n25023 , n20175 );
and ( n25025 , n25019 , n25024 );
and ( n25026 , n25015 , n25024 );
or ( n25027 , n25020 , n25025 , n25026 );
xor ( n25028 , n24565 , n24569 );
xor ( n25029 , n25028 , n24574 );
and ( n25030 , n25027 , n25029 );
xor ( n25031 , n24611 , n24625 );
xor ( n25032 , n25031 , n24630 );
and ( n25033 , n25029 , n25032 );
and ( n25034 , n25027 , n25032 );
or ( n25035 , n25030 , n25033 , n25034 );
and ( n25036 , n22916 , n19805 );
and ( n25037 , n22756 , n19803 );
nor ( n25038 , n25036 , n25037 );
xnor ( n25039 , n25038 , n19750 );
buf ( n25040 , n25039 );
and ( n25041 , n20867 , n20955 );
and ( n25042 , n20803 , n20953 );
nor ( n25043 , n25041 , n25042 );
xnor ( n25044 , n25043 , n20780 );
and ( n25045 , n25040 , n25044 );
and ( n25046 , n21218 , n20674 );
and ( n25047 , n21072 , n20672 );
nor ( n25048 , n25046 , n25047 );
xnor ( n25049 , n25048 , n20542 );
and ( n25050 , n25044 , n25049 );
and ( n25051 , n25040 , n25049 );
or ( n25052 , n25045 , n25050 , n25051 );
xor ( n25053 , n24599 , n24603 );
xor ( n25054 , n25053 , n24608 );
and ( n25055 , n25052 , n25054 );
xor ( n25056 , n24615 , n24619 );
xor ( n25057 , n25056 , n24622 );
and ( n25058 , n25054 , n25057 );
and ( n25059 , n25052 , n25057 );
or ( n25060 , n25055 , n25058 , n25059 );
xor ( n25061 , n24755 , n24759 );
xor ( n25062 , n25061 , n24764 );
and ( n25063 , n25060 , n25062 );
xor ( n25064 , n24842 , n24844 );
xor ( n25065 , n25064 , n24847 );
and ( n25066 , n25062 , n25065 );
and ( n25067 , n25060 , n25065 );
or ( n25068 , n25063 , n25066 , n25067 );
and ( n25069 , n25035 , n25068 );
xor ( n25070 , n24767 , n24769 );
xor ( n25071 , n25070 , n24772 );
and ( n25072 , n25068 , n25071 );
and ( n25073 , n25035 , n25071 );
or ( n25074 , n25069 , n25072 , n25073 );
xor ( n25075 , n24636 , n24667 );
xor ( n25076 , n25075 , n24670 );
and ( n25077 , n25074 , n25076 );
xor ( n25078 , n24856 , n24858 );
xor ( n25079 , n25078 , n24861 );
and ( n25080 , n25076 , n25079 );
and ( n25081 , n25074 , n25079 );
or ( n25082 , n25077 , n25080 , n25081 );
and ( n25083 , n20080 , n22048 );
and ( n25084 , n20004 , n22046 );
nor ( n25085 , n25083 , n25084 );
xnor ( n25086 , n25085 , n21853 );
and ( n25087 , n21704 , n20276 );
and ( n25088 , n21612 , n20274 );
nor ( n25089 , n25087 , n25088 );
xnor ( n25090 , n25089 , n20175 );
and ( n25091 , n25086 , n25090 );
and ( n25092 , n21955 , n20114 );
and ( n25093 , n21876 , n20112 );
nor ( n25094 , n25092 , n25093 );
xnor ( n25095 , n25094 , n19997 );
and ( n25096 , n25090 , n25095 );
and ( n25097 , n25086 , n25095 );
or ( n25098 , n25091 , n25096 , n25097 );
and ( n25099 , n20268 , n21741 );
and ( n25100 , n20182 , n21739 );
nor ( n25101 , n25099 , n25100 );
xnor ( n25102 , n25101 , n21605 );
and ( n25103 , n20452 , n21468 );
and ( n25104 , n20360 , n21466 );
nor ( n25105 , n25103 , n25104 );
xnor ( n25106 , n25105 , n21331 );
and ( n25107 , n25102 , n25106 );
and ( n25108 , n20666 , n21155 );
and ( n25109 , n20618 , n21153 );
nor ( n25110 , n25108 , n25109 );
xnor ( n25111 , n25110 , n20994 );
and ( n25112 , n25106 , n25111 );
and ( n25113 , n25102 , n25111 );
or ( n25114 , n25107 , n25112 , n25113 );
and ( n25115 , n25098 , n25114 );
and ( n25116 , n19418 , n24902 );
and ( n25117 , n19426 , n24900 );
nor ( n25118 , n25116 , n25117 );
xnor ( n25119 , n25118 , n24397 );
and ( n25120 , n19946 , n22381 );
and ( n25121 , n19881 , n22379 );
nor ( n25122 , n25120 , n25121 );
xnor ( n25123 , n25122 , n22228 );
and ( n25124 , n25119 , n25123 );
and ( n25125 , n21451 , n20460 );
and ( n25126 , n21302 , n20458 );
nor ( n25127 , n25125 , n25126 );
xnor ( n25128 , n25127 , n20337 );
and ( n25129 , n25123 , n25128 );
and ( n25130 , n25119 , n25128 );
or ( n25131 , n25124 , n25129 , n25130 );
and ( n25132 , n25114 , n25131 );
and ( n25133 , n25098 , n25131 );
or ( n25134 , n25115 , n25132 , n25133 );
and ( n25135 , n19510 , n23944 );
and ( n25136 , n19496 , n23942 );
nor ( n25137 , n25135 , n25136 );
xnor ( n25138 , n25137 , n23550 );
and ( n25139 , n19605 , n23641 );
and ( n25140 , n19588 , n23639 );
nor ( n25141 , n25139 , n25140 );
xnor ( n25142 , n25141 , n23213 );
and ( n25143 , n25138 , n25142 );
and ( n25144 , n19721 , n23230 );
and ( n25145 , n19637 , n23228 );
nor ( n25146 , n25144 , n25145 );
xnor ( n25147 , n25146 , n22842 );
and ( n25148 , n25142 , n25147 );
and ( n25149 , n25138 , n25147 );
or ( n25150 , n25143 , n25148 , n25149 );
and ( n25151 , n23271 , n19688 );
and ( n25152 , n23141 , n19686 );
nor ( n25153 , n25151 , n25152 );
xnor ( n25154 , n25153 , n19655 );
and ( n25155 , n23573 , n19596 );
and ( n25156 , n23381 , n19594 );
nor ( n25157 , n25155 , n25156 );
xnor ( n25158 , n25157 , n19545 );
and ( n25159 , n25154 , n25158 );
and ( n25160 , n24131 , n19518 );
and ( n25161 , n23968 , n19516 );
nor ( n25162 , n25160 , n25161 );
xnor ( n25163 , n25162 , n19489 );
and ( n25164 , n25158 , n25163 );
and ( n25165 , n25154 , n25163 );
or ( n25166 , n25159 , n25164 , n25165 );
and ( n25167 , n19469 , n24376 );
and ( n25168 , n19434 , n24374 );
nor ( n25169 , n25167 , n25168 );
xnor ( n25170 , n25169 , n23927 );
and ( n25171 , n25166 , n25170 );
and ( n25172 , n19825 , n22859 );
and ( n25173 , n19811 , n22857 );
nor ( n25174 , n25172 , n25173 );
xnor ( n25175 , n25174 , n22418 );
and ( n25176 , n25170 , n25175 );
and ( n25177 , n25166 , n25175 );
or ( n25178 , n25171 , n25176 , n25177 );
and ( n25179 , n25150 , n25178 );
xor ( n25180 , n24828 , n24832 );
xor ( n25181 , n25180 , n24834 );
and ( n25182 , n25178 , n25181 );
and ( n25183 , n25150 , n25181 );
or ( n25184 , n25179 , n25182 , n25183 );
and ( n25185 , n25134 , n25184 );
xor ( n25186 , n24807 , n24823 );
xor ( n25187 , n25186 , n24837 );
and ( n25188 , n25184 , n25187 );
and ( n25189 , n25134 , n25187 );
or ( n25190 , n25185 , n25188 , n25189 );
xor ( n25191 , n24840 , n24850 );
xor ( n25192 , n25191 , n24853 );
and ( n25193 , n25190 , n25192 );
xor ( n25194 , n24955 , n24965 );
xor ( n25195 , n25194 , n24968 );
and ( n25196 , n25192 , n25195 );
and ( n25197 , n25190 , n25195 );
or ( n25198 , n25193 , n25196 , n25197 );
xor ( n25199 , n24775 , n24777 );
xor ( n25200 , n25199 , n24780 );
and ( n25201 , n25198 , n25200 );
xor ( n25202 , n24971 , n24981 );
xor ( n25203 , n25202 , n24984 );
and ( n25204 , n25200 , n25203 );
and ( n25205 , n25198 , n25203 );
or ( n25206 , n25201 , n25204 , n25205 );
and ( n25207 , n25082 , n25206 );
xor ( n25208 , n24783 , n24785 );
xor ( n25209 , n25208 , n24788 );
and ( n25210 , n25206 , n25209 );
and ( n25211 , n25082 , n25209 );
or ( n25212 , n25207 , n25210 , n25211 );
xor ( n25213 , n24679 , n24681 );
xor ( n25214 , n25213 , n24720 );
and ( n25215 , n25212 , n25214 );
xor ( n25216 , n24791 , n24993 );
xor ( n25217 , n25216 , n24996 );
and ( n25218 , n25214 , n25217 );
and ( n25219 , n25212 , n25217 );
or ( n25220 , n25215 , n25218 , n25219 );
and ( n25221 , n25011 , n25220 );
xor ( n25222 , n25011 , n25220 );
xor ( n25223 , n25212 , n25214 );
xor ( n25224 , n25223 , n25217 );
and ( n25225 , n22425 , n19894 );
and ( n25226 , n22198 , n19892 );
nor ( n25227 , n25225 , n25226 );
xnor ( n25228 , n25227 , n19858 );
and ( n25229 , n24527 , n19459 );
and ( n25230 , n24521 , n19457 );
nor ( n25231 , n25229 , n25230 );
xnor ( n25232 , n25231 , n19416 );
and ( n25233 , n25228 , n25232 );
and ( n25234 , n24940 , n19424 );
and ( n25235 , n24621 , n19422 );
nor ( n25236 , n25234 , n25235 );
xnor ( n25237 , n25236 , n19431 );
and ( n25238 , n25232 , n25237 );
and ( n25239 , n25228 , n25237 );
or ( n25240 , n25233 , n25238 , n25239 );
xor ( n25241 , n24886 , n24890 );
xor ( n25242 , n25241 , n24895 );
and ( n25243 , n25240 , n25242 );
xor ( n25244 , n24934 , n24938 );
xor ( n25245 , n25244 , n24941 );
and ( n25246 , n25242 , n25245 );
and ( n25247 , n25240 , n25245 );
or ( n25248 , n25243 , n25246 , n25247 );
xor ( n25249 , n25015 , n25019 );
xor ( n25250 , n25249 , n25024 );
and ( n25251 , n25248 , n25250 );
xor ( n25252 , n24930 , n24944 );
xor ( n25253 , n25252 , n24949 );
and ( n25254 , n25250 , n25253 );
and ( n25255 , n25248 , n25253 );
or ( n25256 , n25251 , n25254 , n25255 );
xor ( n25257 , n24880 , n24913 );
xor ( n25258 , n25257 , n24952 );
and ( n25259 , n25256 , n25258 );
xor ( n25260 , n24957 , n24959 );
xor ( n25261 , n25260 , n24962 );
and ( n25262 , n25258 , n25261 );
and ( n25263 , n25256 , n25261 );
or ( n25264 , n25259 , n25262 , n25263 );
xor ( n25265 , n24795 , n24799 );
xor ( n25266 , n25265 , n24804 );
xor ( n25267 , n24811 , n24815 );
xor ( n25268 , n25267 , n24820 );
and ( n25269 , n25266 , n25268 );
xor ( n25270 , n24898 , n24905 );
xor ( n25271 , n25270 , n24910 );
and ( n25272 , n25268 , n25271 );
and ( n25273 , n25266 , n25271 );
or ( n25274 , n25269 , n25272 , n25273 );
and ( n25275 , n21876 , n20276 );
and ( n25276 , n21704 , n20274 );
nor ( n25277 , n25275 , n25276 );
xnor ( n25278 , n25277 , n20175 );
and ( n25279 , n22235 , n20114 );
and ( n25280 , n21955 , n20112 );
nor ( n25281 , n25279 , n25280 );
xnor ( n25282 , n25281 , n19997 );
and ( n25283 , n25278 , n25282 );
buf ( n25284 , n19330 );
and ( n25285 , n25284 , n19419 );
and ( n25286 , n25282 , n25285 );
and ( n25287 , n25278 , n25285 );
or ( n25288 , n25283 , n25286 , n25287 );
and ( n25289 , n20182 , n22048 );
and ( n25290 , n20080 , n22046 );
nor ( n25291 , n25289 , n25290 );
xnor ( n25292 , n25291 , n21853 );
and ( n25293 , n20360 , n21741 );
and ( n25294 , n20268 , n21739 );
nor ( n25295 , n25293 , n25294 );
xnor ( n25296 , n25295 , n21605 );
and ( n25297 , n25292 , n25296 );
and ( n25298 , n20618 , n21468 );
and ( n25299 , n20452 , n21466 );
nor ( n25300 , n25298 , n25299 );
xnor ( n25301 , n25300 , n21331 );
and ( n25302 , n25296 , n25301 );
and ( n25303 , n25292 , n25301 );
or ( n25304 , n25297 , n25302 , n25303 );
and ( n25305 , n25288 , n25304 );
xor ( n25306 , n24918 , n24922 );
xor ( n25307 , n25306 , n24927 );
and ( n25308 , n25304 , n25307 );
and ( n25309 , n25288 , n25307 );
or ( n25310 , n25305 , n25308 , n25309 );
xor ( n25311 , n24868 , n24872 );
xor ( n25312 , n25311 , n24877 );
and ( n25313 , n25310 , n25312 );
xor ( n25314 , n25052 , n25054 );
xor ( n25315 , n25314 , n25057 );
and ( n25316 , n25312 , n25315 );
and ( n25317 , n25310 , n25315 );
or ( n25318 , n25313 , n25316 , n25317 );
and ( n25319 , n25274 , n25318 );
xor ( n25320 , n25027 , n25029 );
xor ( n25321 , n25320 , n25032 );
and ( n25322 , n25318 , n25321 );
and ( n25323 , n25274 , n25321 );
or ( n25324 , n25319 , n25322 , n25323 );
and ( n25325 , n25264 , n25324 );
xor ( n25326 , n24973 , n24975 );
xor ( n25327 , n25326 , n24978 );
and ( n25328 , n25324 , n25327 );
and ( n25329 , n25264 , n25327 );
or ( n25330 , n25325 , n25328 , n25329 );
and ( n25331 , n20004 , n22381 );
and ( n25332 , n19946 , n22379 );
nor ( n25333 , n25331 , n25332 );
xnor ( n25334 , n25333 , n22228 );
and ( n25335 , n21302 , n20674 );
and ( n25336 , n21218 , n20672 );
nor ( n25337 , n25335 , n25336 );
xnor ( n25338 , n25337 , n20542 );
and ( n25339 , n25334 , n25338 );
and ( n25340 , n21612 , n20460 );
and ( n25341 , n21451 , n20458 );
nor ( n25342 , n25340 , n25341 );
xnor ( n25343 , n25342 , n20337 );
and ( n25344 , n25338 , n25343 );
and ( n25345 , n25334 , n25343 );
or ( n25346 , n25339 , n25344 , n25345 );
and ( n25347 , n19434 , n24902 );
and ( n25348 , n19418 , n24900 );
nor ( n25349 , n25347 , n25348 );
xnor ( n25350 , n25349 , n24397 );
and ( n25351 , n19588 , n23944 );
and ( n25352 , n19510 , n23942 );
nor ( n25353 , n25351 , n25352 );
xnor ( n25354 , n25353 , n23550 );
and ( n25355 , n25350 , n25354 );
and ( n25356 , n19637 , n23641 );
and ( n25357 , n19605 , n23639 );
nor ( n25358 , n25356 , n25357 );
xnor ( n25359 , n25358 , n23213 );
and ( n25360 , n25354 , n25359 );
and ( n25361 , n25350 , n25359 );
or ( n25362 , n25355 , n25360 , n25361 );
and ( n25363 , n25346 , n25362 );
and ( n25364 , n20803 , n21155 );
and ( n25365 , n20666 , n21153 );
nor ( n25366 , n25364 , n25365 );
xnor ( n25367 , n25366 , n20994 );
and ( n25368 , n21072 , n20955 );
and ( n25369 , n20867 , n20953 );
nor ( n25370 , n25368 , n25369 );
xnor ( n25371 , n25370 , n20780 );
and ( n25372 , n25367 , n25371 );
not ( n25373 , n25039 );
and ( n25374 , n25371 , n25373 );
and ( n25375 , n25367 , n25373 );
or ( n25376 , n25372 , n25374 , n25375 );
and ( n25377 , n25362 , n25376 );
and ( n25378 , n25346 , n25376 );
or ( n25379 , n25363 , n25377 , n25378 );
xor ( n25380 , n24394 , n24881 );
xor ( n25381 , n24881 , n24882 );
not ( n25382 , n25381 );
and ( n25383 , n25380 , n25382 );
and ( n25384 , n19426 , n25383 );
not ( n25385 , n25384 );
xnor ( n25386 , n25385 , n24885 );
and ( n25387 , n19496 , n24376 );
and ( n25388 , n19469 , n24374 );
nor ( n25389 , n25387 , n25388 );
xnor ( n25390 , n25389 , n23927 );
and ( n25391 , n25386 , n25390 );
and ( n25392 , n19811 , n23230 );
and ( n25393 , n19721 , n23228 );
nor ( n25394 , n25392 , n25393 );
xnor ( n25395 , n25394 , n22842 );
and ( n25396 , n25390 , n25395 );
and ( n25397 , n25386 , n25395 );
or ( n25398 , n25391 , n25396 , n25397 );
xor ( n25399 , n25086 , n25090 );
xor ( n25400 , n25399 , n25095 );
and ( n25401 , n25398 , n25400 );
xor ( n25402 , n25040 , n25044 );
xor ( n25403 , n25402 , n25049 );
and ( n25404 , n25400 , n25403 );
and ( n25405 , n25398 , n25403 );
or ( n25406 , n25401 , n25404 , n25405 );
and ( n25407 , n25379 , n25406 );
xor ( n25408 , n25098 , n25114 );
xor ( n25409 , n25408 , n25131 );
and ( n25410 , n25406 , n25409 );
and ( n25411 , n25379 , n25409 );
or ( n25412 , n25407 , n25410 , n25411 );
xor ( n25413 , n25134 , n25184 );
xor ( n25414 , n25413 , n25187 );
and ( n25415 , n25412 , n25414 );
xor ( n25416 , n25060 , n25062 );
xor ( n25417 , n25416 , n25065 );
and ( n25418 , n25414 , n25417 );
and ( n25419 , n25412 , n25417 );
or ( n25420 , n25415 , n25418 , n25419 );
xor ( n25421 , n25035 , n25068 );
xor ( n25422 , n25421 , n25071 );
and ( n25423 , n25420 , n25422 );
xor ( n25424 , n25190 , n25192 );
xor ( n25425 , n25424 , n25195 );
and ( n25426 , n25422 , n25425 );
and ( n25427 , n25420 , n25425 );
or ( n25428 , n25423 , n25426 , n25427 );
and ( n25429 , n25330 , n25428 );
xor ( n25430 , n25074 , n25076 );
xor ( n25431 , n25430 , n25079 );
and ( n25432 , n25428 , n25431 );
and ( n25433 , n25330 , n25431 );
or ( n25434 , n25429 , n25432 , n25433 );
xor ( n25435 , n24864 , n24987 );
xor ( n25436 , n25435 , n24990 );
and ( n25437 , n25434 , n25436 );
xor ( n25438 , n25082 , n25206 );
xor ( n25439 , n25438 , n25209 );
and ( n25440 , n25436 , n25439 );
and ( n25441 , n25434 , n25439 );
or ( n25442 , n25437 , n25440 , n25441 );
and ( n25443 , n25224 , n25442 );
xor ( n25444 , n25224 , n25442 );
xor ( n25445 , n25434 , n25436 );
xor ( n25446 , n25445 , n25439 );
and ( n25447 , n24521 , n19518 );
and ( n25448 , n24131 , n19516 );
nor ( n25449 , n25447 , n25448 );
xnor ( n25450 , n25449 , n19489 );
and ( n25451 , n24621 , n19459 );
and ( n25452 , n24527 , n19457 );
nor ( n25453 , n25451 , n25452 );
xnor ( n25454 , n25453 , n19416 );
and ( n25455 , n25450 , n25454 );
and ( n25456 , n25284 , n19424 );
and ( n25457 , n24940 , n19422 );
nor ( n25458 , n25456 , n25457 );
xnor ( n25459 , n25458 , n19431 );
and ( n25460 , n25454 , n25459 );
and ( n25461 , n25450 , n25459 );
or ( n25462 , n25455 , n25460 , n25461 );
xor ( n25463 , n25154 , n25158 );
xor ( n25464 , n25463 , n25163 );
and ( n25465 , n25462 , n25464 );
xor ( n25466 , n25228 , n25232 );
xor ( n25467 , n25466 , n25237 );
and ( n25468 , n25464 , n25467 );
and ( n25469 , n25462 , n25467 );
or ( n25470 , n25465 , n25468 , n25469 );
xor ( n25471 , n25138 , n25142 );
xor ( n25472 , n25471 , n25147 );
and ( n25473 , n25470 , n25472 );
xor ( n25474 , n25166 , n25170 );
xor ( n25475 , n25474 , n25175 );
and ( n25476 , n25472 , n25475 );
and ( n25477 , n25470 , n25475 );
or ( n25478 , n25473 , n25476 , n25477 );
xor ( n25479 , n25150 , n25178 );
xor ( n25480 , n25479 , n25181 );
and ( n25481 , n25478 , n25480 );
xor ( n25482 , n25266 , n25268 );
xor ( n25483 , n25482 , n25271 );
and ( n25484 , n25480 , n25483 );
and ( n25485 , n25478 , n25483 );
or ( n25486 , n25481 , n25484 , n25485 );
xor ( n25487 , n25256 , n25258 );
xor ( n25488 , n25487 , n25261 );
and ( n25489 , n25486 , n25488 );
xor ( n25490 , n25274 , n25318 );
xor ( n25491 , n25490 , n25321 );
and ( n25492 , n25488 , n25491 );
and ( n25493 , n25486 , n25491 );
or ( n25494 , n25489 , n25492 , n25493 );
buf ( n25495 , n19396 );
buf ( n25496 , n19397 );
and ( n25497 , n25495 , n25496 );
not ( n25498 , n25497 );
and ( n25499 , n24882 , n25498 );
not ( n25500 , n25499 );
and ( n25501 , n22198 , n20114 );
and ( n25502 , n22235 , n20112 );
nor ( n25503 , n25501 , n25502 );
xnor ( n25504 , n25503 , n19997 );
and ( n25505 , n25500 , n25504 );
and ( n25506 , n22756 , n19894 );
and ( n25507 , n22425 , n19892 );
nor ( n25508 , n25506 , n25507 );
xnor ( n25509 , n25508 , n19858 );
and ( n25510 , n25504 , n25509 );
and ( n25511 , n25500 , n25509 );
or ( n25512 , n25505 , n25510 , n25511 );
and ( n25513 , n23141 , n19805 );
and ( n25514 , n22916 , n19803 );
nor ( n25515 , n25513 , n25514 );
xnor ( n25516 , n25515 , n19750 );
and ( n25517 , n23381 , n19688 );
and ( n25518 , n23271 , n19686 );
nor ( n25519 , n25517 , n25518 );
xnor ( n25520 , n25519 , n19655 );
and ( n25521 , n25516 , n25520 );
and ( n25522 , n23968 , n19596 );
and ( n25523 , n23573 , n19594 );
nor ( n25524 , n25522 , n25523 );
xnor ( n25525 , n25524 , n19545 );
and ( n25526 , n25520 , n25525 );
and ( n25527 , n25516 , n25525 );
or ( n25528 , n25521 , n25526 , n25527 );
and ( n25529 , n25512 , n25528 );
and ( n25530 , n19881 , n22859 );
and ( n25531 , n19825 , n22857 );
nor ( n25532 , n25530 , n25531 );
xnor ( n25533 , n25532 , n22418 );
and ( n25534 , n25528 , n25533 );
and ( n25535 , n25512 , n25533 );
or ( n25536 , n25529 , n25534 , n25535 );
xor ( n25537 , n25102 , n25106 );
xor ( n25538 , n25537 , n25111 );
and ( n25539 , n25536 , n25538 );
xor ( n25540 , n25119 , n25123 );
xor ( n25541 , n25540 , n25128 );
and ( n25542 , n25538 , n25541 );
and ( n25543 , n25536 , n25541 );
or ( n25544 , n25539 , n25542 , n25543 );
and ( n25545 , n20080 , n22381 );
and ( n25546 , n20004 , n22379 );
nor ( n25547 , n25545 , n25546 );
xnor ( n25548 , n25547 , n22228 );
and ( n25549 , n21955 , n20276 );
and ( n25550 , n21876 , n20274 );
nor ( n25551 , n25549 , n25550 );
xnor ( n25552 , n25551 , n20175 );
and ( n25553 , n25548 , n25552 );
buf ( n25554 , n19331 );
and ( n25555 , n25554 , n19419 );
and ( n25556 , n25552 , n25555 );
and ( n25557 , n25548 , n25555 );
or ( n25558 , n25553 , n25556 , n25557 );
and ( n25559 , n22916 , n19894 );
and ( n25560 , n22756 , n19892 );
nor ( n25561 , n25559 , n25560 );
xnor ( n25562 , n25561 , n19858 );
buf ( n25563 , n25562 );
and ( n25564 , n20666 , n21468 );
and ( n25565 , n20618 , n21466 );
nor ( n25566 , n25564 , n25565 );
xnor ( n25567 , n25566 , n21331 );
and ( n25568 , n25563 , n25567 );
and ( n25569 , n20867 , n21155 );
and ( n25570 , n20803 , n21153 );
nor ( n25571 , n25569 , n25570 );
xnor ( n25572 , n25571 , n20994 );
and ( n25573 , n25567 , n25572 );
and ( n25574 , n25563 , n25572 );
or ( n25575 , n25568 , n25573 , n25574 );
and ( n25576 , n25558 , n25575 );
xor ( n25577 , n25278 , n25282 );
xor ( n25578 , n25577 , n25285 );
and ( n25579 , n25575 , n25578 );
and ( n25580 , n25558 , n25578 );
or ( n25581 , n25576 , n25579 , n25580 );
xor ( n25582 , n25288 , n25304 );
xor ( n25583 , n25582 , n25307 );
and ( n25584 , n25581 , n25583 );
xor ( n25585 , n25240 , n25242 );
xor ( n25586 , n25585 , n25245 );
and ( n25587 , n25583 , n25586 );
and ( n25588 , n25581 , n25586 );
or ( n25589 , n25584 , n25587 , n25588 );
and ( n25590 , n25544 , n25589 );
xor ( n25591 , n25248 , n25250 );
xor ( n25592 , n25591 , n25253 );
and ( n25593 , n25589 , n25592 );
and ( n25594 , n25544 , n25592 );
or ( n25595 , n25590 , n25593 , n25594 );
and ( n25596 , n19946 , n22859 );
and ( n25597 , n19881 , n22857 );
nor ( n25598 , n25596 , n25597 );
xnor ( n25599 , n25598 , n22418 );
and ( n25600 , n21218 , n20955 );
and ( n25601 , n21072 , n20953 );
nor ( n25602 , n25600 , n25601 );
xnor ( n25603 , n25602 , n20780 );
and ( n25604 , n25599 , n25603 );
and ( n25605 , n21451 , n20674 );
and ( n25606 , n21302 , n20672 );
nor ( n25607 , n25605 , n25606 );
xnor ( n25608 , n25607 , n20542 );
and ( n25609 , n25603 , n25608 );
and ( n25610 , n25599 , n25608 );
or ( n25611 , n25604 , n25609 , n25610 );
and ( n25612 , n20268 , n22048 );
and ( n25613 , n20182 , n22046 );
nor ( n25614 , n25612 , n25613 );
xnor ( n25615 , n25614 , n21853 );
and ( n25616 , n20452 , n21741 );
and ( n25617 , n20360 , n21739 );
nor ( n25618 , n25616 , n25617 );
xnor ( n25619 , n25618 , n21605 );
and ( n25620 , n25615 , n25619 );
and ( n25621 , n21704 , n20460 );
and ( n25622 , n21612 , n20458 );
nor ( n25623 , n25621 , n25622 );
xnor ( n25624 , n25623 , n20337 );
and ( n25625 , n25619 , n25624 );
and ( n25626 , n25615 , n25624 );
or ( n25627 , n25620 , n25625 , n25626 );
and ( n25628 , n25611 , n25627 );
and ( n25629 , n19418 , n25383 );
and ( n25630 , n19426 , n25381 );
nor ( n25631 , n25629 , n25630 );
xnor ( n25632 , n25631 , n24885 );
and ( n25633 , n19510 , n24376 );
and ( n25634 , n19496 , n24374 );
nor ( n25635 , n25633 , n25634 );
xnor ( n25636 , n25635 , n23927 );
and ( n25637 , n25632 , n25636 );
and ( n25638 , n19605 , n23944 );
and ( n25639 , n19588 , n23942 );
nor ( n25640 , n25638 , n25639 );
xnor ( n25641 , n25640 , n23550 );
and ( n25642 , n25636 , n25641 );
and ( n25643 , n25632 , n25641 );
or ( n25644 , n25637 , n25642 , n25643 );
and ( n25645 , n25627 , n25644 );
and ( n25646 , n25611 , n25644 );
or ( n25647 , n25628 , n25645 , n25646 );
xor ( n25648 , n25334 , n25338 );
xor ( n25649 , n25648 , n25343 );
xor ( n25650 , n25292 , n25296 );
xor ( n25651 , n25650 , n25301 );
and ( n25652 , n25649 , n25651 );
xor ( n25653 , n25367 , n25371 );
xor ( n25654 , n25653 , n25373 );
and ( n25655 , n25651 , n25654 );
and ( n25656 , n25649 , n25654 );
or ( n25657 , n25652 , n25655 , n25656 );
and ( n25658 , n25647 , n25657 );
and ( n25659 , n23271 , n19805 );
and ( n25660 , n23141 , n19803 );
nor ( n25661 , n25659 , n25660 );
xnor ( n25662 , n25661 , n19750 );
and ( n25663 , n23573 , n19688 );
and ( n25664 , n23381 , n19686 );
nor ( n25665 , n25663 , n25664 );
xnor ( n25666 , n25665 , n19655 );
and ( n25667 , n25662 , n25666 );
and ( n25668 , n24131 , n19596 );
and ( n25669 , n23968 , n19594 );
nor ( n25670 , n25668 , n25669 );
xnor ( n25671 , n25670 , n19545 );
and ( n25672 , n25666 , n25671 );
and ( n25673 , n25662 , n25671 );
or ( n25674 , n25667 , n25672 , n25673 );
and ( n25675 , n22425 , n20114 );
and ( n25676 , n22198 , n20112 );
nor ( n25677 , n25675 , n25676 );
xnor ( n25678 , n25677 , n19997 );
and ( n25679 , n24527 , n19518 );
and ( n25680 , n24521 , n19516 );
nor ( n25681 , n25679 , n25680 );
xnor ( n25682 , n25681 , n19489 );
and ( n25683 , n25678 , n25682 );
and ( n25684 , n24940 , n19459 );
and ( n25685 , n24621 , n19457 );
nor ( n25686 , n25684 , n25685 );
xnor ( n25687 , n25686 , n19416 );
and ( n25688 , n25682 , n25687 );
and ( n25689 , n25678 , n25687 );
or ( n25690 , n25683 , n25688 , n25689 );
and ( n25691 , n25674 , n25690 );
xor ( n25692 , n25500 , n25504 );
xor ( n25693 , n25692 , n25509 );
and ( n25694 , n25690 , n25693 );
and ( n25695 , n25674 , n25693 );
or ( n25696 , n25691 , n25694 , n25695 );
xor ( n25697 , n25350 , n25354 );
xor ( n25698 , n25697 , n25359 );
and ( n25699 , n25696 , n25698 );
xor ( n25700 , n25386 , n25390 );
xor ( n25701 , n25700 , n25395 );
and ( n25702 , n25698 , n25701 );
and ( n25703 , n25696 , n25701 );
or ( n25704 , n25699 , n25702 , n25703 );
and ( n25705 , n25657 , n25704 );
and ( n25706 , n25647 , n25704 );
or ( n25707 , n25658 , n25705 , n25706 );
xor ( n25708 , n25379 , n25406 );
xor ( n25709 , n25708 , n25409 );
and ( n25710 , n25707 , n25709 );
xor ( n25711 , n25310 , n25312 );
xor ( n25712 , n25711 , n25315 );
and ( n25713 , n25709 , n25712 );
and ( n25714 , n25707 , n25712 );
or ( n25715 , n25710 , n25713 , n25714 );
and ( n25716 , n25595 , n25715 );
xor ( n25717 , n25412 , n25414 );
xor ( n25718 , n25717 , n25417 );
and ( n25719 , n25715 , n25718 );
and ( n25720 , n25595 , n25718 );
or ( n25721 , n25716 , n25719 , n25720 );
and ( n25722 , n25494 , n25721 );
xor ( n25723 , n25264 , n25324 );
xor ( n25724 , n25723 , n25327 );
and ( n25725 , n25721 , n25724 );
and ( n25726 , n25494 , n25724 );
or ( n25727 , n25722 , n25725 , n25726 );
xor ( n25728 , n25198 , n25200 );
xor ( n25729 , n25728 , n25203 );
and ( n25730 , n25727 , n25729 );
xor ( n25731 , n25330 , n25428 );
xor ( n25732 , n25731 , n25431 );
and ( n25733 , n25729 , n25732 );
and ( n25734 , n25727 , n25732 );
or ( n25735 , n25730 , n25733 , n25734 );
and ( n25736 , n25446 , n25735 );
xor ( n25737 , n25446 , n25735 );
xor ( n25738 , n25727 , n25729 );
xor ( n25739 , n25738 , n25732 );
and ( n25740 , n19469 , n24902 );
and ( n25741 , n19434 , n24900 );
nor ( n25742 , n25740 , n25741 );
xnor ( n25743 , n25742 , n24397 );
and ( n25744 , n19721 , n23641 );
and ( n25745 , n19637 , n23639 );
nor ( n25746 , n25744 , n25745 );
xnor ( n25747 , n25746 , n23213 );
and ( n25748 , n25743 , n25747 );
and ( n25749 , n19825 , n23230 );
and ( n25750 , n19811 , n23228 );
nor ( n25751 , n25749 , n25750 );
xnor ( n25752 , n25751 , n22842 );
and ( n25753 , n25747 , n25752 );
and ( n25754 , n25743 , n25752 );
or ( n25755 , n25748 , n25753 , n25754 );
and ( n25756 , n22235 , n20276 );
and ( n25757 , n21955 , n20274 );
nor ( n25758 , n25756 , n25757 );
xnor ( n25759 , n25758 , n20175 );
and ( n25760 , n25554 , n19424 );
and ( n25761 , n25284 , n19422 );
nor ( n25762 , n25760 , n25761 );
xnor ( n25763 , n25762 , n19431 );
and ( n25764 , n25759 , n25763 );
buf ( n25765 , n19332 );
and ( n25766 , n25765 , n19419 );
and ( n25767 , n25763 , n25766 );
and ( n25768 , n25759 , n25766 );
or ( n25769 , n25764 , n25767 , n25768 );
xor ( n25770 , n25516 , n25520 );
xor ( n25771 , n25770 , n25525 );
and ( n25772 , n25769 , n25771 );
xor ( n25773 , n25450 , n25454 );
xor ( n25774 , n25773 , n25459 );
and ( n25775 , n25771 , n25774 );
and ( n25776 , n25769 , n25774 );
or ( n25777 , n25772 , n25775 , n25776 );
and ( n25778 , n25755 , n25777 );
xor ( n25779 , n25512 , n25528 );
xor ( n25780 , n25779 , n25533 );
and ( n25781 , n25777 , n25780 );
and ( n25782 , n25755 , n25780 );
or ( n25783 , n25778 , n25781 , n25782 );
xor ( n25784 , n25398 , n25400 );
xor ( n25785 , n25784 , n25403 );
and ( n25786 , n25783 , n25785 );
xor ( n25787 , n25536 , n25538 );
xor ( n25788 , n25787 , n25541 );
and ( n25789 , n25785 , n25788 );
and ( n25790 , n25783 , n25788 );
or ( n25791 , n25786 , n25789 , n25790 );
xor ( n25792 , n25346 , n25362 );
xor ( n25793 , n25792 , n25376 );
xor ( n25794 , n25470 , n25472 );
xor ( n25795 , n25794 , n25475 );
and ( n25796 , n25793 , n25795 );
xor ( n25797 , n25581 , n25583 );
xor ( n25798 , n25797 , n25586 );
and ( n25799 , n25795 , n25798 );
and ( n25800 , n25793 , n25798 );
or ( n25801 , n25796 , n25799 , n25800 );
and ( n25802 , n25791 , n25801 );
xor ( n25803 , n25478 , n25480 );
xor ( n25804 , n25803 , n25483 );
and ( n25805 , n25801 , n25804 );
and ( n25806 , n25791 , n25804 );
or ( n25807 , n25802 , n25805 , n25806 );
and ( n25808 , n20618 , n21741 );
and ( n25809 , n20452 , n21739 );
nor ( n25810 , n25808 , n25809 );
xnor ( n25811 , n25810 , n21605 );
and ( n25812 , n20803 , n21468 );
and ( n25813 , n20666 , n21466 );
nor ( n25814 , n25812 , n25813 );
xnor ( n25815 , n25814 , n21331 );
and ( n25816 , n25811 , n25815 );
and ( n25817 , n21072 , n21155 );
and ( n25818 , n20867 , n21153 );
nor ( n25819 , n25817 , n25818 );
xnor ( n25820 , n25819 , n20994 );
and ( n25821 , n25815 , n25820 );
and ( n25822 , n25811 , n25820 );
or ( n25823 , n25816 , n25821 , n25822 );
and ( n25824 , n20182 , n22381 );
and ( n25825 , n20080 , n22379 );
nor ( n25826 , n25824 , n25825 );
xnor ( n25827 , n25826 , n22228 );
and ( n25828 , n20360 , n22048 );
and ( n25829 , n20268 , n22046 );
nor ( n25830 , n25828 , n25829 );
xnor ( n25831 , n25830 , n21853 );
and ( n25832 , n25827 , n25831 );
and ( n25833 , n21876 , n20460 );
and ( n25834 , n21704 , n20458 );
nor ( n25835 , n25833 , n25834 );
xnor ( n25836 , n25835 , n20337 );
and ( n25837 , n25831 , n25836 );
and ( n25838 , n25827 , n25836 );
or ( n25839 , n25832 , n25837 , n25838 );
and ( n25840 , n25823 , n25839 );
and ( n25841 , n21302 , n20955 );
and ( n25842 , n21218 , n20953 );
nor ( n25843 , n25841 , n25842 );
xnor ( n25844 , n25843 , n20780 );
and ( n25845 , n21612 , n20674 );
and ( n25846 , n21451 , n20672 );
nor ( n25847 , n25845 , n25846 );
xnor ( n25848 , n25847 , n20542 );
and ( n25849 , n25844 , n25848 );
not ( n25850 , n25562 );
and ( n25851 , n25848 , n25850 );
and ( n25852 , n25844 , n25850 );
or ( n25853 , n25849 , n25851 , n25852 );
and ( n25854 , n25839 , n25853 );
and ( n25855 , n25823 , n25853 );
or ( n25856 , n25840 , n25854 , n25855 );
xor ( n25857 , n25615 , n25619 );
xor ( n25858 , n25857 , n25624 );
xor ( n25859 , n25548 , n25552 );
xor ( n25860 , n25859 , n25555 );
and ( n25861 , n25858 , n25860 );
xor ( n25862 , n25563 , n25567 );
xor ( n25863 , n25862 , n25572 );
and ( n25864 , n25860 , n25863 );
and ( n25865 , n25858 , n25863 );
or ( n25866 , n25861 , n25864 , n25865 );
and ( n25867 , n25856 , n25866 );
xor ( n25868 , n25462 , n25464 );
xor ( n25869 , n25868 , n25467 );
and ( n25870 , n25866 , n25869 );
and ( n25871 , n25856 , n25869 );
or ( n25872 , n25867 , n25870 , n25871 );
and ( n25873 , n19434 , n25383 );
and ( n25874 , n19418 , n25381 );
nor ( n25875 , n25873 , n25874 );
xnor ( n25876 , n25875 , n24885 );
and ( n25877 , n19588 , n24376 );
and ( n25878 , n19510 , n24374 );
nor ( n25879 , n25877 , n25878 );
xnor ( n25880 , n25879 , n23927 );
and ( n25881 , n25876 , n25880 );
and ( n25882 , n20004 , n22859 );
and ( n25883 , n19946 , n22857 );
nor ( n25884 , n25882 , n25883 );
xnor ( n25885 , n25884 , n22418 );
and ( n25886 , n25880 , n25885 );
and ( n25887 , n25876 , n25885 );
or ( n25888 , n25881 , n25886 , n25887 );
buf ( n25889 , n19398 );
buf ( n25890 , n19399 );
and ( n25891 , n25889 , n25890 );
not ( n25892 , n25891 );
and ( n25893 , n25496 , n25892 );
not ( n25894 , n25893 );
and ( n25895 , n22198 , n20276 );
and ( n25896 , n22235 , n20274 );
nor ( n25897 , n25895 , n25896 );
xnor ( n25898 , n25897 , n20175 );
and ( n25899 , n25894 , n25898 );
and ( n25900 , n22756 , n20114 );
and ( n25901 , n22425 , n20112 );
nor ( n25902 , n25900 , n25901 );
xnor ( n25903 , n25902 , n19997 );
and ( n25904 , n25898 , n25903 );
and ( n25905 , n25894 , n25903 );
or ( n25906 , n25899 , n25904 , n25905 );
and ( n25907 , n19811 , n23641 );
and ( n25908 , n19721 , n23639 );
nor ( n25909 , n25907 , n25908 );
xnor ( n25910 , n25909 , n23213 );
and ( n25911 , n25906 , n25910 );
and ( n25912 , n19881 , n23230 );
and ( n25913 , n19825 , n23228 );
nor ( n25914 , n25912 , n25913 );
xnor ( n25915 , n25914 , n22842 );
and ( n25916 , n25910 , n25915 );
and ( n25917 , n25906 , n25915 );
or ( n25918 , n25911 , n25916 , n25917 );
and ( n25919 , n25888 , n25918 );
xor ( n25920 , n25599 , n25603 );
xor ( n25921 , n25920 , n25608 );
and ( n25922 , n25918 , n25921 );
and ( n25923 , n25888 , n25921 );
or ( n25924 , n25919 , n25922 , n25923 );
xor ( n25925 , n25611 , n25627 );
xor ( n25926 , n25925 , n25644 );
and ( n25927 , n25924 , n25926 );
xor ( n25928 , n25558 , n25575 );
xor ( n25929 , n25928 , n25578 );
and ( n25930 , n25926 , n25929 );
and ( n25931 , n25924 , n25929 );
or ( n25932 , n25927 , n25930 , n25931 );
and ( n25933 , n25872 , n25932 );
xor ( n25934 , n25647 , n25657 );
xor ( n25935 , n25934 , n25704 );
and ( n25936 , n25932 , n25935 );
and ( n25937 , n25872 , n25935 );
or ( n25938 , n25933 , n25936 , n25937 );
xor ( n25939 , n25544 , n25589 );
xor ( n25940 , n25939 , n25592 );
and ( n25941 , n25938 , n25940 );
xor ( n25942 , n25707 , n25709 );
xor ( n25943 , n25942 , n25712 );
and ( n25944 , n25940 , n25943 );
and ( n25945 , n25938 , n25943 );
or ( n25946 , n25941 , n25944 , n25945 );
and ( n25947 , n25807 , n25946 );
xor ( n25948 , n25486 , n25488 );
xor ( n25949 , n25948 , n25491 );
and ( n25950 , n25946 , n25949 );
and ( n25951 , n25807 , n25949 );
or ( n25952 , n25947 , n25950 , n25951 );
xor ( n25953 , n25420 , n25422 );
xor ( n25954 , n25953 , n25425 );
and ( n25955 , n25952 , n25954 );
xor ( n25956 , n25494 , n25721 );
xor ( n25957 , n25956 , n25724 );
and ( n25958 , n25954 , n25957 );
and ( n25959 , n25952 , n25957 );
or ( n25960 , n25955 , n25958 , n25959 );
and ( n25961 , n25739 , n25960 );
xor ( n25962 , n25739 , n25960 );
xor ( n25963 , n25952 , n25954 );
xor ( n25964 , n25963 , n25957 );
and ( n25965 , n21955 , n20460 );
and ( n25966 , n21876 , n20458 );
nor ( n25967 , n25965 , n25966 );
xnor ( n25968 , n25967 , n20337 );
and ( n25969 , n25765 , n19424 );
and ( n25970 , n25554 , n19422 );
nor ( n25971 , n25969 , n25970 );
xnor ( n25972 , n25971 , n19431 );
and ( n25973 , n25968 , n25972 );
buf ( n25974 , n19333 );
and ( n25975 , n25974 , n19419 );
and ( n25976 , n25972 , n25975 );
and ( n25977 , n25968 , n25975 );
or ( n25978 , n25973 , n25976 , n25977 );
and ( n25979 , n20452 , n22048 );
and ( n25980 , n20360 , n22046 );
nor ( n25981 , n25979 , n25980 );
xnor ( n25982 , n25981 , n21853 );
and ( n25983 , n20666 , n21741 );
and ( n25984 , n20618 , n21739 );
nor ( n25985 , n25983 , n25984 );
xnor ( n25986 , n25985 , n21605 );
and ( n25987 , n25982 , n25986 );
and ( n25988 , n20867 , n21468 );
and ( n25989 , n20803 , n21466 );
nor ( n25990 , n25988 , n25989 );
xnor ( n25991 , n25990 , n21331 );
and ( n25992 , n25986 , n25991 );
and ( n25993 , n25982 , n25991 );
or ( n25994 , n25987 , n25992 , n25993 );
and ( n25995 , n25978 , n25994 );
and ( n25996 , n22916 , n20114 );
and ( n25997 , n22756 , n20112 );
nor ( n25998 , n25996 , n25997 );
xnor ( n25999 , n25998 , n19997 );
buf ( n26000 , n25999 );
and ( n26001 , n21218 , n21155 );
and ( n26002 , n21072 , n21153 );
nor ( n26003 , n26001 , n26002 );
xnor ( n26004 , n26003 , n20994 );
and ( n26005 , n26000 , n26004 );
and ( n26006 , n21451 , n20955 );
and ( n26007 , n21302 , n20953 );
nor ( n26008 , n26006 , n26007 );
xnor ( n26009 , n26008 , n20780 );
and ( n26010 , n26004 , n26009 );
and ( n26011 , n26000 , n26009 );
or ( n26012 , n26005 , n26010 , n26011 );
and ( n26013 , n25994 , n26012 );
and ( n26014 , n25978 , n26012 );
or ( n26015 , n25995 , n26013 , n26014 );
xor ( n26016 , n25743 , n25747 );
xor ( n26017 , n26016 , n25752 );
and ( n26018 , n26015 , n26017 );
xor ( n26019 , n25632 , n25636 );
xor ( n26020 , n26019 , n25641 );
and ( n26021 , n26017 , n26020 );
and ( n26022 , n26015 , n26020 );
or ( n26023 , n26018 , n26021 , n26022 );
xor ( n26024 , n24882 , n25495 );
xor ( n26025 , n25495 , n25496 );
not ( n26026 , n26025 );
and ( n26027 , n26024 , n26026 );
and ( n26028 , n19426 , n26027 );
not ( n26029 , n26028 );
xnor ( n26030 , n26029 , n25499 );
and ( n26031 , n19496 , n24902 );
and ( n26032 , n19469 , n24900 );
nor ( n26033 , n26031 , n26032 );
xnor ( n26034 , n26033 , n24397 );
and ( n26035 , n26030 , n26034 );
and ( n26036 , n19637 , n23944 );
and ( n26037 , n19605 , n23942 );
nor ( n26038 , n26036 , n26037 );
xnor ( n26039 , n26038 , n23550 );
and ( n26040 , n26034 , n26039 );
and ( n26041 , n26030 , n26039 );
or ( n26042 , n26035 , n26040 , n26041 );
and ( n26043 , n23141 , n19894 );
and ( n26044 , n22916 , n19892 );
nor ( n26045 , n26043 , n26044 );
xnor ( n26046 , n26045 , n19858 );
and ( n26047 , n23381 , n19805 );
and ( n26048 , n23271 , n19803 );
nor ( n26049 , n26047 , n26048 );
xnor ( n26050 , n26049 , n19750 );
and ( n26051 , n26046 , n26050 );
and ( n26052 , n23968 , n19688 );
and ( n26053 , n23573 , n19686 );
nor ( n26054 , n26052 , n26053 );
xnor ( n26055 , n26054 , n19655 );
and ( n26056 , n26050 , n26055 );
and ( n26057 , n26046 , n26055 );
or ( n26058 , n26051 , n26056 , n26057 );
and ( n26059 , n24521 , n19596 );
and ( n26060 , n24131 , n19594 );
nor ( n26061 , n26059 , n26060 );
xnor ( n26062 , n26061 , n19545 );
and ( n26063 , n24621 , n19518 );
and ( n26064 , n24527 , n19516 );
nor ( n26065 , n26063 , n26064 );
xnor ( n26066 , n26065 , n19489 );
and ( n26067 , n26062 , n26066 );
and ( n26068 , n25284 , n19459 );
and ( n26069 , n24940 , n19457 );
nor ( n26070 , n26068 , n26069 );
xnor ( n26071 , n26070 , n19416 );
and ( n26072 , n26066 , n26071 );
and ( n26073 , n26062 , n26071 );
or ( n26074 , n26067 , n26072 , n26073 );
and ( n26075 , n26058 , n26074 );
xor ( n26076 , n25759 , n25763 );
xor ( n26077 , n26076 , n25766 );
and ( n26078 , n26074 , n26077 );
and ( n26079 , n26058 , n26077 );
or ( n26080 , n26075 , n26078 , n26079 );
and ( n26081 , n26042 , n26080 );
xor ( n26082 , n25674 , n25690 );
xor ( n26083 , n26082 , n25693 );
and ( n26084 , n26080 , n26083 );
and ( n26085 , n26042 , n26083 );
or ( n26086 , n26081 , n26084 , n26085 );
and ( n26087 , n26023 , n26086 );
xor ( n26088 , n25649 , n25651 );
xor ( n26089 , n26088 , n25654 );
and ( n26090 , n26086 , n26089 );
and ( n26091 , n26023 , n26089 );
or ( n26092 , n26087 , n26090 , n26091 );
and ( n26093 , n20080 , n22859 );
and ( n26094 , n20004 , n22857 );
nor ( n26095 , n26093 , n26094 );
xnor ( n26096 , n26095 , n22418 );
and ( n26097 , n20268 , n22381 );
and ( n26098 , n20182 , n22379 );
nor ( n26099 , n26097 , n26098 );
xnor ( n26100 , n26099 , n22228 );
and ( n26101 , n26096 , n26100 );
and ( n26102 , n21704 , n20674 );
and ( n26103 , n21612 , n20672 );
nor ( n26104 , n26102 , n26103 );
xnor ( n26105 , n26104 , n20542 );
and ( n26106 , n26100 , n26105 );
and ( n26107 , n26096 , n26105 );
or ( n26108 , n26101 , n26106 , n26107 );
xor ( n26109 , n25662 , n25666 );
xor ( n26110 , n26109 , n25671 );
and ( n26111 , n26108 , n26110 );
xor ( n26112 , n25678 , n25682 );
xor ( n26113 , n26112 , n25687 );
and ( n26114 , n26110 , n26113 );
and ( n26115 , n26108 , n26113 );
or ( n26116 , n26111 , n26114 , n26115 );
and ( n26117 , n19469 , n25383 );
and ( n26118 , n19434 , n25381 );
nor ( n26119 , n26117 , n26118 );
xnor ( n26120 , n26119 , n24885 );
and ( n26121 , n19605 , n24376 );
and ( n26122 , n19588 , n24374 );
nor ( n26123 , n26121 , n26122 );
xnor ( n26124 , n26123 , n23927 );
and ( n26125 , n26120 , n26124 );
and ( n26126 , n19721 , n23944 );
and ( n26127 , n19637 , n23942 );
nor ( n26128 , n26126 , n26127 );
xnor ( n26129 , n26128 , n23550 );
and ( n26130 , n26124 , n26129 );
and ( n26131 , n26120 , n26129 );
or ( n26132 , n26125 , n26130 , n26131 );
and ( n26133 , n23271 , n19894 );
and ( n26134 , n23141 , n19892 );
nor ( n26135 , n26133 , n26134 );
xnor ( n26136 , n26135 , n19858 );
and ( n26137 , n23573 , n19805 );
and ( n26138 , n23381 , n19803 );
nor ( n26139 , n26137 , n26138 );
xnor ( n26140 , n26139 , n19750 );
and ( n26141 , n26136 , n26140 );
and ( n26142 , n24131 , n19688 );
and ( n26143 , n23968 , n19686 );
nor ( n26144 , n26142 , n26143 );
xnor ( n26145 , n26144 , n19655 );
and ( n26146 , n26140 , n26145 );
and ( n26147 , n26136 , n26145 );
or ( n26148 , n26141 , n26146 , n26147 );
and ( n26149 , n22425 , n20276 );
and ( n26150 , n22198 , n20274 );
nor ( n26151 , n26149 , n26150 );
xnor ( n26152 , n26151 , n20175 );
and ( n26153 , n24527 , n19596 );
and ( n26154 , n24521 , n19594 );
nor ( n26155 , n26153 , n26154 );
xnor ( n26156 , n26155 , n19545 );
and ( n26157 , n26152 , n26156 );
and ( n26158 , n25554 , n19459 );
and ( n26159 , n25284 , n19457 );
nor ( n26160 , n26158 , n26159 );
xnor ( n26161 , n26160 , n19416 );
and ( n26162 , n26156 , n26161 );
and ( n26163 , n26152 , n26161 );
or ( n26164 , n26157 , n26162 , n26163 );
and ( n26165 , n26148 , n26164 );
and ( n26166 , n19825 , n23641 );
and ( n26167 , n19811 , n23639 );
nor ( n26168 , n26166 , n26167 );
xnor ( n26169 , n26168 , n23213 );
and ( n26170 , n26164 , n26169 );
and ( n26171 , n26148 , n26169 );
or ( n26172 , n26165 , n26170 , n26171 );
and ( n26173 , n26132 , n26172 );
xor ( n26174 , n25811 , n25815 );
xor ( n26175 , n26174 , n25820 );
and ( n26176 , n26172 , n26175 );
and ( n26177 , n26132 , n26175 );
or ( n26178 , n26173 , n26176 , n26177 );
and ( n26179 , n26116 , n26178 );
xor ( n26180 , n25769 , n25771 );
xor ( n26181 , n26180 , n25774 );
and ( n26182 , n26178 , n26181 );
and ( n26183 , n26116 , n26181 );
or ( n26184 , n26179 , n26182 , n26183 );
xor ( n26185 , n25755 , n25777 );
xor ( n26186 , n26185 , n25780 );
and ( n26187 , n26184 , n26186 );
xor ( n26188 , n25696 , n25698 );
xor ( n26189 , n26188 , n25701 );
and ( n26190 , n26186 , n26189 );
and ( n26191 , n26184 , n26189 );
or ( n26192 , n26187 , n26190 , n26191 );
and ( n26193 , n26092 , n26192 );
xor ( n26194 , n25783 , n25785 );
xor ( n26195 , n26194 , n25788 );
and ( n26196 , n26192 , n26195 );
and ( n26197 , n26092 , n26195 );
or ( n26198 , n26193 , n26196 , n26197 );
xor ( n26199 , n25791 , n25801 );
xor ( n26200 , n26199 , n25804 );
and ( n26201 , n26198 , n26200 );
xor ( n26202 , n25938 , n25940 );
xor ( n26203 , n26202 , n25943 );
and ( n26204 , n26200 , n26203 );
and ( n26205 , n26198 , n26203 );
or ( n26206 , n26201 , n26204 , n26205 );
xor ( n26207 , n25595 , n25715 );
xor ( n26208 , n26207 , n25718 );
and ( n26209 , n26206 , n26208 );
xor ( n26210 , n25807 , n25946 );
xor ( n26211 , n26210 , n25949 );
and ( n26212 , n26208 , n26211 );
and ( n26213 , n26206 , n26211 );
or ( n26214 , n26209 , n26212 , n26213 );
and ( n26215 , n25964 , n26214 );
xor ( n26216 , n25964 , n26214 );
xor ( n26217 , n26206 , n26208 );
xor ( n26218 , n26217 , n26211 );
and ( n26219 , n19418 , n26027 );
and ( n26220 , n19426 , n26025 );
nor ( n26221 , n26219 , n26220 );
xnor ( n26222 , n26221 , n25499 );
and ( n26223 , n19510 , n24902 );
and ( n26224 , n19496 , n24900 );
nor ( n26225 , n26223 , n26224 );
xnor ( n26226 , n26225 , n24397 );
and ( n26227 , n26222 , n26226 );
and ( n26228 , n19946 , n23230 );
and ( n26229 , n19881 , n23228 );
nor ( n26230 , n26228 , n26229 );
xnor ( n26231 , n26230 , n22842 );
and ( n26232 , n26226 , n26231 );
and ( n26233 , n26222 , n26231 );
or ( n26234 , n26227 , n26232 , n26233 );
xor ( n26235 , n25827 , n25831 );
xor ( n26236 , n26235 , n25836 );
and ( n26237 , n26234 , n26236 );
xor ( n26238 , n25844 , n25848 );
xor ( n26239 , n26238 , n25850 );
and ( n26240 , n26236 , n26239 );
and ( n26241 , n26234 , n26239 );
or ( n26242 , n26237 , n26240 , n26241 );
xor ( n26243 , n25823 , n25839 );
xor ( n26244 , n26243 , n25853 );
and ( n26245 , n26242 , n26244 );
xor ( n26246 , n25858 , n25860 );
xor ( n26247 , n26246 , n25863 );
and ( n26248 , n26244 , n26247 );
and ( n26249 , n26242 , n26247 );
or ( n26250 , n26245 , n26248 , n26249 );
xor ( n26251 , n25856 , n25866 );
xor ( n26252 , n26251 , n25869 );
and ( n26253 , n26250 , n26252 );
xor ( n26254 , n25924 , n25926 );
xor ( n26255 , n26254 , n25929 );
and ( n26256 , n26252 , n26255 );
and ( n26257 , n26250 , n26255 );
or ( n26258 , n26253 , n26256 , n26257 );
xor ( n26259 , n25872 , n25932 );
xor ( n26260 , n26259 , n25935 );
and ( n26261 , n26258 , n26260 );
xor ( n26262 , n25793 , n25795 );
xor ( n26263 , n26262 , n25798 );
and ( n26264 , n26260 , n26263 );
and ( n26265 , n26258 , n26263 );
or ( n26266 , n26261 , n26264 , n26265 );
and ( n26267 , n20182 , n22859 );
and ( n26268 , n20080 , n22857 );
nor ( n26269 , n26267 , n26268 );
xnor ( n26270 , n26269 , n22418 );
and ( n26271 , n21876 , n20674 );
and ( n26272 , n21704 , n20672 );
nor ( n26273 , n26271 , n26272 );
xnor ( n26274 , n26273 , n20542 );
and ( n26275 , n26270 , n26274 );
and ( n26276 , n22235 , n20460 );
and ( n26277 , n21955 , n20458 );
nor ( n26278 , n26276 , n26277 );
xnor ( n26279 , n26278 , n20337 );
and ( n26280 , n26274 , n26279 );
and ( n26281 , n26270 , n26279 );
or ( n26282 , n26275 , n26280 , n26281 );
and ( n26283 , n20360 , n22381 );
and ( n26284 , n20268 , n22379 );
nor ( n26285 , n26283 , n26284 );
xnor ( n26286 , n26285 , n22228 );
and ( n26287 , n20618 , n22048 );
and ( n26288 , n20452 , n22046 );
nor ( n26289 , n26287 , n26288 );
xnor ( n26290 , n26289 , n21853 );
and ( n26291 , n26286 , n26290 );
not ( n26292 , n25999 );
and ( n26293 , n26290 , n26292 );
and ( n26294 , n26286 , n26292 );
or ( n26295 , n26291 , n26293 , n26294 );
and ( n26296 , n26282 , n26295 );
xor ( n26297 , n26046 , n26050 );
xor ( n26298 , n26297 , n26055 );
and ( n26299 , n26295 , n26298 );
and ( n26300 , n26282 , n26298 );
or ( n26301 , n26296 , n26299 , n26300 );
xor ( n26302 , n26030 , n26034 );
xor ( n26303 , n26302 , n26039 );
and ( n26304 , n26301 , n26303 );
xor ( n26305 , n25906 , n25910 );
xor ( n26306 , n26305 , n25915 );
and ( n26307 , n26303 , n26306 );
and ( n26308 , n26301 , n26306 );
or ( n26309 , n26304 , n26307 , n26308 );
and ( n26310 , n24940 , n19518 );
and ( n26311 , n24621 , n19516 );
nor ( n26312 , n26310 , n26311 );
xnor ( n26313 , n26312 , n19489 );
and ( n26314 , n25974 , n19424 );
and ( n26315 , n25765 , n19422 );
nor ( n26316 , n26314 , n26315 );
xnor ( n26317 , n26316 , n19431 );
and ( n26318 , n26313 , n26317 );
buf ( n26319 , n19334 );
and ( n26320 , n26319 , n19419 );
and ( n26321 , n26317 , n26320 );
and ( n26322 , n26313 , n26320 );
or ( n26323 , n26318 , n26321 , n26322 );
xor ( n26324 , n25894 , n25898 );
xor ( n26325 , n26324 , n25903 );
and ( n26326 , n26323 , n26325 );
xor ( n26327 , n26062 , n26066 );
xor ( n26328 , n26327 , n26071 );
and ( n26329 , n26325 , n26328 );
and ( n26330 , n26323 , n26328 );
or ( n26331 , n26326 , n26329 , n26330 );
xor ( n26332 , n25876 , n25880 );
xor ( n26333 , n26332 , n25885 );
and ( n26334 , n26331 , n26333 );
xor ( n26335 , n26058 , n26074 );
xor ( n26336 , n26335 , n26077 );
and ( n26337 , n26333 , n26336 );
and ( n26338 , n26331 , n26336 );
or ( n26339 , n26334 , n26337 , n26338 );
and ( n26340 , n26309 , n26339 );
xor ( n26341 , n25888 , n25918 );
xor ( n26342 , n26341 , n25921 );
and ( n26343 , n26339 , n26342 );
and ( n26344 , n26309 , n26342 );
or ( n26345 , n26340 , n26343 , n26344 );
xor ( n26346 , n25496 , n25889 );
xor ( n26347 , n25889 , n25890 );
not ( n26348 , n26347 );
and ( n26349 , n26346 , n26348 );
and ( n26350 , n19426 , n26349 );
not ( n26351 , n26350 );
xnor ( n26352 , n26351 , n25893 );
and ( n26353 , n19496 , n25383 );
and ( n26354 , n19469 , n25381 );
nor ( n26355 , n26353 , n26354 );
xnor ( n26356 , n26355 , n24885 );
and ( n26357 , n26352 , n26356 );
and ( n26358 , n19811 , n23944 );
and ( n26359 , n19721 , n23942 );
nor ( n26360 , n26358 , n26359 );
xnor ( n26361 , n26360 , n23550 );
and ( n26362 , n26356 , n26361 );
and ( n26363 , n26352 , n26361 );
or ( n26364 , n26357 , n26362 , n26363 );
buf ( n26365 , n19400 );
buf ( n26366 , n19401 );
and ( n26367 , n26365 , n26366 );
not ( n26368 , n26367 );
and ( n26369 , n25890 , n26368 );
not ( n26370 , n26369 );
and ( n26371 , n22198 , n20460 );
and ( n26372 , n22235 , n20458 );
nor ( n26373 , n26371 , n26372 );
xnor ( n26374 , n26373 , n20337 );
and ( n26375 , n26370 , n26374 );
and ( n26376 , n22756 , n20276 );
and ( n26377 , n22425 , n20274 );
nor ( n26378 , n26376 , n26377 );
xnor ( n26379 , n26378 , n20175 );
and ( n26380 , n26374 , n26379 );
and ( n26381 , n26370 , n26379 );
or ( n26382 , n26375 , n26380 , n26381 );
and ( n26383 , n23141 , n20114 );
and ( n26384 , n22916 , n20112 );
nor ( n26385 , n26383 , n26384 );
xnor ( n26386 , n26385 , n19997 );
and ( n26387 , n23381 , n19894 );
and ( n26388 , n23271 , n19892 );
nor ( n26389 , n26387 , n26388 );
xnor ( n26390 , n26389 , n19858 );
and ( n26391 , n26386 , n26390 );
and ( n26392 , n23968 , n19805 );
and ( n26393 , n23573 , n19803 );
nor ( n26394 , n26392 , n26393 );
xnor ( n26395 , n26394 , n19750 );
and ( n26396 , n26390 , n26395 );
and ( n26397 , n26386 , n26395 );
or ( n26398 , n26391 , n26396 , n26397 );
and ( n26399 , n26382 , n26398 );
and ( n26400 , n19881 , n23641 );
and ( n26401 , n19825 , n23639 );
nor ( n26402 , n26400 , n26401 );
xnor ( n26403 , n26402 , n23213 );
and ( n26404 , n26398 , n26403 );
and ( n26405 , n26382 , n26403 );
or ( n26406 , n26399 , n26404 , n26405 );
and ( n26407 , n26364 , n26406 );
xor ( n26408 , n25982 , n25986 );
xor ( n26409 , n26408 , n25991 );
and ( n26410 , n26406 , n26409 );
and ( n26411 , n26364 , n26409 );
or ( n26412 , n26407 , n26410 , n26411 );
and ( n26413 , n25765 , n19459 );
and ( n26414 , n25554 , n19457 );
nor ( n26415 , n26413 , n26414 );
xnor ( n26416 , n26415 , n19416 );
and ( n26417 , n26319 , n19424 );
and ( n26418 , n25974 , n19422 );
nor ( n26419 , n26417 , n26418 );
xnor ( n26420 , n26419 , n19431 );
and ( n26421 , n26416 , n26420 );
buf ( n26422 , n19335 );
and ( n26423 , n26422 , n19419 );
and ( n26424 , n26420 , n26423 );
and ( n26425 , n26416 , n26423 );
or ( n26426 , n26421 , n26424 , n26425 );
and ( n26427 , n20004 , n23230 );
and ( n26428 , n19946 , n23228 );
nor ( n26429 , n26427 , n26428 );
xnor ( n26430 , n26429 , n22842 );
and ( n26431 , n26426 , n26430 );
and ( n26432 , n21612 , n20955 );
and ( n26433 , n21451 , n20953 );
nor ( n26434 , n26432 , n26433 );
xnor ( n26435 , n26434 , n20780 );
and ( n26436 , n26430 , n26435 );
and ( n26437 , n26426 , n26435 );
or ( n26438 , n26431 , n26436 , n26437 );
xor ( n26439 , n26096 , n26100 );
xor ( n26440 , n26439 , n26105 );
and ( n26441 , n26438 , n26440 );
xor ( n26442 , n26000 , n26004 );
xor ( n26443 , n26442 , n26009 );
and ( n26444 , n26440 , n26443 );
and ( n26445 , n26438 , n26443 );
or ( n26446 , n26441 , n26444 , n26445 );
and ( n26447 , n26412 , n26446 );
xor ( n26448 , n26108 , n26110 );
xor ( n26449 , n26448 , n26113 );
and ( n26450 , n26446 , n26449 );
and ( n26451 , n26412 , n26449 );
or ( n26452 , n26447 , n26450 , n26451 );
xor ( n26453 , n26015 , n26017 );
xor ( n26454 , n26453 , n26020 );
and ( n26455 , n26452 , n26454 );
xor ( n26456 , n26042 , n26080 );
xor ( n26457 , n26456 , n26083 );
and ( n26458 , n26454 , n26457 );
and ( n26459 , n26452 , n26457 );
or ( n26460 , n26455 , n26458 , n26459 );
and ( n26461 , n26345 , n26460 );
xor ( n26462 , n26023 , n26086 );
xor ( n26463 , n26462 , n26089 );
and ( n26464 , n26460 , n26463 );
and ( n26465 , n26345 , n26463 );
or ( n26466 , n26461 , n26464 , n26465 );
and ( n26467 , n20803 , n21741 );
and ( n26468 , n20666 , n21739 );
nor ( n26469 , n26467 , n26468 );
xnor ( n26470 , n26469 , n21605 );
and ( n26471 , n21072 , n21468 );
and ( n26472 , n20867 , n21466 );
nor ( n26473 , n26471 , n26472 );
xnor ( n26474 , n26473 , n21331 );
and ( n26475 , n26470 , n26474 );
and ( n26476 , n21302 , n21155 );
and ( n26477 , n21218 , n21153 );
nor ( n26478 , n26476 , n26477 );
xnor ( n26479 , n26478 , n20994 );
and ( n26480 , n26474 , n26479 );
and ( n26481 , n26470 , n26479 );
or ( n26482 , n26475 , n26480 , n26481 );
and ( n26483 , n19434 , n26027 );
and ( n26484 , n19418 , n26025 );
nor ( n26485 , n26483 , n26484 );
xnor ( n26486 , n26485 , n25499 );
and ( n26487 , n19588 , n24902 );
and ( n26488 , n19510 , n24900 );
nor ( n26489 , n26487 , n26488 );
xnor ( n26490 , n26489 , n24397 );
and ( n26491 , n26486 , n26490 );
and ( n26492 , n19637 , n24376 );
and ( n26493 , n19605 , n24374 );
nor ( n26494 , n26492 , n26493 );
xnor ( n26495 , n26494 , n23927 );
and ( n26496 , n26490 , n26495 );
and ( n26497 , n26486 , n26495 );
or ( n26498 , n26491 , n26496 , n26497 );
and ( n26499 , n26482 , n26498 );
xor ( n26500 , n25968 , n25972 );
xor ( n26501 , n26500 , n25975 );
and ( n26502 , n26498 , n26501 );
and ( n26503 , n26482 , n26501 );
or ( n26504 , n26499 , n26502 , n26503 );
and ( n26505 , n24521 , n19688 );
and ( n26506 , n24131 , n19686 );
nor ( n26507 , n26505 , n26506 );
xnor ( n26508 , n26507 , n19655 );
and ( n26509 , n24621 , n19596 );
and ( n26510 , n24527 , n19594 );
nor ( n26511 , n26509 , n26510 );
xnor ( n26512 , n26511 , n19545 );
and ( n26513 , n26508 , n26512 );
and ( n26514 , n25284 , n19518 );
and ( n26515 , n24940 , n19516 );
nor ( n26516 , n26514 , n26515 );
xnor ( n26517 , n26516 , n19489 );
and ( n26518 , n26512 , n26517 );
and ( n26519 , n26508 , n26517 );
or ( n26520 , n26513 , n26518 , n26519 );
xor ( n26521 , n26152 , n26156 );
xor ( n26522 , n26521 , n26161 );
and ( n26523 , n26520 , n26522 );
xor ( n26524 , n26313 , n26317 );
xor ( n26525 , n26524 , n26320 );
and ( n26526 , n26522 , n26525 );
and ( n26527 , n26520 , n26525 );
or ( n26528 , n26523 , n26526 , n26527 );
xor ( n26529 , n26222 , n26226 );
xor ( n26530 , n26529 , n26231 );
and ( n26531 , n26528 , n26530 );
xor ( n26532 , n26148 , n26164 );
xor ( n26533 , n26532 , n26169 );
and ( n26534 , n26530 , n26533 );
and ( n26535 , n26528 , n26533 );
or ( n26536 , n26531 , n26534 , n26535 );
and ( n26537 , n26504 , n26536 );
xor ( n26538 , n25978 , n25994 );
xor ( n26539 , n26538 , n26012 );
and ( n26540 , n26536 , n26539 );
and ( n26541 , n26504 , n26539 );
or ( n26542 , n26537 , n26540 , n26541 );
xor ( n26543 , n26116 , n26178 );
xor ( n26544 , n26543 , n26181 );
and ( n26545 , n26542 , n26544 );
xor ( n26546 , n26242 , n26244 );
xor ( n26547 , n26546 , n26247 );
and ( n26548 , n26544 , n26547 );
and ( n26549 , n26542 , n26547 );
or ( n26550 , n26545 , n26548 , n26549 );
xor ( n26551 , n26184 , n26186 );
xor ( n26552 , n26551 , n26189 );
and ( n26553 , n26550 , n26552 );
xor ( n26554 , n26250 , n26252 );
xor ( n26555 , n26554 , n26255 );
and ( n26556 , n26552 , n26555 );
and ( n26557 , n26550 , n26555 );
or ( n26558 , n26553 , n26556 , n26557 );
and ( n26559 , n26466 , n26558 );
xor ( n26560 , n26092 , n26192 );
xor ( n26561 , n26560 , n26195 );
and ( n26562 , n26558 , n26561 );
and ( n26563 , n26466 , n26561 );
or ( n26564 , n26559 , n26562 , n26563 );
and ( n26565 , n26266 , n26564 );
xor ( n26566 , n26198 , n26200 );
xor ( n26567 , n26566 , n26203 );
and ( n26568 , n26564 , n26567 );
and ( n26569 , n26266 , n26567 );
or ( n26570 , n26565 , n26568 , n26569 );
and ( n26571 , n26218 , n26570 );
xor ( n26572 , n26218 , n26570 );
xor ( n26573 , n26266 , n26564 );
xor ( n26574 , n26573 , n26567 );
xor ( n26575 , n26234 , n26236 );
xor ( n26576 , n26575 , n26239 );
xor ( n26577 , n26132 , n26172 );
xor ( n26578 , n26577 , n26175 );
and ( n26579 , n26576 , n26578 );
xor ( n26580 , n26301 , n26303 );
xor ( n26581 , n26580 , n26306 );
and ( n26582 , n26578 , n26581 );
and ( n26583 , n26576 , n26581 );
or ( n26584 , n26579 , n26582 , n26583 );
xor ( n26585 , n26309 , n26339 );
xor ( n26586 , n26585 , n26342 );
and ( n26587 , n26584 , n26586 );
xor ( n26588 , n26452 , n26454 );
xor ( n26589 , n26588 , n26457 );
and ( n26590 , n26586 , n26589 );
and ( n26591 , n26584 , n26589 );
or ( n26592 , n26587 , n26590 , n26591 );
and ( n26593 , n20268 , n22859 );
and ( n26594 , n20182 , n22857 );
nor ( n26595 , n26593 , n26594 );
xnor ( n26596 , n26595 , n22418 );
and ( n26597 , n20452 , n22381 );
and ( n26598 , n20360 , n22379 );
nor ( n26599 , n26597 , n26598 );
xnor ( n26600 , n26599 , n22228 );
and ( n26601 , n26596 , n26600 );
and ( n26602 , n20666 , n22048 );
and ( n26603 , n20618 , n22046 );
nor ( n26604 , n26602 , n26603 );
xnor ( n26605 , n26604 , n21853 );
and ( n26606 , n26600 , n26605 );
and ( n26607 , n26596 , n26605 );
or ( n26608 , n26601 , n26606 , n26607 );
and ( n26609 , n20080 , n23230 );
and ( n26610 , n20004 , n23228 );
nor ( n26611 , n26609 , n26610 );
xnor ( n26612 , n26611 , n22842 );
and ( n26613 , n21704 , n20955 );
and ( n26614 , n21612 , n20953 );
nor ( n26615 , n26613 , n26614 );
xnor ( n26616 , n26615 , n20780 );
and ( n26617 , n26612 , n26616 );
and ( n26618 , n21955 , n20674 );
and ( n26619 , n21876 , n20672 );
nor ( n26620 , n26618 , n26619 );
xnor ( n26621 , n26620 , n20542 );
and ( n26622 , n26616 , n26621 );
and ( n26623 , n26612 , n26621 );
or ( n26624 , n26617 , n26622 , n26623 );
and ( n26625 , n26608 , n26624 );
xor ( n26626 , n26136 , n26140 );
xor ( n26627 , n26626 , n26145 );
and ( n26628 , n26624 , n26627 );
and ( n26629 , n26608 , n26627 );
or ( n26630 , n26625 , n26628 , n26629 );
xor ( n26631 , n26120 , n26124 );
xor ( n26632 , n26631 , n26129 );
and ( n26633 , n26630 , n26632 );
xor ( n26634 , n26323 , n26325 );
xor ( n26635 , n26634 , n26328 );
and ( n26636 , n26632 , n26635 );
and ( n26637 , n26630 , n26635 );
or ( n26638 , n26633 , n26636 , n26637 );
and ( n26639 , n19418 , n26349 );
and ( n26640 , n19426 , n26347 );
nor ( n26641 , n26639 , n26640 );
xnor ( n26642 , n26641 , n25893 );
and ( n26643 , n19510 , n25383 );
and ( n26644 , n19496 , n25381 );
nor ( n26645 , n26643 , n26644 );
xnor ( n26646 , n26645 , n24885 );
and ( n26647 , n26642 , n26646 );
and ( n26648 , n19605 , n24902 );
and ( n26649 , n19588 , n24900 );
nor ( n26650 , n26648 , n26649 );
xnor ( n26651 , n26650 , n24397 );
and ( n26652 , n26646 , n26651 );
and ( n26653 , n26642 , n26651 );
or ( n26654 , n26647 , n26652 , n26653 );
and ( n26655 , n22916 , n20276 );
and ( n26656 , n22756 , n20274 );
nor ( n26657 , n26655 , n26656 );
xnor ( n26658 , n26657 , n20175 );
buf ( n26659 , n26658 );
and ( n26660 , n20867 , n21741 );
and ( n26661 , n20803 , n21739 );
nor ( n26662 , n26660 , n26661 );
xnor ( n26663 , n26662 , n21605 );
and ( n26664 , n26659 , n26663 );
and ( n26665 , n21218 , n21468 );
and ( n26666 , n21072 , n21466 );
nor ( n26667 , n26665 , n26666 );
xnor ( n26668 , n26667 , n21331 );
and ( n26669 , n26663 , n26668 );
and ( n26670 , n26659 , n26668 );
or ( n26671 , n26664 , n26669 , n26670 );
and ( n26672 , n26654 , n26671 );
and ( n26673 , n24940 , n19596 );
and ( n26674 , n24621 , n19594 );
nor ( n26675 , n26673 , n26674 );
xnor ( n26676 , n26675 , n19545 );
and ( n26677 , n25974 , n19459 );
and ( n26678 , n25765 , n19457 );
nor ( n26679 , n26677 , n26678 );
xnor ( n26680 , n26679 , n19416 );
and ( n26681 , n26676 , n26680 );
and ( n26682 , n26422 , n19424 );
and ( n26683 , n26319 , n19422 );
nor ( n26684 , n26682 , n26683 );
xnor ( n26685 , n26684 , n19431 );
and ( n26686 , n26680 , n26685 );
and ( n26687 , n26676 , n26685 );
or ( n26688 , n26681 , n26686 , n26687 );
and ( n26689 , n19946 , n23641 );
and ( n26690 , n19881 , n23639 );
nor ( n26691 , n26689 , n26690 );
xnor ( n26692 , n26691 , n23213 );
and ( n26693 , n26688 , n26692 );
and ( n26694 , n21451 , n21155 );
and ( n26695 , n21302 , n21153 );
nor ( n26696 , n26694 , n26695 );
xnor ( n26697 , n26696 , n20994 );
and ( n26698 , n26692 , n26697 );
and ( n26699 , n26688 , n26697 );
or ( n26700 , n26693 , n26698 , n26699 );
and ( n26701 , n26671 , n26700 );
and ( n26702 , n26654 , n26700 );
or ( n26703 , n26672 , n26701 , n26702 );
and ( n26704 , n19469 , n26027 );
and ( n26705 , n19434 , n26025 );
nor ( n26706 , n26704 , n26705 );
xnor ( n26707 , n26706 , n25499 );
and ( n26708 , n19721 , n24376 );
and ( n26709 , n19637 , n24374 );
nor ( n26710 , n26708 , n26709 );
xnor ( n26711 , n26710 , n23927 );
and ( n26712 , n26707 , n26711 );
and ( n26713 , n19825 , n23944 );
and ( n26714 , n19811 , n23942 );
nor ( n26715 , n26713 , n26714 );
xnor ( n26716 , n26715 , n23550 );
and ( n26717 , n26711 , n26716 );
and ( n26718 , n26707 , n26716 );
or ( n26719 , n26712 , n26717 , n26718 );
xor ( n26720 , n26470 , n26474 );
xor ( n26721 , n26720 , n26479 );
and ( n26722 , n26719 , n26721 );
xor ( n26723 , n26286 , n26290 );
xor ( n26724 , n26723 , n26292 );
and ( n26725 , n26721 , n26724 );
and ( n26726 , n26719 , n26724 );
or ( n26727 , n26722 , n26725 , n26726 );
and ( n26728 , n26703 , n26727 );
xor ( n26729 , n26482 , n26498 );
xor ( n26730 , n26729 , n26501 );
and ( n26731 , n26727 , n26730 );
and ( n26732 , n26703 , n26730 );
or ( n26733 , n26728 , n26731 , n26732 );
and ( n26734 , n26638 , n26733 );
xor ( n26735 , n26331 , n26333 );
xor ( n26736 , n26735 , n26336 );
and ( n26737 , n26733 , n26736 );
and ( n26738 , n26638 , n26736 );
or ( n26739 , n26734 , n26737 , n26738 );
and ( n26740 , n23271 , n20114 );
and ( n26741 , n23141 , n20112 );
nor ( n26742 , n26740 , n26741 );
xnor ( n26743 , n26742 , n19997 );
and ( n26744 , n23573 , n19894 );
and ( n26745 , n23381 , n19892 );
nor ( n26746 , n26744 , n26745 );
xnor ( n26747 , n26746 , n19858 );
and ( n26748 , n26743 , n26747 );
and ( n26749 , n24131 , n19805 );
and ( n26750 , n23968 , n19803 );
nor ( n26751 , n26749 , n26750 );
xnor ( n26752 , n26751 , n19750 );
and ( n26753 , n26747 , n26752 );
and ( n26754 , n26743 , n26752 );
or ( n26755 , n26748 , n26753 , n26754 );
and ( n26756 , n22425 , n20460 );
and ( n26757 , n22198 , n20458 );
nor ( n26758 , n26756 , n26757 );
xnor ( n26759 , n26758 , n20337 );
and ( n26760 , n24527 , n19688 );
and ( n26761 , n24521 , n19686 );
nor ( n26762 , n26760 , n26761 );
xnor ( n26763 , n26762 , n19655 );
and ( n26764 , n26759 , n26763 );
and ( n26765 , n25554 , n19518 );
and ( n26766 , n25284 , n19516 );
nor ( n26767 , n26765 , n26766 );
xnor ( n26768 , n26767 , n19489 );
and ( n26769 , n26763 , n26768 );
and ( n26770 , n26759 , n26768 );
or ( n26771 , n26764 , n26769 , n26770 );
and ( n26772 , n26755 , n26771 );
xor ( n26773 , n26370 , n26374 );
xor ( n26774 , n26773 , n26379 );
and ( n26775 , n26771 , n26774 );
and ( n26776 , n26755 , n26774 );
or ( n26777 , n26772 , n26775 , n26776 );
xor ( n26778 , n26270 , n26274 );
xor ( n26779 , n26778 , n26279 );
and ( n26780 , n26777 , n26779 );
xor ( n26781 , n26382 , n26398 );
xor ( n26782 , n26781 , n26403 );
and ( n26783 , n26779 , n26782 );
and ( n26784 , n26777 , n26782 );
or ( n26785 , n26780 , n26783 , n26784 );
xor ( n26786 , n26386 , n26390 );
xor ( n26787 , n26786 , n26395 );
xor ( n26788 , n26416 , n26420 );
xor ( n26789 , n26788 , n26423 );
and ( n26790 , n26787 , n26789 );
xor ( n26791 , n26508 , n26512 );
xor ( n26792 , n26791 , n26517 );
and ( n26793 , n26789 , n26792 );
and ( n26794 , n26787 , n26792 );
or ( n26795 , n26790 , n26793 , n26794 );
xor ( n26796 , n26486 , n26490 );
xor ( n26797 , n26796 , n26495 );
and ( n26798 , n26795 , n26797 );
xor ( n26799 , n26426 , n26430 );
xor ( n26800 , n26799 , n26435 );
and ( n26801 , n26797 , n26800 );
and ( n26802 , n26795 , n26800 );
or ( n26803 , n26798 , n26801 , n26802 );
and ( n26804 , n26785 , n26803 );
xor ( n26805 , n26282 , n26295 );
xor ( n26806 , n26805 , n26298 );
and ( n26807 , n26803 , n26806 );
and ( n26808 , n26785 , n26806 );
or ( n26809 , n26804 , n26807 , n26808 );
xor ( n26810 , n26504 , n26536 );
xor ( n26811 , n26810 , n26539 );
and ( n26812 , n26809 , n26811 );
xor ( n26813 , n26412 , n26446 );
xor ( n26814 , n26813 , n26449 );
and ( n26815 , n26811 , n26814 );
and ( n26816 , n26809 , n26814 );
or ( n26817 , n26812 , n26815 , n26816 );
and ( n26818 , n26739 , n26817 );
xor ( n26819 , n26542 , n26544 );
xor ( n26820 , n26819 , n26547 );
and ( n26821 , n26817 , n26820 );
and ( n26822 , n26739 , n26820 );
or ( n26823 , n26818 , n26821 , n26822 );
and ( n26824 , n26592 , n26823 );
xor ( n26825 , n26345 , n26460 );
xor ( n26826 , n26825 , n26463 );
and ( n26827 , n26823 , n26826 );
and ( n26828 , n26592 , n26826 );
or ( n26829 , n26824 , n26827 , n26828 );
xor ( n26830 , n26258 , n26260 );
xor ( n26831 , n26830 , n26263 );
and ( n26832 , n26829 , n26831 );
xor ( n26833 , n26466 , n26558 );
xor ( n26834 , n26833 , n26561 );
and ( n26835 , n26831 , n26834 );
and ( n26836 , n26829 , n26834 );
or ( n26837 , n26832 , n26835 , n26836 );
and ( n26838 , n26574 , n26837 );
xor ( n26839 , n26574 , n26837 );
xor ( n26840 , n26829 , n26831 );
xor ( n26841 , n26840 , n26834 );
and ( n26842 , n21876 , n20955 );
and ( n26843 , n21704 , n20953 );
nor ( n26844 , n26842 , n26843 );
xnor ( n26845 , n26844 , n20780 );
and ( n26846 , n22235 , n20674 );
and ( n26847 , n21955 , n20672 );
nor ( n26848 , n26846 , n26847 );
xnor ( n26849 , n26848 , n20542 );
and ( n26850 , n26845 , n26849 );
buf ( n26851 , n19336 );
and ( n26852 , n26851 , n19419 );
and ( n26853 , n26849 , n26852 );
and ( n26854 , n26845 , n26852 );
or ( n26855 , n26850 , n26853 , n26854 );
and ( n26856 , n20182 , n23230 );
and ( n26857 , n20080 , n23228 );
nor ( n26858 , n26856 , n26857 );
xnor ( n26859 , n26858 , n22842 );
and ( n26860 , n20360 , n22859 );
and ( n26861 , n20268 , n22857 );
nor ( n26862 , n26860 , n26861 );
xnor ( n26863 , n26862 , n22418 );
and ( n26864 , n26859 , n26863 );
and ( n26865 , n20618 , n22381 );
and ( n26866 , n20452 , n22379 );
nor ( n26867 , n26865 , n26866 );
xnor ( n26868 , n26867 , n22228 );
and ( n26869 , n26863 , n26868 );
and ( n26870 , n26859 , n26868 );
or ( n26871 , n26864 , n26869 , n26870 );
and ( n26872 , n26855 , n26871 );
and ( n26873 , n20803 , n22048 );
and ( n26874 , n20666 , n22046 );
nor ( n26875 , n26873 , n26874 );
xnor ( n26876 , n26875 , n21853 );
and ( n26877 , n21072 , n21741 );
and ( n26878 , n20867 , n21739 );
nor ( n26879 , n26877 , n26878 );
xnor ( n26880 , n26879 , n21605 );
and ( n26881 , n26876 , n26880 );
not ( n26882 , n26658 );
and ( n26883 , n26880 , n26882 );
and ( n26884 , n26876 , n26882 );
or ( n26885 , n26881 , n26883 , n26884 );
and ( n26886 , n26871 , n26885 );
and ( n26887 , n26855 , n26885 );
or ( n26888 , n26872 , n26886 , n26887 );
xor ( n26889 , n26352 , n26356 );
xor ( n26890 , n26889 , n26361 );
and ( n26891 , n26888 , n26890 );
xor ( n26892 , n26520 , n26522 );
xor ( n26893 , n26892 , n26525 );
and ( n26894 , n26890 , n26893 );
and ( n26895 , n26888 , n26893 );
or ( n26896 , n26891 , n26894 , n26895 );
xor ( n26897 , n26364 , n26406 );
xor ( n26898 , n26897 , n26409 );
and ( n26899 , n26896 , n26898 );
xor ( n26900 , n26438 , n26440 );
xor ( n26901 , n26900 , n26443 );
and ( n26902 , n26898 , n26901 );
and ( n26903 , n26896 , n26901 );
or ( n26904 , n26899 , n26902 , n26903 );
xor ( n26905 , n26576 , n26578 );
xor ( n26906 , n26905 , n26581 );
and ( n26907 , n26904 , n26906 );
xor ( n26908 , n26638 , n26733 );
xor ( n26909 , n26908 , n26736 );
and ( n26910 , n26906 , n26909 );
and ( n26911 , n26904 , n26909 );
or ( n26912 , n26907 , n26910 , n26911 );
and ( n26913 , n20004 , n23641 );
and ( n26914 , n19946 , n23639 );
nor ( n26915 , n26913 , n26914 );
xnor ( n26916 , n26915 , n23213 );
and ( n26917 , n21302 , n21468 );
and ( n26918 , n21218 , n21466 );
nor ( n26919 , n26917 , n26918 );
xnor ( n26920 , n26919 , n21331 );
and ( n26921 , n26916 , n26920 );
and ( n26922 , n21612 , n21155 );
and ( n26923 , n21451 , n21153 );
nor ( n26924 , n26922 , n26923 );
xnor ( n26925 , n26924 , n20994 );
and ( n26926 , n26920 , n26925 );
and ( n26927 , n26916 , n26925 );
or ( n26928 , n26921 , n26926 , n26927 );
and ( n26929 , n19588 , n25383 );
and ( n26930 , n19510 , n25381 );
nor ( n26931 , n26929 , n26930 );
xnor ( n26932 , n26931 , n24885 );
and ( n26933 , n19637 , n24902 );
and ( n26934 , n19605 , n24900 );
nor ( n26935 , n26933 , n26934 );
xnor ( n26936 , n26935 , n24397 );
and ( n26937 , n26932 , n26936 );
and ( n26938 , n19881 , n23944 );
and ( n26939 , n19825 , n23942 );
nor ( n26940 , n26938 , n26939 );
xnor ( n26941 , n26940 , n23550 );
and ( n26942 , n26936 , n26941 );
and ( n26943 , n26932 , n26941 );
or ( n26944 , n26937 , n26942 , n26943 );
and ( n26945 , n26928 , n26944 );
and ( n26946 , n25765 , n19518 );
and ( n26947 , n25554 , n19516 );
nor ( n26948 , n26946 , n26947 );
xnor ( n26949 , n26948 , n19489 );
and ( n26950 , n26319 , n19459 );
and ( n26951 , n25974 , n19457 );
nor ( n26952 , n26950 , n26951 );
xnor ( n26953 , n26952 , n19416 );
and ( n26954 , n26949 , n26953 );
and ( n26955 , n26851 , n19424 );
and ( n26956 , n26422 , n19422 );
nor ( n26957 , n26955 , n26956 );
xnor ( n26958 , n26957 , n19431 );
and ( n26959 , n26953 , n26958 );
and ( n26960 , n26949 , n26958 );
or ( n26961 , n26954 , n26959 , n26960 );
and ( n26962 , n24521 , n19805 );
and ( n26963 , n24131 , n19803 );
nor ( n26964 , n26962 , n26963 );
xnor ( n26965 , n26964 , n19750 );
and ( n26966 , n24621 , n19688 );
and ( n26967 , n24527 , n19686 );
nor ( n26968 , n26966 , n26967 );
xnor ( n26969 , n26968 , n19655 );
and ( n26970 , n26965 , n26969 );
and ( n26971 , n25284 , n19596 );
and ( n26972 , n24940 , n19594 );
nor ( n26973 , n26971 , n26972 );
xnor ( n26974 , n26973 , n19545 );
and ( n26975 , n26969 , n26974 );
and ( n26976 , n26965 , n26974 );
or ( n26977 , n26970 , n26975 , n26976 );
and ( n26978 , n26961 , n26977 );
and ( n26979 , n19434 , n26349 );
and ( n26980 , n19418 , n26347 );
nor ( n26981 , n26979 , n26980 );
xnor ( n26982 , n26981 , n25893 );
and ( n26983 , n26977 , n26982 );
and ( n26984 , n26961 , n26982 );
or ( n26985 , n26978 , n26983 , n26984 );
and ( n26986 , n26944 , n26985 );
and ( n26987 , n26928 , n26985 );
or ( n26988 , n26945 , n26986 , n26987 );
xor ( n26989 , n25890 , n26365 );
xor ( n26990 , n26365 , n26366 );
not ( n26991 , n26990 );
and ( n26992 , n26989 , n26991 );
and ( n26993 , n19426 , n26992 );
not ( n26994 , n26993 );
xnor ( n26995 , n26994 , n26369 );
and ( n26996 , n19496 , n26027 );
and ( n26997 , n19469 , n26025 );
nor ( n26998 , n26996 , n26997 );
xnor ( n26999 , n26998 , n25499 );
and ( n27000 , n26995 , n26999 );
and ( n27001 , n19811 , n24376 );
and ( n27002 , n19721 , n24374 );
nor ( n27003 , n27001 , n27002 );
xnor ( n27004 , n27003 , n23927 );
and ( n27005 , n26999 , n27004 );
and ( n27006 , n26995 , n27004 );
or ( n27007 , n27000 , n27005 , n27006 );
xor ( n27008 , n26596 , n26600 );
xor ( n27009 , n27008 , n26605 );
and ( n27010 , n27007 , n27009 );
xor ( n27011 , n26659 , n26663 );
xor ( n27012 , n27011 , n26668 );
and ( n27013 , n27009 , n27012 );
and ( n27014 , n27007 , n27012 );
or ( n27015 , n27010 , n27013 , n27014 );
and ( n27016 , n26988 , n27015 );
xor ( n27017 , n26608 , n26624 );
xor ( n27018 , n27017 , n26627 );
and ( n27019 , n27015 , n27018 );
and ( n27020 , n26988 , n27018 );
or ( n27021 , n27016 , n27019 , n27020 );
xor ( n27022 , n26528 , n26530 );
xor ( n27023 , n27022 , n26533 );
and ( n27024 , n27021 , n27023 );
xor ( n27025 , n26630 , n26632 );
xor ( n27026 , n27025 , n26635 );
and ( n27027 , n27023 , n27026 );
and ( n27028 , n27021 , n27026 );
or ( n27029 , n27024 , n27027 , n27028 );
buf ( n27030 , n19402 );
buf ( n27031 , n19403 );
and ( n27032 , n27030 , n27031 );
not ( n27033 , n27032 );
and ( n27034 , n26366 , n27033 );
not ( n27035 , n27034 );
and ( n27036 , n22198 , n20674 );
and ( n27037 , n22235 , n20672 );
nor ( n27038 , n27036 , n27037 );
xnor ( n27039 , n27038 , n20542 );
and ( n27040 , n27035 , n27039 );
and ( n27041 , n22756 , n20460 );
and ( n27042 , n22425 , n20458 );
nor ( n27043 , n27041 , n27042 );
xnor ( n27044 , n27043 , n20337 );
and ( n27045 , n27039 , n27044 );
and ( n27046 , n27035 , n27044 );
or ( n27047 , n27040 , n27045 , n27046 );
and ( n27048 , n23141 , n20276 );
and ( n27049 , n22916 , n20274 );
nor ( n27050 , n27048 , n27049 );
xnor ( n27051 , n27050 , n20175 );
and ( n27052 , n23381 , n20114 );
and ( n27053 , n23271 , n20112 );
nor ( n27054 , n27052 , n27053 );
xnor ( n27055 , n27054 , n19997 );
and ( n27056 , n27051 , n27055 );
and ( n27057 , n23968 , n19894 );
and ( n27058 , n23573 , n19892 );
nor ( n27059 , n27057 , n27058 );
xnor ( n27060 , n27059 , n19858 );
and ( n27061 , n27055 , n27060 );
and ( n27062 , n27051 , n27060 );
or ( n27063 , n27056 , n27061 , n27062 );
and ( n27064 , n27047 , n27063 );
xor ( n27065 , n26676 , n26680 );
xor ( n27066 , n27065 , n26685 );
and ( n27067 , n27063 , n27066 );
and ( n27068 , n27047 , n27066 );
or ( n27069 , n27064 , n27067 , n27068 );
xor ( n27070 , n26707 , n26711 );
xor ( n27071 , n27070 , n26716 );
and ( n27072 , n27069 , n27071 );
xor ( n27073 , n26642 , n26646 );
xor ( n27074 , n27073 , n26651 );
and ( n27075 , n27071 , n27074 );
and ( n27076 , n27069 , n27074 );
or ( n27077 , n27072 , n27075 , n27076 );
xor ( n27078 , n26612 , n26616 );
xor ( n27079 , n27078 , n26621 );
xor ( n27080 , n26688 , n26692 );
xor ( n27081 , n27080 , n26697 );
and ( n27082 , n27079 , n27081 );
xor ( n27083 , n26755 , n26771 );
xor ( n27084 , n27083 , n26774 );
and ( n27085 , n27081 , n27084 );
and ( n27086 , n27079 , n27084 );
or ( n27087 , n27082 , n27085 , n27086 );
and ( n27088 , n27077 , n27087 );
xor ( n27089 , n26654 , n26671 );
xor ( n27090 , n27089 , n26700 );
and ( n27091 , n27087 , n27090 );
and ( n27092 , n27077 , n27090 );
or ( n27093 , n27088 , n27091 , n27092 );
xor ( n27094 , n26703 , n26727 );
xor ( n27095 , n27094 , n26730 );
and ( n27096 , n27093 , n27095 );
xor ( n27097 , n26785 , n26803 );
xor ( n27098 , n27097 , n26806 );
and ( n27099 , n27095 , n27098 );
and ( n27100 , n27093 , n27098 );
or ( n27101 , n27096 , n27099 , n27100 );
and ( n27102 , n27029 , n27101 );
xor ( n27103 , n26809 , n26811 );
xor ( n27104 , n27103 , n26814 );
and ( n27105 , n27101 , n27104 );
and ( n27106 , n27029 , n27104 );
or ( n27107 , n27102 , n27105 , n27106 );
and ( n27108 , n26912 , n27107 );
xor ( n27109 , n26584 , n26586 );
xor ( n27110 , n27109 , n26589 );
and ( n27111 , n27107 , n27110 );
and ( n27112 , n26912 , n27110 );
or ( n27113 , n27108 , n27111 , n27112 );
xor ( n27114 , n26550 , n26552 );
xor ( n27115 , n27114 , n26555 );
and ( n27116 , n27113 , n27115 );
xor ( n27117 , n26592 , n26823 );
xor ( n27118 , n27117 , n26826 );
and ( n27119 , n27115 , n27118 );
and ( n27120 , n27113 , n27118 );
or ( n27121 , n27116 , n27119 , n27120 );
and ( n27122 , n26841 , n27121 );
xor ( n27123 , n26841 , n27121 );
xor ( n27124 , n27113 , n27115 );
xor ( n27125 , n27124 , n27118 );
and ( n27126 , n20080 , n23641 );
and ( n27127 , n20004 , n23639 );
nor ( n27128 , n27126 , n27127 );
xnor ( n27129 , n27128 , n23213 );
and ( n27130 , n21955 , n20955 );
and ( n27131 , n21876 , n20953 );
nor ( n27132 , n27130 , n27131 );
xnor ( n27133 , n27132 , n20780 );
and ( n27134 , n27129 , n27133 );
buf ( n27135 , n19337 );
and ( n27136 , n27135 , n19419 );
and ( n27137 , n27133 , n27136 );
and ( n27138 , n27129 , n27136 );
or ( n27139 , n27134 , n27137 , n27138 );
xor ( n27140 , n26743 , n26747 );
xor ( n27141 , n27140 , n26752 );
and ( n27142 , n27139 , n27141 );
xor ( n27143 , n26759 , n26763 );
xor ( n27144 , n27143 , n26768 );
and ( n27145 , n27141 , n27144 );
and ( n27146 , n27139 , n27144 );
or ( n27147 , n27142 , n27145 , n27146 );
and ( n27148 , n20666 , n22381 );
and ( n27149 , n20618 , n22379 );
nor ( n27150 , n27148 , n27149 );
xnor ( n27151 , n27150 , n22228 );
and ( n27152 , n20867 , n22048 );
and ( n27153 , n20803 , n22046 );
nor ( n27154 , n27152 , n27153 );
xnor ( n27155 , n27154 , n21853 );
and ( n27156 , n27151 , n27155 );
and ( n27157 , n21218 , n21741 );
and ( n27158 , n21072 , n21739 );
nor ( n27159 , n27157 , n27158 );
xnor ( n27160 , n27159 , n21605 );
and ( n27161 , n27155 , n27160 );
and ( n27162 , n27151 , n27160 );
or ( n27163 , n27156 , n27161 , n27162 );
and ( n27164 , n20268 , n23230 );
and ( n27165 , n20182 , n23228 );
nor ( n27166 , n27164 , n27165 );
xnor ( n27167 , n27166 , n22842 );
and ( n27168 , n20452 , n22859 );
and ( n27169 , n20360 , n22857 );
nor ( n27170 , n27168 , n27169 );
xnor ( n27171 , n27170 , n22418 );
and ( n27172 , n27167 , n27171 );
and ( n27173 , n21704 , n21155 );
and ( n27174 , n21612 , n21153 );
nor ( n27175 , n27173 , n27174 );
xnor ( n27176 , n27175 , n20994 );
and ( n27177 , n27171 , n27176 );
and ( n27178 , n27167 , n27176 );
or ( n27179 , n27172 , n27177 , n27178 );
and ( n27180 , n27163 , n27179 );
xor ( n27181 , n26845 , n26849 );
xor ( n27182 , n27181 , n26852 );
and ( n27183 , n27179 , n27182 );
and ( n27184 , n27163 , n27182 );
or ( n27185 , n27180 , n27183 , n27184 );
and ( n27186 , n27147 , n27185 );
xor ( n27187 , n26787 , n26789 );
xor ( n27188 , n27187 , n26792 );
and ( n27189 , n27185 , n27188 );
and ( n27190 , n27147 , n27188 );
or ( n27191 , n27186 , n27189 , n27190 );
xor ( n27192 , n26719 , n26721 );
xor ( n27193 , n27192 , n26724 );
and ( n27194 , n27191 , n27193 );
xor ( n27195 , n26795 , n26797 );
xor ( n27196 , n27195 , n26800 );
and ( n27197 , n27193 , n27196 );
and ( n27198 , n27191 , n27196 );
or ( n27199 , n27194 , n27197 , n27198 );
and ( n27200 , n19510 , n26027 );
and ( n27201 , n19496 , n26025 );
nor ( n27202 , n27200 , n27201 );
xnor ( n27203 , n27202 , n25499 );
and ( n27204 , n19605 , n25383 );
and ( n27205 , n19588 , n25381 );
nor ( n27206 , n27204 , n27205 );
xnor ( n27207 , n27206 , n24885 );
and ( n27208 , n27203 , n27207 );
and ( n27209 , n19721 , n24902 );
and ( n27210 , n19637 , n24900 );
nor ( n27211 , n27209 , n27210 );
xnor ( n27212 , n27211 , n24397 );
and ( n27213 , n27207 , n27212 );
and ( n27214 , n27203 , n27212 );
or ( n27215 , n27208 , n27213 , n27214 );
and ( n27216 , n22916 , n20460 );
and ( n27217 , n22756 , n20458 );
nor ( n27218 , n27216 , n27217 );
xnor ( n27219 , n27218 , n20337 );
buf ( n27220 , n27219 );
and ( n27221 , n19946 , n23944 );
and ( n27222 , n19881 , n23942 );
nor ( n27223 , n27221 , n27222 );
xnor ( n27224 , n27223 , n23550 );
and ( n27225 , n27220 , n27224 );
and ( n27226 , n21451 , n21468 );
and ( n27227 , n21302 , n21466 );
nor ( n27228 , n27226 , n27227 );
xnor ( n27229 , n27228 , n21331 );
and ( n27230 , n27224 , n27229 );
and ( n27231 , n27220 , n27229 );
or ( n27232 , n27225 , n27230 , n27231 );
and ( n27233 , n27215 , n27232 );
and ( n27234 , n22425 , n20674 );
and ( n27235 , n22198 , n20672 );
nor ( n27236 , n27234 , n27235 );
xnor ( n27237 , n27236 , n20542 );
and ( n27238 , n24527 , n19805 );
and ( n27239 , n24521 , n19803 );
nor ( n27240 , n27238 , n27239 );
xnor ( n27241 , n27240 , n19750 );
and ( n27242 , n27237 , n27241 );
and ( n27243 , n25554 , n19596 );
and ( n27244 , n25284 , n19594 );
nor ( n27245 , n27243 , n27244 );
xnor ( n27246 , n27245 , n19545 );
and ( n27247 , n27241 , n27246 );
and ( n27248 , n27237 , n27246 );
or ( n27249 , n27242 , n27247 , n27248 );
and ( n27250 , n24940 , n19688 );
and ( n27251 , n24621 , n19686 );
nor ( n27252 , n27250 , n27251 );
xnor ( n27253 , n27252 , n19655 );
and ( n27254 , n25974 , n19518 );
and ( n27255 , n25765 , n19516 );
nor ( n27256 , n27254 , n27255 );
xnor ( n27257 , n27256 , n19489 );
and ( n27258 , n27253 , n27257 );
and ( n27259 , n26422 , n19459 );
and ( n27260 , n26319 , n19457 );
nor ( n27261 , n27259 , n27260 );
xnor ( n27262 , n27261 , n19416 );
and ( n27263 , n27257 , n27262 );
and ( n27264 , n27253 , n27262 );
or ( n27265 , n27258 , n27263 , n27264 );
and ( n27266 , n27249 , n27265 );
and ( n27267 , n19418 , n26992 );
and ( n27268 , n19426 , n26990 );
nor ( n27269 , n27267 , n27268 );
xnor ( n27270 , n27269 , n26369 );
and ( n27271 , n27265 , n27270 );
and ( n27272 , n27249 , n27270 );
or ( n27273 , n27266 , n27271 , n27272 );
and ( n27274 , n27232 , n27273 );
and ( n27275 , n27215 , n27273 );
or ( n27276 , n27233 , n27274 , n27275 );
and ( n27277 , n23271 , n20276 );
and ( n27278 , n23141 , n20274 );
nor ( n27279 , n27277 , n27278 );
xnor ( n27280 , n27279 , n20175 );
and ( n27281 , n23573 , n20114 );
and ( n27282 , n23381 , n20112 );
nor ( n27283 , n27281 , n27282 );
xnor ( n27284 , n27283 , n19997 );
and ( n27285 , n27280 , n27284 );
and ( n27286 , n24131 , n19894 );
and ( n27287 , n23968 , n19892 );
nor ( n27288 , n27286 , n27287 );
xnor ( n27289 , n27288 , n19858 );
and ( n27290 , n27284 , n27289 );
and ( n27291 , n27280 , n27289 );
or ( n27292 , n27285 , n27290 , n27291 );
and ( n27293 , n19469 , n26349 );
and ( n27294 , n19434 , n26347 );
nor ( n27295 , n27293 , n27294 );
xnor ( n27296 , n27295 , n25893 );
and ( n27297 , n27292 , n27296 );
and ( n27298 , n19825 , n24376 );
and ( n27299 , n19811 , n24374 );
nor ( n27300 , n27298 , n27299 );
xnor ( n27301 , n27300 , n23927 );
and ( n27302 , n27296 , n27301 );
and ( n27303 , n27292 , n27301 );
or ( n27304 , n27297 , n27302 , n27303 );
xor ( n27305 , n26916 , n26920 );
xor ( n27306 , n27305 , n26925 );
and ( n27307 , n27304 , n27306 );
xor ( n27308 , n26859 , n26863 );
xor ( n27309 , n27308 , n26868 );
and ( n27310 , n27306 , n27309 );
and ( n27311 , n27304 , n27309 );
or ( n27312 , n27307 , n27310 , n27311 );
and ( n27313 , n27276 , n27312 );
xor ( n27314 , n26855 , n26871 );
xor ( n27315 , n27314 , n26885 );
and ( n27316 , n27312 , n27315 );
and ( n27317 , n27276 , n27315 );
or ( n27318 , n27313 , n27316 , n27317 );
xor ( n27319 , n26777 , n26779 );
xor ( n27320 , n27319 , n26782 );
and ( n27321 , n27318 , n27320 );
xor ( n27322 , n26888 , n26890 );
xor ( n27323 , n27322 , n26893 );
and ( n27324 , n27320 , n27323 );
and ( n27325 , n27318 , n27323 );
or ( n27326 , n27321 , n27324 , n27325 );
and ( n27327 , n27199 , n27326 );
xor ( n27328 , n26896 , n26898 );
xor ( n27329 , n27328 , n26901 );
and ( n27330 , n27326 , n27329 );
and ( n27331 , n27199 , n27329 );
or ( n27332 , n27327 , n27330 , n27331 );
xor ( n27333 , n26932 , n26936 );
xor ( n27334 , n27333 , n26941 );
xor ( n27335 , n26995 , n26999 );
xor ( n27336 , n27335 , n27004 );
and ( n27337 , n27334 , n27336 );
xor ( n27338 , n26961 , n26977 );
xor ( n27339 , n27338 , n26982 );
and ( n27340 , n27336 , n27339 );
and ( n27341 , n27334 , n27339 );
or ( n27342 , n27337 , n27340 , n27341 );
and ( n27343 , n22235 , n20955 );
and ( n27344 , n21955 , n20953 );
nor ( n27345 , n27343 , n27344 );
xnor ( n27346 , n27345 , n20780 );
and ( n27347 , n27135 , n19424 );
and ( n27348 , n26851 , n19422 );
nor ( n27349 , n27347 , n27348 );
xnor ( n27350 , n27349 , n19431 );
and ( n27351 , n27346 , n27350 );
buf ( n27352 , n19338 );
and ( n27353 , n27352 , n19419 );
and ( n27354 , n27350 , n27353 );
and ( n27355 , n27346 , n27353 );
or ( n27356 , n27351 , n27354 , n27355 );
xor ( n27357 , n27035 , n27039 );
xor ( n27358 , n27357 , n27044 );
and ( n27359 , n27356 , n27358 );
xor ( n27360 , n26949 , n26953 );
xor ( n27361 , n27360 , n26958 );
and ( n27362 , n27358 , n27361 );
and ( n27363 , n27356 , n27361 );
or ( n27364 , n27359 , n27362 , n27363 );
xor ( n27365 , n26876 , n26880 );
xor ( n27366 , n27365 , n26882 );
and ( n27367 , n27364 , n27366 );
xor ( n27368 , n27047 , n27063 );
xor ( n27369 , n27368 , n27066 );
and ( n27370 , n27366 , n27369 );
and ( n27371 , n27364 , n27369 );
or ( n27372 , n27367 , n27370 , n27371 );
and ( n27373 , n27342 , n27372 );
xor ( n27374 , n26928 , n26944 );
xor ( n27375 , n27374 , n26985 );
and ( n27376 , n27372 , n27375 );
and ( n27377 , n27342 , n27375 );
or ( n27378 , n27373 , n27376 , n27377 );
xor ( n27379 , n27077 , n27087 );
xor ( n27380 , n27379 , n27090 );
and ( n27381 , n27378 , n27380 );
xor ( n27382 , n26988 , n27015 );
xor ( n27383 , n27382 , n27018 );
and ( n27384 , n27380 , n27383 );
and ( n27385 , n27378 , n27383 );
or ( n27386 , n27381 , n27384 , n27385 );
xor ( n27387 , n27021 , n27023 );
xor ( n27388 , n27387 , n27026 );
and ( n27389 , n27386 , n27388 );
xor ( n27390 , n27093 , n27095 );
xor ( n27391 , n27390 , n27098 );
and ( n27392 , n27388 , n27391 );
and ( n27393 , n27386 , n27391 );
or ( n27394 , n27389 , n27392 , n27393 );
and ( n27395 , n27332 , n27394 );
xor ( n27396 , n26904 , n26906 );
xor ( n27397 , n27396 , n26909 );
and ( n27398 , n27394 , n27397 );
and ( n27399 , n27332 , n27397 );
or ( n27400 , n27395 , n27398 , n27399 );
xor ( n27401 , n26739 , n26817 );
xor ( n27402 , n27401 , n26820 );
and ( n27403 , n27400 , n27402 );
xor ( n27404 , n26912 , n27107 );
xor ( n27405 , n27404 , n27110 );
and ( n27406 , n27402 , n27405 );
and ( n27407 , n27400 , n27405 );
or ( n27408 , n27403 , n27406 , n27407 );
and ( n27409 , n27125 , n27408 );
xor ( n27410 , n27125 , n27408 );
xor ( n27411 , n27400 , n27402 );
xor ( n27412 , n27411 , n27405 );
xor ( n27413 , n27007 , n27009 );
xor ( n27414 , n27413 , n27012 );
xor ( n27415 , n27069 , n27071 );
xor ( n27416 , n27415 , n27074 );
and ( n27417 , n27414 , n27416 );
xor ( n27418 , n27079 , n27081 );
xor ( n27419 , n27418 , n27084 );
and ( n27420 , n27416 , n27419 );
and ( n27421 , n27414 , n27419 );
or ( n27422 , n27417 , n27420 , n27421 );
and ( n27423 , n21072 , n22048 );
and ( n27424 , n20867 , n22046 );
nor ( n27425 , n27423 , n27424 );
xnor ( n27426 , n27425 , n21853 );
and ( n27427 , n21302 , n21741 );
and ( n27428 , n21218 , n21739 );
nor ( n27429 , n27427 , n27428 );
xnor ( n27430 , n27429 , n21605 );
and ( n27431 , n27426 , n27430 );
and ( n27432 , n21612 , n21468 );
and ( n27433 , n21451 , n21466 );
nor ( n27434 , n27432 , n27433 );
xnor ( n27435 , n27434 , n21331 );
and ( n27436 , n27430 , n27435 );
and ( n27437 , n27426 , n27435 );
or ( n27438 , n27431 , n27436 , n27437 );
and ( n27439 , n23141 , n20460 );
and ( n27440 , n22916 , n20458 );
nor ( n27441 , n27439 , n27440 );
xnor ( n27442 , n27441 , n20337 );
and ( n27443 , n23381 , n20276 );
and ( n27444 , n23271 , n20274 );
nor ( n27445 , n27443 , n27444 );
xnor ( n27446 , n27445 , n20175 );
and ( n27447 , n27442 , n27446 );
and ( n27448 , n23968 , n20114 );
and ( n27449 , n23573 , n20112 );
nor ( n27450 , n27448 , n27449 );
xnor ( n27451 , n27450 , n19997 );
and ( n27452 , n27446 , n27451 );
and ( n27453 , n27442 , n27451 );
or ( n27454 , n27447 , n27452 , n27453 );
and ( n27455 , n24521 , n19894 );
and ( n27456 , n24131 , n19892 );
nor ( n27457 , n27455 , n27456 );
xnor ( n27458 , n27457 , n19858 );
and ( n27459 , n24621 , n19805 );
and ( n27460 , n24527 , n19803 );
nor ( n27461 , n27459 , n27460 );
xnor ( n27462 , n27461 , n19750 );
and ( n27463 , n27458 , n27462 );
and ( n27464 , n25284 , n19688 );
and ( n27465 , n24940 , n19686 );
nor ( n27466 , n27464 , n27465 );
xnor ( n27467 , n27466 , n19655 );
and ( n27468 , n27462 , n27467 );
and ( n27469 , n27458 , n27467 );
or ( n27470 , n27463 , n27468 , n27469 );
and ( n27471 , n27454 , n27470 );
and ( n27472 , n20004 , n23944 );
and ( n27473 , n19946 , n23942 );
nor ( n27474 , n27472 , n27473 );
xnor ( n27475 , n27474 , n23550 );
and ( n27476 , n27470 , n27475 );
and ( n27477 , n27454 , n27475 );
or ( n27478 , n27471 , n27476 , n27477 );
and ( n27479 , n27438 , n27478 );
and ( n27480 , n20618 , n22859 );
and ( n27481 , n20452 , n22857 );
nor ( n27482 , n27480 , n27481 );
xnor ( n27483 , n27482 , n22418 );
and ( n27484 , n20803 , n22381 );
and ( n27485 , n20666 , n22379 );
nor ( n27486 , n27484 , n27485 );
xnor ( n27487 , n27486 , n22228 );
and ( n27488 , n27483 , n27487 );
not ( n27489 , n27219 );
and ( n27490 , n27487 , n27489 );
and ( n27491 , n27483 , n27489 );
or ( n27492 , n27488 , n27490 , n27491 );
and ( n27493 , n27478 , n27492 );
and ( n27494 , n27438 , n27492 );
or ( n27495 , n27479 , n27493 , n27494 );
and ( n27496 , n20182 , n23641 );
and ( n27497 , n20080 , n23639 );
nor ( n27498 , n27496 , n27497 );
xnor ( n27499 , n27498 , n23213 );
and ( n27500 , n20360 , n23230 );
and ( n27501 , n20268 , n23228 );
nor ( n27502 , n27500 , n27501 );
xnor ( n27503 , n27502 , n22842 );
and ( n27504 , n27499 , n27503 );
and ( n27505 , n21876 , n21155 );
and ( n27506 , n21704 , n21153 );
nor ( n27507 , n27505 , n27506 );
xnor ( n27508 , n27507 , n20994 );
and ( n27509 , n27503 , n27508 );
and ( n27510 , n27499 , n27508 );
or ( n27511 , n27504 , n27509 , n27510 );
xor ( n27512 , n27051 , n27055 );
xor ( n27513 , n27512 , n27060 );
and ( n27514 , n27511 , n27513 );
xor ( n27515 , n26965 , n26969 );
xor ( n27516 , n27515 , n26974 );
and ( n27517 , n27513 , n27516 );
and ( n27518 , n27511 , n27516 );
or ( n27519 , n27514 , n27517 , n27518 );
and ( n27520 , n27495 , n27519 );
xor ( n27521 , n27139 , n27141 );
xor ( n27522 , n27521 , n27144 );
and ( n27523 , n27519 , n27522 );
and ( n27524 , n27495 , n27522 );
or ( n27525 , n27520 , n27523 , n27524 );
xor ( n27526 , n26366 , n27030 );
xor ( n27527 , n27030 , n27031 );
not ( n27528 , n27527 );
and ( n27529 , n27526 , n27528 );
and ( n27530 , n19426 , n27529 );
not ( n27531 , n27530 );
xnor ( n27532 , n27531 , n27034 );
and ( n27533 , n19637 , n25383 );
and ( n27534 , n19605 , n25381 );
nor ( n27535 , n27533 , n27534 );
xnor ( n27536 , n27535 , n24885 );
and ( n27537 , n27532 , n27536 );
and ( n27538 , n19811 , n24902 );
and ( n27539 , n19721 , n24900 );
nor ( n27540 , n27538 , n27539 );
xnor ( n27541 , n27540 , n24397 );
and ( n27542 , n27536 , n27541 );
and ( n27543 , n27532 , n27541 );
or ( n27544 , n27537 , n27542 , n27543 );
buf ( n27545 , n19404 );
buf ( n27546 , n19405 );
and ( n27547 , n27545 , n27546 );
not ( n27548 , n27547 );
and ( n27549 , n27031 , n27548 );
not ( n27550 , n27549 );
and ( n27551 , n22198 , n20955 );
and ( n27552 , n22235 , n20953 );
nor ( n27553 , n27551 , n27552 );
xnor ( n27554 , n27553 , n20780 );
and ( n27555 , n27550 , n27554 );
and ( n27556 , n22756 , n20674 );
and ( n27557 , n22425 , n20672 );
nor ( n27558 , n27556 , n27557 );
xnor ( n27559 , n27558 , n20542 );
and ( n27560 , n27554 , n27559 );
and ( n27561 , n27550 , n27559 );
or ( n27562 , n27555 , n27560 , n27561 );
and ( n27563 , n19496 , n26349 );
and ( n27564 , n19469 , n26347 );
nor ( n27565 , n27563 , n27564 );
xnor ( n27566 , n27565 , n25893 );
and ( n27567 , n27562 , n27566 );
and ( n27568 , n19881 , n24376 );
and ( n27569 , n19825 , n24374 );
nor ( n27570 , n27568 , n27569 );
xnor ( n27571 , n27570 , n23927 );
and ( n27572 , n27566 , n27571 );
and ( n27573 , n27562 , n27571 );
or ( n27574 , n27567 , n27572 , n27573 );
and ( n27575 , n27544 , n27574 );
xor ( n27576 , n27220 , n27224 );
xor ( n27577 , n27576 , n27229 );
and ( n27578 , n27574 , n27577 );
and ( n27579 , n27544 , n27577 );
or ( n27580 , n27575 , n27578 , n27579 );
and ( n27581 , n25765 , n19596 );
and ( n27582 , n25554 , n19594 );
nor ( n27583 , n27581 , n27582 );
xnor ( n27584 , n27583 , n19545 );
and ( n27585 , n26319 , n19518 );
and ( n27586 , n25974 , n19516 );
nor ( n27587 , n27585 , n27586 );
xnor ( n27588 , n27587 , n19489 );
and ( n27589 , n27584 , n27588 );
and ( n27590 , n26851 , n19459 );
and ( n27591 , n26422 , n19457 );
nor ( n27592 , n27590 , n27591 );
xnor ( n27593 , n27592 , n19416 );
and ( n27594 , n27588 , n27593 );
and ( n27595 , n27584 , n27593 );
or ( n27596 , n27589 , n27594 , n27595 );
and ( n27597 , n19434 , n26992 );
and ( n27598 , n19418 , n26990 );
nor ( n27599 , n27597 , n27598 );
xnor ( n27600 , n27599 , n26369 );
and ( n27601 , n27596 , n27600 );
and ( n27602 , n19588 , n26027 );
and ( n27603 , n19510 , n26025 );
nor ( n27604 , n27602 , n27603 );
xnor ( n27605 , n27604 , n25499 );
and ( n27606 , n27600 , n27605 );
and ( n27607 , n27596 , n27605 );
or ( n27608 , n27601 , n27606 , n27607 );
xor ( n27609 , n27151 , n27155 );
xor ( n27610 , n27609 , n27160 );
and ( n27611 , n27608 , n27610 );
xor ( n27612 , n27167 , n27171 );
xor ( n27613 , n27612 , n27176 );
and ( n27614 , n27610 , n27613 );
and ( n27615 , n27608 , n27613 );
or ( n27616 , n27611 , n27614 , n27615 );
and ( n27617 , n27580 , n27616 );
xor ( n27618 , n27163 , n27179 );
xor ( n27619 , n27618 , n27182 );
and ( n27620 , n27616 , n27619 );
and ( n27621 , n27580 , n27619 );
or ( n27622 , n27617 , n27620 , n27621 );
and ( n27623 , n27525 , n27622 );
xor ( n27624 , n27147 , n27185 );
xor ( n27625 , n27624 , n27188 );
and ( n27626 , n27622 , n27625 );
and ( n27627 , n27525 , n27625 );
or ( n27628 , n27623 , n27626 , n27627 );
and ( n27629 , n27422 , n27628 );
xor ( n27630 , n27191 , n27193 );
xor ( n27631 , n27630 , n27196 );
and ( n27632 , n27628 , n27631 );
and ( n27633 , n27422 , n27631 );
or ( n27634 , n27629 , n27632 , n27633 );
xor ( n27635 , n27129 , n27133 );
xor ( n27636 , n27635 , n27136 );
xor ( n27637 , n27292 , n27296 );
xor ( n27638 , n27637 , n27301 );
and ( n27639 , n27636 , n27638 );
xor ( n27640 , n27249 , n27265 );
xor ( n27641 , n27640 , n27270 );
and ( n27642 , n27638 , n27641 );
and ( n27643 , n27636 , n27641 );
or ( n27644 , n27639 , n27642 , n27643 );
xor ( n27645 , n27215 , n27232 );
xor ( n27646 , n27645 , n27273 );
and ( n27647 , n27644 , n27646 );
xor ( n27648 , n27304 , n27306 );
xor ( n27649 , n27648 , n27309 );
and ( n27650 , n27646 , n27649 );
and ( n27651 , n27644 , n27649 );
or ( n27652 , n27647 , n27650 , n27651 );
xor ( n27653 , n27276 , n27312 );
xor ( n27654 , n27653 , n27315 );
and ( n27655 , n27652 , n27654 );
xor ( n27656 , n27342 , n27372 );
xor ( n27657 , n27656 , n27375 );
and ( n27658 , n27654 , n27657 );
and ( n27659 , n27652 , n27657 );
or ( n27660 , n27655 , n27658 , n27659 );
xor ( n27661 , n27318 , n27320 );
xor ( n27662 , n27661 , n27323 );
and ( n27663 , n27660 , n27662 );
xor ( n27664 , n27378 , n27380 );
xor ( n27665 , n27664 , n27383 );
and ( n27666 , n27662 , n27665 );
and ( n27667 , n27660 , n27665 );
or ( n27668 , n27663 , n27666 , n27667 );
and ( n27669 , n27634 , n27668 );
xor ( n27670 , n27199 , n27326 );
xor ( n27671 , n27670 , n27329 );
and ( n27672 , n27668 , n27671 );
and ( n27673 , n27634 , n27671 );
or ( n27674 , n27669 , n27672 , n27673 );
xor ( n27675 , n27029 , n27101 );
xor ( n27676 , n27675 , n27104 );
and ( n27677 , n27674 , n27676 );
xor ( n27678 , n27332 , n27394 );
xor ( n27679 , n27678 , n27397 );
and ( n27680 , n27676 , n27679 );
and ( n27681 , n27674 , n27679 );
or ( n27682 , n27677 , n27680 , n27681 );
and ( n27683 , n27412 , n27682 );
xor ( n27684 , n27412 , n27682 );
xor ( n27685 , n27674 , n27676 );
xor ( n27686 , n27685 , n27679 );
xor ( n27687 , n27280 , n27284 );
xor ( n27688 , n27687 , n27289 );
xor ( n27689 , n27346 , n27350 );
xor ( n27690 , n27689 , n27353 );
and ( n27691 , n27688 , n27690 );
xor ( n27692 , n27253 , n27257 );
xor ( n27693 , n27692 , n27262 );
and ( n27694 , n27690 , n27693 );
and ( n27695 , n27688 , n27693 );
or ( n27696 , n27691 , n27694 , n27695 );
xor ( n27697 , n27203 , n27207 );
xor ( n27698 , n27697 , n27212 );
and ( n27699 , n27696 , n27698 );
xor ( n27700 , n27511 , n27513 );
xor ( n27701 , n27700 , n27516 );
and ( n27702 , n27698 , n27701 );
and ( n27703 , n27696 , n27701 );
or ( n27704 , n27699 , n27702 , n27703 );
xor ( n27705 , n27334 , n27336 );
xor ( n27706 , n27705 , n27339 );
and ( n27707 , n27704 , n27706 );
xor ( n27708 , n27364 , n27366 );
xor ( n27709 , n27708 , n27369 );
and ( n27710 , n27706 , n27709 );
and ( n27711 , n27704 , n27709 );
or ( n27712 , n27707 , n27710 , n27711 );
and ( n27713 , n20452 , n23230 );
and ( n27714 , n20360 , n23228 );
nor ( n27715 , n27713 , n27714 );
xnor ( n27716 , n27715 , n22842 );
and ( n27717 , n20666 , n22859 );
and ( n27718 , n20618 , n22857 );
nor ( n27719 , n27717 , n27718 );
xnor ( n27720 , n27719 , n22418 );
and ( n27721 , n27716 , n27720 );
and ( n27722 , n20867 , n22381 );
and ( n27723 , n20803 , n22379 );
nor ( n27724 , n27722 , n27723 );
xnor ( n27725 , n27724 , n22228 );
and ( n27726 , n27720 , n27725 );
and ( n27727 , n27716 , n27725 );
or ( n27728 , n27721 , n27726 , n27727 );
and ( n27729 , n22916 , n20674 );
and ( n27730 , n22756 , n20672 );
nor ( n27731 , n27729 , n27730 );
xnor ( n27732 , n27731 , n20542 );
buf ( n27733 , n27732 );
and ( n27734 , n21218 , n22048 );
and ( n27735 , n21072 , n22046 );
nor ( n27736 , n27734 , n27735 );
xnor ( n27737 , n27736 , n21853 );
and ( n27738 , n27733 , n27737 );
and ( n27739 , n21451 , n21741 );
and ( n27740 , n21302 , n21739 );
nor ( n27741 , n27739 , n27740 );
xnor ( n27742 , n27741 , n21605 );
and ( n27743 , n27737 , n27742 );
and ( n27744 , n27733 , n27742 );
or ( n27745 , n27738 , n27743 , n27744 );
and ( n27746 , n27728 , n27745 );
and ( n27747 , n27135 , n19459 );
and ( n27748 , n26851 , n19457 );
nor ( n27749 , n27747 , n27748 );
xnor ( n27750 , n27749 , n19416 );
buf ( n27751 , n19339 );
and ( n27752 , n27751 , n19424 );
and ( n27753 , n27352 , n19422 );
nor ( n27754 , n27752 , n27753 );
xnor ( n27755 , n27754 , n19431 );
and ( n27756 , n27750 , n27755 );
buf ( n27757 , n19340 );
and ( n27758 , n27757 , n19419 );
and ( n27759 , n27755 , n27758 );
and ( n27760 , n27750 , n27758 );
or ( n27761 , n27756 , n27759 , n27760 );
and ( n27762 , n24940 , n19805 );
and ( n27763 , n24621 , n19803 );
nor ( n27764 , n27762 , n27763 );
xnor ( n27765 , n27764 , n19750 );
and ( n27766 , n25974 , n19596 );
and ( n27767 , n25765 , n19594 );
nor ( n27768 , n27766 , n27767 );
xnor ( n27769 , n27768 , n19545 );
and ( n27770 , n27765 , n27769 );
and ( n27771 , n26422 , n19518 );
and ( n27772 , n26319 , n19516 );
nor ( n27773 , n27771 , n27772 );
xnor ( n27774 , n27773 , n19489 );
and ( n27775 , n27769 , n27774 );
and ( n27776 , n27765 , n27774 );
or ( n27777 , n27770 , n27775 , n27776 );
and ( n27778 , n27761 , n27777 );
and ( n27779 , n19418 , n27529 );
and ( n27780 , n19426 , n27527 );
nor ( n27781 , n27779 , n27780 );
xnor ( n27782 , n27781 , n27034 );
and ( n27783 , n27777 , n27782 );
and ( n27784 , n27761 , n27782 );
or ( n27785 , n27778 , n27783 , n27784 );
and ( n27786 , n27745 , n27785 );
and ( n27787 , n27728 , n27785 );
or ( n27788 , n27746 , n27786 , n27787 );
and ( n27789 , n19510 , n26349 );
and ( n27790 , n19496 , n26347 );
nor ( n27791 , n27789 , n27790 );
xnor ( n27792 , n27791 , n25893 );
and ( n27793 , n19605 , n26027 );
and ( n27794 , n19588 , n26025 );
nor ( n27795 , n27793 , n27794 );
xnor ( n27796 , n27795 , n25499 );
and ( n27797 , n27792 , n27796 );
and ( n27798 , n19721 , n25383 );
and ( n27799 , n19637 , n25381 );
nor ( n27800 , n27798 , n27799 );
xnor ( n27801 , n27800 , n24885 );
and ( n27802 , n27796 , n27801 );
and ( n27803 , n27792 , n27801 );
or ( n27804 , n27797 , n27802 , n27803 );
xor ( n27805 , n27426 , n27430 );
xor ( n27806 , n27805 , n27435 );
and ( n27807 , n27804 , n27806 );
xor ( n27808 , n27483 , n27487 );
xor ( n27809 , n27808 , n27489 );
and ( n27810 , n27806 , n27809 );
and ( n27811 , n27804 , n27809 );
or ( n27812 , n27807 , n27810 , n27811 );
and ( n27813 , n27788 , n27812 );
xor ( n27814 , n27442 , n27446 );
xor ( n27815 , n27814 , n27451 );
xor ( n27816 , n27584 , n27588 );
xor ( n27817 , n27816 , n27593 );
and ( n27818 , n27815 , n27817 );
xor ( n27819 , n27458 , n27462 );
xor ( n27820 , n27819 , n27467 );
and ( n27821 , n27817 , n27820 );
and ( n27822 , n27815 , n27820 );
or ( n27823 , n27818 , n27821 , n27822 );
xor ( n27824 , n27562 , n27566 );
xor ( n27825 , n27824 , n27571 );
and ( n27826 , n27823 , n27825 );
xor ( n27827 , n27596 , n27600 );
xor ( n27828 , n27827 , n27605 );
and ( n27829 , n27825 , n27828 );
and ( n27830 , n27823 , n27828 );
or ( n27831 , n27826 , n27829 , n27830 );
and ( n27832 , n27812 , n27831 );
and ( n27833 , n27788 , n27831 );
or ( n27834 , n27813 , n27832 , n27833 );
and ( n27835 , n21955 , n21155 );
and ( n27836 , n21876 , n21153 );
nor ( n27837 , n27835 , n27836 );
xnor ( n27838 , n27837 , n20994 );
and ( n27839 , n27352 , n19424 );
and ( n27840 , n27135 , n19422 );
nor ( n27841 , n27839 , n27840 );
xnor ( n27842 , n27841 , n19431 );
and ( n27843 , n27838 , n27842 );
and ( n27844 , n27751 , n19419 );
and ( n27845 , n27842 , n27844 );
and ( n27846 , n27838 , n27844 );
or ( n27847 , n27843 , n27845 , n27846 );
and ( n27848 , n20080 , n23944 );
and ( n27849 , n20004 , n23942 );
nor ( n27850 , n27848 , n27849 );
xnor ( n27851 , n27850 , n23550 );
and ( n27852 , n20268 , n23641 );
and ( n27853 , n20182 , n23639 );
nor ( n27854 , n27852 , n27853 );
xnor ( n27855 , n27854 , n23213 );
and ( n27856 , n27851 , n27855 );
and ( n27857 , n21704 , n21468 );
and ( n27858 , n21612 , n21466 );
nor ( n27859 , n27857 , n27858 );
xnor ( n27860 , n27859 , n21331 );
and ( n27861 , n27855 , n27860 );
and ( n27862 , n27851 , n27860 );
or ( n27863 , n27856 , n27861 , n27862 );
and ( n27864 , n27847 , n27863 );
xor ( n27865 , n27237 , n27241 );
xor ( n27866 , n27865 , n27246 );
and ( n27867 , n27863 , n27866 );
and ( n27868 , n27847 , n27866 );
or ( n27869 , n27864 , n27867 , n27868 );
xor ( n27870 , n27438 , n27478 );
xor ( n27871 , n27870 , n27492 );
and ( n27872 , n27869 , n27871 );
xor ( n27873 , n27356 , n27358 );
xor ( n27874 , n27873 , n27361 );
and ( n27875 , n27871 , n27874 );
and ( n27876 , n27869 , n27874 );
or ( n27877 , n27872 , n27875 , n27876 );
and ( n27878 , n27834 , n27877 );
xor ( n27879 , n27495 , n27519 );
xor ( n27880 , n27879 , n27522 );
and ( n27881 , n27877 , n27880 );
and ( n27882 , n27834 , n27880 );
or ( n27883 , n27878 , n27881 , n27882 );
and ( n27884 , n27712 , n27883 );
xor ( n27885 , n27414 , n27416 );
xor ( n27886 , n27885 , n27419 );
and ( n27887 , n27883 , n27886 );
and ( n27888 , n27712 , n27886 );
or ( n27889 , n27884 , n27887 , n27888 );
and ( n27890 , n23271 , n20460 );
and ( n27891 , n23141 , n20458 );
nor ( n27892 , n27890 , n27891 );
xnor ( n27893 , n27892 , n20337 );
and ( n27894 , n23573 , n20276 );
and ( n27895 , n23381 , n20274 );
nor ( n27896 , n27894 , n27895 );
xnor ( n27897 , n27896 , n20175 );
and ( n27898 , n27893 , n27897 );
and ( n27899 , n24131 , n20114 );
and ( n27900 , n23968 , n20112 );
nor ( n27901 , n27899 , n27900 );
xnor ( n27902 , n27901 , n19997 );
and ( n27903 , n27897 , n27902 );
and ( n27904 , n27893 , n27902 );
or ( n27905 , n27898 , n27903 , n27904 );
and ( n27906 , n22425 , n20955 );
and ( n27907 , n22198 , n20953 );
nor ( n27908 , n27906 , n27907 );
xnor ( n27909 , n27908 , n20780 );
and ( n27910 , n24527 , n19894 );
and ( n27911 , n24521 , n19892 );
nor ( n27912 , n27910 , n27911 );
xnor ( n27913 , n27912 , n19858 );
and ( n27914 , n27909 , n27913 );
and ( n27915 , n25554 , n19688 );
and ( n27916 , n25284 , n19686 );
nor ( n27917 , n27915 , n27916 );
xnor ( n27918 , n27917 , n19655 );
and ( n27919 , n27913 , n27918 );
and ( n27920 , n27909 , n27918 );
or ( n27921 , n27914 , n27919 , n27920 );
and ( n27922 , n27905 , n27921 );
and ( n27923 , n19946 , n24376 );
and ( n27924 , n19881 , n24374 );
nor ( n27925 , n27923 , n27924 );
xnor ( n27926 , n27925 , n23927 );
and ( n27927 , n27921 , n27926 );
and ( n27928 , n27905 , n27926 );
or ( n27929 , n27922 , n27927 , n27928 );
xor ( n27930 , n27499 , n27503 );
xor ( n27931 , n27930 , n27508 );
and ( n27932 , n27929 , n27931 );
xor ( n27933 , n27454 , n27470 );
xor ( n27934 , n27933 , n27475 );
and ( n27935 , n27931 , n27934 );
and ( n27936 , n27929 , n27934 );
or ( n27937 , n27932 , n27935 , n27936 );
xor ( n27938 , n27544 , n27574 );
xor ( n27939 , n27938 , n27577 );
and ( n27940 , n27937 , n27939 );
xor ( n27941 , n27608 , n27610 );
xor ( n27942 , n27941 , n27613 );
and ( n27943 , n27939 , n27942 );
and ( n27944 , n27937 , n27942 );
or ( n27945 , n27940 , n27943 , n27944 );
xor ( n27946 , n27580 , n27616 );
xor ( n27947 , n27946 , n27619 );
and ( n27948 , n27945 , n27947 );
xor ( n27949 , n27644 , n27646 );
xor ( n27950 , n27949 , n27649 );
and ( n27951 , n27947 , n27950 );
and ( n27952 , n27945 , n27950 );
or ( n27953 , n27948 , n27951 , n27952 );
xor ( n27954 , n27652 , n27654 );
xor ( n27955 , n27954 , n27657 );
and ( n27956 , n27953 , n27955 );
xor ( n27957 , n27525 , n27622 );
xor ( n27958 , n27957 , n27625 );
and ( n27959 , n27955 , n27958 );
and ( n27960 , n27953 , n27958 );
or ( n27961 , n27956 , n27959 , n27960 );
and ( n27962 , n27889 , n27961 );
xor ( n27963 , n27422 , n27628 );
xor ( n27964 , n27963 , n27631 );
and ( n27965 , n27961 , n27964 );
and ( n27966 , n27889 , n27964 );
or ( n27967 , n27962 , n27965 , n27966 );
xor ( n27968 , n27386 , n27388 );
xor ( n27969 , n27968 , n27391 );
and ( n27970 , n27967 , n27969 );
xor ( n27971 , n27634 , n27668 );
xor ( n27972 , n27971 , n27671 );
and ( n27973 , n27969 , n27972 );
and ( n27974 , n27967 , n27972 );
or ( n27975 , n27970 , n27973 , n27974 );
and ( n27976 , n27686 , n27975 );
xor ( n27977 , n27686 , n27975 );
xor ( n27978 , n27967 , n27969 );
xor ( n27979 , n27978 , n27972 );
and ( n27980 , n19469 , n26992 );
and ( n27981 , n19434 , n26990 );
nor ( n27982 , n27980 , n27981 );
xnor ( n27983 , n27982 , n26369 );
and ( n27984 , n19825 , n24902 );
and ( n27985 , n19811 , n24900 );
nor ( n27986 , n27984 , n27985 );
xnor ( n27987 , n27986 , n24397 );
and ( n27988 , n27983 , n27987 );
xor ( n27989 , n27550 , n27554 );
xor ( n27990 , n27989 , n27559 );
and ( n27991 , n27987 , n27990 );
and ( n27992 , n27983 , n27990 );
or ( n27993 , n27988 , n27991 , n27992 );
xor ( n27994 , n27532 , n27536 );
xor ( n27995 , n27994 , n27541 );
and ( n27996 , n27993 , n27995 );
xor ( n27997 , n27688 , n27690 );
xor ( n27998 , n27997 , n27693 );
and ( n27999 , n27995 , n27998 );
and ( n28000 , n27993 , n27998 );
or ( n28001 , n27996 , n27999 , n28000 );
xor ( n28002 , n27636 , n27638 );
xor ( n28003 , n28002 , n27641 );
and ( n28004 , n28001 , n28003 );
xor ( n28005 , n27696 , n27698 );
xor ( n28006 , n28005 , n27701 );
and ( n28007 , n28003 , n28006 );
and ( n28008 , n28001 , n28006 );
or ( n28009 , n28004 , n28007 , n28008 );
and ( n28010 , n20803 , n22859 );
and ( n28011 , n20666 , n22857 );
nor ( n28012 , n28010 , n28011 );
xnor ( n28013 , n28012 , n22418 );
and ( n28014 , n21072 , n22381 );
and ( n28015 , n20867 , n22379 );
nor ( n28016 , n28014 , n28015 );
xnor ( n28017 , n28016 , n22228 );
and ( n28018 , n28013 , n28017 );
and ( n28019 , n21302 , n22048 );
and ( n28020 , n21218 , n22046 );
nor ( n28021 , n28019 , n28020 );
xnor ( n28022 , n28021 , n21853 );
and ( n28023 , n28017 , n28022 );
and ( n28024 , n28013 , n28022 );
or ( n28025 , n28018 , n28023 , n28024 );
and ( n28026 , n20182 , n23944 );
and ( n28027 , n20080 , n23942 );
nor ( n28028 , n28026 , n28027 );
xnor ( n28029 , n28028 , n23550 );
and ( n28030 , n21876 , n21468 );
and ( n28031 , n21704 , n21466 );
nor ( n28032 , n28030 , n28031 );
xnor ( n28033 , n28032 , n21331 );
and ( n28034 , n28029 , n28033 );
and ( n28035 , n22235 , n21155 );
and ( n28036 , n21955 , n21153 );
nor ( n28037 , n28035 , n28036 );
xnor ( n28038 , n28037 , n20994 );
and ( n28039 , n28033 , n28038 );
and ( n28040 , n28029 , n28038 );
or ( n28041 , n28034 , n28039 , n28040 );
and ( n28042 , n28025 , n28041 );
and ( n28043 , n20360 , n23641 );
and ( n28044 , n20268 , n23639 );
nor ( n28045 , n28043 , n28044 );
xnor ( n28046 , n28045 , n23213 );
and ( n28047 , n20618 , n23230 );
and ( n28048 , n20452 , n23228 );
nor ( n28049 , n28047 , n28048 );
xnor ( n28050 , n28049 , n22842 );
and ( n28051 , n28046 , n28050 );
not ( n28052 , n27732 );
and ( n28053 , n28050 , n28052 );
and ( n28054 , n28046 , n28052 );
or ( n28055 , n28051 , n28053 , n28054 );
and ( n28056 , n28041 , n28055 );
and ( n28057 , n28025 , n28055 );
or ( n28058 , n28042 , n28056 , n28057 );
xor ( n28059 , n27031 , n27545 );
xor ( n28060 , n27545 , n27546 );
not ( n28061 , n28060 );
and ( n28062 , n28059 , n28061 );
and ( n28063 , n19426 , n28062 );
not ( n28064 , n28063 );
xnor ( n28065 , n28064 , n27549 );
and ( n28066 , n19637 , n26027 );
and ( n28067 , n19605 , n26025 );
nor ( n28068 , n28066 , n28067 );
xnor ( n28069 , n28068 , n25499 );
and ( n28070 , n28065 , n28069 );
and ( n28071 , n19811 , n25383 );
and ( n28072 , n19721 , n25381 );
nor ( n28073 , n28071 , n28072 );
xnor ( n28074 , n28073 , n24885 );
and ( n28075 , n28069 , n28074 );
and ( n28076 , n28065 , n28074 );
or ( n28077 , n28070 , n28075 , n28076 );
xor ( n28078 , n27716 , n27720 );
xor ( n28079 , n28078 , n27725 );
and ( n28080 , n28077 , n28079 );
xor ( n28081 , n27733 , n27737 );
xor ( n28082 , n28081 , n27742 );
and ( n28083 , n28079 , n28082 );
and ( n28084 , n28077 , n28082 );
or ( n28085 , n28080 , n28083 , n28084 );
and ( n28086 , n28058 , n28085 );
xor ( n28087 , n27847 , n27863 );
xor ( n28088 , n28087 , n27866 );
and ( n28089 , n28085 , n28088 );
and ( n28090 , n28058 , n28088 );
or ( n28091 , n28086 , n28089 , n28090 );
buf ( n28092 , n19406 );
buf ( n28093 , n19407 );
and ( n28094 , n28092 , n28093 );
not ( n28095 , n28094 );
and ( n28096 , n27546 , n28095 );
not ( n28097 , n28096 );
and ( n28098 , n22198 , n21155 );
and ( n28099 , n22235 , n21153 );
nor ( n28100 , n28098 , n28099 );
xnor ( n28101 , n28100 , n20994 );
and ( n28102 , n28097 , n28101 );
and ( n28103 , n22756 , n20955 );
and ( n28104 , n22425 , n20953 );
nor ( n28105 , n28103 , n28104 );
xnor ( n28106 , n28105 , n20780 );
and ( n28107 , n28101 , n28106 );
and ( n28108 , n28097 , n28106 );
or ( n28109 , n28102 , n28107 , n28108 );
and ( n28110 , n20004 , n24376 );
and ( n28111 , n19946 , n24374 );
nor ( n28112 , n28110 , n28111 );
xnor ( n28113 , n28112 , n23927 );
and ( n28114 , n28109 , n28113 );
and ( n28115 , n21612 , n21741 );
and ( n28116 , n21451 , n21739 );
nor ( n28117 , n28115 , n28116 );
xnor ( n28118 , n28117 , n21605 );
and ( n28119 , n28113 , n28118 );
and ( n28120 , n28109 , n28118 );
or ( n28121 , n28114 , n28119 , n28120 );
and ( n28122 , n19496 , n26992 );
and ( n28123 , n19469 , n26990 );
nor ( n28124 , n28122 , n28123 );
xnor ( n28125 , n28124 , n26369 );
and ( n28126 , n19881 , n24902 );
and ( n28127 , n19825 , n24900 );
nor ( n28128 , n28126 , n28127 );
xnor ( n28129 , n28128 , n24397 );
and ( n28130 , n28125 , n28129 );
xor ( n28131 , n27750 , n27755 );
xor ( n28132 , n28131 , n27758 );
and ( n28133 , n28129 , n28132 );
and ( n28134 , n28125 , n28132 );
or ( n28135 , n28130 , n28133 , n28134 );
and ( n28136 , n28121 , n28135 );
xor ( n28137 , n27851 , n27855 );
xor ( n28138 , n28137 , n27860 );
and ( n28139 , n28135 , n28138 );
and ( n28140 , n28121 , n28138 );
or ( n28141 , n28136 , n28139 , n28140 );
xor ( n28142 , n27804 , n27806 );
xor ( n28143 , n28142 , n27809 );
and ( n28144 , n28141 , n28143 );
xor ( n28145 , n27929 , n27931 );
xor ( n28146 , n28145 , n27934 );
and ( n28147 , n28143 , n28146 );
and ( n28148 , n28141 , n28146 );
or ( n28149 , n28144 , n28147 , n28148 );
and ( n28150 , n28091 , n28149 );
xor ( n28151 , n27869 , n27871 );
xor ( n28152 , n28151 , n27874 );
and ( n28153 , n28149 , n28152 );
and ( n28154 , n28091 , n28152 );
or ( n28155 , n28150 , n28153 , n28154 );
and ( n28156 , n28009 , n28155 );
xor ( n28157 , n27704 , n27706 );
xor ( n28158 , n28157 , n27709 );
and ( n28159 , n28155 , n28158 );
and ( n28160 , n28009 , n28158 );
or ( n28161 , n28156 , n28159 , n28160 );
and ( n28162 , n23141 , n20674 );
and ( n28163 , n22916 , n20672 );
nor ( n28164 , n28162 , n28163 );
xnor ( n28165 , n28164 , n20542 );
and ( n28166 , n23381 , n20460 );
and ( n28167 , n23271 , n20458 );
nor ( n28168 , n28166 , n28167 );
xnor ( n28169 , n28168 , n20337 );
and ( n28170 , n28165 , n28169 );
and ( n28171 , n23968 , n20276 );
and ( n28172 , n23573 , n20274 );
nor ( n28173 , n28171 , n28172 );
xnor ( n28174 , n28173 , n20175 );
and ( n28175 , n28169 , n28174 );
and ( n28176 , n28165 , n28174 );
or ( n28177 , n28170 , n28175 , n28176 );
and ( n28178 , n24521 , n20114 );
and ( n28179 , n24131 , n20112 );
nor ( n28180 , n28178 , n28179 );
xnor ( n28181 , n28180 , n19997 );
and ( n28182 , n24621 , n19894 );
and ( n28183 , n24527 , n19892 );
nor ( n28184 , n28182 , n28183 );
xnor ( n28185 , n28184 , n19858 );
and ( n28186 , n28181 , n28185 );
and ( n28187 , n25284 , n19805 );
and ( n28188 , n24940 , n19803 );
nor ( n28189 , n28187 , n28188 );
xnor ( n28190 , n28189 , n19750 );
and ( n28191 , n28185 , n28190 );
and ( n28192 , n28181 , n28190 );
or ( n28193 , n28186 , n28191 , n28192 );
and ( n28194 , n28177 , n28193 );
and ( n28195 , n19434 , n27529 );
and ( n28196 , n19418 , n27527 );
nor ( n28197 , n28195 , n28196 );
xnor ( n28198 , n28197 , n27034 );
and ( n28199 , n28193 , n28198 );
and ( n28200 , n28177 , n28198 );
or ( n28201 , n28194 , n28199 , n28200 );
and ( n28202 , n27352 , n19459 );
and ( n28203 , n27135 , n19457 );
nor ( n28204 , n28202 , n28203 );
xnor ( n28205 , n28204 , n19416 );
and ( n28206 , n27757 , n19424 );
and ( n28207 , n27751 , n19422 );
nor ( n28208 , n28206 , n28207 );
xnor ( n28209 , n28208 , n19431 );
and ( n28210 , n28205 , n28209 );
buf ( n28211 , n19341 );
and ( n28212 , n28211 , n19419 );
and ( n28213 , n28209 , n28212 );
and ( n28214 , n28205 , n28212 );
or ( n28215 , n28210 , n28213 , n28214 );
and ( n28216 , n25765 , n19688 );
and ( n28217 , n25554 , n19686 );
nor ( n28218 , n28216 , n28217 );
xnor ( n28219 , n28218 , n19655 );
and ( n28220 , n26319 , n19596 );
and ( n28221 , n25974 , n19594 );
nor ( n28222 , n28220 , n28221 );
xnor ( n28223 , n28222 , n19545 );
and ( n28224 , n28219 , n28223 );
and ( n28225 , n26851 , n19518 );
and ( n28226 , n26422 , n19516 );
nor ( n28227 , n28225 , n28226 );
xnor ( n28228 , n28227 , n19489 );
and ( n28229 , n28223 , n28228 );
and ( n28230 , n28219 , n28228 );
or ( n28231 , n28224 , n28229 , n28230 );
and ( n28232 , n28215 , n28231 );
and ( n28233 , n19588 , n26349 );
and ( n28234 , n19510 , n26347 );
nor ( n28235 , n28233 , n28234 );
xnor ( n28236 , n28235 , n25893 );
and ( n28237 , n28231 , n28236 );
and ( n28238 , n28215 , n28236 );
or ( n28239 , n28232 , n28237 , n28238 );
and ( n28240 , n28201 , n28239 );
xor ( n28241 , n27838 , n27842 );
xor ( n28242 , n28241 , n27844 );
and ( n28243 , n28239 , n28242 );
and ( n28244 , n28201 , n28242 );
or ( n28245 , n28240 , n28243 , n28244 );
xor ( n28246 , n27893 , n27897 );
xor ( n28247 , n28246 , n27902 );
xor ( n28248 , n27909 , n27913 );
xor ( n28249 , n28248 , n27918 );
and ( n28250 , n28247 , n28249 );
xor ( n28251 , n27765 , n27769 );
xor ( n28252 , n28251 , n27774 );
and ( n28253 , n28249 , n28252 );
and ( n28254 , n28247 , n28252 );
or ( n28255 , n28250 , n28253 , n28254 );
xor ( n28256 , n27905 , n27921 );
xor ( n28257 , n28256 , n27926 );
and ( n28258 , n28255 , n28257 );
xor ( n28259 , n27761 , n27777 );
xor ( n28260 , n28259 , n27782 );
and ( n28261 , n28257 , n28260 );
and ( n28262 , n28255 , n28260 );
or ( n28263 , n28258 , n28261 , n28262 );
and ( n28264 , n28245 , n28263 );
xor ( n28265 , n27728 , n27745 );
xor ( n28266 , n28265 , n27785 );
and ( n28267 , n28263 , n28266 );
and ( n28268 , n28245 , n28266 );
or ( n28269 , n28264 , n28267 , n28268 );
xor ( n28270 , n27788 , n27812 );
xor ( n28271 , n28270 , n27831 );
and ( n28272 , n28269 , n28271 );
xor ( n28273 , n27937 , n27939 );
xor ( n28274 , n28273 , n27942 );
and ( n28275 , n28271 , n28274 );
and ( n28276 , n28269 , n28274 );
or ( n28277 , n28272 , n28275 , n28276 );
xor ( n28278 , n27834 , n27877 );
xor ( n28279 , n28278 , n27880 );
and ( n28280 , n28277 , n28279 );
xor ( n28281 , n27945 , n27947 );
xor ( n28282 , n28281 , n27950 );
and ( n28283 , n28279 , n28282 );
and ( n28284 , n28277 , n28282 );
or ( n28285 , n28280 , n28283 , n28284 );
and ( n28286 , n28161 , n28285 );
xor ( n28287 , n27712 , n27883 );
xor ( n28288 , n28287 , n27886 );
and ( n28289 , n28285 , n28288 );
and ( n28290 , n28161 , n28288 );
or ( n28291 , n28286 , n28289 , n28290 );
xor ( n28292 , n27660 , n27662 );
xor ( n28293 , n28292 , n27665 );
and ( n28294 , n28291 , n28293 );
xor ( n28295 , n27889 , n27961 );
xor ( n28296 , n28295 , n27964 );
and ( n28297 , n28293 , n28296 );
and ( n28298 , n28291 , n28296 );
or ( n28299 , n28294 , n28297 , n28298 );
and ( n28300 , n27979 , n28299 );
xor ( n28301 , n27979 , n28299 );
xor ( n28302 , n28291 , n28293 );
xor ( n28303 , n28302 , n28296 );
and ( n28304 , n20666 , n23230 );
and ( n28305 , n20618 , n23228 );
nor ( n28306 , n28304 , n28305 );
xnor ( n28307 , n28306 , n22842 );
and ( n28308 , n20867 , n22859 );
and ( n28309 , n20803 , n22857 );
nor ( n28310 , n28308 , n28309 );
xnor ( n28311 , n28310 , n22418 );
and ( n28312 , n28307 , n28311 );
and ( n28313 , n21218 , n22381 );
and ( n28314 , n21072 , n22379 );
nor ( n28315 , n28313 , n28314 );
xnor ( n28316 , n28315 , n22228 );
and ( n28317 , n28311 , n28316 );
and ( n28318 , n28307 , n28316 );
or ( n28319 , n28312 , n28317 , n28318 );
and ( n28320 , n20268 , n23944 );
and ( n28321 , n20182 , n23942 );
nor ( n28322 , n28320 , n28321 );
xnor ( n28323 , n28322 , n23550 );
and ( n28324 , n20452 , n23641 );
and ( n28325 , n20360 , n23639 );
nor ( n28326 , n28324 , n28325 );
xnor ( n28327 , n28326 , n23213 );
and ( n28328 , n28323 , n28327 );
and ( n28329 , n21704 , n21741 );
and ( n28330 , n21612 , n21739 );
nor ( n28331 , n28329 , n28330 );
xnor ( n28332 , n28331 , n21605 );
and ( n28333 , n28327 , n28332 );
and ( n28334 , n28323 , n28332 );
or ( n28335 , n28328 , n28333 , n28334 );
and ( n28336 , n28319 , n28335 );
and ( n28337 , n22425 , n21155 );
and ( n28338 , n22198 , n21153 );
nor ( n28339 , n28337 , n28338 );
xnor ( n28340 , n28339 , n20994 );
buf ( n28341 , n28340 );
and ( n28342 , n20080 , n24376 );
and ( n28343 , n20004 , n24374 );
nor ( n28344 , n28342 , n28343 );
xnor ( n28345 , n28344 , n23927 );
and ( n28346 , n28341 , n28345 );
and ( n28347 , n21955 , n21468 );
and ( n28348 , n21876 , n21466 );
nor ( n28349 , n28347 , n28348 );
xnor ( n28350 , n28349 , n21331 );
and ( n28351 , n28345 , n28350 );
and ( n28352 , n28341 , n28350 );
or ( n28353 , n28346 , n28351 , n28352 );
and ( n28354 , n28335 , n28353 );
and ( n28355 , n28319 , n28353 );
or ( n28356 , n28336 , n28354 , n28355 );
and ( n28357 , n19469 , n27529 );
and ( n28358 , n19434 , n27527 );
nor ( n28359 , n28357 , n28358 );
xnor ( n28360 , n28359 , n27034 );
and ( n28361 , n19721 , n26027 );
and ( n28362 , n19637 , n26025 );
nor ( n28363 , n28361 , n28362 );
xnor ( n28364 , n28363 , n25499 );
and ( n28365 , n28360 , n28364 );
and ( n28366 , n19825 , n25383 );
and ( n28367 , n19811 , n25381 );
nor ( n28368 , n28366 , n28367 );
xnor ( n28369 , n28368 , n24885 );
and ( n28370 , n28364 , n28369 );
and ( n28371 , n28360 , n28369 );
or ( n28372 , n28365 , n28370 , n28371 );
and ( n28373 , n24131 , n20276 );
and ( n28374 , n23968 , n20274 );
nor ( n28375 , n28373 , n28374 );
xnor ( n28376 , n28375 , n20175 );
and ( n28377 , n24527 , n20114 );
and ( n28378 , n24521 , n20112 );
nor ( n28379 , n28377 , n28378 );
xnor ( n28380 , n28379 , n19997 );
and ( n28381 , n28376 , n28380 );
and ( n28382 , n24940 , n19894 );
and ( n28383 , n24621 , n19892 );
nor ( n28384 , n28382 , n28383 );
xnor ( n28385 , n28384 , n19858 );
and ( n28386 , n28380 , n28385 );
and ( n28387 , n28376 , n28385 );
or ( n28388 , n28381 , n28386 , n28387 );
and ( n28389 , n25554 , n19805 );
and ( n28390 , n25284 , n19803 );
nor ( n28391 , n28389 , n28390 );
xnor ( n28392 , n28391 , n19750 );
and ( n28393 , n25974 , n19688 );
and ( n28394 , n25765 , n19686 );
nor ( n28395 , n28393 , n28394 );
xnor ( n28396 , n28395 , n19655 );
and ( n28397 , n28392 , n28396 );
and ( n28398 , n26422 , n19596 );
and ( n28399 , n26319 , n19594 );
nor ( n28400 , n28398 , n28399 );
xnor ( n28401 , n28400 , n19545 );
and ( n28402 , n28396 , n28401 );
and ( n28403 , n28392 , n28401 );
or ( n28404 , n28397 , n28402 , n28403 );
and ( n28405 , n28388 , n28404 );
and ( n28406 , n19418 , n28062 );
and ( n28407 , n19426 , n28060 );
nor ( n28408 , n28406 , n28407 );
xnor ( n28409 , n28408 , n27549 );
and ( n28410 , n28404 , n28409 );
and ( n28411 , n28388 , n28409 );
or ( n28412 , n28405 , n28410 , n28411 );
and ( n28413 , n28372 , n28412 );
and ( n28414 , n22916 , n20955 );
and ( n28415 , n22756 , n20953 );
nor ( n28416 , n28414 , n28415 );
xnor ( n28417 , n28416 , n20780 );
and ( n28418 , n23271 , n20674 );
and ( n28419 , n23141 , n20672 );
nor ( n28420 , n28418 , n28419 );
xnor ( n28421 , n28420 , n20542 );
and ( n28422 , n28417 , n28421 );
and ( n28423 , n23573 , n20460 );
and ( n28424 , n23381 , n20458 );
nor ( n28425 , n28423 , n28424 );
xnor ( n28426 , n28425 , n20337 );
and ( n28427 , n28421 , n28426 );
and ( n28428 , n28417 , n28426 );
or ( n28429 , n28422 , n28427 , n28428 );
and ( n28430 , n19946 , n24902 );
and ( n28431 , n19881 , n24900 );
nor ( n28432 , n28430 , n28431 );
xnor ( n28433 , n28432 , n24397 );
and ( n28434 , n28429 , n28433 );
and ( n28435 , n21451 , n22048 );
and ( n28436 , n21302 , n22046 );
nor ( n28437 , n28435 , n28436 );
xnor ( n28438 , n28437 , n21853 );
and ( n28439 , n28433 , n28438 );
and ( n28440 , n28429 , n28438 );
or ( n28441 , n28434 , n28439 , n28440 );
and ( n28442 , n28412 , n28441 );
and ( n28443 , n28372 , n28441 );
or ( n28444 , n28413 , n28442 , n28443 );
and ( n28445 , n28356 , n28444 );
xor ( n28446 , n28025 , n28041 );
xor ( n28447 , n28446 , n28055 );
and ( n28448 , n28444 , n28447 );
and ( n28449 , n28356 , n28447 );
or ( n28450 , n28445 , n28448 , n28449 );
and ( n28451 , n27135 , n19518 );
and ( n28452 , n26851 , n19516 );
nor ( n28453 , n28451 , n28452 );
xnor ( n28454 , n28453 , n19489 );
and ( n28455 , n27751 , n19459 );
and ( n28456 , n27352 , n19457 );
nor ( n28457 , n28455 , n28456 );
xnor ( n28458 , n28457 , n19416 );
and ( n28459 , n28454 , n28458 );
and ( n28460 , n28211 , n19424 );
and ( n28461 , n27757 , n19422 );
nor ( n28462 , n28460 , n28461 );
xnor ( n28463 , n28462 , n19431 );
and ( n28464 , n28458 , n28463 );
and ( n28465 , n28454 , n28463 );
or ( n28466 , n28459 , n28464 , n28465 );
and ( n28467 , n19510 , n26992 );
and ( n28468 , n19496 , n26990 );
nor ( n28469 , n28467 , n28468 );
xnor ( n28470 , n28469 , n26369 );
and ( n28471 , n28466 , n28470 );
and ( n28472 , n19605 , n26349 );
and ( n28473 , n19588 , n26347 );
nor ( n28474 , n28472 , n28473 );
xnor ( n28475 , n28474 , n25893 );
and ( n28476 , n28470 , n28475 );
and ( n28477 , n28466 , n28475 );
or ( n28478 , n28471 , n28476 , n28477 );
xor ( n28479 , n28013 , n28017 );
xor ( n28480 , n28479 , n28022 );
and ( n28481 , n28478 , n28480 );
xor ( n28482 , n28029 , n28033 );
xor ( n28483 , n28482 , n28038 );
and ( n28484 , n28480 , n28483 );
and ( n28485 , n28478 , n28483 );
or ( n28486 , n28481 , n28484 , n28485 );
xor ( n28487 , n28097 , n28101 );
xor ( n28488 , n28487 , n28106 );
xor ( n28489 , n28165 , n28169 );
xor ( n28490 , n28489 , n28174 );
and ( n28491 , n28488 , n28490 );
xor ( n28492 , n28205 , n28209 );
xor ( n28493 , n28492 , n28212 );
and ( n28494 , n28490 , n28493 );
and ( n28495 , n28488 , n28493 );
or ( n28496 , n28491 , n28494 , n28495 );
xor ( n28497 , n28065 , n28069 );
xor ( n28498 , n28497 , n28074 );
and ( n28499 , n28496 , n28498 );
xor ( n28500 , n28215 , n28231 );
xor ( n28501 , n28500 , n28236 );
and ( n28502 , n28498 , n28501 );
and ( n28503 , n28496 , n28501 );
or ( n28504 , n28499 , n28502 , n28503 );
and ( n28505 , n28486 , n28504 );
xor ( n28506 , n28121 , n28135 );
xor ( n28507 , n28506 , n28138 );
and ( n28508 , n28504 , n28507 );
and ( n28509 , n28486 , n28507 );
or ( n28510 , n28505 , n28508 , n28509 );
and ( n28511 , n28450 , n28510 );
xor ( n28512 , n28109 , n28113 );
xor ( n28513 , n28512 , n28118 );
xor ( n28514 , n28177 , n28193 );
xor ( n28515 , n28514 , n28198 );
and ( n28516 , n28513 , n28515 );
xor ( n28517 , n28046 , n28050 );
xor ( n28518 , n28517 , n28052 );
and ( n28519 , n28515 , n28518 );
and ( n28520 , n28513 , n28518 );
or ( n28521 , n28516 , n28519 , n28520 );
xor ( n28522 , n28201 , n28239 );
xor ( n28523 , n28522 , n28242 );
and ( n28524 , n28521 , n28523 );
xor ( n28525 , n28077 , n28079 );
xor ( n28526 , n28525 , n28082 );
and ( n28527 , n28523 , n28526 );
and ( n28528 , n28521 , n28526 );
or ( n28529 , n28524 , n28527 , n28528 );
and ( n28530 , n28510 , n28529 );
and ( n28531 , n28450 , n28529 );
or ( n28532 , n28511 , n28530 , n28531 );
xor ( n28533 , n27792 , n27796 );
xor ( n28534 , n28533 , n27801 );
xor ( n28535 , n27983 , n27987 );
xor ( n28536 , n28535 , n27990 );
and ( n28537 , n28534 , n28536 );
xor ( n28538 , n27815 , n27817 );
xor ( n28539 , n28538 , n27820 );
and ( n28540 , n28536 , n28539 );
and ( n28541 , n28534 , n28539 );
or ( n28542 , n28537 , n28540 , n28541 );
xor ( n28543 , n27823 , n27825 );
xor ( n28544 , n28543 , n27828 );
and ( n28545 , n28542 , n28544 );
xor ( n28546 , n27993 , n27995 );
xor ( n28547 , n28546 , n27998 );
and ( n28548 , n28544 , n28547 );
and ( n28549 , n28542 , n28547 );
or ( n28550 , n28545 , n28548 , n28549 );
and ( n28551 , n28532 , n28550 );
xor ( n28552 , n28001 , n28003 );
xor ( n28553 , n28552 , n28006 );
and ( n28554 , n28550 , n28553 );
and ( n28555 , n28532 , n28553 );
or ( n28556 , n28551 , n28554 , n28555 );
xor ( n28557 , n28245 , n28263 );
xor ( n28558 , n28557 , n28266 );
xor ( n28559 , n28058 , n28085 );
xor ( n28560 , n28559 , n28088 );
and ( n28561 , n28558 , n28560 );
xor ( n28562 , n28141 , n28143 );
xor ( n28563 , n28562 , n28146 );
and ( n28564 , n28560 , n28563 );
and ( n28565 , n28558 , n28563 );
or ( n28566 , n28561 , n28564 , n28565 );
xor ( n28567 , n28091 , n28149 );
xor ( n28568 , n28567 , n28152 );
and ( n28569 , n28566 , n28568 );
xor ( n28570 , n28269 , n28271 );
xor ( n28571 , n28570 , n28274 );
and ( n28572 , n28568 , n28571 );
and ( n28573 , n28566 , n28571 );
or ( n28574 , n28569 , n28572 , n28573 );
and ( n28575 , n28556 , n28574 );
xor ( n28576 , n28009 , n28155 );
xor ( n28577 , n28576 , n28158 );
and ( n28578 , n28574 , n28577 );
and ( n28579 , n28556 , n28577 );
or ( n28580 , n28575 , n28578 , n28579 );
xor ( n28581 , n27953 , n27955 );
xor ( n28582 , n28581 , n27958 );
and ( n28583 , n28580 , n28582 );
xor ( n28584 , n28161 , n28285 );
xor ( n28585 , n28584 , n28288 );
and ( n28586 , n28582 , n28585 );
and ( n28587 , n28580 , n28585 );
or ( n28588 , n28583 , n28586 , n28587 );
and ( n28589 , n28303 , n28588 );
xor ( n28590 , n28303 , n28588 );
xor ( n28591 , n28580 , n28582 );
xor ( n28592 , n28591 , n28585 );
and ( n28593 , n20182 , n24376 );
and ( n28594 , n20080 , n24374 );
nor ( n28595 , n28593 , n28594 );
xnor ( n28596 , n28595 , n23927 );
and ( n28597 , n20360 , n23944 );
and ( n28598 , n20268 , n23942 );
nor ( n28599 , n28597 , n28598 );
xnor ( n28600 , n28599 , n23550 );
and ( n28601 , n28596 , n28600 );
and ( n28602 , n20618 , n23641 );
and ( n28603 , n20452 , n23639 );
nor ( n28604 , n28602 , n28603 );
xnor ( n28605 , n28604 , n23213 );
and ( n28606 , n28600 , n28605 );
and ( n28607 , n28596 , n28605 );
or ( n28608 , n28601 , n28606 , n28607 );
and ( n28609 , n26851 , n19596 );
and ( n28610 , n26422 , n19594 );
nor ( n28611 , n28609 , n28610 );
xnor ( n28612 , n28611 , n19545 );
and ( n28613 , n27352 , n19518 );
and ( n28614 , n27135 , n19516 );
nor ( n28615 , n28613 , n28614 );
xnor ( n28616 , n28615 , n19489 );
and ( n28617 , n28612 , n28616 );
and ( n28618 , n27757 , n19459 );
and ( n28619 , n27751 , n19457 );
nor ( n28620 , n28618 , n28619 );
xnor ( n28621 , n28620 , n19416 );
and ( n28622 , n28616 , n28621 );
and ( n28623 , n28612 , n28621 );
or ( n28624 , n28617 , n28622 , n28623 );
xor ( n28625 , n27546 , n28092 );
xor ( n28626 , n28092 , n28093 );
not ( n28627 , n28626 );
and ( n28628 , n28625 , n28627 );
and ( n28629 , n19426 , n28628 );
not ( n28630 , n28629 );
xnor ( n28631 , n28630 , n28096 );
and ( n28632 , n28624 , n28631 );
and ( n28633 , n19637 , n26349 );
and ( n28634 , n19605 , n26347 );
nor ( n28635 , n28633 , n28634 );
xnor ( n28636 , n28635 , n25893 );
and ( n28637 , n28631 , n28636 );
and ( n28638 , n28624 , n28636 );
or ( n28639 , n28632 , n28637 , n28638 );
and ( n28640 , n28608 , n28639 );
and ( n28641 , n20803 , n23230 );
and ( n28642 , n20666 , n23228 );
nor ( n28643 , n28641 , n28642 );
xnor ( n28644 , n28643 , n22842 );
and ( n28645 , n21072 , n22859 );
and ( n28646 , n20867 , n22857 );
nor ( n28647 , n28645 , n28646 );
xnor ( n28648 , n28647 , n22418 );
and ( n28649 , n28644 , n28648 );
not ( n28650 , n28340 );
and ( n28651 , n28648 , n28650 );
and ( n28652 , n28644 , n28650 );
or ( n28653 , n28649 , n28651 , n28652 );
and ( n28654 , n28639 , n28653 );
and ( n28655 , n28608 , n28653 );
or ( n28656 , n28640 , n28654 , n28655 );
and ( n28657 , n20004 , n24902 );
and ( n28658 , n19946 , n24900 );
nor ( n28659 , n28657 , n28658 );
xnor ( n28660 , n28659 , n24397 );
and ( n28661 , n21302 , n22381 );
and ( n28662 , n21218 , n22379 );
nor ( n28663 , n28661 , n28662 );
xnor ( n28664 , n28663 , n22228 );
and ( n28665 , n28660 , n28664 );
and ( n28666 , n21612 , n22048 );
and ( n28667 , n21451 , n22046 );
nor ( n28668 , n28666 , n28667 );
xnor ( n28669 , n28668 , n21853 );
and ( n28670 , n28664 , n28669 );
and ( n28671 , n28660 , n28669 );
or ( n28672 , n28665 , n28670 , n28671 );
buf ( n28673 , n19408 );
buf ( n28674 , n19409 );
and ( n28675 , n28673 , n28674 );
not ( n28676 , n28675 );
and ( n28677 , n28093 , n28676 );
not ( n28678 , n28677 );
and ( n28679 , n22198 , n21468 );
and ( n28680 , n22235 , n21466 );
nor ( n28681 , n28679 , n28680 );
xnor ( n28682 , n28681 , n21331 );
and ( n28683 , n28678 , n28682 );
and ( n28684 , n22756 , n21155 );
and ( n28685 , n22425 , n21153 );
nor ( n28686 , n28684 , n28685 );
xnor ( n28687 , n28686 , n20994 );
and ( n28688 , n28682 , n28687 );
and ( n28689 , n28678 , n28687 );
or ( n28690 , n28683 , n28688 , n28689 );
and ( n28691 , n23141 , n20955 );
and ( n28692 , n22916 , n20953 );
nor ( n28693 , n28691 , n28692 );
xnor ( n28694 , n28693 , n20780 );
and ( n28695 , n23381 , n20674 );
and ( n28696 , n23271 , n20672 );
nor ( n28697 , n28695 , n28696 );
xnor ( n28698 , n28697 , n20542 );
and ( n28699 , n28694 , n28698 );
buf ( n28700 , n19343 );
and ( n28701 , n28700 , n19419 );
and ( n28702 , n28698 , n28701 );
and ( n28703 , n28694 , n28701 );
or ( n28704 , n28699 , n28702 , n28703 );
and ( n28705 , n28690 , n28704 );
and ( n28706 , n19434 , n28062 );
and ( n28707 , n19418 , n28060 );
nor ( n28708 , n28706 , n28707 );
xnor ( n28709 , n28708 , n27549 );
and ( n28710 , n28704 , n28709 );
and ( n28711 , n28690 , n28709 );
or ( n28712 , n28705 , n28710 , n28711 );
and ( n28713 , n28672 , n28712 );
and ( n28714 , n23968 , n20460 );
and ( n28715 , n23573 , n20458 );
nor ( n28716 , n28714 , n28715 );
xnor ( n28717 , n28716 , n20337 );
and ( n28718 , n24521 , n20276 );
and ( n28719 , n24131 , n20274 );
nor ( n28720 , n28718 , n28719 );
xnor ( n28721 , n28720 , n20175 );
and ( n28722 , n28717 , n28721 );
and ( n28723 , n24621 , n20114 );
and ( n28724 , n24527 , n20112 );
nor ( n28725 , n28723 , n28724 );
xnor ( n28726 , n28725 , n19997 );
and ( n28727 , n28721 , n28726 );
and ( n28728 , n28717 , n28726 );
or ( n28729 , n28722 , n28727 , n28728 );
and ( n28730 , n25284 , n19894 );
and ( n28731 , n24940 , n19892 );
nor ( n28732 , n28730 , n28731 );
xnor ( n28733 , n28732 , n19858 );
and ( n28734 , n25765 , n19805 );
and ( n28735 , n25554 , n19803 );
nor ( n28736 , n28734 , n28735 );
xnor ( n28737 , n28736 , n19750 );
and ( n28738 , n28733 , n28737 );
and ( n28739 , n26319 , n19688 );
and ( n28740 , n25974 , n19686 );
nor ( n28741 , n28739 , n28740 );
xnor ( n28742 , n28741 , n19655 );
and ( n28743 , n28737 , n28742 );
and ( n28744 , n28733 , n28742 );
or ( n28745 , n28738 , n28743 , n28744 );
and ( n28746 , n28729 , n28745 );
and ( n28747 , n19588 , n26992 );
and ( n28748 , n19510 , n26990 );
nor ( n28749 , n28747 , n28748 );
xnor ( n28750 , n28749 , n26369 );
and ( n28751 , n28745 , n28750 );
and ( n28752 , n28729 , n28750 );
or ( n28753 , n28746 , n28751 , n28752 );
and ( n28754 , n28712 , n28753 );
and ( n28755 , n28672 , n28753 );
or ( n28756 , n28713 , n28754 , n28755 );
and ( n28757 , n28656 , n28756 );
xor ( n28758 , n28319 , n28335 );
xor ( n28759 , n28758 , n28353 );
and ( n28760 , n28756 , n28759 );
and ( n28761 , n28656 , n28759 );
or ( n28762 , n28757 , n28760 , n28761 );
and ( n28763 , n19496 , n27529 );
and ( n28764 , n19469 , n27527 );
nor ( n28765 , n28763 , n28764 );
xnor ( n28766 , n28765 , n27034 );
and ( n28767 , n19811 , n26027 );
and ( n28768 , n19721 , n26025 );
nor ( n28769 , n28767 , n28768 );
xnor ( n28770 , n28769 , n25499 );
and ( n28771 , n28766 , n28770 );
and ( n28772 , n19881 , n25383 );
and ( n28773 , n19825 , n25381 );
nor ( n28774 , n28772 , n28773 );
xnor ( n28775 , n28774 , n24885 );
and ( n28776 , n28770 , n28775 );
and ( n28777 , n28766 , n28775 );
or ( n28778 , n28771 , n28776 , n28777 );
xor ( n28779 , n28307 , n28311 );
xor ( n28780 , n28779 , n28316 );
and ( n28781 , n28778 , n28780 );
xor ( n28782 , n28341 , n28345 );
xor ( n28783 , n28782 , n28350 );
and ( n28784 , n28780 , n28783 );
and ( n28785 , n28778 , n28783 );
or ( n28786 , n28781 , n28784 , n28785 );
xor ( n28787 , n28372 , n28412 );
xor ( n28788 , n28787 , n28441 );
and ( n28789 , n28786 , n28788 );
xor ( n28790 , n28478 , n28480 );
xor ( n28791 , n28790 , n28483 );
and ( n28792 , n28788 , n28791 );
and ( n28793 , n28786 , n28791 );
or ( n28794 , n28789 , n28792 , n28793 );
and ( n28795 , n28762 , n28794 );
xor ( n28796 , n28356 , n28444 );
xor ( n28797 , n28796 , n28447 );
and ( n28798 , n28794 , n28797 );
and ( n28799 , n28762 , n28797 );
or ( n28800 , n28795 , n28798 , n28799 );
and ( n28801 , n21876 , n21741 );
and ( n28802 , n21704 , n21739 );
nor ( n28803 , n28801 , n28802 );
xnor ( n28804 , n28803 , n21605 );
and ( n28805 , n22235 , n21468 );
and ( n28806 , n21955 , n21466 );
nor ( n28807 , n28805 , n28806 );
xnor ( n28808 , n28807 , n21331 );
and ( n28809 , n28804 , n28808 );
buf ( n28810 , n19342 );
and ( n28811 , n28810 , n19419 );
and ( n28812 , n28808 , n28811 );
and ( n28813 , n28804 , n28811 );
or ( n28814 , n28809 , n28812 , n28813 );
xor ( n28815 , n28219 , n28223 );
xor ( n28816 , n28815 , n28228 );
and ( n28817 , n28814 , n28816 );
xor ( n28818 , n28181 , n28185 );
xor ( n28819 , n28818 , n28190 );
and ( n28820 , n28816 , n28819 );
and ( n28821 , n28814 , n28819 );
or ( n28822 , n28817 , n28820 , n28821 );
xor ( n28823 , n28125 , n28129 );
xor ( n28824 , n28823 , n28132 );
and ( n28825 , n28822 , n28824 );
xor ( n28826 , n28247 , n28249 );
xor ( n28827 , n28826 , n28252 );
and ( n28828 , n28824 , n28827 );
and ( n28829 , n28822 , n28827 );
or ( n28830 , n28825 , n28828 , n28829 );
xor ( n28831 , n28255 , n28257 );
xor ( n28832 , n28831 , n28260 );
and ( n28833 , n28830 , n28832 );
xor ( n28834 , n28534 , n28536 );
xor ( n28835 , n28834 , n28539 );
and ( n28836 , n28832 , n28835 );
and ( n28837 , n28830 , n28835 );
or ( n28838 , n28833 , n28836 , n28837 );
and ( n28839 , n28800 , n28838 );
xor ( n28840 , n28542 , n28544 );
xor ( n28841 , n28840 , n28547 );
and ( n28842 , n28838 , n28841 );
and ( n28843 , n28800 , n28841 );
or ( n28844 , n28839 , n28842 , n28843 );
xor ( n28845 , n28417 , n28421 );
xor ( n28846 , n28845 , n28426 );
xor ( n28847 , n28376 , n28380 );
xor ( n28848 , n28847 , n28385 );
and ( n28849 , n28846 , n28848 );
xor ( n28850 , n28454 , n28458 );
xor ( n28851 , n28850 , n28463 );
and ( n28852 , n28848 , n28851 );
and ( n28853 , n28846 , n28851 );
or ( n28854 , n28849 , n28852 , n28853 );
xor ( n28855 , n28360 , n28364 );
xor ( n28856 , n28855 , n28369 );
and ( n28857 , n28854 , n28856 );
xor ( n28858 , n28323 , n28327 );
xor ( n28859 , n28858 , n28332 );
and ( n28860 , n28856 , n28859 );
and ( n28861 , n28854 , n28859 );
or ( n28862 , n28857 , n28860 , n28861 );
xor ( n28863 , n28466 , n28470 );
xor ( n28864 , n28863 , n28475 );
xor ( n28865 , n28388 , n28404 );
xor ( n28866 , n28865 , n28409 );
and ( n28867 , n28864 , n28866 );
xor ( n28868 , n28429 , n28433 );
xor ( n28869 , n28868 , n28438 );
and ( n28870 , n28866 , n28869 );
and ( n28871 , n28864 , n28869 );
or ( n28872 , n28867 , n28870 , n28871 );
and ( n28873 , n28862 , n28872 );
and ( n28874 , n20080 , n24902 );
and ( n28875 , n20004 , n24900 );
nor ( n28876 , n28874 , n28875 );
xnor ( n28877 , n28876 , n24397 );
and ( n28878 , n20268 , n24376 );
and ( n28879 , n20182 , n24374 );
nor ( n28880 , n28878 , n28879 );
xnor ( n28881 , n28880 , n23927 );
and ( n28882 , n28877 , n28881 );
and ( n28883 , n21704 , n22048 );
and ( n28884 , n21612 , n22046 );
nor ( n28885 , n28883 , n28884 );
xnor ( n28886 , n28885 , n21853 );
and ( n28887 , n28881 , n28886 );
and ( n28888 , n28877 , n28886 );
or ( n28889 , n28882 , n28887 , n28888 );
and ( n28890 , n22425 , n21468 );
and ( n28891 , n22198 , n21466 );
nor ( n28892 , n28890 , n28891 );
xnor ( n28893 , n28892 , n21331 );
buf ( n28894 , n28893 );
and ( n28895 , n21955 , n21741 );
and ( n28896 , n21876 , n21739 );
nor ( n28897 , n28895 , n28896 );
xnor ( n28898 , n28897 , n21605 );
and ( n28899 , n28894 , n28898 );
and ( n28900 , n28810 , n19424 );
and ( n28901 , n28211 , n19422 );
nor ( n28902 , n28900 , n28901 );
xnor ( n28903 , n28902 , n19431 );
and ( n28904 , n28898 , n28903 );
and ( n28905 , n28894 , n28903 );
or ( n28906 , n28899 , n28904 , n28905 );
and ( n28907 , n28889 , n28906 );
xor ( n28908 , n28392 , n28396 );
xor ( n28909 , n28908 , n28401 );
and ( n28910 , n28906 , n28909 );
and ( n28911 , n28889 , n28909 );
or ( n28912 , n28907 , n28910 , n28911 );
xor ( n28913 , n28488 , n28490 );
xor ( n28914 , n28913 , n28493 );
and ( n28915 , n28912 , n28914 );
xor ( n28916 , n28814 , n28816 );
xor ( n28917 , n28916 , n28819 );
and ( n28918 , n28914 , n28917 );
and ( n28919 , n28912 , n28917 );
or ( n28920 , n28915 , n28918 , n28919 );
and ( n28921 , n28872 , n28920 );
and ( n28922 , n28862 , n28920 );
or ( n28923 , n28873 , n28921 , n28922 );
xor ( n28924 , n28486 , n28504 );
xor ( n28925 , n28924 , n28507 );
and ( n28926 , n28923 , n28925 );
xor ( n28927 , n28521 , n28523 );
xor ( n28928 , n28927 , n28526 );
and ( n28929 , n28925 , n28928 );
and ( n28930 , n28923 , n28928 );
or ( n28931 , n28926 , n28929 , n28930 );
xor ( n28932 , n28450 , n28510 );
xor ( n28933 , n28932 , n28529 );
and ( n28934 , n28931 , n28933 );
xor ( n28935 , n28558 , n28560 );
xor ( n28936 , n28935 , n28563 );
and ( n28937 , n28933 , n28936 );
and ( n28938 , n28931 , n28936 );
or ( n28939 , n28934 , n28937 , n28938 );
and ( n28940 , n28844 , n28939 );
xor ( n28941 , n28532 , n28550 );
xor ( n28942 , n28941 , n28553 );
and ( n28943 , n28939 , n28942 );
and ( n28944 , n28844 , n28942 );
or ( n28945 , n28940 , n28943 , n28944 );
xor ( n28946 , n28277 , n28279 );
xor ( n28947 , n28946 , n28282 );
and ( n28948 , n28945 , n28947 );
xor ( n28949 , n28556 , n28574 );
xor ( n28950 , n28949 , n28577 );
and ( n28951 , n28947 , n28950 );
and ( n28952 , n28945 , n28950 );
or ( n28953 , n28948 , n28951 , n28952 );
and ( n28954 , n28592 , n28953 );
xor ( n28955 , n28592 , n28953 );
xor ( n28956 , n28945 , n28947 );
xor ( n28957 , n28956 , n28950 );
xor ( n28958 , n28660 , n28664 );
xor ( n28959 , n28958 , n28669 );
xor ( n28960 , n28596 , n28600 );
xor ( n28961 , n28960 , n28605 );
and ( n28962 , n28959 , n28961 );
xor ( n28963 , n28644 , n28648 );
xor ( n28964 , n28963 , n28650 );
and ( n28965 , n28961 , n28964 );
and ( n28966 , n28959 , n28964 );
or ( n28967 , n28962 , n28965 , n28966 );
and ( n28968 , n20452 , n23944 );
and ( n28969 , n20360 , n23942 );
nor ( n28970 , n28968 , n28969 );
xnor ( n28971 , n28970 , n23550 );
and ( n28972 , n20666 , n23641 );
and ( n28973 , n20618 , n23639 );
nor ( n28974 , n28972 , n28973 );
xnor ( n28975 , n28974 , n23213 );
and ( n28976 , n28971 , n28975 );
and ( n28977 , n20867 , n23230 );
and ( n28978 , n20803 , n23228 );
nor ( n28979 , n28977 , n28978 );
xnor ( n28980 , n28979 , n22842 );
and ( n28981 , n28975 , n28980 );
and ( n28982 , n28971 , n28980 );
or ( n28983 , n28976 , n28981 , n28982 );
and ( n28984 , n26422 , n19688 );
and ( n28985 , n26319 , n19686 );
nor ( n28986 , n28984 , n28985 );
xnor ( n28987 , n28986 , n19655 );
and ( n28988 , n27135 , n19596 );
and ( n28989 , n26851 , n19594 );
nor ( n28990 , n28988 , n28989 );
xnor ( n28991 , n28990 , n19545 );
and ( n28992 , n28987 , n28991 );
and ( n28993 , n27751 , n19518 );
and ( n28994 , n27352 , n19516 );
nor ( n28995 , n28993 , n28994 );
xnor ( n28996 , n28995 , n19489 );
and ( n28997 , n28991 , n28996 );
and ( n28998 , n28987 , n28996 );
or ( n28999 , n28992 , n28997 , n28998 );
and ( n29000 , n24940 , n20114 );
and ( n29001 , n24621 , n20112 );
nor ( n29002 , n29000 , n29001 );
xnor ( n29003 , n29002 , n19997 );
and ( n29004 , n25554 , n19894 );
and ( n29005 , n25284 , n19892 );
nor ( n29006 , n29004 , n29005 );
xnor ( n29007 , n29006 , n19858 );
and ( n29008 , n29003 , n29007 );
and ( n29009 , n25974 , n19805 );
and ( n29010 , n25765 , n19803 );
nor ( n29011 , n29009 , n29010 );
xnor ( n29012 , n29011 , n19750 );
and ( n29013 , n29007 , n29012 );
and ( n29014 , n29003 , n29012 );
or ( n29015 , n29008 , n29013 , n29014 );
and ( n29016 , n28999 , n29015 );
and ( n29017 , n19510 , n27529 );
and ( n29018 , n19496 , n27527 );
nor ( n29019 , n29017 , n29018 );
xnor ( n29020 , n29019 , n27034 );
and ( n29021 , n29015 , n29020 );
and ( n29022 , n28999 , n29020 );
or ( n29023 , n29016 , n29021 , n29022 );
and ( n29024 , n28983 , n29023 );
xor ( n29025 , n28804 , n28808 );
xor ( n29026 , n29025 , n28811 );
and ( n29027 , n29023 , n29026 );
and ( n29028 , n28983 , n29026 );
or ( n29029 , n29024 , n29027 , n29028 );
and ( n29030 , n28967 , n29029 );
xor ( n29031 , n28608 , n28639 );
xor ( n29032 , n29031 , n28653 );
and ( n29033 , n29029 , n29032 );
and ( n29034 , n28967 , n29032 );
or ( n29035 , n29030 , n29033 , n29034 );
and ( n29036 , n19469 , n28062 );
and ( n29037 , n19434 , n28060 );
nor ( n29038 , n29036 , n29037 );
xnor ( n29039 , n29038 , n27549 );
and ( n29040 , n19605 , n26992 );
and ( n29041 , n19588 , n26990 );
nor ( n29042 , n29040 , n29041 );
xnor ( n29043 , n29042 , n26369 );
and ( n29044 , n29039 , n29043 );
and ( n29045 , n19721 , n26349 );
and ( n29046 , n19637 , n26347 );
nor ( n29047 , n29045 , n29046 );
xnor ( n29048 , n29047 , n25893 );
and ( n29049 , n29043 , n29048 );
and ( n29050 , n29039 , n29048 );
or ( n29051 , n29044 , n29049 , n29050 );
and ( n29052 , n19946 , n25383 );
and ( n29053 , n19881 , n25381 );
nor ( n29054 , n29052 , n29053 );
xnor ( n29055 , n29054 , n24885 );
and ( n29056 , n21218 , n22859 );
and ( n29057 , n21072 , n22857 );
nor ( n29058 , n29056 , n29057 );
xnor ( n29059 , n29058 , n22418 );
and ( n29060 , n29055 , n29059 );
and ( n29061 , n21451 , n22381 );
and ( n29062 , n21302 , n22379 );
nor ( n29063 , n29061 , n29062 );
xnor ( n29064 , n29063 , n22228 );
and ( n29065 , n29059 , n29064 );
and ( n29066 , n29055 , n29064 );
or ( n29067 , n29060 , n29065 , n29066 );
and ( n29068 , n29051 , n29067 );
and ( n29069 , n22916 , n21155 );
and ( n29070 , n22756 , n21153 );
nor ( n29071 , n29069 , n29070 );
xnor ( n29072 , n29071 , n20994 );
and ( n29073 , n23271 , n20955 );
and ( n29074 , n23141 , n20953 );
nor ( n29075 , n29073 , n29074 );
xnor ( n29076 , n29075 , n20780 );
and ( n29077 , n29072 , n29076 );
buf ( n29078 , n19344 );
and ( n29079 , n29078 , n19419 );
and ( n29080 , n29076 , n29079 );
and ( n29081 , n29072 , n29079 );
or ( n29082 , n29077 , n29080 , n29081 );
and ( n29083 , n23573 , n20674 );
and ( n29084 , n23381 , n20672 );
nor ( n29085 , n29083 , n29084 );
xnor ( n29086 , n29085 , n20542 );
and ( n29087 , n24131 , n20460 );
and ( n29088 , n23968 , n20458 );
nor ( n29089 , n29087 , n29088 );
xnor ( n29090 , n29089 , n20337 );
and ( n29091 , n29086 , n29090 );
and ( n29092 , n24527 , n20276 );
and ( n29093 , n24521 , n20274 );
nor ( n29094 , n29092 , n29093 );
xnor ( n29095 , n29094 , n20175 );
and ( n29096 , n29090 , n29095 );
and ( n29097 , n29086 , n29095 );
or ( n29098 , n29091 , n29096 , n29097 );
and ( n29099 , n29082 , n29098 );
and ( n29100 , n19418 , n28628 );
and ( n29101 , n19426 , n28626 );
nor ( n29102 , n29100 , n29101 );
xnor ( n29103 , n29102 , n28096 );
and ( n29104 , n29098 , n29103 );
and ( n29105 , n29082 , n29103 );
or ( n29106 , n29099 , n29104 , n29105 );
and ( n29107 , n29067 , n29106 );
and ( n29108 , n29051 , n29106 );
or ( n29109 , n29068 , n29107 , n29108 );
xor ( n29110 , n28766 , n28770 );
xor ( n29111 , n29110 , n28775 );
xor ( n29112 , n28624 , n28631 );
xor ( n29113 , n29112 , n28636 );
and ( n29114 , n29111 , n29113 );
xor ( n29115 , n28729 , n28745 );
xor ( n29116 , n29115 , n28750 );
and ( n29117 , n29113 , n29116 );
and ( n29118 , n29111 , n29116 );
or ( n29119 , n29114 , n29117 , n29118 );
and ( n29120 , n29109 , n29119 );
xor ( n29121 , n28672 , n28712 );
xor ( n29122 , n29121 , n28753 );
and ( n29123 , n29119 , n29122 );
and ( n29124 , n29109 , n29122 );
or ( n29125 , n29120 , n29123 , n29124 );
and ( n29126 , n29035 , n29125 );
xor ( n29127 , n28656 , n28756 );
xor ( n29128 , n29127 , n28759 );
and ( n29129 , n29125 , n29128 );
and ( n29130 , n29035 , n29128 );
or ( n29131 , n29126 , n29129 , n29130 );
xor ( n29132 , n28513 , n28515 );
xor ( n29133 , n29132 , n28518 );
xor ( n29134 , n28496 , n28498 );
xor ( n29135 , n29134 , n28501 );
and ( n29136 , n29133 , n29135 );
xor ( n29137 , n28822 , n28824 );
xor ( n29138 , n29137 , n28827 );
and ( n29139 , n29135 , n29138 );
and ( n29140 , n29133 , n29138 );
or ( n29141 , n29136 , n29139 , n29140 );
and ( n29142 , n29131 , n29141 );
xor ( n29143 , n28830 , n28832 );
xor ( n29144 , n29143 , n28835 );
and ( n29145 , n29141 , n29144 );
and ( n29146 , n29131 , n29144 );
or ( n29147 , n29142 , n29145 , n29146 );
and ( n29148 , n22235 , n21741 );
and ( n29149 , n21955 , n21739 );
nor ( n29150 , n29148 , n29149 );
xnor ( n29151 , n29150 , n21605 );
and ( n29152 , n28211 , n19459 );
and ( n29153 , n27757 , n19457 );
nor ( n29154 , n29152 , n29153 );
xnor ( n29155 , n29154 , n19416 );
and ( n29156 , n29151 , n29155 );
and ( n29157 , n28700 , n19424 );
and ( n29158 , n28810 , n19422 );
nor ( n29159 , n29157 , n29158 );
xnor ( n29160 , n29159 , n19431 );
and ( n29161 , n29155 , n29160 );
and ( n29162 , n29151 , n29160 );
or ( n29163 , n29156 , n29161 , n29162 );
and ( n29164 , n19825 , n26027 );
and ( n29165 , n19811 , n26025 );
nor ( n29166 , n29164 , n29165 );
xnor ( n29167 , n29166 , n25499 );
and ( n29168 , n29163 , n29167 );
xor ( n29169 , n28694 , n28698 );
xor ( n29170 , n29169 , n28701 );
and ( n29171 , n29167 , n29170 );
and ( n29172 , n29163 , n29170 );
or ( n29173 , n29168 , n29171 , n29172 );
xor ( n29174 , n28678 , n28682 );
xor ( n29175 , n29174 , n28687 );
xor ( n29176 , n28717 , n28721 );
xor ( n29177 , n29176 , n28726 );
and ( n29178 , n29175 , n29177 );
xor ( n29179 , n28612 , n28616 );
xor ( n29180 , n29179 , n28621 );
and ( n29181 , n29177 , n29180 );
and ( n29182 , n29175 , n29180 );
or ( n29183 , n29178 , n29181 , n29182 );
and ( n29184 , n29173 , n29183 );
xor ( n29185 , n28690 , n28704 );
xor ( n29186 , n29185 , n28709 );
and ( n29187 , n29183 , n29186 );
and ( n29188 , n29173 , n29186 );
or ( n29189 , n29184 , n29187 , n29188 );
xor ( n29190 , n28778 , n28780 );
xor ( n29191 , n29190 , n28783 );
and ( n29192 , n29189 , n29191 );
xor ( n29193 , n28864 , n28866 );
xor ( n29194 , n29193 , n28869 );
and ( n29195 , n29191 , n29194 );
and ( n29196 , n29189 , n29194 );
or ( n29197 , n29192 , n29195 , n29196 );
xor ( n29198 , n28862 , n28872 );
xor ( n29199 , n29198 , n28920 );
and ( n29200 , n29197 , n29199 );
xor ( n29201 , n28786 , n28788 );
xor ( n29202 , n29201 , n28791 );
and ( n29203 , n29199 , n29202 );
and ( n29204 , n29197 , n29202 );
or ( n29205 , n29200 , n29203 , n29204 );
xor ( n29206 , n28762 , n28794 );
xor ( n29207 , n29206 , n28797 );
and ( n29208 , n29205 , n29207 );
xor ( n29209 , n28923 , n28925 );
xor ( n29210 , n29209 , n28928 );
and ( n29211 , n29207 , n29210 );
and ( n29212 , n29205 , n29210 );
or ( n29213 , n29208 , n29211 , n29212 );
and ( n29214 , n29147 , n29213 );
xor ( n29215 , n28800 , n28838 );
xor ( n29216 , n29215 , n28841 );
and ( n29217 , n29213 , n29216 );
and ( n29218 , n29147 , n29216 );
or ( n29219 , n29214 , n29217 , n29218 );
xor ( n29220 , n28566 , n28568 );
xor ( n29221 , n29220 , n28571 );
and ( n29222 , n29219 , n29221 );
xor ( n29223 , n28844 , n28939 );
xor ( n29224 , n29223 , n28942 );
and ( n29225 , n29221 , n29224 );
and ( n29226 , n29219 , n29224 );
or ( n29227 , n29222 , n29225 , n29226 );
and ( n29228 , n28957 , n29227 );
xor ( n29229 , n28957 , n29227 );
xor ( n29230 , n29219 , n29221 );
xor ( n29231 , n29230 , n29224 );
and ( n29232 , n20182 , n24902 );
and ( n29233 , n20080 , n24900 );
nor ( n29234 , n29232 , n29233 );
xnor ( n29235 , n29234 , n24397 );
and ( n29236 , n20360 , n24376 );
and ( n29237 , n20268 , n24374 );
nor ( n29238 , n29236 , n29237 );
xnor ( n29239 , n29238 , n23927 );
and ( n29240 , n29235 , n29239 );
and ( n29241 , n20618 , n23944 );
and ( n29242 , n20452 , n23942 );
nor ( n29243 , n29241 , n29242 );
xnor ( n29244 , n29243 , n23550 );
and ( n29245 , n29239 , n29244 );
and ( n29246 , n29235 , n29244 );
or ( n29247 , n29240 , n29245 , n29246 );
not ( n29248 , n28674 );
buf ( n29249 , n29248 );
and ( n29250 , n21876 , n22048 );
and ( n29251 , n21704 , n22046 );
nor ( n29252 , n29250 , n29251 );
xnor ( n29253 , n29252 , n21853 );
and ( n29254 , n29249 , n29253 );
not ( n29255 , n28893 );
and ( n29256 , n29253 , n29255 );
and ( n29257 , n29249 , n29255 );
or ( n29258 , n29254 , n29256 , n29257 );
and ( n29259 , n29247 , n29258 );
xor ( n29260 , n28733 , n28737 );
xor ( n29261 , n29260 , n28742 );
and ( n29262 , n29258 , n29261 );
and ( n29263 , n29247 , n29261 );
or ( n29264 , n29259 , n29262 , n29263 );
xor ( n29265 , n28846 , n28848 );
xor ( n29266 , n29265 , n28851 );
and ( n29267 , n29264 , n29266 );
xor ( n29268 , n28983 , n29023 );
xor ( n29269 , n29268 , n29026 );
and ( n29270 , n29266 , n29269 );
and ( n29271 , n29264 , n29269 );
or ( n29272 , n29267 , n29270 , n29271 );
xor ( n29273 , n28093 , n28673 );
xor ( n29274 , n28673 , n28674 );
not ( n29275 , n29274 );
and ( n29276 , n29273 , n29275 );
and ( n29277 , n19426 , n29276 );
not ( n29278 , n29277 );
xnor ( n29279 , n29278 , n28677 );
and ( n29280 , n19811 , n26349 );
and ( n29281 , n19721 , n26347 );
nor ( n29282 , n29280 , n29281 );
xnor ( n29283 , n29282 , n25893 );
and ( n29284 , n29279 , n29283 );
and ( n29285 , n20004 , n25383 );
and ( n29286 , n19946 , n25381 );
nor ( n29287 , n29285 , n29286 );
xnor ( n29288 , n29287 , n24885 );
and ( n29289 , n29283 , n29288 );
and ( n29290 , n29279 , n29288 );
or ( n29291 , n29284 , n29289 , n29290 );
and ( n29292 , n20803 , n23641 );
and ( n29293 , n20666 , n23639 );
nor ( n29294 , n29292 , n29293 );
xnor ( n29295 , n29294 , n23213 );
and ( n29296 , n21072 , n23230 );
and ( n29297 , n20867 , n23228 );
nor ( n29298 , n29296 , n29297 );
xnor ( n29299 , n29298 , n22842 );
and ( n29300 , n29295 , n29299 );
and ( n29301 , n21302 , n22859 );
and ( n29302 , n21218 , n22857 );
nor ( n29303 , n29301 , n29302 );
xnor ( n29304 , n29303 , n22418 );
and ( n29305 , n29299 , n29304 );
and ( n29306 , n29295 , n29304 );
or ( n29307 , n29300 , n29305 , n29306 );
and ( n29308 , n29291 , n29307 );
and ( n29309 , n22198 , n21741 );
and ( n29310 , n22235 , n21739 );
nor ( n29311 , n29309 , n29310 );
xnor ( n29312 , n29311 , n21605 );
and ( n29313 , n22756 , n21468 );
and ( n29314 , n22425 , n21466 );
nor ( n29315 , n29313 , n29314 );
xnor ( n29316 , n29315 , n21331 );
and ( n29317 , n29312 , n29316 );
buf ( n29318 , n19345 );
and ( n29319 , n29318 , n19419 );
and ( n29320 , n29316 , n29319 );
and ( n29321 , n29312 , n29319 );
or ( n29322 , n29317 , n29320 , n29321 );
and ( n29323 , n19434 , n28628 );
and ( n29324 , n19418 , n28626 );
nor ( n29325 , n29323 , n29324 );
xnor ( n29326 , n29325 , n28096 );
and ( n29327 , n29322 , n29326 );
and ( n29328 , n21612 , n22381 );
and ( n29329 , n21451 , n22379 );
nor ( n29330 , n29328 , n29329 );
xnor ( n29331 , n29330 , n22228 );
and ( n29332 , n29326 , n29331 );
and ( n29333 , n29322 , n29331 );
or ( n29334 , n29327 , n29332 , n29333 );
and ( n29335 , n29307 , n29334 );
and ( n29336 , n29291 , n29334 );
or ( n29337 , n29308 , n29335 , n29336 );
xor ( n29338 , n28971 , n28975 );
xor ( n29339 , n29338 , n28980 );
xor ( n29340 , n28877 , n28881 );
xor ( n29341 , n29340 , n28886 );
and ( n29342 , n29339 , n29341 );
xor ( n29343 , n28894 , n28898 );
xor ( n29344 , n29343 , n28903 );
and ( n29345 , n29341 , n29344 );
and ( n29346 , n29339 , n29344 );
or ( n29347 , n29342 , n29345 , n29346 );
and ( n29348 , n29337 , n29347 );
xor ( n29349 , n28889 , n28906 );
xor ( n29350 , n29349 , n28909 );
and ( n29351 , n29347 , n29350 );
and ( n29352 , n29337 , n29350 );
or ( n29353 , n29348 , n29351 , n29352 );
and ( n29354 , n29272 , n29353 );
xor ( n29355 , n28854 , n28856 );
xor ( n29356 , n29355 , n28859 );
and ( n29357 , n29353 , n29356 );
and ( n29358 , n29272 , n29356 );
or ( n29359 , n29354 , n29357 , n29358 );
and ( n29360 , n26851 , n19688 );
and ( n29361 , n26422 , n19686 );
nor ( n29362 , n29360 , n29361 );
xnor ( n29363 , n29362 , n19655 );
and ( n29364 , n27352 , n19596 );
and ( n29365 , n27135 , n19594 );
nor ( n29366 , n29364 , n29365 );
xnor ( n29367 , n29366 , n19545 );
and ( n29368 , n29363 , n29367 );
and ( n29369 , n27757 , n19518 );
and ( n29370 , n27751 , n19516 );
nor ( n29371 , n29369 , n29370 );
xnor ( n29372 , n29371 , n19489 );
and ( n29373 , n29367 , n29372 );
and ( n29374 , n29363 , n29372 );
or ( n29375 , n29368 , n29373 , n29374 );
and ( n29376 , n25284 , n20114 );
and ( n29377 , n24940 , n20112 );
nor ( n29378 , n29376 , n29377 );
xnor ( n29379 , n29378 , n19997 );
and ( n29380 , n25765 , n19894 );
and ( n29381 , n25554 , n19892 );
nor ( n29382 , n29380 , n29381 );
xnor ( n29383 , n29382 , n19858 );
and ( n29384 , n29379 , n29383 );
and ( n29385 , n26319 , n19805 );
and ( n29386 , n25974 , n19803 );
nor ( n29387 , n29385 , n29386 );
xnor ( n29388 , n29387 , n19750 );
and ( n29389 , n29383 , n29388 );
and ( n29390 , n29379 , n29388 );
or ( n29391 , n29384 , n29389 , n29390 );
and ( n29392 , n29375 , n29391 );
and ( n29393 , n19637 , n26992 );
and ( n29394 , n19605 , n26990 );
nor ( n29395 , n29393 , n29394 );
xnor ( n29396 , n29395 , n26369 );
and ( n29397 , n29391 , n29396 );
and ( n29398 , n29375 , n29396 );
or ( n29399 , n29392 , n29397 , n29398 );
and ( n29400 , n23141 , n21155 );
and ( n29401 , n22916 , n21153 );
nor ( n29402 , n29400 , n29401 );
xnor ( n29403 , n29402 , n20994 );
and ( n29404 , n23381 , n20955 );
and ( n29405 , n23271 , n20953 );
nor ( n29406 , n29404 , n29405 );
xnor ( n29407 , n29406 , n20780 );
and ( n29408 , n29403 , n29407 );
and ( n29409 , n29078 , n19424 );
and ( n29410 , n28700 , n19422 );
nor ( n29411 , n29409 , n29410 );
xnor ( n29412 , n29411 , n19431 );
and ( n29413 , n29407 , n29412 );
and ( n29414 , n29403 , n29412 );
or ( n29415 , n29408 , n29413 , n29414 );
and ( n29416 , n23968 , n20674 );
and ( n29417 , n23573 , n20672 );
nor ( n29418 , n29416 , n29417 );
xnor ( n29419 , n29418 , n20542 );
and ( n29420 , n24521 , n20460 );
and ( n29421 , n24131 , n20458 );
nor ( n29422 , n29420 , n29421 );
xnor ( n29423 , n29422 , n20337 );
and ( n29424 , n29419 , n29423 );
and ( n29425 , n24621 , n20276 );
and ( n29426 , n24527 , n20274 );
nor ( n29427 , n29425 , n29426 );
xnor ( n29428 , n29427 , n20175 );
and ( n29429 , n29423 , n29428 );
and ( n29430 , n29419 , n29428 );
or ( n29431 , n29424 , n29429 , n29430 );
and ( n29432 , n29415 , n29431 );
and ( n29433 , n19588 , n27529 );
and ( n29434 , n19510 , n27527 );
nor ( n29435 , n29433 , n29434 );
xnor ( n29436 , n29435 , n27034 );
and ( n29437 , n29431 , n29436 );
and ( n29438 , n29415 , n29436 );
or ( n29439 , n29432 , n29437 , n29438 );
and ( n29440 , n29399 , n29439 );
xor ( n29441 , n29055 , n29059 );
xor ( n29442 , n29441 , n29064 );
and ( n29443 , n29439 , n29442 );
and ( n29444 , n29399 , n29442 );
or ( n29445 , n29440 , n29443 , n29444 );
xor ( n29446 , n29086 , n29090 );
xor ( n29447 , n29446 , n29095 );
xor ( n29448 , n29151 , n29155 );
xor ( n29449 , n29448 , n29160 );
and ( n29450 , n29447 , n29449 );
xor ( n29451 , n28987 , n28991 );
xor ( n29452 , n29451 , n28996 );
and ( n29453 , n29449 , n29452 );
and ( n29454 , n29447 , n29452 );
or ( n29455 , n29450 , n29453 , n29454 );
xor ( n29456 , n29039 , n29043 );
xor ( n29457 , n29456 , n29048 );
and ( n29458 , n29455 , n29457 );
xor ( n29459 , n29082 , n29098 );
xor ( n29460 , n29459 , n29103 );
and ( n29461 , n29457 , n29460 );
and ( n29462 , n29455 , n29460 );
or ( n29463 , n29458 , n29461 , n29462 );
and ( n29464 , n29445 , n29463 );
xor ( n29465 , n29051 , n29067 );
xor ( n29466 , n29465 , n29106 );
and ( n29467 , n29463 , n29466 );
and ( n29468 , n29445 , n29466 );
or ( n29469 , n29464 , n29467 , n29468 );
xor ( n29470 , n28967 , n29029 );
xor ( n29471 , n29470 , n29032 );
and ( n29472 , n29469 , n29471 );
xor ( n29473 , n28912 , n28914 );
xor ( n29474 , n29473 , n28917 );
and ( n29475 , n29471 , n29474 );
and ( n29476 , n29469 , n29474 );
or ( n29477 , n29472 , n29475 , n29476 );
and ( n29478 , n29359 , n29477 );
xor ( n29479 , n29133 , n29135 );
xor ( n29480 , n29479 , n29138 );
and ( n29481 , n29477 , n29480 );
and ( n29482 , n29359 , n29480 );
or ( n29483 , n29478 , n29481 , n29482 );
and ( n29484 , n19496 , n28062 );
and ( n29485 , n19469 , n28060 );
nor ( n29486 , n29484 , n29485 );
xnor ( n29487 , n29486 , n27549 );
and ( n29488 , n19881 , n26027 );
and ( n29489 , n19825 , n26025 );
nor ( n29490 , n29488 , n29489 );
xnor ( n29491 , n29490 , n25499 );
and ( n29492 , n29487 , n29491 );
xor ( n29493 , n29072 , n29076 );
xor ( n29494 , n29493 , n29079 );
and ( n29495 , n29491 , n29494 );
and ( n29496 , n29487 , n29494 );
or ( n29497 , n29492 , n29495 , n29496 );
xor ( n29498 , n28999 , n29015 );
xor ( n29499 , n29498 , n29020 );
and ( n29500 , n29497 , n29499 );
xor ( n29501 , n29163 , n29167 );
xor ( n29502 , n29501 , n29170 );
and ( n29503 , n29499 , n29502 );
and ( n29504 , n29497 , n29502 );
or ( n29505 , n29500 , n29503 , n29504 );
xor ( n29506 , n28959 , n28961 );
xor ( n29507 , n29506 , n28964 );
and ( n29508 , n29505 , n29507 );
xor ( n29509 , n29111 , n29113 );
xor ( n29510 , n29509 , n29116 );
and ( n29511 , n29507 , n29510 );
and ( n29512 , n29505 , n29510 );
or ( n29513 , n29508 , n29511 , n29512 );
xor ( n29514 , n29109 , n29119 );
xor ( n29515 , n29514 , n29122 );
and ( n29516 , n29513 , n29515 );
xor ( n29517 , n29189 , n29191 );
xor ( n29518 , n29517 , n29194 );
and ( n29519 , n29515 , n29518 );
and ( n29520 , n29513 , n29518 );
or ( n29521 , n29516 , n29519 , n29520 );
xor ( n29522 , n29035 , n29125 );
xor ( n29523 , n29522 , n29128 );
and ( n29524 , n29521 , n29523 );
xor ( n29525 , n29197 , n29199 );
xor ( n29526 , n29525 , n29202 );
and ( n29527 , n29523 , n29526 );
and ( n29528 , n29521 , n29526 );
or ( n29529 , n29524 , n29527 , n29528 );
and ( n29530 , n29483 , n29529 );
xor ( n29531 , n29131 , n29141 );
xor ( n29532 , n29531 , n29144 );
and ( n29533 , n29529 , n29532 );
and ( n29534 , n29483 , n29532 );
or ( n29535 , n29530 , n29533 , n29534 );
xor ( n29536 , n28931 , n28933 );
xor ( n29537 , n29536 , n28936 );
and ( n29538 , n29535 , n29537 );
xor ( n29539 , n29147 , n29213 );
xor ( n29540 , n29539 , n29216 );
and ( n29541 , n29537 , n29540 );
and ( n29542 , n29535 , n29540 );
or ( n29543 , n29538 , n29541 , n29542 );
and ( n29544 , n29231 , n29543 );
xor ( n29545 , n29231 , n29543 );
xor ( n29546 , n29535 , n29537 );
xor ( n29547 , n29546 , n29540 );
and ( n29548 , n20080 , n25383 );
and ( n29549 , n20004 , n25381 );
nor ( n29550 , n29548 , n29549 );
xnor ( n29551 , n29550 , n24885 );
and ( n29552 , n20268 , n24902 );
and ( n29553 , n20182 , n24900 );
nor ( n29554 , n29552 , n29553 );
xnor ( n29555 , n29554 , n24397 );
and ( n29556 , n29551 , n29555 );
and ( n29557 , n21704 , n22381 );
and ( n29558 , n21612 , n22379 );
nor ( n29559 , n29557 , n29558 );
xnor ( n29560 , n29559 , n22228 );
and ( n29561 , n29555 , n29560 );
and ( n29562 , n29551 , n29560 );
or ( n29563 , n29556 , n29561 , n29562 );
and ( n29564 , n21955 , n22048 );
and ( n29565 , n21876 , n22046 );
nor ( n29566 , n29564 , n29565 );
xnor ( n29567 , n29566 , n21853 );
and ( n29568 , n28674 , n29567 );
and ( n29569 , n28810 , n19459 );
and ( n29570 , n28211 , n19457 );
nor ( n29571 , n29569 , n29570 );
xnor ( n29572 , n29571 , n19416 );
and ( n29573 , n29567 , n29572 );
and ( n29574 , n28674 , n29572 );
or ( n29575 , n29568 , n29573 , n29574 );
and ( n29576 , n29563 , n29575 );
xor ( n29577 , n29003 , n29007 );
xor ( n29578 , n29577 , n29012 );
and ( n29579 , n29575 , n29578 );
and ( n29580 , n29563 , n29578 );
or ( n29581 , n29576 , n29579 , n29580 );
xor ( n29582 , n29175 , n29177 );
xor ( n29583 , n29582 , n29180 );
and ( n29584 , n29581 , n29583 );
xor ( n29585 , n29247 , n29258 );
xor ( n29586 , n29585 , n29261 );
and ( n29587 , n29583 , n29586 );
and ( n29588 , n29581 , n29586 );
or ( n29589 , n29584 , n29587 , n29588 );
xor ( n29590 , n29173 , n29183 );
xor ( n29591 , n29590 , n29186 );
and ( n29592 , n29589 , n29591 );
xor ( n29593 , n29264 , n29266 );
xor ( n29594 , n29593 , n29269 );
and ( n29595 , n29591 , n29594 );
and ( n29596 , n29589 , n29594 );
or ( n29597 , n29592 , n29595 , n29596 );
and ( n29598 , n19946 , n26027 );
and ( n29599 , n19881 , n26025 );
nor ( n29600 , n29598 , n29599 );
xnor ( n29601 , n29600 , n25499 );
and ( n29602 , n21218 , n23230 );
and ( n29603 , n21072 , n23228 );
nor ( n29604 , n29602 , n29603 );
xnor ( n29605 , n29604 , n22842 );
and ( n29606 , n29601 , n29605 );
and ( n29607 , n21451 , n22859 );
and ( n29608 , n21302 , n22857 );
nor ( n29609 , n29607 , n29608 );
xnor ( n29610 , n29609 , n22418 );
and ( n29611 , n29605 , n29610 );
and ( n29612 , n29601 , n29610 );
or ( n29613 , n29606 , n29611 , n29612 );
and ( n29614 , n22425 , n21741 );
and ( n29615 , n22198 , n21739 );
nor ( n29616 , n29614 , n29615 );
xnor ( n29617 , n29616 , n21605 );
and ( n29618 , n22916 , n21468 );
and ( n29619 , n22756 , n21466 );
nor ( n29620 , n29618 , n29619 );
xnor ( n29621 , n29620 , n21331 );
and ( n29622 , n29617 , n29621 );
buf ( n29623 , n19346 );
and ( n29624 , n29623 , n19419 );
and ( n29625 , n29621 , n29624 );
and ( n29626 , n29617 , n29624 );
or ( n29627 , n29622 , n29625 , n29626 );
and ( n29628 , n19418 , n29276 );
and ( n29629 , n19426 , n29274 );
nor ( n29630 , n29628 , n29629 );
xnor ( n29631 , n29630 , n28677 );
and ( n29632 , n29627 , n29631 );
and ( n29633 , n19510 , n28062 );
and ( n29634 , n19496 , n28060 );
nor ( n29635 , n29633 , n29634 );
xnor ( n29636 , n29635 , n27549 );
and ( n29637 , n29631 , n29636 );
and ( n29638 , n29627 , n29636 );
or ( n29639 , n29632 , n29637 , n29638 );
and ( n29640 , n29613 , n29639 );
and ( n29641 , n27135 , n19688 );
and ( n29642 , n26851 , n19686 );
nor ( n29643 , n29641 , n29642 );
xnor ( n29644 , n29643 , n19655 );
and ( n29645 , n27751 , n19596 );
and ( n29646 , n27352 , n19594 );
nor ( n29647 , n29645 , n29646 );
xnor ( n29648 , n29647 , n19545 );
and ( n29649 , n29644 , n29648 );
and ( n29650 , n28211 , n19518 );
and ( n29651 , n27757 , n19516 );
nor ( n29652 , n29650 , n29651 );
xnor ( n29653 , n29652 , n19489 );
and ( n29654 , n29648 , n29653 );
and ( n29655 , n29644 , n29653 );
or ( n29656 , n29649 , n29654 , n29655 );
and ( n29657 , n19605 , n27529 );
and ( n29658 , n19588 , n27527 );
nor ( n29659 , n29657 , n29658 );
xnor ( n29660 , n29659 , n27034 );
and ( n29661 , n29656 , n29660 );
and ( n29662 , n19721 , n26992 );
and ( n29663 , n19637 , n26990 );
nor ( n29664 , n29662 , n29663 );
xnor ( n29665 , n29664 , n26369 );
and ( n29666 , n29660 , n29665 );
and ( n29667 , n29656 , n29665 );
or ( n29668 , n29661 , n29666 , n29667 );
and ( n29669 , n29639 , n29668 );
and ( n29670 , n29613 , n29668 );
or ( n29671 , n29640 , n29669 , n29670 );
and ( n29672 , n20452 , n24376 );
and ( n29673 , n20360 , n24374 );
nor ( n29674 , n29672 , n29673 );
xnor ( n29675 , n29674 , n23927 );
and ( n29676 , n20666 , n23944 );
and ( n29677 , n20618 , n23942 );
nor ( n29678 , n29676 , n29677 );
xnor ( n29679 , n29678 , n23550 );
and ( n29680 , n29675 , n29679 );
and ( n29681 , n20867 , n23641 );
and ( n29682 , n20803 , n23639 );
nor ( n29683 , n29681 , n29682 );
xnor ( n29684 , n29683 , n23213 );
and ( n29685 , n29679 , n29684 );
and ( n29686 , n29675 , n29684 );
or ( n29687 , n29680 , n29685 , n29686 );
and ( n29688 , n23271 , n21155 );
and ( n29689 , n23141 , n21153 );
nor ( n29690 , n29688 , n29689 );
xnor ( n29691 , n29690 , n20994 );
and ( n29692 , n23573 , n20955 );
and ( n29693 , n23381 , n20953 );
nor ( n29694 , n29692 , n29693 );
xnor ( n29695 , n29694 , n20780 );
and ( n29696 , n29691 , n29695 );
and ( n29697 , n29318 , n19424 );
and ( n29698 , n29078 , n19422 );
nor ( n29699 , n29697 , n29698 );
xnor ( n29700 , n29699 , n19431 );
and ( n29701 , n29695 , n29700 );
and ( n29702 , n29691 , n29700 );
or ( n29703 , n29696 , n29701 , n29702 );
and ( n29704 , n24131 , n20674 );
and ( n29705 , n23968 , n20672 );
nor ( n29706 , n29704 , n29705 );
xnor ( n29707 , n29706 , n20542 );
and ( n29708 , n24527 , n20460 );
and ( n29709 , n24521 , n20458 );
nor ( n29710 , n29708 , n29709 );
xnor ( n29711 , n29710 , n20337 );
and ( n29712 , n29707 , n29711 );
and ( n29713 , n24940 , n20276 );
and ( n29714 , n24621 , n20274 );
nor ( n29715 , n29713 , n29714 );
xnor ( n29716 , n29715 , n20175 );
and ( n29717 , n29711 , n29716 );
and ( n29718 , n29707 , n29716 );
or ( n29719 , n29712 , n29717 , n29718 );
and ( n29720 , n29703 , n29719 );
and ( n29721 , n25554 , n20114 );
and ( n29722 , n25284 , n20112 );
nor ( n29723 , n29721 , n29722 );
xnor ( n29724 , n29723 , n19997 );
and ( n29725 , n25974 , n19894 );
and ( n29726 , n25765 , n19892 );
nor ( n29727 , n29725 , n29726 );
xnor ( n29728 , n29727 , n19858 );
and ( n29729 , n29724 , n29728 );
and ( n29730 , n26422 , n19805 );
and ( n29731 , n26319 , n19803 );
nor ( n29732 , n29730 , n29731 );
xnor ( n29733 , n29732 , n19750 );
and ( n29734 , n29728 , n29733 );
and ( n29735 , n29724 , n29733 );
or ( n29736 , n29729 , n29734 , n29735 );
and ( n29737 , n29719 , n29736 );
and ( n29738 , n29703 , n29736 );
or ( n29739 , n29720 , n29737 , n29738 );
and ( n29740 , n29687 , n29739 );
xor ( n29741 , n29249 , n29253 );
xor ( n29742 , n29741 , n29255 );
and ( n29743 , n29739 , n29742 );
and ( n29744 , n29687 , n29742 );
or ( n29745 , n29740 , n29743 , n29744 );
and ( n29746 , n29671 , n29745 );
xor ( n29747 , n29312 , n29316 );
xor ( n29748 , n29747 , n29319 );
xor ( n29749 , n29419 , n29423 );
xor ( n29750 , n29749 , n29428 );
and ( n29751 , n29748 , n29750 );
xor ( n29752 , n29363 , n29367 );
xor ( n29753 , n29752 , n29372 );
and ( n29754 , n29750 , n29753 );
and ( n29755 , n29748 , n29753 );
or ( n29756 , n29751 , n29754 , n29755 );
xor ( n29757 , n29279 , n29283 );
xor ( n29758 , n29757 , n29288 );
and ( n29759 , n29756 , n29758 );
xor ( n29760 , n29322 , n29326 );
xor ( n29761 , n29760 , n29331 );
and ( n29762 , n29758 , n29761 );
and ( n29763 , n29756 , n29761 );
or ( n29764 , n29759 , n29762 , n29763 );
and ( n29765 , n29745 , n29764 );
and ( n29766 , n29671 , n29764 );
or ( n29767 , n29746 , n29765 , n29766 );
xor ( n29768 , n29375 , n29391 );
xor ( n29769 , n29768 , n29396 );
xor ( n29770 , n29415 , n29431 );
xor ( n29771 , n29770 , n29436 );
and ( n29772 , n29769 , n29771 );
xor ( n29773 , n29487 , n29491 );
xor ( n29774 , n29773 , n29494 );
and ( n29775 , n29771 , n29774 );
and ( n29776 , n29769 , n29774 );
or ( n29777 , n29772 , n29775 , n29776 );
xor ( n29778 , n29291 , n29307 );
xor ( n29779 , n29778 , n29334 );
and ( n29780 , n29777 , n29779 );
xor ( n29781 , n29399 , n29439 );
xor ( n29782 , n29781 , n29442 );
and ( n29783 , n29779 , n29782 );
and ( n29784 , n29777 , n29782 );
or ( n29785 , n29780 , n29783 , n29784 );
and ( n29786 , n29767 , n29785 );
xor ( n29787 , n29337 , n29347 );
xor ( n29788 , n29787 , n29350 );
and ( n29789 , n29785 , n29788 );
and ( n29790 , n29767 , n29788 );
or ( n29791 , n29786 , n29789 , n29790 );
and ( n29792 , n29597 , n29791 );
xor ( n29793 , n29272 , n29353 );
xor ( n29794 , n29793 , n29356 );
and ( n29795 , n29791 , n29794 );
and ( n29796 , n29597 , n29794 );
or ( n29797 , n29792 , n29795 , n29796 );
xor ( n29798 , n29359 , n29477 );
xor ( n29799 , n29798 , n29480 );
and ( n29800 , n29797 , n29799 );
xor ( n29801 , n29521 , n29523 );
xor ( n29802 , n29801 , n29526 );
and ( n29803 , n29799 , n29802 );
and ( n29804 , n29797 , n29802 );
or ( n29805 , n29800 , n29803 , n29804 );
xor ( n29806 , n29205 , n29207 );
xor ( n29807 , n29806 , n29210 );
and ( n29808 , n29805 , n29807 );
xor ( n29809 , n29483 , n29529 );
xor ( n29810 , n29809 , n29532 );
and ( n29811 , n29807 , n29810 );
and ( n29812 , n29805 , n29810 );
or ( n29813 , n29808 , n29811 , n29812 );
and ( n29814 , n29547 , n29813 );
xor ( n29815 , n29547 , n29813 );
xor ( n29816 , n29805 , n29807 );
xor ( n29817 , n29816 , n29810 );
and ( n29818 , n19469 , n28628 );
and ( n29819 , n19434 , n28626 );
nor ( n29820 , n29818 , n29819 );
xnor ( n29821 , n29820 , n28096 );
and ( n29822 , n19825 , n26349 );
and ( n29823 , n19811 , n26347 );
nor ( n29824 , n29822 , n29823 );
xnor ( n29825 , n29824 , n25893 );
and ( n29826 , n29821 , n29825 );
xor ( n29827 , n29403 , n29407 );
xor ( n29828 , n29827 , n29412 );
and ( n29829 , n29825 , n29828 );
and ( n29830 , n29821 , n29828 );
or ( n29831 , n29826 , n29829 , n29830 );
xor ( n29832 , n29235 , n29239 );
xor ( n29833 , n29832 , n29244 );
and ( n29834 , n29831 , n29833 );
xor ( n29835 , n29295 , n29299 );
xor ( n29836 , n29835 , n29304 );
and ( n29837 , n29833 , n29836 );
and ( n29838 , n29831 , n29836 );
or ( n29839 , n29834 , n29837 , n29838 );
xor ( n29840 , n29455 , n29457 );
xor ( n29841 , n29840 , n29460 );
and ( n29842 , n29839 , n29841 );
xor ( n29843 , n29339 , n29341 );
xor ( n29844 , n29843 , n29344 );
and ( n29845 , n29841 , n29844 );
and ( n29846 , n29839 , n29844 );
or ( n29847 , n29842 , n29845 , n29846 );
xor ( n29848 , n29445 , n29463 );
xor ( n29849 , n29848 , n29466 );
and ( n29850 , n29847 , n29849 );
xor ( n29851 , n29505 , n29507 );
xor ( n29852 , n29851 , n29510 );
and ( n29853 , n29849 , n29852 );
and ( n29854 , n29847 , n29852 );
or ( n29855 , n29850 , n29853 , n29854 );
xor ( n29856 , n29513 , n29515 );
xor ( n29857 , n29856 , n29518 );
and ( n29858 , n29855 , n29857 );
xor ( n29859 , n29469 , n29471 );
xor ( n29860 , n29859 , n29474 );
and ( n29861 , n29857 , n29860 );
and ( n29862 , n29855 , n29860 );
or ( n29863 , n29858 , n29861 , n29862 );
and ( n29864 , n21876 , n22381 );
and ( n29865 , n21704 , n22379 );
nor ( n29866 , n29864 , n29865 );
xnor ( n29867 , n29866 , n22228 );
and ( n29868 , n22235 , n22048 );
and ( n29869 , n21955 , n22046 );
nor ( n29870 , n29868 , n29869 );
xnor ( n29871 , n29870 , n21853 );
and ( n29872 , n29867 , n29871 );
and ( n29873 , n28700 , n19459 );
and ( n29874 , n28810 , n19457 );
nor ( n29875 , n29873 , n29874 );
xnor ( n29876 , n29875 , n19416 );
and ( n29877 , n29871 , n29876 );
and ( n29878 , n29867 , n29876 );
or ( n29879 , n29872 , n29877 , n29878 );
and ( n29880 , n20618 , n24376 );
and ( n29881 , n20452 , n24374 );
nor ( n29882 , n29880 , n29881 );
xnor ( n29883 , n29882 , n23927 );
and ( n29884 , n20803 , n23944 );
and ( n29885 , n20666 , n23942 );
nor ( n29886 , n29884 , n29885 );
xnor ( n29887 , n29886 , n23550 );
and ( n29888 , n29883 , n29887 );
and ( n29889 , n21072 , n23641 );
and ( n29890 , n20867 , n23639 );
nor ( n29891 , n29889 , n29890 );
xnor ( n29892 , n29891 , n23213 );
and ( n29893 , n29887 , n29892 );
and ( n29894 , n29883 , n29892 );
or ( n29895 , n29888 , n29893 , n29894 );
and ( n29896 , n29879 , n29895 );
xor ( n29897 , n29379 , n29383 );
xor ( n29898 , n29897 , n29388 );
and ( n29899 , n29895 , n29898 );
and ( n29900 , n29879 , n29898 );
or ( n29901 , n29896 , n29899 , n29900 );
and ( n29902 , n20004 , n26027 );
and ( n29903 , n19946 , n26025 );
nor ( n29904 , n29902 , n29903 );
xnor ( n29905 , n29904 , n25499 );
and ( n29906 , n21302 , n23230 );
and ( n29907 , n21218 , n23228 );
nor ( n29908 , n29906 , n29907 );
xnor ( n29909 , n29908 , n22842 );
and ( n29910 , n29905 , n29909 );
and ( n29911 , n21612 , n22859 );
and ( n29912 , n21451 , n22857 );
nor ( n29913 , n29911 , n29912 );
xnor ( n29914 , n29913 , n22418 );
and ( n29915 , n29909 , n29914 );
and ( n29916 , n29905 , n29914 );
or ( n29917 , n29910 , n29915 , n29916 );
and ( n29918 , n22756 , n21741 );
and ( n29919 , n22425 , n21739 );
nor ( n29920 , n29918 , n29919 );
xnor ( n29921 , n29920 , n21605 );
and ( n29922 , n23141 , n21468 );
and ( n29923 , n22916 , n21466 );
nor ( n29924 , n29922 , n29923 );
xnor ( n29925 , n29924 , n21331 );
and ( n29926 , n29921 , n29925 );
and ( n29927 , n29623 , n19424 );
and ( n29928 , n29318 , n19422 );
nor ( n29929 , n29927 , n29928 );
xnor ( n29930 , n29929 , n19431 );
and ( n29931 , n29925 , n29930 );
and ( n29932 , n29921 , n29930 );
or ( n29933 , n29926 , n29931 , n29932 );
and ( n29934 , n19434 , n29276 );
and ( n29935 , n19418 , n29274 );
nor ( n29936 , n29934 , n29935 );
xnor ( n29937 , n29936 , n28677 );
and ( n29938 , n29933 , n29937 );
and ( n29939 , n19588 , n28062 );
and ( n29940 , n19510 , n28060 );
nor ( n29941 , n29939 , n29940 );
xnor ( n29942 , n29941 , n27549 );
and ( n29943 , n29937 , n29942 );
and ( n29944 , n29933 , n29942 );
or ( n29945 , n29938 , n29943 , n29944 );
and ( n29946 , n29917 , n29945 );
xor ( n29947 , n29601 , n29605 );
xor ( n29948 , n29947 , n29610 );
and ( n29949 , n29945 , n29948 );
and ( n29950 , n29917 , n29948 );
or ( n29951 , n29946 , n29949 , n29950 );
and ( n29952 , n29901 , n29951 );
xor ( n29953 , n29447 , n29449 );
xor ( n29954 , n29953 , n29452 );
and ( n29955 , n29951 , n29954 );
and ( n29956 , n29901 , n29954 );
or ( n29957 , n29952 , n29955 , n29956 );
and ( n29958 , n27757 , n19596 );
and ( n29959 , n27751 , n19594 );
nor ( n29960 , n29958 , n29959 );
xnor ( n29961 , n29960 , n19545 );
and ( n29962 , n28810 , n19518 );
and ( n29963 , n28211 , n19516 );
nor ( n29964 , n29962 , n29963 );
xnor ( n29965 , n29964 , n19489 );
and ( n29966 , n29961 , n29965 );
and ( n29967 , n29078 , n19459 );
and ( n29968 , n28700 , n19457 );
nor ( n29969 , n29967 , n29968 );
xnor ( n29970 , n29969 , n19416 );
and ( n29971 , n29965 , n29970 );
and ( n29972 , n29961 , n29970 );
or ( n29973 , n29966 , n29971 , n29972 );
buf ( n29974 , n19410 );
xor ( n29975 , n28674 , n29974 );
not ( n29976 , n29974 );
and ( n29977 , n29975 , n29976 );
and ( n29978 , n19426 , n29977 );
not ( n29979 , n29978 );
xnor ( n29980 , n29979 , n28674 );
and ( n29981 , n29973 , n29980 );
and ( n29982 , n19637 , n27529 );
and ( n29983 , n19605 , n27527 );
nor ( n29984 , n29982 , n29983 );
xnor ( n29985 , n29984 , n27034 );
and ( n29986 , n29980 , n29985 );
and ( n29987 , n29973 , n29985 );
or ( n29988 , n29981 , n29986 , n29987 );
and ( n29989 , n22198 , n22048 );
and ( n29990 , n22235 , n22046 );
nor ( n29991 , n29989 , n29990 );
xnor ( n29992 , n29991 , n21853 );
and ( n29993 , n29623 , n19422 );
not ( n29994 , n29993 );
and ( n29995 , n29994 , n19431 );
and ( n29996 , n29992 , n29995 );
and ( n29997 , n20182 , n25383 );
and ( n29998 , n20080 , n25381 );
nor ( n29999 , n29997 , n29998 );
xnor ( n30000 , n29999 , n24885 );
and ( n30001 , n29996 , n30000 );
and ( n30002 , n20360 , n24902 );
and ( n30003 , n20268 , n24900 );
nor ( n30004 , n30002 , n30003 );
xnor ( n30005 , n30004 , n24397 );
and ( n30006 , n30000 , n30005 );
and ( n30007 , n29996 , n30005 );
or ( n30008 , n30001 , n30006 , n30007 );
and ( n30009 , n29988 , n30008 );
xor ( n30010 , n28674 , n29567 );
xor ( n30011 , n30010 , n29572 );
and ( n30012 , n30008 , n30011 );
and ( n30013 , n29988 , n30011 );
or ( n30014 , n30009 , n30012 , n30013 );
and ( n30015 , n19496 , n28628 );
and ( n30016 , n19469 , n28626 );
nor ( n30017 , n30015 , n30016 );
xnor ( n30018 , n30017 , n28096 );
and ( n30019 , n19811 , n26992 );
and ( n30020 , n19721 , n26990 );
nor ( n30021 , n30019 , n30020 );
xnor ( n30022 , n30021 , n26369 );
and ( n30023 , n30018 , n30022 );
and ( n30024 , n19881 , n26349 );
and ( n30025 , n19825 , n26347 );
nor ( n30026 , n30024 , n30025 );
xnor ( n30027 , n30026 , n25893 );
and ( n30028 , n30022 , n30027 );
and ( n30029 , n30018 , n30027 );
or ( n30030 , n30023 , n30028 , n30029 );
and ( n30031 , n23381 , n21155 );
and ( n30032 , n23271 , n21153 );
nor ( n30033 , n30031 , n30032 );
xnor ( n30034 , n30033 , n20994 );
and ( n30035 , n23968 , n20955 );
and ( n30036 , n23573 , n20953 );
nor ( n30037 , n30035 , n30036 );
xnor ( n30038 , n30037 , n20780 );
and ( n30039 , n30034 , n30038 );
and ( n30040 , n24521 , n20674 );
and ( n30041 , n24131 , n20672 );
nor ( n30042 , n30040 , n30041 );
xnor ( n30043 , n30042 , n20542 );
and ( n30044 , n30038 , n30043 );
and ( n30045 , n30034 , n30043 );
or ( n30046 , n30039 , n30044 , n30045 );
and ( n30047 , n26319 , n19894 );
and ( n30048 , n25974 , n19892 );
nor ( n30049 , n30047 , n30048 );
xnor ( n30050 , n30049 , n19858 );
and ( n30051 , n26851 , n19805 );
and ( n30052 , n26422 , n19803 );
nor ( n30053 , n30051 , n30052 );
xnor ( n30054 , n30053 , n19750 );
and ( n30055 , n30050 , n30054 );
and ( n30056 , n27352 , n19688 );
and ( n30057 , n27135 , n19686 );
nor ( n30058 , n30056 , n30057 );
xnor ( n30059 , n30058 , n19655 );
and ( n30060 , n30054 , n30059 );
and ( n30061 , n30050 , n30059 );
or ( n30062 , n30055 , n30060 , n30061 );
and ( n30063 , n30046 , n30062 );
and ( n30064 , n24621 , n20460 );
and ( n30065 , n24527 , n20458 );
nor ( n30066 , n30064 , n30065 );
xnor ( n30067 , n30066 , n20337 );
and ( n30068 , n25284 , n20276 );
and ( n30069 , n24940 , n20274 );
nor ( n30070 , n30068 , n30069 );
xnor ( n30071 , n30070 , n20175 );
and ( n30072 , n30067 , n30071 );
and ( n30073 , n25765 , n20114 );
and ( n30074 , n25554 , n20112 );
nor ( n30075 , n30073 , n30074 );
xnor ( n30076 , n30075 , n19997 );
and ( n30077 , n30071 , n30076 );
and ( n30078 , n30067 , n30076 );
or ( n30079 , n30072 , n30077 , n30078 );
and ( n30080 , n30062 , n30079 );
and ( n30081 , n30046 , n30079 );
or ( n30082 , n30063 , n30080 , n30081 );
and ( n30083 , n30030 , n30082 );
xor ( n30084 , n29551 , n29555 );
xor ( n30085 , n30084 , n29560 );
and ( n30086 , n30082 , n30085 );
and ( n30087 , n30030 , n30085 );
or ( n30088 , n30083 , n30086 , n30087 );
and ( n30089 , n30014 , n30088 );
xor ( n30090 , n29563 , n29575 );
xor ( n30091 , n30090 , n29578 );
and ( n30092 , n30088 , n30091 );
and ( n30093 , n30014 , n30091 );
or ( n30094 , n30089 , n30092 , n30093 );
and ( n30095 , n29957 , n30094 );
xor ( n30096 , n29497 , n29499 );
xor ( n30097 , n30096 , n29502 );
and ( n30098 , n30094 , n30097 );
and ( n30099 , n29957 , n30097 );
or ( n30100 , n30095 , n30098 , n30099 );
xor ( n30101 , n29617 , n29621 );
xor ( n30102 , n30101 , n29624 );
xor ( n30103 , n29691 , n29695 );
xor ( n30104 , n30103 , n29700 );
and ( n30105 , n30102 , n30104 );
xor ( n30106 , n29707 , n29711 );
xor ( n30107 , n30106 , n29716 );
and ( n30108 , n30104 , n30107 );
and ( n30109 , n30102 , n30107 );
or ( n30110 , n30105 , n30108 , n30109 );
xor ( n30111 , n29656 , n29660 );
xor ( n30112 , n30111 , n29665 );
and ( n30113 , n30110 , n30112 );
xor ( n30114 , n29821 , n29825 );
xor ( n30115 , n30114 , n29828 );
and ( n30116 , n30112 , n30115 );
and ( n30117 , n30110 , n30115 );
or ( n30118 , n30113 , n30116 , n30117 );
xor ( n30119 , n29613 , n29639 );
xor ( n30120 , n30119 , n29668 );
and ( n30121 , n30118 , n30120 );
xor ( n30122 , n29687 , n29739 );
xor ( n30123 , n30122 , n29742 );
and ( n30124 , n30120 , n30123 );
and ( n30125 , n30118 , n30123 );
or ( n30126 , n30121 , n30124 , n30125 );
xor ( n30127 , n29671 , n29745 );
xor ( n30128 , n30127 , n29764 );
and ( n30129 , n30126 , n30128 );
xor ( n30130 , n29581 , n29583 );
xor ( n30131 , n30130 , n29586 );
and ( n30132 , n30128 , n30131 );
and ( n30133 , n30126 , n30131 );
or ( n30134 , n30129 , n30132 , n30133 );
and ( n30135 , n30100 , n30134 );
xor ( n30136 , n29589 , n29591 );
xor ( n30137 , n30136 , n29594 );
and ( n30138 , n30134 , n30137 );
and ( n30139 , n30100 , n30137 );
or ( n30140 , n30135 , n30138 , n30139 );
xor ( n30141 , n29675 , n29679 );
xor ( n30142 , n30141 , n29684 );
xor ( n30143 , n29627 , n29631 );
xor ( n30144 , n30143 , n29636 );
and ( n30145 , n30142 , n30144 );
xor ( n30146 , n29703 , n29719 );
xor ( n30147 , n30146 , n29736 );
and ( n30148 , n30144 , n30147 );
and ( n30149 , n30142 , n30147 );
or ( n30150 , n30145 , n30148 , n30149 );
xor ( n30151 , n29831 , n29833 );
xor ( n30152 , n30151 , n29836 );
and ( n30153 , n30150 , n30152 );
xor ( n30154 , n29769 , n29771 );
xor ( n30155 , n30154 , n29774 );
and ( n30156 , n30152 , n30155 );
and ( n30157 , n30150 , n30155 );
or ( n30158 , n30153 , n30156 , n30157 );
xor ( n30159 , n29777 , n29779 );
xor ( n30160 , n30159 , n29782 );
and ( n30161 , n30158 , n30160 );
xor ( n30162 , n29839 , n29841 );
xor ( n30163 , n30162 , n29844 );
and ( n30164 , n30160 , n30163 );
and ( n30165 , n30158 , n30163 );
or ( n30166 , n30161 , n30164 , n30165 );
xor ( n30167 , n29767 , n29785 );
xor ( n30168 , n30167 , n29788 );
and ( n30169 , n30166 , n30168 );
xor ( n30170 , n29847 , n29849 );
xor ( n30171 , n30170 , n29852 );
and ( n30172 , n30168 , n30171 );
and ( n30173 , n30166 , n30171 );
or ( n30174 , n30169 , n30172 , n30173 );
and ( n30175 , n30140 , n30174 );
xor ( n30176 , n29597 , n29791 );
xor ( n30177 , n30176 , n29794 );
and ( n30178 , n30174 , n30177 );
and ( n30179 , n30140 , n30177 );
or ( n30180 , n30175 , n30178 , n30179 );
and ( n30181 , n29863 , n30180 );
xor ( n30182 , n29797 , n29799 );
xor ( n30183 , n30182 , n29802 );
and ( n30184 , n30180 , n30183 );
and ( n30185 , n29863 , n30183 );
or ( n30186 , n30181 , n30184 , n30185 );
and ( n30187 , n29817 , n30186 );
xor ( n30188 , n29817 , n30186 );
and ( n30189 , n20867 , n23944 );
and ( n30190 , n20803 , n23942 );
nor ( n30191 , n30189 , n30190 );
xnor ( n30192 , n30191 , n23550 );
and ( n30193 , n21218 , n23641 );
and ( n30194 , n21072 , n23639 );
nor ( n30195 , n30193 , n30194 );
xnor ( n30196 , n30195 , n23213 );
and ( n30197 , n30192 , n30196 );
and ( n30198 , n21451 , n23230 );
and ( n30199 , n21302 , n23228 );
nor ( n30200 , n30198 , n30199 );
xnor ( n30201 , n30200 , n22842 );
and ( n30202 , n30196 , n30201 );
and ( n30203 , n30192 , n30201 );
or ( n30204 , n30197 , n30202 , n30203 );
and ( n30205 , n20268 , n25383 );
and ( n30206 , n20182 , n25381 );
nor ( n30207 , n30205 , n30206 );
xnor ( n30208 , n30207 , n24885 );
and ( n30209 , n20452 , n24902 );
and ( n30210 , n20360 , n24900 );
nor ( n30211 , n30209 , n30210 );
xnor ( n30212 , n30211 , n24397 );
and ( n30213 , n30208 , n30212 );
and ( n30214 , n20666 , n24376 );
and ( n30215 , n20618 , n24374 );
nor ( n30216 , n30214 , n30215 );
xnor ( n30217 , n30216 , n23927 );
and ( n30218 , n30212 , n30217 );
and ( n30219 , n30208 , n30217 );
or ( n30220 , n30213 , n30218 , n30219 );
and ( n30221 , n30204 , n30220 );
xor ( n30222 , n29867 , n29871 );
xor ( n30223 , n30222 , n29876 );
and ( n30224 , n30220 , n30223 );
and ( n30225 , n30204 , n30223 );
or ( n30226 , n30221 , n30224 , n30225 );
xor ( n30227 , n29992 , n29995 );
and ( n30228 , n20080 , n26027 );
and ( n30229 , n20004 , n26025 );
nor ( n30230 , n30228 , n30229 );
xnor ( n30231 , n30230 , n25499 );
and ( n30232 , n30227 , n30231 );
and ( n30233 , n21955 , n22381 );
and ( n30234 , n21876 , n22379 );
nor ( n30235 , n30233 , n30234 );
xnor ( n30236 , n30235 , n22228 );
and ( n30237 , n30231 , n30236 );
and ( n30238 , n30227 , n30236 );
or ( n30239 , n30232 , n30237 , n30238 );
xor ( n30240 , n29644 , n29648 );
xor ( n30241 , n30240 , n29653 );
and ( n30242 , n30239 , n30241 );
xor ( n30243 , n29724 , n29728 );
xor ( n30244 , n30243 , n29733 );
and ( n30245 , n30241 , n30244 );
and ( n30246 , n30239 , n30244 );
or ( n30247 , n30242 , n30245 , n30246 );
and ( n30248 , n30226 , n30247 );
xor ( n30249 , n29748 , n29750 );
xor ( n30250 , n30249 , n29753 );
and ( n30251 , n30247 , n30250 );
and ( n30252 , n30226 , n30250 );
or ( n30253 , n30248 , n30251 , n30252 );
xor ( n30254 , n29756 , n29758 );
xor ( n30255 , n30254 , n29761 );
and ( n30256 , n30253 , n30255 );
xor ( n30257 , n29901 , n29951 );
xor ( n30258 , n30257 , n29954 );
and ( n30259 , n30255 , n30258 );
and ( n30260 , n30253 , n30258 );
or ( n30261 , n30256 , n30259 , n30260 );
and ( n30262 , n24527 , n20674 );
and ( n30263 , n24521 , n20672 );
nor ( n30264 , n30262 , n30263 );
xnor ( n30265 , n30264 , n20542 );
and ( n30266 , n24940 , n20460 );
and ( n30267 , n24621 , n20458 );
nor ( n30268 , n30266 , n30267 );
xnor ( n30269 , n30268 , n20337 );
and ( n30270 , n30265 , n30269 );
and ( n30271 , n25554 , n20276 );
and ( n30272 , n25284 , n20274 );
nor ( n30273 , n30271 , n30272 );
xnor ( n30274 , n30273 , n20175 );
and ( n30275 , n30269 , n30274 );
and ( n30276 , n30265 , n30274 );
or ( n30277 , n30270 , n30275 , n30276 );
and ( n30278 , n27751 , n19688 );
and ( n30279 , n27352 , n19686 );
nor ( n30280 , n30278 , n30279 );
xnor ( n30281 , n30280 , n19655 );
and ( n30282 , n28211 , n19596 );
and ( n30283 , n27757 , n19594 );
nor ( n30284 , n30282 , n30283 );
xnor ( n30285 , n30284 , n19545 );
and ( n30286 , n30281 , n30285 );
and ( n30287 , n28700 , n19518 );
and ( n30288 , n28810 , n19516 );
nor ( n30289 , n30287 , n30288 );
xnor ( n30290 , n30289 , n19489 );
and ( n30291 , n30285 , n30290 );
and ( n30292 , n30281 , n30290 );
or ( n30293 , n30286 , n30291 , n30292 );
and ( n30294 , n30277 , n30293 );
and ( n30295 , n25974 , n20114 );
and ( n30296 , n25765 , n20112 );
nor ( n30297 , n30295 , n30296 );
xnor ( n30298 , n30297 , n19997 );
and ( n30299 , n26422 , n19894 );
and ( n30300 , n26319 , n19892 );
nor ( n30301 , n30299 , n30300 );
xnor ( n30302 , n30301 , n19858 );
and ( n30303 , n30298 , n30302 );
and ( n30304 , n27135 , n19805 );
and ( n30305 , n26851 , n19803 );
nor ( n30306 , n30304 , n30305 );
xnor ( n30307 , n30306 , n19750 );
and ( n30308 , n30302 , n30307 );
and ( n30309 , n30298 , n30307 );
or ( n30310 , n30303 , n30308 , n30309 );
and ( n30311 , n30293 , n30310 );
and ( n30312 , n30277 , n30310 );
or ( n30313 , n30294 , n30311 , n30312 );
and ( n30314 , n22425 , n22048 );
and ( n30315 , n22198 , n22046 );
nor ( n30316 , n30314 , n30315 );
xnor ( n30317 , n30316 , n21853 );
and ( n30318 , n22916 , n21741 );
and ( n30319 , n22756 , n21739 );
nor ( n30320 , n30318 , n30319 );
xnor ( n30321 , n30320 , n21605 );
and ( n30322 , n30317 , n30321 );
and ( n30323 , n30321 , n29993 );
and ( n30324 , n30317 , n29993 );
or ( n30325 , n30322 , n30323 , n30324 );
and ( n30326 , n23271 , n21468 );
and ( n30327 , n23141 , n21466 );
nor ( n30328 , n30326 , n30327 );
xnor ( n30329 , n30328 , n21331 );
and ( n30330 , n23573 , n21155 );
and ( n30331 , n23381 , n21153 );
nor ( n30332 , n30330 , n30331 );
xnor ( n30333 , n30332 , n20994 );
and ( n30334 , n30329 , n30333 );
and ( n30335 , n24131 , n20955 );
and ( n30336 , n23968 , n20953 );
nor ( n30337 , n30335 , n30336 );
xnor ( n30338 , n30337 , n20780 );
and ( n30339 , n30333 , n30338 );
and ( n30340 , n30329 , n30338 );
or ( n30341 , n30334 , n30339 , n30340 );
and ( n30342 , n30325 , n30341 );
and ( n30343 , n19469 , n29276 );
and ( n30344 , n19434 , n29274 );
nor ( n30345 , n30343 , n30344 );
xnor ( n30346 , n30345 , n28677 );
and ( n30347 , n30341 , n30346 );
and ( n30348 , n30325 , n30346 );
or ( n30349 , n30342 , n30347 , n30348 );
and ( n30350 , n30313 , n30349 );
xor ( n30351 , n29883 , n29887 );
xor ( n30352 , n30351 , n29892 );
and ( n30353 , n30349 , n30352 );
and ( n30354 , n30313 , n30352 );
or ( n30355 , n30350 , n30353 , n30354 );
xor ( n30356 , n29879 , n29895 );
xor ( n30357 , n30356 , n29898 );
and ( n30358 , n30355 , n30357 );
xor ( n30359 , n29988 , n30008 );
xor ( n30360 , n30359 , n30011 );
and ( n30361 , n30357 , n30360 );
and ( n30362 , n30355 , n30360 );
or ( n30363 , n30358 , n30361 , n30362 );
and ( n30364 , n19510 , n28628 );
and ( n30365 , n19496 , n28626 );
nor ( n30366 , n30364 , n30365 );
xnor ( n30367 , n30366 , n28096 );
and ( n30368 , n19721 , n27529 );
and ( n30369 , n19637 , n27527 );
nor ( n30370 , n30368 , n30369 );
xnor ( n30371 , n30370 , n27034 );
and ( n30372 , n30367 , n30371 );
and ( n30373 , n19825 , n26992 );
and ( n30374 , n19811 , n26990 );
nor ( n30375 , n30373 , n30374 );
xnor ( n30376 , n30375 , n26369 );
and ( n30377 , n30371 , n30376 );
and ( n30378 , n30367 , n30376 );
or ( n30379 , n30372 , n30377 , n30378 );
and ( n30380 , n19418 , n29977 );
and ( n30381 , n19426 , n29974 );
nor ( n30382 , n30380 , n30381 );
xnor ( n30383 , n30382 , n28674 );
and ( n30384 , n19605 , n28062 );
and ( n30385 , n19588 , n28060 );
nor ( n30386 , n30384 , n30385 );
xnor ( n30387 , n30386 , n27549 );
and ( n30388 , n30383 , n30387 );
and ( n30389 , n21704 , n22859 );
and ( n30390 , n21612 , n22857 );
nor ( n30391 , n30389 , n30390 );
xnor ( n30392 , n30391 , n22418 );
and ( n30393 , n30387 , n30392 );
and ( n30394 , n30383 , n30392 );
or ( n30395 , n30388 , n30393 , n30394 );
and ( n30396 , n30379 , n30395 );
xor ( n30397 , n29905 , n29909 );
xor ( n30398 , n30397 , n29914 );
and ( n30399 , n30395 , n30398 );
and ( n30400 , n30379 , n30398 );
or ( n30401 , n30396 , n30399 , n30400 );
and ( n30402 , n22198 , n22381 );
and ( n30403 , n22235 , n22379 );
nor ( n30404 , n30402 , n30403 );
xnor ( n30405 , n30404 , n22228 );
and ( n30406 , n29623 , n19457 );
not ( n30407 , n30406 );
and ( n30408 , n30407 , n19416 );
and ( n30409 , n30405 , n30408 );
and ( n30410 , n22235 , n22381 );
and ( n30411 , n21955 , n22379 );
nor ( n30412 , n30410 , n30411 );
xnor ( n30413 , n30412 , n22228 );
and ( n30414 , n30409 , n30413 );
and ( n30415 , n29318 , n19459 );
and ( n30416 , n29078 , n19457 );
nor ( n30417 , n30415 , n30416 );
xnor ( n30418 , n30417 , n19416 );
and ( n30419 , n30413 , n30418 );
and ( n30420 , n30409 , n30418 );
or ( n30421 , n30414 , n30419 , n30420 );
and ( n30422 , n19946 , n26349 );
and ( n30423 , n19881 , n26347 );
nor ( n30424 , n30422 , n30423 );
xnor ( n30425 , n30424 , n25893 );
and ( n30426 , n30421 , n30425 );
xor ( n30427 , n29921 , n29925 );
xor ( n30428 , n30427 , n29930 );
and ( n30429 , n30425 , n30428 );
and ( n30430 , n30421 , n30428 );
or ( n30431 , n30426 , n30429 , n30430 );
xor ( n30432 , n30018 , n30022 );
xor ( n30433 , n30432 , n30027 );
and ( n30434 , n30431 , n30433 );
xor ( n30435 , n29996 , n30000 );
xor ( n30436 , n30435 , n30005 );
and ( n30437 , n30433 , n30436 );
and ( n30438 , n30431 , n30436 );
or ( n30439 , n30434 , n30437 , n30438 );
and ( n30440 , n30401 , n30439 );
xor ( n30441 , n30030 , n30082 );
xor ( n30442 , n30441 , n30085 );
and ( n30443 , n30439 , n30442 );
and ( n30444 , n30401 , n30442 );
or ( n30445 , n30440 , n30443 , n30444 );
and ( n30446 , n30363 , n30445 );
xor ( n30447 , n30014 , n30088 );
xor ( n30448 , n30447 , n30091 );
and ( n30449 , n30445 , n30448 );
and ( n30450 , n30363 , n30448 );
or ( n30451 , n30446 , n30449 , n30450 );
and ( n30452 , n30261 , n30451 );
xor ( n30453 , n29957 , n30094 );
xor ( n30454 , n30453 , n30097 );
and ( n30455 , n30451 , n30454 );
and ( n30456 , n30261 , n30454 );
or ( n30457 , n30452 , n30455 , n30456 );
xor ( n30458 , n30034 , n30038 );
xor ( n30459 , n30458 , n30043 );
xor ( n30460 , n29961 , n29965 );
xor ( n30461 , n30460 , n29970 );
and ( n30462 , n30459 , n30461 );
xor ( n30463 , n30050 , n30054 );
xor ( n30464 , n30463 , n30059 );
and ( n30465 , n30461 , n30464 );
and ( n30466 , n30459 , n30464 );
or ( n30467 , n30462 , n30465 , n30466 );
xor ( n30468 , n30046 , n30062 );
xor ( n30469 , n30468 , n30079 );
and ( n30470 , n30467 , n30469 );
xor ( n30471 , n29933 , n29937 );
xor ( n30472 , n30471 , n29942 );
and ( n30473 , n30469 , n30472 );
and ( n30474 , n30467 , n30472 );
or ( n30475 , n30470 , n30473 , n30474 );
xor ( n30476 , n29973 , n29980 );
xor ( n30477 , n30476 , n29985 );
xor ( n30478 , n30102 , n30104 );
xor ( n30479 , n30478 , n30107 );
and ( n30480 , n30477 , n30479 );
xor ( n30481 , n30239 , n30241 );
xor ( n30482 , n30481 , n30244 );
and ( n30483 , n30479 , n30482 );
and ( n30484 , n30477 , n30482 );
or ( n30485 , n30480 , n30483 , n30484 );
and ( n30486 , n30475 , n30485 );
xor ( n30487 , n29917 , n29945 );
xor ( n30488 , n30487 , n29948 );
and ( n30489 , n30485 , n30488 );
and ( n30490 , n30475 , n30488 );
or ( n30491 , n30486 , n30489 , n30490 );
xor ( n30492 , n30118 , n30120 );
xor ( n30493 , n30492 , n30123 );
and ( n30494 , n30491 , n30493 );
xor ( n30495 , n30150 , n30152 );
xor ( n30496 , n30495 , n30155 );
and ( n30497 , n30493 , n30496 );
and ( n30498 , n30491 , n30496 );
or ( n30499 , n30494 , n30497 , n30498 );
xor ( n30500 , n30126 , n30128 );
xor ( n30501 , n30500 , n30131 );
and ( n30502 , n30499 , n30501 );
xor ( n30503 , n30158 , n30160 );
xor ( n30504 , n30503 , n30163 );
and ( n30505 , n30501 , n30504 );
and ( n30506 , n30499 , n30504 );
or ( n30507 , n30502 , n30505 , n30506 );
and ( n30508 , n30457 , n30507 );
xor ( n30509 , n30100 , n30134 );
xor ( n30510 , n30509 , n30137 );
and ( n30511 , n30507 , n30510 );
and ( n30512 , n30457 , n30510 );
or ( n30513 , n30508 , n30511 , n30512 );
xor ( n30514 , n29855 , n29857 );
xor ( n30515 , n30514 , n29860 );
and ( n30516 , n30513 , n30515 );
xor ( n30517 , n30140 , n30174 );
xor ( n30518 , n30517 , n30177 );
and ( n30519 , n30515 , n30518 );
and ( n30520 , n30513 , n30518 );
or ( n30521 , n30516 , n30519 , n30520 );
xor ( n30522 , n29863 , n30180 );
xor ( n30523 , n30522 , n30183 );
and ( n30524 , n30521 , n30523 );
xor ( n30525 , n30521 , n30523 );
xor ( n30526 , n30513 , n30515 );
xor ( n30527 , n30526 , n30518 );
and ( n30528 , n20182 , n26027 );
and ( n30529 , n20080 , n26025 );
nor ( n30530 , n30528 , n30529 );
xnor ( n30531 , n30530 , n25499 );
and ( n30532 , n20360 , n25383 );
and ( n30533 , n20268 , n25381 );
nor ( n30534 , n30532 , n30533 );
xnor ( n30535 , n30534 , n24885 );
and ( n30536 , n30531 , n30535 );
and ( n30537 , n20618 , n24902 );
and ( n30538 , n20452 , n24900 );
nor ( n30539 , n30537 , n30538 );
xnor ( n30540 , n30539 , n24397 );
and ( n30541 , n30535 , n30540 );
and ( n30542 , n30531 , n30540 );
or ( n30543 , n30536 , n30541 , n30542 );
and ( n30544 , n20803 , n24376 );
and ( n30545 , n20666 , n24374 );
nor ( n30546 , n30544 , n30545 );
xnor ( n30547 , n30546 , n23927 );
and ( n30548 , n21072 , n23944 );
and ( n30549 , n20867 , n23942 );
nor ( n30550 , n30548 , n30549 );
xnor ( n30551 , n30550 , n23550 );
and ( n30552 , n30547 , n30551 );
and ( n30553 , n21302 , n23641 );
and ( n30554 , n21218 , n23639 );
nor ( n30555 , n30553 , n30554 );
xnor ( n30556 , n30555 , n23213 );
and ( n30557 , n30551 , n30556 );
and ( n30558 , n30547 , n30556 );
or ( n30559 , n30552 , n30557 , n30558 );
and ( n30560 , n30543 , n30559 );
xor ( n30561 , n30067 , n30071 );
xor ( n30562 , n30561 , n30076 );
and ( n30563 , n30559 , n30562 );
and ( n30564 , n30543 , n30562 );
or ( n30565 , n30560 , n30563 , n30564 );
and ( n30566 , n26851 , n19894 );
and ( n30567 , n26422 , n19892 );
nor ( n30568 , n30566 , n30567 );
xnor ( n30569 , n30568 , n19858 );
and ( n30570 , n27352 , n19805 );
and ( n30571 , n27135 , n19803 );
nor ( n30572 , n30570 , n30571 );
xnor ( n30573 , n30572 , n19750 );
and ( n30574 , n30569 , n30573 );
and ( n30575 , n27757 , n19688 );
and ( n30576 , n27751 , n19686 );
nor ( n30577 , n30575 , n30576 );
xnor ( n30578 , n30577 , n19655 );
and ( n30579 , n30573 , n30578 );
and ( n30580 , n30569 , n30578 );
or ( n30581 , n30574 , n30579 , n30580 );
and ( n30582 , n25284 , n20460 );
and ( n30583 , n24940 , n20458 );
nor ( n30584 , n30582 , n30583 );
xnor ( n30585 , n30584 , n20337 );
and ( n30586 , n25765 , n20276 );
and ( n30587 , n25554 , n20274 );
nor ( n30588 , n30586 , n30587 );
xnor ( n30589 , n30588 , n20175 );
and ( n30590 , n30585 , n30589 );
and ( n30591 , n26319 , n20114 );
and ( n30592 , n25974 , n20112 );
nor ( n30593 , n30591 , n30592 );
xnor ( n30594 , n30593 , n19997 );
and ( n30595 , n30589 , n30594 );
and ( n30596 , n30585 , n30594 );
or ( n30597 , n30590 , n30595 , n30596 );
and ( n30598 , n30581 , n30597 );
and ( n30599 , n19496 , n29276 );
and ( n30600 , n19469 , n29274 );
nor ( n30601 , n30599 , n30600 );
xnor ( n30602 , n30601 , n28677 );
and ( n30603 , n30597 , n30602 );
and ( n30604 , n30581 , n30602 );
or ( n30605 , n30598 , n30603 , n30604 );
xor ( n30606 , n30192 , n30196 );
xor ( n30607 , n30606 , n30201 );
and ( n30608 , n30605 , n30607 );
xor ( n30609 , n30227 , n30231 );
xor ( n30610 , n30609 , n30236 );
and ( n30611 , n30607 , n30610 );
and ( n30612 , n30605 , n30610 );
or ( n30613 , n30608 , n30611 , n30612 );
and ( n30614 , n30565 , n30613 );
xor ( n30615 , n30204 , n30220 );
xor ( n30616 , n30615 , n30223 );
and ( n30617 , n30613 , n30616 );
and ( n30618 , n30565 , n30616 );
or ( n30619 , n30614 , n30617 , n30618 );
xor ( n30620 , n30142 , n30144 );
xor ( n30621 , n30620 , n30147 );
and ( n30622 , n30619 , n30621 );
xor ( n30623 , n30110 , n30112 );
xor ( n30624 , n30623 , n30115 );
and ( n30625 , n30621 , n30624 );
and ( n30626 , n30619 , n30624 );
or ( n30627 , n30622 , n30625 , n30626 );
and ( n30628 , n19637 , n28062 );
and ( n30629 , n19605 , n28060 );
nor ( n30630 , n30628 , n30629 );
xnor ( n30631 , n30630 , n27549 );
and ( n30632 , n21612 , n23230 );
and ( n30633 , n21451 , n23228 );
nor ( n30634 , n30632 , n30633 );
xnor ( n30635 , n30634 , n22842 );
and ( n30636 , n30631 , n30635 );
and ( n30637 , n21876 , n22859 );
and ( n30638 , n21704 , n22857 );
nor ( n30639 , n30637 , n30638 );
xnor ( n30640 , n30639 , n22418 );
and ( n30641 , n30635 , n30640 );
and ( n30642 , n30631 , n30640 );
or ( n30643 , n30636 , n30641 , n30642 );
and ( n30644 , n28810 , n19596 );
and ( n30645 , n28211 , n19594 );
nor ( n30646 , n30644 , n30645 );
xnor ( n30647 , n30646 , n19545 );
and ( n30648 , n29078 , n19518 );
and ( n30649 , n28700 , n19516 );
nor ( n30650 , n30648 , n30649 );
xnor ( n30651 , n30650 , n19489 );
and ( n30652 , n30647 , n30651 );
and ( n30653 , n29623 , n19459 );
and ( n30654 , n29318 , n19457 );
nor ( n30655 , n30653 , n30654 );
xnor ( n30656 , n30655 , n19416 );
and ( n30657 , n30651 , n30656 );
and ( n30658 , n30647 , n30656 );
or ( n30659 , n30652 , n30657 , n30658 );
and ( n30660 , n19811 , n27529 );
and ( n30661 , n19721 , n27527 );
nor ( n30662 , n30660 , n30661 );
xnor ( n30663 , n30662 , n27034 );
and ( n30664 , n30659 , n30663 );
and ( n30665 , n19881 , n26992 );
and ( n30666 , n19825 , n26990 );
nor ( n30667 , n30665 , n30666 );
xnor ( n30668 , n30667 , n26369 );
and ( n30669 , n30663 , n30668 );
and ( n30670 , n30659 , n30668 );
or ( n30671 , n30664 , n30669 , n30670 );
and ( n30672 , n30643 , n30671 );
and ( n30673 , n22756 , n22048 );
and ( n30674 , n22425 , n22046 );
nor ( n30675 , n30673 , n30674 );
xnor ( n30676 , n30675 , n21853 );
and ( n30677 , n23141 , n21741 );
and ( n30678 , n22916 , n21739 );
nor ( n30679 , n30677 , n30678 );
xnor ( n30680 , n30679 , n21605 );
and ( n30681 , n30676 , n30680 );
and ( n30682 , n23381 , n21468 );
and ( n30683 , n23271 , n21466 );
nor ( n30684 , n30682 , n30683 );
xnor ( n30685 , n30684 , n21331 );
and ( n30686 , n30680 , n30685 );
and ( n30687 , n30676 , n30685 );
or ( n30688 , n30681 , n30686 , n30687 );
and ( n30689 , n23968 , n21155 );
and ( n30690 , n23573 , n21153 );
nor ( n30691 , n30689 , n30690 );
xnor ( n30692 , n30691 , n20994 );
and ( n30693 , n24521 , n20955 );
and ( n30694 , n24131 , n20953 );
nor ( n30695 , n30693 , n30694 );
xnor ( n30696 , n30695 , n20780 );
and ( n30697 , n30692 , n30696 );
and ( n30698 , n24621 , n20674 );
and ( n30699 , n24527 , n20672 );
nor ( n30700 , n30698 , n30699 );
xnor ( n30701 , n30700 , n20542 );
and ( n30702 , n30696 , n30701 );
and ( n30703 , n30692 , n30701 );
or ( n30704 , n30697 , n30702 , n30703 );
and ( n30705 , n30688 , n30704 );
and ( n30706 , n19434 , n29977 );
and ( n30707 , n19418 , n29974 );
nor ( n30708 , n30706 , n30707 );
xnor ( n30709 , n30708 , n28674 );
and ( n30710 , n30704 , n30709 );
and ( n30711 , n30688 , n30709 );
or ( n30712 , n30705 , n30710 , n30711 );
and ( n30713 , n30671 , n30712 );
and ( n30714 , n30643 , n30712 );
or ( n30715 , n30672 , n30713 , n30714 );
and ( n30716 , n19588 , n28628 );
and ( n30717 , n19510 , n28626 );
nor ( n30718 , n30716 , n30717 );
xnor ( n30719 , n30718 , n28096 );
and ( n30720 , n20004 , n26349 );
and ( n30721 , n19946 , n26347 );
nor ( n30722 , n30720 , n30721 );
xnor ( n30723 , n30722 , n25893 );
and ( n30724 , n30719 , n30723 );
xor ( n30725 , n30329 , n30333 );
xor ( n30726 , n30725 , n30338 );
and ( n30727 , n30723 , n30726 );
and ( n30728 , n30719 , n30726 );
or ( n30729 , n30724 , n30727 , n30728 );
xor ( n30730 , n30208 , n30212 );
xor ( n30731 , n30730 , n30217 );
and ( n30732 , n30729 , n30731 );
xor ( n30733 , n30383 , n30387 );
xor ( n30734 , n30733 , n30392 );
and ( n30735 , n30731 , n30734 );
and ( n30736 , n30729 , n30734 );
or ( n30737 , n30732 , n30735 , n30736 );
and ( n30738 , n30715 , n30737 );
xor ( n30739 , n30379 , n30395 );
xor ( n30740 , n30739 , n30398 );
and ( n30741 , n30737 , n30740 );
and ( n30742 , n30715 , n30740 );
or ( n30743 , n30738 , n30741 , n30742 );
xor ( n30744 , n30226 , n30247 );
xor ( n30745 , n30744 , n30250 );
and ( n30746 , n30743 , n30745 );
xor ( n30747 , n30355 , n30357 );
xor ( n30748 , n30747 , n30360 );
and ( n30749 , n30745 , n30748 );
and ( n30750 , n30743 , n30748 );
or ( n30751 , n30746 , n30749 , n30750 );
and ( n30752 , n30627 , n30751 );
xor ( n30753 , n30253 , n30255 );
xor ( n30754 , n30753 , n30258 );
and ( n30755 , n30751 , n30754 );
and ( n30756 , n30627 , n30754 );
or ( n30757 , n30752 , n30755 , n30756 );
xor ( n30758 , n30261 , n30451 );
xor ( n30759 , n30758 , n30454 );
and ( n30760 , n30757 , n30759 );
xor ( n30761 , n30499 , n30501 );
xor ( n30762 , n30761 , n30504 );
and ( n30763 , n30759 , n30762 );
and ( n30764 , n30757 , n30762 );
or ( n30765 , n30760 , n30763 , n30764 );
xor ( n30766 , n30166 , n30168 );
xor ( n30767 , n30766 , n30171 );
and ( n30768 , n30765 , n30767 );
xor ( n30769 , n30457 , n30507 );
xor ( n30770 , n30769 , n30510 );
and ( n30771 , n30767 , n30770 );
and ( n30772 , n30765 , n30770 );
or ( n30773 , n30768 , n30771 , n30772 );
and ( n30774 , n30527 , n30773 );
xor ( n30775 , n30527 , n30773 );
xor ( n30776 , n30765 , n30767 );
xor ( n30777 , n30776 , n30770 );
xor ( n30778 , n30367 , n30371 );
xor ( n30779 , n30778 , n30376 );
xor ( n30780 , n30277 , n30293 );
xor ( n30781 , n30780 , n30310 );
and ( n30782 , n30779 , n30781 );
xor ( n30783 , n30325 , n30341 );
xor ( n30784 , n30783 , n30346 );
and ( n30785 , n30781 , n30784 );
and ( n30786 , n30779 , n30784 );
or ( n30787 , n30782 , n30785 , n30786 );
xor ( n30788 , n30317 , n30321 );
xor ( n30789 , n30788 , n29993 );
xor ( n30790 , n30265 , n30269 );
xor ( n30791 , n30790 , n30274 );
and ( n30792 , n30789 , n30791 );
xor ( n30793 , n30281 , n30285 );
xor ( n30794 , n30793 , n30290 );
and ( n30795 , n30791 , n30794 );
and ( n30796 , n30789 , n30794 );
or ( n30797 , n30792 , n30795 , n30796 );
xor ( n30798 , n30459 , n30461 );
xor ( n30799 , n30798 , n30464 );
and ( n30800 , n30797 , n30799 );
xor ( n30801 , n30421 , n30425 );
xor ( n30802 , n30801 , n30428 );
and ( n30803 , n30799 , n30802 );
and ( n30804 , n30797 , n30802 );
or ( n30805 , n30800 , n30803 , n30804 );
and ( n30806 , n30787 , n30805 );
xor ( n30807 , n30313 , n30349 );
xor ( n30808 , n30807 , n30352 );
and ( n30809 , n30805 , n30808 );
and ( n30810 , n30787 , n30808 );
or ( n30811 , n30806 , n30809 , n30810 );
xor ( n30812 , n30401 , n30439 );
xor ( n30813 , n30812 , n30442 );
and ( n30814 , n30811 , n30813 );
xor ( n30815 , n30475 , n30485 );
xor ( n30816 , n30815 , n30488 );
and ( n30817 , n30813 , n30816 );
and ( n30818 , n30811 , n30816 );
or ( n30819 , n30814 , n30817 , n30818 );
xor ( n30820 , n30363 , n30445 );
xor ( n30821 , n30820 , n30448 );
and ( n30822 , n30819 , n30821 );
xor ( n30823 , n30491 , n30493 );
xor ( n30824 , n30823 , n30496 );
and ( n30825 , n30821 , n30824 );
and ( n30826 , n30819 , n30824 );
or ( n30827 , n30822 , n30825 , n30826 );
and ( n30828 , n22235 , n22859 );
and ( n30829 , n21955 , n22857 );
nor ( n30830 , n30828 , n30829 );
xnor ( n30831 , n30830 , n22418 );
and ( n30832 , n28211 , n19688 );
and ( n30833 , n27757 , n19686 );
nor ( n30834 , n30832 , n30833 );
xnor ( n30835 , n30834 , n19655 );
and ( n30836 , n30831 , n30835 );
and ( n30837 , n29318 , n19518 );
and ( n30838 , n29078 , n19516 );
nor ( n30839 , n30837 , n30838 );
xnor ( n30840 , n30839 , n19489 );
and ( n30841 , n30835 , n30840 );
and ( n30842 , n30831 , n30840 );
or ( n30843 , n30836 , n30841 , n30842 );
xor ( n30844 , n30676 , n30680 );
xor ( n30845 , n30844 , n30685 );
and ( n30846 , n30843 , n30845 );
xor ( n30847 , n30647 , n30651 );
xor ( n30848 , n30847 , n30656 );
and ( n30849 , n30845 , n30848 );
and ( n30850 , n30843 , n30848 );
or ( n30851 , n30846 , n30849 , n30850 );
xor ( n30852 , n30692 , n30696 );
xor ( n30853 , n30852 , n30701 );
xor ( n30854 , n30569 , n30573 );
xor ( n30855 , n30854 , n30578 );
and ( n30856 , n30853 , n30855 );
xor ( n30857 , n30585 , n30589 );
xor ( n30858 , n30857 , n30594 );
and ( n30859 , n30855 , n30858 );
and ( n30860 , n30853 , n30858 );
or ( n30861 , n30856 , n30859 , n30860 );
and ( n30862 , n30851 , n30861 );
xor ( n30863 , n30659 , n30663 );
xor ( n30864 , n30863 , n30668 );
and ( n30865 , n30861 , n30864 );
and ( n30866 , n30851 , n30864 );
or ( n30867 , n30862 , n30865 , n30866 );
xor ( n30868 , n30581 , n30597 );
xor ( n30869 , n30868 , n30602 );
xor ( n30870 , n30688 , n30704 );
xor ( n30871 , n30870 , n30709 );
and ( n30872 , n30869 , n30871 );
xor ( n30873 , n30719 , n30723 );
xor ( n30874 , n30873 , n30726 );
and ( n30875 , n30871 , n30874 );
and ( n30876 , n30869 , n30874 );
or ( n30877 , n30872 , n30875 , n30876 );
and ( n30878 , n30867 , n30877 );
xor ( n30879 , n30643 , n30671 );
xor ( n30880 , n30879 , n30712 );
and ( n30881 , n30877 , n30880 );
and ( n30882 , n30867 , n30880 );
or ( n30883 , n30878 , n30881 , n30882 );
and ( n30884 , n20080 , n26349 );
and ( n30885 , n20004 , n26347 );
nor ( n30886 , n30884 , n30885 );
xnor ( n30887 , n30886 , n25893 );
and ( n30888 , n20452 , n25383 );
and ( n30889 , n20360 , n25381 );
nor ( n30890 , n30888 , n30889 );
xnor ( n30891 , n30890 , n24885 );
and ( n30892 , n30887 , n30891 );
and ( n30893 , n20666 , n24902 );
and ( n30894 , n20618 , n24900 );
nor ( n30895 , n30893 , n30894 );
xnor ( n30896 , n30895 , n24397 );
and ( n30897 , n30891 , n30896 );
and ( n30898 , n30887 , n30896 );
or ( n30899 , n30892 , n30897 , n30898 );
xor ( n30900 , n30405 , n30408 );
and ( n30901 , n20268 , n26027 );
and ( n30902 , n20182 , n26025 );
nor ( n30903 , n30901 , n30902 );
xnor ( n30904 , n30903 , n25499 );
and ( n30905 , n30900 , n30904 );
and ( n30906 , n21955 , n22859 );
and ( n30907 , n21876 , n22857 );
nor ( n30908 , n30906 , n30907 );
xnor ( n30909 , n30908 , n22418 );
and ( n30910 , n30904 , n30909 );
and ( n30911 , n30900 , n30909 );
or ( n30912 , n30905 , n30910 , n30911 );
and ( n30913 , n30899 , n30912 );
xor ( n30914 , n30298 , n30302 );
xor ( n30915 , n30914 , n30307 );
and ( n30916 , n30912 , n30915 );
and ( n30917 , n30899 , n30915 );
or ( n30918 , n30913 , n30916 , n30917 );
and ( n30919 , n25974 , n20276 );
and ( n30920 , n25765 , n20274 );
nor ( n30921 , n30919 , n30920 );
xnor ( n30922 , n30921 , n20175 );
and ( n30923 , n27751 , n19805 );
and ( n30924 , n27352 , n19803 );
nor ( n30925 , n30923 , n30924 );
xnor ( n30926 , n30925 , n19750 );
and ( n30927 , n30922 , n30926 );
and ( n30928 , n28700 , n19596 );
and ( n30929 , n28810 , n19594 );
nor ( n30930 , n30928 , n30929 );
xnor ( n30931 , n30930 , n19545 );
and ( n30932 , n30926 , n30931 );
and ( n30933 , n30922 , n30931 );
or ( n30934 , n30927 , n30932 , n30933 );
and ( n30935 , n25554 , n20460 );
and ( n30936 , n25284 , n20458 );
nor ( n30937 , n30935 , n30936 );
xnor ( n30938 , n30937 , n20337 );
and ( n30939 , n26422 , n20114 );
and ( n30940 , n26319 , n20112 );
nor ( n30941 , n30939 , n30940 );
xnor ( n30942 , n30941 , n19997 );
and ( n30943 , n30938 , n30942 );
and ( n30944 , n27135 , n19894 );
and ( n30945 , n26851 , n19892 );
nor ( n30946 , n30944 , n30945 );
xnor ( n30947 , n30946 , n19858 );
and ( n30948 , n30942 , n30947 );
and ( n30949 , n30938 , n30947 );
or ( n30950 , n30943 , n30948 , n30949 );
and ( n30951 , n30934 , n30950 );
and ( n30952 , n19825 , n27529 );
and ( n30953 , n19811 , n27527 );
nor ( n30954 , n30952 , n30953 );
xnor ( n30955 , n30954 , n27034 );
and ( n30956 , n30950 , n30955 );
and ( n30957 , n30934 , n30955 );
or ( n30958 , n30951 , n30956 , n30957 );
xor ( n30959 , n30531 , n30535 );
xor ( n30960 , n30959 , n30540 );
and ( n30961 , n30958 , n30960 );
xor ( n30962 , n30547 , n30551 );
xor ( n30963 , n30962 , n30556 );
and ( n30964 , n30960 , n30963 );
and ( n30965 , n30958 , n30963 );
or ( n30966 , n30961 , n30964 , n30965 );
and ( n30967 , n30918 , n30966 );
xor ( n30968 , n30543 , n30559 );
xor ( n30969 , n30968 , n30562 );
and ( n30970 , n30966 , n30969 );
and ( n30971 , n30918 , n30969 );
or ( n30972 , n30967 , n30970 , n30971 );
and ( n30973 , n30883 , n30972 );
and ( n30974 , n19469 , n29977 );
and ( n30975 , n19434 , n29974 );
nor ( n30976 , n30974 , n30975 );
xnor ( n30977 , n30976 , n28674 );
and ( n30978 , n19605 , n28628 );
and ( n30979 , n19588 , n28626 );
nor ( n30980 , n30978 , n30979 );
xnor ( n30981 , n30980 , n28096 );
and ( n30982 , n30977 , n30981 );
and ( n30983 , n19946 , n26992 );
and ( n30984 , n19881 , n26990 );
nor ( n30985 , n30983 , n30984 );
xnor ( n30986 , n30985 , n26369 );
and ( n30987 , n30981 , n30986 );
and ( n30988 , n30977 , n30986 );
or ( n30989 , n30982 , n30987 , n30988 );
and ( n30990 , n20867 , n24376 );
and ( n30991 , n20803 , n24374 );
nor ( n30992 , n30990 , n30991 );
xnor ( n30993 , n30992 , n23927 );
and ( n30994 , n21218 , n23944 );
and ( n30995 , n21072 , n23942 );
nor ( n30996 , n30994 , n30995 );
xnor ( n30997 , n30996 , n23550 );
and ( n30998 , n30993 , n30997 );
and ( n30999 , n21451 , n23641 );
and ( n31000 , n21302 , n23639 );
nor ( n31001 , n30999 , n31000 );
xnor ( n31002 , n31001 , n23213 );
and ( n31003 , n30997 , n31002 );
and ( n31004 , n30993 , n31002 );
or ( n31005 , n30998 , n31003 , n31004 );
and ( n31006 , n30989 , n31005 );
xor ( n31007 , n30409 , n30413 );
xor ( n31008 , n31007 , n30418 );
and ( n31009 , n31005 , n31008 );
and ( n31010 , n30989 , n31008 );
or ( n31011 , n31006 , n31009 , n31010 );
and ( n31012 , n22425 , n22381 );
and ( n31013 , n22198 , n22379 );
nor ( n31014 , n31012 , n31013 );
xnor ( n31015 , n31014 , n22228 );
and ( n31016 , n22916 , n22048 );
and ( n31017 , n22756 , n22046 );
nor ( n31018 , n31016 , n31017 );
xnor ( n31019 , n31018 , n21853 );
and ( n31020 , n31015 , n31019 );
and ( n31021 , n31019 , n30406 );
and ( n31022 , n31015 , n30406 );
or ( n31023 , n31020 , n31021 , n31022 );
and ( n31024 , n19721 , n28062 );
and ( n31025 , n19637 , n28060 );
nor ( n31026 , n31024 , n31025 );
xnor ( n31027 , n31026 , n27549 );
and ( n31028 , n31023 , n31027 );
and ( n31029 , n21704 , n23230 );
and ( n31030 , n21612 , n23228 );
nor ( n31031 , n31029 , n31030 );
xnor ( n31032 , n31031 , n22842 );
and ( n31033 , n31027 , n31032 );
and ( n31034 , n31023 , n31032 );
or ( n31035 , n31028 , n31033 , n31034 );
and ( n31036 , n24131 , n21155 );
and ( n31037 , n23968 , n21153 );
nor ( n31038 , n31036 , n31037 );
xnor ( n31039 , n31038 , n20994 );
and ( n31040 , n24527 , n20955 );
and ( n31041 , n24521 , n20953 );
nor ( n31042 , n31040 , n31041 );
xnor ( n31043 , n31042 , n20780 );
and ( n31044 , n31039 , n31043 );
and ( n31045 , n24940 , n20674 );
and ( n31046 , n24621 , n20672 );
nor ( n31047 , n31045 , n31046 );
xnor ( n31048 , n31047 , n20542 );
and ( n31049 , n31043 , n31048 );
and ( n31050 , n31039 , n31048 );
or ( n31051 , n31044 , n31049 , n31050 );
and ( n31052 , n22756 , n22381 );
and ( n31053 , n22425 , n22379 );
nor ( n31054 , n31052 , n31053 );
xnor ( n31055 , n31054 , n22228 );
and ( n31056 , n29623 , n19516 );
not ( n31057 , n31056 );
and ( n31058 , n31057 , n19489 );
and ( n31059 , n31055 , n31058 );
and ( n31060 , n23271 , n21741 );
and ( n31061 , n23141 , n21739 );
nor ( n31062 , n31060 , n31061 );
xnor ( n31063 , n31062 , n21605 );
and ( n31064 , n31059 , n31063 );
and ( n31065 , n23573 , n21468 );
and ( n31066 , n23381 , n21466 );
nor ( n31067 , n31065 , n31066 );
xnor ( n31068 , n31067 , n21331 );
and ( n31069 , n31063 , n31068 );
and ( n31070 , n31059 , n31068 );
or ( n31071 , n31064 , n31069 , n31070 );
and ( n31072 , n31051 , n31071 );
and ( n31073 , n19510 , n29276 );
and ( n31074 , n19496 , n29274 );
nor ( n31075 , n31073 , n31074 );
xnor ( n31076 , n31075 , n28677 );
and ( n31077 , n31071 , n31076 );
and ( n31078 , n31051 , n31076 );
or ( n31079 , n31072 , n31077 , n31078 );
and ( n31080 , n31035 , n31079 );
xor ( n31081 , n30631 , n30635 );
xor ( n31082 , n31081 , n30640 );
and ( n31083 , n31079 , n31082 );
and ( n31084 , n31035 , n31082 );
or ( n31085 , n31080 , n31083 , n31084 );
and ( n31086 , n31011 , n31085 );
xor ( n31087 , n30605 , n30607 );
xor ( n31088 , n31087 , n30610 );
and ( n31089 , n31085 , n31088 );
and ( n31090 , n31011 , n31088 );
or ( n31091 , n31086 , n31089 , n31090 );
and ( n31092 , n30972 , n31091 );
and ( n31093 , n30883 , n31091 );
or ( n31094 , n30973 , n31092 , n31093 );
xor ( n31095 , n30467 , n30469 );
xor ( n31096 , n31095 , n30472 );
xor ( n31097 , n30431 , n30433 );
xor ( n31098 , n31097 , n30436 );
and ( n31099 , n31096 , n31098 );
xor ( n31100 , n30477 , n30479 );
xor ( n31101 , n31100 , n30482 );
and ( n31102 , n31098 , n31101 );
and ( n31103 , n31096 , n31101 );
or ( n31104 , n31099 , n31102 , n31103 );
and ( n31105 , n31094 , n31104 );
xor ( n31106 , n30619 , n30621 );
xor ( n31107 , n31106 , n30624 );
and ( n31108 , n31104 , n31107 );
and ( n31109 , n31094 , n31107 );
or ( n31110 , n31105 , n31108 , n31109 );
xor ( n31111 , n30565 , n30613 );
xor ( n31112 , n31111 , n30616 );
xor ( n31113 , n30715 , n30737 );
xor ( n31114 , n31113 , n30740 );
and ( n31115 , n31112 , n31114 );
xor ( n31116 , n30787 , n30805 );
xor ( n31117 , n31116 , n30808 );
and ( n31118 , n31114 , n31117 );
and ( n31119 , n31112 , n31117 );
or ( n31120 , n31115 , n31118 , n31119 );
xor ( n31121 , n30743 , n30745 );
xor ( n31122 , n31121 , n30748 );
and ( n31123 , n31120 , n31122 );
xor ( n31124 , n30811 , n30813 );
xor ( n31125 , n31124 , n30816 );
and ( n31126 , n31122 , n31125 );
and ( n31127 , n31120 , n31125 );
or ( n31128 , n31123 , n31126 , n31127 );
and ( n31129 , n31110 , n31128 );
xor ( n31130 , n30627 , n30751 );
xor ( n31131 , n31130 , n30754 );
and ( n31132 , n31128 , n31131 );
and ( n31133 , n31110 , n31131 );
or ( n31134 , n31129 , n31132 , n31133 );
and ( n31135 , n30827 , n31134 );
xor ( n31136 , n30757 , n30759 );
xor ( n31137 , n31136 , n30762 );
and ( n31138 , n31134 , n31137 );
and ( n31139 , n30827 , n31137 );
or ( n31140 , n31135 , n31138 , n31139 );
and ( n31141 , n30777 , n31140 );
xor ( n31142 , n30777 , n31140 );
xor ( n31143 , n30827 , n31134 );
xor ( n31144 , n31143 , n31137 );
xor ( n31145 , n31055 , n31058 );
and ( n31146 , n28810 , n19688 );
and ( n31147 , n28211 , n19686 );
nor ( n31148 , n31146 , n31147 );
xnor ( n31149 , n31148 , n19655 );
and ( n31150 , n31145 , n31149 );
and ( n31151 , n29078 , n19596 );
and ( n31152 , n28700 , n19594 );
nor ( n31153 , n31151 , n31152 );
xnor ( n31154 , n31153 , n19545 );
and ( n31155 , n31149 , n31154 );
and ( n31156 , n31145 , n31154 );
or ( n31157 , n31150 , n31155 , n31156 );
and ( n31158 , n19881 , n27529 );
and ( n31159 , n19825 , n27527 );
nor ( n31160 , n31158 , n31159 );
xnor ( n31161 , n31160 , n27034 );
and ( n31162 , n31157 , n31161 );
and ( n31163 , n20004 , n26992 );
and ( n31164 , n19946 , n26990 );
nor ( n31165 , n31163 , n31164 );
xnor ( n31166 , n31165 , n26369 );
and ( n31167 , n31161 , n31166 );
and ( n31168 , n31157 , n31166 );
or ( n31169 , n31162 , n31167 , n31168 );
xor ( n31170 , n30887 , n30891 );
xor ( n31171 , n31170 , n30896 );
and ( n31172 , n31169 , n31171 );
xor ( n31173 , n30900 , n30904 );
xor ( n31174 , n31173 , n30909 );
and ( n31175 , n31171 , n31174 );
and ( n31176 , n31169 , n31174 );
or ( n31177 , n31172 , n31175 , n31176 );
xor ( n31178 , n30789 , n30791 );
xor ( n31179 , n31178 , n30794 );
and ( n31180 , n31177 , n31179 );
xor ( n31181 , n30899 , n30912 );
xor ( n31182 , n31181 , n30915 );
and ( n31183 , n31179 , n31182 );
and ( n31184 , n31177 , n31182 );
or ( n31185 , n31180 , n31183 , n31184 );
xor ( n31186 , n30729 , n30731 );
xor ( n31187 , n31186 , n30734 );
and ( n31188 , n31185 , n31187 );
xor ( n31189 , n30779 , n30781 );
xor ( n31190 , n31189 , n30784 );
and ( n31191 , n31187 , n31190 );
and ( n31192 , n31185 , n31190 );
or ( n31193 , n31188 , n31191 , n31192 );
and ( n31194 , n20182 , n26349 );
and ( n31195 , n20080 , n26347 );
nor ( n31196 , n31194 , n31195 );
xnor ( n31197 , n31196 , n25893 );
and ( n31198 , n21072 , n24376 );
and ( n31199 , n20867 , n24374 );
nor ( n31200 , n31198 , n31199 );
xnor ( n31201 , n31200 , n23927 );
and ( n31202 , n31197 , n31201 );
and ( n31203 , n21612 , n23641 );
and ( n31204 , n21451 , n23639 );
nor ( n31205 , n31203 , n31204 );
xnor ( n31206 , n31205 , n23213 );
and ( n31207 , n31201 , n31206 );
and ( n31208 , n31197 , n31206 );
or ( n31209 , n31202 , n31207 , n31208 );
and ( n31210 , n20360 , n26027 );
and ( n31211 , n20268 , n26025 );
nor ( n31212 , n31210 , n31211 );
xnor ( n31213 , n31212 , n25499 );
and ( n31214 , n20618 , n25383 );
and ( n31215 , n20452 , n25381 );
nor ( n31216 , n31214 , n31215 );
xnor ( n31217 , n31216 , n24885 );
and ( n31218 , n31213 , n31217 );
and ( n31219 , n20803 , n24902 );
and ( n31220 , n20666 , n24900 );
nor ( n31221 , n31219 , n31220 );
xnor ( n31222 , n31221 , n24397 );
and ( n31223 , n31217 , n31222 );
and ( n31224 , n31213 , n31222 );
or ( n31225 , n31218 , n31223 , n31224 );
and ( n31226 , n31209 , n31225 );
and ( n31227 , n26319 , n20276 );
and ( n31228 , n25974 , n20274 );
nor ( n31229 , n31227 , n31228 );
xnor ( n31230 , n31229 , n20175 );
and ( n31231 , n27352 , n19894 );
and ( n31232 , n27135 , n19892 );
nor ( n31233 , n31231 , n31232 );
xnor ( n31234 , n31233 , n19858 );
and ( n31235 , n31230 , n31234 );
and ( n31236 , n27757 , n19805 );
and ( n31237 , n27751 , n19803 );
nor ( n31238 , n31236 , n31237 );
xnor ( n31239 , n31238 , n19750 );
and ( n31240 , n31234 , n31239 );
and ( n31241 , n31230 , n31239 );
or ( n31242 , n31235 , n31240 , n31241 );
and ( n31243 , n19588 , n29276 );
and ( n31244 , n19510 , n29274 );
nor ( n31245 , n31243 , n31244 );
xnor ( n31246 , n31245 , n28677 );
and ( n31247 , n31242 , n31246 );
xor ( n31248 , n31015 , n31019 );
xor ( n31249 , n31248 , n30406 );
and ( n31250 , n31246 , n31249 );
and ( n31251 , n31242 , n31249 );
or ( n31252 , n31247 , n31250 , n31251 );
and ( n31253 , n31225 , n31252 );
and ( n31254 , n31209 , n31252 );
or ( n31255 , n31226 , n31253 , n31254 );
and ( n31256 , n19811 , n28062 );
and ( n31257 , n19721 , n28060 );
nor ( n31258 , n31256 , n31257 );
xnor ( n31259 , n31258 , n27549 );
and ( n31260 , n21302 , n23944 );
and ( n31261 , n21218 , n23942 );
nor ( n31262 , n31260 , n31261 );
xnor ( n31263 , n31262 , n23550 );
and ( n31264 , n31259 , n31263 );
and ( n31265 , n21876 , n23230 );
and ( n31266 , n21704 , n23228 );
nor ( n31267 , n31265 , n31266 );
xnor ( n31268 , n31267 , n22842 );
and ( n31269 , n31263 , n31268 );
and ( n31270 , n31259 , n31268 );
or ( n31271 , n31264 , n31269 , n31270 );
and ( n31272 , n22198 , n22859 );
and ( n31273 , n22235 , n22857 );
nor ( n31274 , n31272 , n31273 );
xnor ( n31275 , n31274 , n22418 );
and ( n31276 , n23141 , n22048 );
and ( n31277 , n22916 , n22046 );
nor ( n31278 , n31276 , n31277 );
xnor ( n31279 , n31278 , n21853 );
and ( n31280 , n31275 , n31279 );
and ( n31281 , n23381 , n21741 );
and ( n31282 , n23271 , n21739 );
nor ( n31283 , n31281 , n31282 );
xnor ( n31284 , n31283 , n21605 );
and ( n31285 , n31279 , n31284 );
and ( n31286 , n31275 , n31284 );
or ( n31287 , n31280 , n31285 , n31286 );
and ( n31288 , n23968 , n21468 );
and ( n31289 , n23573 , n21466 );
nor ( n31290 , n31288 , n31289 );
xnor ( n31291 , n31290 , n21331 );
and ( n31292 , n24521 , n21155 );
and ( n31293 , n24131 , n21153 );
nor ( n31294 , n31292 , n31293 );
xnor ( n31295 , n31294 , n20994 );
and ( n31296 , n31291 , n31295 );
and ( n31297 , n24621 , n20955 );
and ( n31298 , n24527 , n20953 );
nor ( n31299 , n31297 , n31298 );
xnor ( n31300 , n31299 , n20780 );
and ( n31301 , n31295 , n31300 );
and ( n31302 , n31291 , n31300 );
or ( n31303 , n31296 , n31301 , n31302 );
and ( n31304 , n31287 , n31303 );
and ( n31305 , n25284 , n20674 );
and ( n31306 , n24940 , n20672 );
nor ( n31307 , n31305 , n31306 );
xnor ( n31308 , n31307 , n20542 );
and ( n31309 , n25765 , n20460 );
and ( n31310 , n25554 , n20458 );
nor ( n31311 , n31309 , n31310 );
xnor ( n31312 , n31311 , n20337 );
and ( n31313 , n31308 , n31312 );
and ( n31314 , n26851 , n20114 );
and ( n31315 , n26422 , n20112 );
nor ( n31316 , n31314 , n31315 );
xnor ( n31317 , n31316 , n19997 );
and ( n31318 , n31312 , n31317 );
and ( n31319 , n31308 , n31317 );
or ( n31320 , n31313 , n31318 , n31319 );
and ( n31321 , n31303 , n31320 );
and ( n31322 , n31287 , n31320 );
or ( n31323 , n31304 , n31321 , n31322 );
and ( n31324 , n31271 , n31323 );
xor ( n31325 , n30993 , n30997 );
xor ( n31326 , n31325 , n31002 );
and ( n31327 , n31323 , n31326 );
and ( n31328 , n31271 , n31326 );
or ( n31329 , n31324 , n31327 , n31328 );
and ( n31330 , n31255 , n31329 );
xor ( n31331 , n30989 , n31005 );
xor ( n31332 , n31331 , n31008 );
and ( n31333 , n31329 , n31332 );
and ( n31334 , n31255 , n31332 );
or ( n31335 , n31330 , n31333 , n31334 );
xor ( n31336 , n30797 , n30799 );
xor ( n31337 , n31336 , n30802 );
and ( n31338 , n31335 , n31337 );
xor ( n31339 , n31011 , n31085 );
xor ( n31340 , n31339 , n31088 );
and ( n31341 , n31337 , n31340 );
and ( n31342 , n31335 , n31340 );
or ( n31343 , n31338 , n31341 , n31342 );
and ( n31344 , n31193 , n31343 );
xor ( n31345 , n31096 , n31098 );
xor ( n31346 , n31345 , n31101 );
and ( n31347 , n31343 , n31346 );
and ( n31348 , n31193 , n31346 );
or ( n31349 , n31344 , n31347 , n31348 );
xor ( n31350 , n31094 , n31104 );
xor ( n31351 , n31350 , n31107 );
and ( n31352 , n31349 , n31351 );
xor ( n31353 , n31120 , n31122 );
xor ( n31354 , n31353 , n31125 );
and ( n31355 , n31351 , n31354 );
and ( n31356 , n31349 , n31354 );
or ( n31357 , n31352 , n31355 , n31356 );
xor ( n31358 , n30819 , n30821 );
xor ( n31359 , n31358 , n30824 );
and ( n31360 , n31357 , n31359 );
xor ( n31361 , n31110 , n31128 );
xor ( n31362 , n31361 , n31131 );
and ( n31363 , n31359 , n31362 );
and ( n31364 , n31357 , n31362 );
or ( n31365 , n31360 , n31363 , n31364 );
and ( n31366 , n31144 , n31365 );
xor ( n31367 , n31144 , n31365 );
xor ( n31368 , n31357 , n31359 );
xor ( n31369 , n31368 , n31362 );
xor ( n31370 , n30977 , n30981 );
xor ( n31371 , n31370 , n30986 );
xor ( n31372 , n30934 , n30950 );
xor ( n31373 , n31372 , n30955 );
and ( n31374 , n31371 , n31373 );
xor ( n31375 , n31023 , n31027 );
xor ( n31376 , n31375 , n31032 );
and ( n31377 , n31373 , n31376 );
and ( n31378 , n31371 , n31376 );
or ( n31379 , n31374 , n31377 , n31378 );
xor ( n31380 , n30831 , n30835 );
xor ( n31381 , n31380 , n30840 );
xor ( n31382 , n30922 , n30926 );
xor ( n31383 , n31382 , n30931 );
and ( n31384 , n31381 , n31383 );
xor ( n31385 , n30938 , n30942 );
xor ( n31386 , n31385 , n30947 );
and ( n31387 , n31383 , n31386 );
and ( n31388 , n31381 , n31386 );
or ( n31389 , n31384 , n31387 , n31388 );
and ( n31390 , n19496 , n29977 );
and ( n31391 , n19469 , n29974 );
nor ( n31392 , n31390 , n31391 );
xnor ( n31393 , n31392 , n28674 );
and ( n31394 , n19637 , n28628 );
and ( n31395 , n19605 , n28626 );
nor ( n31396 , n31394 , n31395 );
xnor ( n31397 , n31396 , n28096 );
and ( n31398 , n31393 , n31397 );
xor ( n31399 , n31059 , n31063 );
xor ( n31400 , n31399 , n31068 );
and ( n31401 , n31397 , n31400 );
and ( n31402 , n31393 , n31400 );
or ( n31403 , n31398 , n31401 , n31402 );
and ( n31404 , n31389 , n31403 );
xor ( n31405 , n31051 , n31071 );
xor ( n31406 , n31405 , n31076 );
and ( n31407 , n31403 , n31406 );
and ( n31408 , n31389 , n31406 );
or ( n31409 , n31404 , n31407 , n31408 );
and ( n31410 , n31379 , n31409 );
xor ( n31411 , n30958 , n30960 );
xor ( n31412 , n31411 , n30963 );
and ( n31413 , n31409 , n31412 );
and ( n31414 , n31379 , n31412 );
or ( n31415 , n31410 , n31413 , n31414 );
xor ( n31416 , n30867 , n30877 );
xor ( n31417 , n31416 , n30880 );
and ( n31418 , n31415 , n31417 );
xor ( n31419 , n30918 , n30966 );
xor ( n31420 , n31419 , n30969 );
and ( n31421 , n31417 , n31420 );
and ( n31422 , n31415 , n31420 );
or ( n31423 , n31418 , n31421 , n31422 );
xor ( n31424 , n30883 , n30972 );
xor ( n31425 , n31424 , n31091 );
and ( n31426 , n31423 , n31425 );
xor ( n31427 , n31112 , n31114 );
xor ( n31428 , n31427 , n31117 );
and ( n31429 , n31425 , n31428 );
and ( n31430 , n31423 , n31428 );
or ( n31431 , n31426 , n31429 , n31430 );
and ( n31432 , n20268 , n26349 );
and ( n31433 , n20182 , n26347 );
nor ( n31434 , n31432 , n31433 );
xnor ( n31435 , n31434 , n25893 );
and ( n31436 , n20666 , n25383 );
and ( n31437 , n20618 , n25381 );
nor ( n31438 , n31436 , n31437 );
xnor ( n31439 , n31438 , n24885 );
and ( n31440 , n31435 , n31439 );
and ( n31441 , n20867 , n24902 );
and ( n31442 , n20803 , n24900 );
nor ( n31443 , n31441 , n31442 );
xnor ( n31444 , n31443 , n24397 );
and ( n31445 , n31439 , n31444 );
and ( n31446 , n31435 , n31444 );
or ( n31447 , n31440 , n31445 , n31446 );
and ( n31448 , n22425 , n22859 );
and ( n31449 , n22198 , n22857 );
nor ( n31450 , n31448 , n31449 );
xnor ( n31451 , n31450 , n22418 );
and ( n31452 , n22916 , n22381 );
and ( n31453 , n22756 , n22379 );
nor ( n31454 , n31452 , n31453 );
xnor ( n31455 , n31454 , n22228 );
and ( n31456 , n31451 , n31455 );
and ( n31457 , n31455 , n31056 );
and ( n31458 , n31451 , n31056 );
or ( n31459 , n31456 , n31457 , n31458 );
and ( n31460 , n20452 , n26027 );
and ( n31461 , n20360 , n26025 );
nor ( n31462 , n31460 , n31461 );
xnor ( n31463 , n31462 , n25499 );
and ( n31464 , n31459 , n31463 );
and ( n31465 , n29623 , n19518 );
and ( n31466 , n29318 , n19516 );
nor ( n31467 , n31465 , n31466 );
xnor ( n31468 , n31467 , n19489 );
and ( n31469 , n31463 , n31468 );
and ( n31470 , n31459 , n31468 );
or ( n31471 , n31464 , n31469 , n31470 );
and ( n31472 , n31447 , n31471 );
xor ( n31473 , n31039 , n31043 );
xor ( n31474 , n31473 , n31048 );
and ( n31475 , n31471 , n31474 );
and ( n31476 , n31447 , n31474 );
or ( n31477 , n31472 , n31475 , n31476 );
xor ( n31478 , n30843 , n30845 );
xor ( n31479 , n31478 , n30848 );
and ( n31480 , n31477 , n31479 );
xor ( n31481 , n30853 , n30855 );
xor ( n31482 , n31481 , n30858 );
and ( n31483 , n31479 , n31482 );
and ( n31484 , n31477 , n31482 );
or ( n31485 , n31480 , n31483 , n31484 );
xor ( n31486 , n30851 , n30861 );
xor ( n31487 , n31486 , n30864 );
and ( n31488 , n31485 , n31487 );
xor ( n31489 , n31035 , n31079 );
xor ( n31490 , n31489 , n31082 );
and ( n31491 , n31487 , n31490 );
and ( n31492 , n31485 , n31490 );
or ( n31493 , n31488 , n31491 , n31492 );
and ( n31494 , n20080 , n26992 );
and ( n31495 , n20004 , n26990 );
nor ( n31496 , n31494 , n31495 );
xnor ( n31497 , n31496 , n26369 );
and ( n31498 , n21218 , n24376 );
and ( n31499 , n21072 , n24374 );
nor ( n31500 , n31498 , n31499 );
xnor ( n31501 , n31500 , n23927 );
and ( n31502 , n31497 , n31501 );
and ( n31503 , n21451 , n23944 );
and ( n31504 , n21302 , n23942 );
nor ( n31505 , n31503 , n31504 );
xnor ( n31506 , n31505 , n23550 );
and ( n31507 , n31501 , n31506 );
and ( n31508 , n31497 , n31506 );
or ( n31509 , n31502 , n31507 , n31508 );
and ( n31510 , n26422 , n20276 );
and ( n31511 , n26319 , n20274 );
nor ( n31512 , n31510 , n31511 );
xnor ( n31513 , n31512 , n20175 );
and ( n31514 , n28211 , n19805 );
and ( n31515 , n27757 , n19803 );
nor ( n31516 , n31514 , n31515 );
xnor ( n31517 , n31516 , n19750 );
and ( n31518 , n31513 , n31517 );
and ( n31519 , n29318 , n19596 );
and ( n31520 , n29078 , n19594 );
nor ( n31521 , n31519 , n31520 );
xnor ( n31522 , n31521 , n19545 );
and ( n31523 , n31517 , n31522 );
and ( n31524 , n31513 , n31522 );
or ( n31525 , n31518 , n31523 , n31524 );
and ( n31526 , n19605 , n29276 );
and ( n31527 , n19588 , n29274 );
nor ( n31528 , n31526 , n31527 );
xnor ( n31529 , n31528 , n28677 );
and ( n31530 , n31525 , n31529 );
and ( n31531 , n19946 , n27529 );
and ( n31532 , n19881 , n27527 );
nor ( n31533 , n31531 , n31532 );
xnor ( n31534 , n31533 , n27034 );
and ( n31535 , n31529 , n31534 );
and ( n31536 , n31525 , n31534 );
or ( n31537 , n31530 , n31535 , n31536 );
and ( n31538 , n31509 , n31537 );
xor ( n31539 , n31259 , n31263 );
xor ( n31540 , n31539 , n31268 );
and ( n31541 , n31537 , n31540 );
and ( n31542 , n31509 , n31540 );
or ( n31543 , n31538 , n31541 , n31542 );
and ( n31544 , n19825 , n28062 );
and ( n31545 , n19811 , n28060 );
nor ( n31546 , n31544 , n31545 );
xnor ( n31547 , n31546 , n27549 );
and ( n31548 , n21704 , n23641 );
and ( n31549 , n21612 , n23639 );
nor ( n31550 , n31548 , n31549 );
xnor ( n31551 , n31550 , n23213 );
and ( n31552 , n31547 , n31551 );
and ( n31553 , n21955 , n23230 );
and ( n31554 , n21876 , n23228 );
nor ( n31555 , n31553 , n31554 );
xnor ( n31556 , n31555 , n22842 );
and ( n31557 , n31551 , n31556 );
and ( n31558 , n31547 , n31556 );
or ( n31559 , n31552 , n31557 , n31558 );
and ( n31560 , n23271 , n22048 );
and ( n31561 , n23141 , n22046 );
nor ( n31562 , n31560 , n31561 );
xnor ( n31563 , n31562 , n21853 );
and ( n31564 , n23573 , n21741 );
and ( n31565 , n23381 , n21739 );
nor ( n31566 , n31564 , n31565 );
xnor ( n31567 , n31566 , n21605 );
and ( n31568 , n31563 , n31567 );
and ( n31569 , n24131 , n21468 );
and ( n31570 , n23968 , n21466 );
nor ( n31571 , n31569 , n31570 );
xnor ( n31572 , n31571 , n21331 );
and ( n31573 , n31567 , n31572 );
and ( n31574 , n31563 , n31572 );
or ( n31575 , n31568 , n31573 , n31574 );
and ( n31576 , n25974 , n20460 );
and ( n31577 , n25765 , n20458 );
nor ( n31578 , n31576 , n31577 );
xnor ( n31579 , n31578 , n20337 );
and ( n31580 , n27135 , n20114 );
and ( n31581 , n26851 , n20112 );
nor ( n31582 , n31580 , n31581 );
xnor ( n31583 , n31582 , n19997 );
and ( n31584 , n31579 , n31583 );
and ( n31585 , n27751 , n19894 );
and ( n31586 , n27352 , n19892 );
nor ( n31587 , n31585 , n31586 );
xnor ( n31588 , n31587 , n19858 );
and ( n31589 , n31583 , n31588 );
and ( n31590 , n31579 , n31588 );
or ( n31591 , n31584 , n31589 , n31590 );
and ( n31592 , n31575 , n31591 );
and ( n31593 , n24527 , n21155 );
and ( n31594 , n24521 , n21153 );
nor ( n31595 , n31593 , n31594 );
xnor ( n31596 , n31595 , n20994 );
and ( n31597 , n24940 , n20955 );
and ( n31598 , n24621 , n20953 );
nor ( n31599 , n31597 , n31598 );
xnor ( n31600 , n31599 , n20780 );
and ( n31601 , n31596 , n31600 );
and ( n31602 , n25554 , n20674 );
and ( n31603 , n25284 , n20672 );
nor ( n31604 , n31602 , n31603 );
xnor ( n31605 , n31604 , n20542 );
and ( n31606 , n31600 , n31605 );
and ( n31607 , n31596 , n31605 );
or ( n31608 , n31601 , n31606 , n31607 );
and ( n31609 , n31591 , n31608 );
and ( n31610 , n31575 , n31608 );
or ( n31611 , n31592 , n31609 , n31610 );
and ( n31612 , n31559 , n31611 );
xor ( n31613 , n31197 , n31201 );
xor ( n31614 , n31613 , n31206 );
and ( n31615 , n31611 , n31614 );
and ( n31616 , n31559 , n31614 );
or ( n31617 , n31612 , n31615 , n31616 );
and ( n31618 , n31543 , n31617 );
xor ( n31619 , n31209 , n31225 );
xor ( n31620 , n31619 , n31252 );
and ( n31621 , n31617 , n31620 );
and ( n31622 , n31543 , n31620 );
or ( n31623 , n31618 , n31621 , n31622 );
xor ( n31624 , n30869 , n30871 );
xor ( n31625 , n31624 , n30874 );
and ( n31626 , n31623 , n31625 );
xor ( n31627 , n31255 , n31329 );
xor ( n31628 , n31627 , n31332 );
and ( n31629 , n31625 , n31628 );
and ( n31630 , n31623 , n31628 );
or ( n31631 , n31626 , n31629 , n31630 );
and ( n31632 , n31493 , n31631 );
xor ( n31633 , n31185 , n31187 );
xor ( n31634 , n31633 , n31190 );
and ( n31635 , n31631 , n31634 );
and ( n31636 , n31493 , n31634 );
or ( n31637 , n31632 , n31635 , n31636 );
xor ( n31638 , n31213 , n31217 );
xor ( n31639 , n31638 , n31222 );
xor ( n31640 , n31287 , n31303 );
xor ( n31641 , n31640 , n31320 );
and ( n31642 , n31639 , n31641 );
xor ( n31643 , n31393 , n31397 );
xor ( n31644 , n31643 , n31400 );
and ( n31645 , n31641 , n31644 );
and ( n31646 , n31639 , n31644 );
or ( n31647 , n31642 , n31645 , n31646 );
and ( n31648 , n22756 , n22859 );
and ( n31649 , n22425 , n22857 );
nor ( n31650 , n31648 , n31649 );
xnor ( n31651 , n31650 , n22418 );
and ( n31652 , n23141 , n22381 );
and ( n31653 , n22916 , n22379 );
nor ( n31654 , n31652 , n31653 );
xnor ( n31655 , n31654 , n22228 );
and ( n31656 , n31651 , n31655 );
and ( n31657 , n22235 , n23230 );
and ( n31658 , n21955 , n23228 );
nor ( n31659 , n31657 , n31658 );
xnor ( n31660 , n31659 , n22842 );
and ( n31661 , n31656 , n31660 );
and ( n31662 , n28700 , n19688 );
and ( n31663 , n28810 , n19686 );
nor ( n31664 , n31662 , n31663 );
xnor ( n31665 , n31664 , n19655 );
and ( n31666 , n31660 , n31665 );
and ( n31667 , n31656 , n31665 );
or ( n31668 , n31661 , n31666 , n31667 );
and ( n31669 , n19510 , n29977 );
and ( n31670 , n19496 , n29974 );
nor ( n31671 , n31669 , n31670 );
xnor ( n31672 , n31671 , n28674 );
and ( n31673 , n31668 , n31672 );
and ( n31674 , n19721 , n28628 );
and ( n31675 , n19637 , n28626 );
nor ( n31676 , n31674 , n31675 );
xnor ( n31677 , n31676 , n28096 );
and ( n31678 , n31672 , n31677 );
and ( n31679 , n31668 , n31677 );
or ( n31680 , n31673 , n31678 , n31679 );
xor ( n31681 , n31157 , n31161 );
xor ( n31682 , n31681 , n31166 );
and ( n31683 , n31680 , n31682 );
xor ( n31684 , n31242 , n31246 );
xor ( n31685 , n31684 , n31249 );
and ( n31686 , n31682 , n31685 );
and ( n31687 , n31680 , n31685 );
or ( n31688 , n31683 , n31686 , n31687 );
and ( n31689 , n31647 , n31688 );
xor ( n31690 , n31271 , n31323 );
xor ( n31691 , n31690 , n31326 );
and ( n31692 , n31688 , n31691 );
and ( n31693 , n31647 , n31691 );
or ( n31694 , n31689 , n31692 , n31693 );
xor ( n31695 , n31177 , n31179 );
xor ( n31696 , n31695 , n31182 );
and ( n31697 , n31694 , n31696 );
xor ( n31698 , n31379 , n31409 );
xor ( n31699 , n31698 , n31412 );
and ( n31700 , n31696 , n31699 );
and ( n31701 , n31694 , n31699 );
or ( n31702 , n31697 , n31700 , n31701 );
xor ( n31703 , n31335 , n31337 );
xor ( n31704 , n31703 , n31340 );
and ( n31705 , n31702 , n31704 );
xor ( n31706 , n31415 , n31417 );
xor ( n31707 , n31706 , n31420 );
and ( n31708 , n31704 , n31707 );
and ( n31709 , n31702 , n31707 );
or ( n31710 , n31705 , n31708 , n31709 );
and ( n31711 , n31637 , n31710 );
xor ( n31712 , n31193 , n31343 );
xor ( n31713 , n31712 , n31346 );
and ( n31714 , n31710 , n31713 );
and ( n31715 , n31637 , n31713 );
or ( n31716 , n31711 , n31714 , n31715 );
and ( n31717 , n31431 , n31716 );
xor ( n31718 , n31349 , n31351 );
xor ( n31719 , n31718 , n31354 );
and ( n31720 , n31716 , n31719 );
and ( n31721 , n31431 , n31719 );
or ( n31722 , n31717 , n31720 , n31721 );
and ( n31723 , n31369 , n31722 );
xor ( n31724 , n31369 , n31722 );
xor ( n31725 , n31431 , n31716 );
xor ( n31726 , n31725 , n31719 );
xor ( n31727 , n31371 , n31373 );
xor ( n31728 , n31727 , n31376 );
xor ( n31729 , n31169 , n31171 );
xor ( n31730 , n31729 , n31174 );
and ( n31731 , n31728 , n31730 );
xor ( n31732 , n31389 , n31403 );
xor ( n31733 , n31732 , n31406 );
and ( n31734 , n31730 , n31733 );
and ( n31735 , n31728 , n31733 );
or ( n31736 , n31731 , n31734 , n31735 );
and ( n31737 , n21302 , n24376 );
and ( n31738 , n21218 , n24374 );
nor ( n31739 , n31737 , n31738 );
xnor ( n31740 , n31739 , n23927 );
and ( n31741 , n21612 , n23944 );
and ( n31742 , n21451 , n23942 );
nor ( n31743 , n31741 , n31742 );
xnor ( n31744 , n31743 , n23550 );
and ( n31745 , n31740 , n31744 );
and ( n31746 , n21876 , n23641 );
and ( n31747 , n21704 , n23639 );
nor ( n31748 , n31746 , n31747 );
xnor ( n31749 , n31748 , n23213 );
and ( n31750 , n31744 , n31749 );
and ( n31751 , n31740 , n31749 );
or ( n31752 , n31745 , n31750 , n31751 );
xor ( n31753 , n31291 , n31295 );
xor ( n31754 , n31753 , n31300 );
and ( n31755 , n31752 , n31754 );
xor ( n31756 , n31308 , n31312 );
xor ( n31757 , n31756 , n31317 );
and ( n31758 , n31754 , n31757 );
and ( n31759 , n31752 , n31757 );
or ( n31760 , n31755 , n31758 , n31759 );
and ( n31761 , n26851 , n20276 );
and ( n31762 , n26422 , n20274 );
nor ( n31763 , n31761 , n31762 );
xnor ( n31764 , n31763 , n20175 );
and ( n31765 , n27352 , n20114 );
and ( n31766 , n27135 , n20112 );
nor ( n31767 , n31765 , n31766 );
xnor ( n31768 , n31767 , n19997 );
and ( n31769 , n31764 , n31768 );
and ( n31770 , n27757 , n19894 );
and ( n31771 , n27751 , n19892 );
nor ( n31772 , n31770 , n31771 );
xnor ( n31773 , n31772 , n19858 );
and ( n31774 , n31768 , n31773 );
and ( n31775 , n31764 , n31773 );
or ( n31776 , n31769 , n31774 , n31775 );
and ( n31777 , n25284 , n20955 );
and ( n31778 , n24940 , n20953 );
nor ( n31779 , n31777 , n31778 );
xnor ( n31780 , n31779 , n20780 );
and ( n31781 , n25765 , n20674 );
and ( n31782 , n25554 , n20672 );
nor ( n31783 , n31781 , n31782 );
xnor ( n31784 , n31783 , n20542 );
and ( n31785 , n31780 , n31784 );
and ( n31786 , n26319 , n20460 );
and ( n31787 , n25974 , n20458 );
nor ( n31788 , n31786 , n31787 );
xnor ( n31789 , n31788 , n20337 );
and ( n31790 , n31784 , n31789 );
and ( n31791 , n31780 , n31789 );
or ( n31792 , n31785 , n31790 , n31791 );
and ( n31793 , n31776 , n31792 );
and ( n31794 , n19588 , n29977 );
and ( n31795 , n19510 , n29974 );
nor ( n31796 , n31794 , n31795 );
xnor ( n31797 , n31796 , n28674 );
and ( n31798 , n31792 , n31797 );
and ( n31799 , n31776 , n31797 );
or ( n31800 , n31793 , n31798 , n31799 );
and ( n31801 , n22198 , n23230 );
and ( n31802 , n22235 , n23228 );
nor ( n31803 , n31801 , n31802 );
xnor ( n31804 , n31803 , n22842 );
and ( n31805 , n23381 , n22048 );
and ( n31806 , n23271 , n22046 );
nor ( n31807 , n31805 , n31806 );
xnor ( n31808 , n31807 , n21853 );
and ( n31809 , n31804 , n31808 );
and ( n31810 , n29623 , n19594 );
not ( n31811 , n31810 );
and ( n31812 , n31811 , n19545 );
and ( n31813 , n31808 , n31812 );
and ( n31814 , n31804 , n31812 );
or ( n31815 , n31809 , n31813 , n31814 );
and ( n31816 , n23968 , n21741 );
and ( n31817 , n23573 , n21739 );
nor ( n31818 , n31816 , n31817 );
xnor ( n31819 , n31818 , n21605 );
and ( n31820 , n24521 , n21468 );
and ( n31821 , n24131 , n21466 );
nor ( n31822 , n31820 , n31821 );
xnor ( n31823 , n31822 , n21331 );
and ( n31824 , n31819 , n31823 );
and ( n31825 , n24621 , n21155 );
and ( n31826 , n24527 , n21153 );
nor ( n31827 , n31825 , n31826 );
xnor ( n31828 , n31827 , n20994 );
and ( n31829 , n31823 , n31828 );
and ( n31830 , n31819 , n31828 );
or ( n31831 , n31824 , n31829 , n31830 );
and ( n31832 , n31815 , n31831 );
and ( n31833 , n19881 , n28062 );
and ( n31834 , n19825 , n28060 );
nor ( n31835 , n31833 , n31834 );
xnor ( n31836 , n31835 , n27549 );
and ( n31837 , n31831 , n31836 );
and ( n31838 , n31815 , n31836 );
or ( n31839 , n31832 , n31837 , n31838 );
and ( n31840 , n31800 , n31839 );
xor ( n31841 , n31547 , n31551 );
xor ( n31842 , n31841 , n31556 );
and ( n31843 , n31839 , n31842 );
and ( n31844 , n31800 , n31842 );
or ( n31845 , n31840 , n31843 , n31844 );
and ( n31846 , n31760 , n31845 );
xor ( n31847 , n31651 , n31655 );
and ( n31848 , n28810 , n19805 );
and ( n31849 , n28211 , n19803 );
nor ( n31850 , n31848 , n31849 );
xnor ( n31851 , n31850 , n19750 );
and ( n31852 , n31847 , n31851 );
and ( n31853 , n29623 , n19596 );
and ( n31854 , n29318 , n19594 );
nor ( n31855 , n31853 , n31854 );
xnor ( n31856 , n31855 , n19545 );
and ( n31857 , n31851 , n31856 );
and ( n31858 , n31847 , n31856 );
or ( n31859 , n31852 , n31857 , n31858 );
and ( n31860 , n19637 , n29276 );
and ( n31861 , n19605 , n29274 );
nor ( n31862 , n31860 , n31861 );
xnor ( n31863 , n31862 , n28677 );
and ( n31864 , n31859 , n31863 );
and ( n31865 , n20004 , n27529 );
and ( n31866 , n19946 , n27527 );
nor ( n31867 , n31865 , n31866 );
xnor ( n31868 , n31867 , n27034 );
and ( n31869 , n31863 , n31868 );
and ( n31870 , n31859 , n31868 );
or ( n31871 , n31864 , n31869 , n31870 );
xor ( n31872 , n31435 , n31439 );
xor ( n31873 , n31872 , n31444 );
and ( n31874 , n31871 , n31873 );
xor ( n31875 , n31497 , n31501 );
xor ( n31876 , n31875 , n31506 );
and ( n31877 , n31873 , n31876 );
and ( n31878 , n31871 , n31876 );
or ( n31879 , n31874 , n31877 , n31878 );
and ( n31880 , n31845 , n31879 );
and ( n31881 , n31760 , n31879 );
or ( n31882 , n31846 , n31880 , n31881 );
xor ( n31883 , n31275 , n31279 );
xor ( n31884 , n31883 , n31284 );
xor ( n31885 , n31230 , n31234 );
xor ( n31886 , n31885 , n31239 );
and ( n31887 , n31884 , n31886 );
xor ( n31888 , n31145 , n31149 );
xor ( n31889 , n31888 , n31154 );
and ( n31890 , n31886 , n31889 );
and ( n31891 , n31884 , n31889 );
or ( n31892 , n31887 , n31890 , n31891 );
and ( n31893 , n20618 , n26027 );
and ( n31894 , n20452 , n26025 );
nor ( n31895 , n31893 , n31894 );
xnor ( n31896 , n31895 , n25499 );
and ( n31897 , n20803 , n25383 );
and ( n31898 , n20666 , n25381 );
nor ( n31899 , n31897 , n31898 );
xnor ( n31900 , n31899 , n24885 );
and ( n31901 , n31896 , n31900 );
and ( n31902 , n21072 , n24902 );
and ( n31903 , n20867 , n24900 );
nor ( n31904 , n31902 , n31903 );
xnor ( n31905 , n31904 , n24397 );
and ( n31906 , n31900 , n31905 );
and ( n31907 , n31896 , n31905 );
or ( n31908 , n31901 , n31906 , n31907 );
and ( n31909 , n20182 , n26992 );
and ( n31910 , n20080 , n26990 );
nor ( n31911 , n31909 , n31910 );
xnor ( n31912 , n31911 , n26369 );
and ( n31913 , n20360 , n26349 );
and ( n31914 , n20268 , n26347 );
nor ( n31915 , n31913 , n31914 );
xnor ( n31916 , n31915 , n25893 );
and ( n31917 , n31912 , n31916 );
xor ( n31918 , n31451 , n31455 );
xor ( n31919 , n31918 , n31056 );
and ( n31920 , n31916 , n31919 );
and ( n31921 , n31912 , n31919 );
or ( n31922 , n31917 , n31920 , n31921 );
and ( n31923 , n31908 , n31922 );
xor ( n31924 , n31459 , n31463 );
xor ( n31925 , n31924 , n31468 );
and ( n31926 , n31922 , n31925 );
and ( n31927 , n31908 , n31925 );
or ( n31928 , n31923 , n31926 , n31927 );
and ( n31929 , n31892 , n31928 );
xor ( n31930 , n31381 , n31383 );
xor ( n31931 , n31930 , n31386 );
and ( n31932 , n31928 , n31931 );
and ( n31933 , n31892 , n31931 );
or ( n31934 , n31929 , n31932 , n31933 );
and ( n31935 , n31882 , n31934 );
xor ( n31936 , n31477 , n31479 );
xor ( n31937 , n31936 , n31482 );
and ( n31938 , n31934 , n31937 );
and ( n31939 , n31882 , n31937 );
or ( n31940 , n31935 , n31938 , n31939 );
and ( n31941 , n31736 , n31940 );
xor ( n31942 , n31485 , n31487 );
xor ( n31943 , n31942 , n31490 );
and ( n31944 , n31940 , n31943 );
and ( n31945 , n31736 , n31943 );
or ( n31946 , n31941 , n31944 , n31945 );
xor ( n31947 , n31563 , n31567 );
xor ( n31948 , n31947 , n31572 );
xor ( n31949 , n31579 , n31583 );
xor ( n31950 , n31949 , n31588 );
and ( n31951 , n31948 , n31950 );
xor ( n31952 , n31596 , n31600 );
xor ( n31953 , n31952 , n31605 );
and ( n31954 , n31950 , n31953 );
and ( n31955 , n31948 , n31953 );
or ( n31956 , n31951 , n31954 , n31955 );
xor ( n31957 , n31575 , n31591 );
xor ( n31958 , n31957 , n31608 );
and ( n31959 , n31956 , n31958 );
xor ( n31960 , n31668 , n31672 );
xor ( n31961 , n31960 , n31677 );
and ( n31962 , n31958 , n31961 );
and ( n31963 , n31956 , n31961 );
or ( n31964 , n31959 , n31962 , n31963 );
xor ( n31965 , n31447 , n31471 );
xor ( n31966 , n31965 , n31474 );
and ( n31967 , n31964 , n31966 );
xor ( n31968 , n31509 , n31537 );
xor ( n31969 , n31968 , n31540 );
and ( n31970 , n31966 , n31969 );
and ( n31971 , n31964 , n31969 );
or ( n31972 , n31967 , n31970 , n31971 );
xor ( n31973 , n31543 , n31617 );
xor ( n31974 , n31973 , n31620 );
and ( n31975 , n31972 , n31974 );
xor ( n31976 , n31647 , n31688 );
xor ( n31977 , n31976 , n31691 );
and ( n31978 , n31974 , n31977 );
and ( n31979 , n31972 , n31977 );
or ( n31980 , n31975 , n31978 , n31979 );
xor ( n31981 , n31623 , n31625 );
xor ( n31982 , n31981 , n31628 );
and ( n31983 , n31980 , n31982 );
xor ( n31984 , n31694 , n31696 );
xor ( n31985 , n31984 , n31699 );
and ( n31986 , n31982 , n31985 );
and ( n31987 , n31980 , n31985 );
or ( n31988 , n31983 , n31986 , n31987 );
and ( n31989 , n31946 , n31988 );
xor ( n31990 , n31493 , n31631 );
xor ( n31991 , n31990 , n31634 );
and ( n31992 , n31988 , n31991 );
and ( n31993 , n31946 , n31991 );
or ( n31994 , n31989 , n31992 , n31993 );
xor ( n31995 , n31423 , n31425 );
xor ( n31996 , n31995 , n31428 );
and ( n31997 , n31994 , n31996 );
xor ( n31998 , n31637 , n31710 );
xor ( n31999 , n31998 , n31713 );
and ( n32000 , n31996 , n31999 );
and ( n32001 , n31994 , n31999 );
or ( n32002 , n31997 , n32000 , n32001 );
and ( n32003 , n31726 , n32002 );
xor ( n32004 , n31726 , n32002 );
xor ( n32005 , n31994 , n31996 );
xor ( n32006 , n32005 , n31999 );
and ( n32007 , n20452 , n26349 );
and ( n32008 , n20360 , n26347 );
nor ( n32009 , n32007 , n32008 );
xnor ( n32010 , n32009 , n25893 );
and ( n32011 , n21704 , n23944 );
and ( n32012 , n21612 , n23942 );
nor ( n32013 , n32011 , n32012 );
xnor ( n32014 , n32013 , n23550 );
and ( n32015 , n32010 , n32014 );
and ( n32016 , n21955 , n23641 );
and ( n32017 , n21876 , n23639 );
nor ( n32018 , n32016 , n32017 );
xnor ( n32019 , n32018 , n23213 );
and ( n32020 , n32014 , n32019 );
and ( n32021 , n32010 , n32019 );
or ( n32022 , n32015 , n32020 , n32021 );
and ( n32023 , n20867 , n25383 );
and ( n32024 , n20803 , n25381 );
nor ( n32025 , n32023 , n32024 );
xnor ( n32026 , n32025 , n24885 );
and ( n32027 , n21218 , n24902 );
and ( n32028 , n21072 , n24900 );
nor ( n32029 , n32027 , n32028 );
xnor ( n32030 , n32029 , n24397 );
and ( n32031 , n32026 , n32030 );
and ( n32032 , n21451 , n24376 );
and ( n32033 , n21302 , n24374 );
nor ( n32034 , n32032 , n32033 );
xnor ( n32035 , n32034 , n23927 );
and ( n32036 , n32030 , n32035 );
and ( n32037 , n32026 , n32035 );
or ( n32038 , n32031 , n32036 , n32037 );
and ( n32039 , n32022 , n32038 );
and ( n32040 , n22425 , n23230 );
and ( n32041 , n22198 , n23228 );
nor ( n32042 , n32040 , n32041 );
xnor ( n32043 , n32042 , n22842 );
and ( n32044 , n22916 , n22859 );
and ( n32045 , n22756 , n22857 );
nor ( n32046 , n32044 , n32045 );
xnor ( n32047 , n32046 , n22418 );
and ( n32048 , n32043 , n32047 );
and ( n32049 , n23271 , n22381 );
and ( n32050 , n23141 , n22379 );
nor ( n32051 , n32049 , n32050 );
xnor ( n32052 , n32051 , n22228 );
and ( n32053 , n32047 , n32052 );
and ( n32054 , n32043 , n32052 );
or ( n32055 , n32048 , n32053 , n32054 );
and ( n32056 , n20666 , n26027 );
and ( n32057 , n20618 , n26025 );
nor ( n32058 , n32056 , n32057 );
xnor ( n32059 , n32058 , n25499 );
and ( n32060 , n32055 , n32059 );
and ( n32061 , n29078 , n19688 );
and ( n32062 , n28700 , n19686 );
nor ( n32063 , n32061 , n32062 );
xnor ( n32064 , n32063 , n19655 );
and ( n32065 , n32059 , n32064 );
and ( n32066 , n32055 , n32064 );
or ( n32067 , n32060 , n32065 , n32066 );
and ( n32068 , n32038 , n32067 );
and ( n32069 , n32022 , n32067 );
or ( n32070 , n32039 , n32068 , n32069 );
and ( n32071 , n19811 , n28628 );
and ( n32072 , n19721 , n28626 );
nor ( n32073 , n32071 , n32072 );
xnor ( n32074 , n32073 , n28096 );
xor ( n32075 , n31513 , n31517 );
xor ( n32076 , n32075 , n31522 );
and ( n32077 , n32074 , n32076 );
xor ( n32078 , n31656 , n31660 );
xor ( n32079 , n32078 , n31665 );
and ( n32080 , n32076 , n32079 );
and ( n32081 , n32074 , n32079 );
or ( n32082 , n32077 , n32080 , n32081 );
and ( n32083 , n32070 , n32082 );
xor ( n32084 , n31525 , n31529 );
xor ( n32085 , n32084 , n31534 );
and ( n32086 , n32082 , n32085 );
and ( n32087 , n32070 , n32085 );
or ( n32088 , n32083 , n32086 , n32087 );
xor ( n32089 , n31559 , n31611 );
xor ( n32090 , n32089 , n31614 );
and ( n32091 , n32088 , n32090 );
xor ( n32092 , n31680 , n31682 );
xor ( n32093 , n32092 , n31685 );
and ( n32094 , n32090 , n32093 );
and ( n32095 , n32088 , n32093 );
or ( n32096 , n32091 , n32094 , n32095 );
and ( n32097 , n27751 , n20114 );
and ( n32098 , n27352 , n20112 );
nor ( n32099 , n32097 , n32098 );
xnor ( n32100 , n32099 , n19997 );
and ( n32101 , n28211 , n19894 );
and ( n32102 , n27757 , n19892 );
nor ( n32103 , n32101 , n32102 );
xnor ( n32104 , n32103 , n19858 );
and ( n32105 , n32100 , n32104 );
and ( n32106 , n28700 , n19805 );
and ( n32107 , n28810 , n19803 );
nor ( n32108 , n32106 , n32107 );
xnor ( n32109 , n32108 , n19750 );
and ( n32110 , n32104 , n32109 );
and ( n32111 , n32100 , n32109 );
or ( n32112 , n32105 , n32110 , n32111 );
and ( n32113 , n19605 , n29977 );
and ( n32114 , n19588 , n29974 );
nor ( n32115 , n32113 , n32114 );
xnor ( n32116 , n32115 , n28674 );
and ( n32117 , n32112 , n32116 );
and ( n32118 , n19721 , n29276 );
and ( n32119 , n19637 , n29274 );
nor ( n32120 , n32118 , n32119 );
xnor ( n32121 , n32120 , n28677 );
and ( n32122 , n32116 , n32121 );
and ( n32123 , n32112 , n32121 );
or ( n32124 , n32117 , n32122 , n32123 );
xor ( n32125 , n31896 , n31900 );
xor ( n32126 , n32125 , n31905 );
and ( n32127 , n32124 , n32126 );
xor ( n32128 , n31740 , n31744 );
xor ( n32129 , n32128 , n31749 );
and ( n32130 , n32126 , n32129 );
and ( n32131 , n32124 , n32129 );
or ( n32132 , n32127 , n32130 , n32131 );
xor ( n32133 , n31752 , n31754 );
xor ( n32134 , n32133 , n31757 );
and ( n32135 , n32132 , n32134 );
xor ( n32136 , n31884 , n31886 );
xor ( n32137 , n32136 , n31889 );
and ( n32138 , n32134 , n32137 );
and ( n32139 , n32132 , n32137 );
or ( n32140 , n32135 , n32138 , n32139 );
xor ( n32141 , n31639 , n31641 );
xor ( n32142 , n32141 , n31644 );
and ( n32143 , n32140 , n32142 );
xor ( n32144 , n31892 , n31928 );
xor ( n32145 , n32144 , n31931 );
and ( n32146 , n32142 , n32145 );
and ( n32147 , n32140 , n32145 );
or ( n32148 , n32143 , n32146 , n32147 );
and ( n32149 , n32096 , n32148 );
xor ( n32150 , n31728 , n31730 );
xor ( n32151 , n32150 , n31733 );
and ( n32152 , n32148 , n32151 );
and ( n32153 , n32096 , n32151 );
or ( n32154 , n32149 , n32152 , n32153 );
and ( n32155 , n19946 , n28062 );
and ( n32156 , n19881 , n28060 );
nor ( n32157 , n32155 , n32156 );
xnor ( n32158 , n32157 , n27549 );
and ( n32159 , n20080 , n27529 );
and ( n32160 , n20004 , n27527 );
nor ( n32161 , n32159 , n32160 );
xnor ( n32162 , n32161 , n27034 );
and ( n32163 , n32158 , n32162 );
and ( n32164 , n20268 , n26992 );
and ( n32165 , n20182 , n26990 );
nor ( n32166 , n32164 , n32165 );
xnor ( n32167 , n32166 , n26369 );
and ( n32168 , n32162 , n32167 );
and ( n32169 , n32158 , n32167 );
or ( n32170 , n32163 , n32168 , n32169 );
and ( n32171 , n23573 , n22048 );
and ( n32172 , n23381 , n22046 );
nor ( n32173 , n32171 , n32172 );
xnor ( n32174 , n32173 , n21853 );
and ( n32175 , n24131 , n21741 );
and ( n32176 , n23968 , n21739 );
nor ( n32177 , n32175 , n32176 );
xnor ( n32178 , n32177 , n21605 );
and ( n32179 , n32174 , n32178 );
and ( n32180 , n32178 , n31810 );
and ( n32181 , n32174 , n31810 );
or ( n32182 , n32179 , n32180 , n32181 );
and ( n32183 , n25974 , n20674 );
and ( n32184 , n25765 , n20672 );
nor ( n32185 , n32183 , n32184 );
xnor ( n32186 , n32185 , n20542 );
and ( n32187 , n26422 , n20460 );
and ( n32188 , n26319 , n20458 );
nor ( n32189 , n32187 , n32188 );
xnor ( n32190 , n32189 , n20337 );
and ( n32191 , n32186 , n32190 );
and ( n32192 , n27135 , n20276 );
and ( n32193 , n26851 , n20274 );
nor ( n32194 , n32192 , n32193 );
xnor ( n32195 , n32194 , n20175 );
and ( n32196 , n32190 , n32195 );
and ( n32197 , n32186 , n32195 );
or ( n32198 , n32191 , n32196 , n32197 );
and ( n32199 , n32182 , n32198 );
and ( n32200 , n24527 , n21468 );
and ( n32201 , n24521 , n21466 );
nor ( n32202 , n32200 , n32201 );
xnor ( n32203 , n32202 , n21331 );
and ( n32204 , n24940 , n21155 );
and ( n32205 , n24621 , n21153 );
nor ( n32206 , n32204 , n32205 );
xnor ( n32207 , n32206 , n20994 );
and ( n32208 , n32203 , n32207 );
and ( n32209 , n25554 , n20955 );
and ( n32210 , n25284 , n20953 );
nor ( n32211 , n32209 , n32210 );
xnor ( n32212 , n32211 , n20780 );
and ( n32213 , n32207 , n32212 );
and ( n32214 , n32203 , n32212 );
or ( n32215 , n32208 , n32213 , n32214 );
and ( n32216 , n32198 , n32215 );
and ( n32217 , n32182 , n32215 );
or ( n32218 , n32199 , n32216 , n32217 );
and ( n32219 , n32170 , n32218 );
xor ( n32220 , n31912 , n31916 );
xor ( n32221 , n32220 , n31919 );
and ( n32222 , n32218 , n32221 );
and ( n32223 , n32170 , n32221 );
or ( n32224 , n32219 , n32222 , n32223 );
xor ( n32225 , n31908 , n31922 );
xor ( n32226 , n32225 , n31925 );
and ( n32227 , n32224 , n32226 );
xor ( n32228 , n31800 , n31839 );
xor ( n32229 , n32228 , n31842 );
and ( n32230 , n32226 , n32229 );
and ( n32231 , n32224 , n32229 );
or ( n32232 , n32227 , n32230 , n32231 );
xor ( n32233 , n31760 , n31845 );
xor ( n32234 , n32233 , n31879 );
and ( n32235 , n32232 , n32234 );
xor ( n32236 , n31964 , n31966 );
xor ( n32237 , n32236 , n31969 );
and ( n32238 , n32234 , n32237 );
and ( n32239 , n32232 , n32237 );
or ( n32240 , n32235 , n32238 , n32239 );
xor ( n32241 , n31882 , n31934 );
xor ( n32242 , n32241 , n31937 );
and ( n32243 , n32240 , n32242 );
xor ( n32244 , n31972 , n31974 );
xor ( n32245 , n32244 , n31977 );
and ( n32246 , n32242 , n32245 );
and ( n32247 , n32240 , n32245 );
or ( n32248 , n32243 , n32246 , n32247 );
and ( n32249 , n32154 , n32248 );
xor ( n32250 , n31736 , n31940 );
xor ( n32251 , n32250 , n31943 );
and ( n32252 , n32248 , n32251 );
and ( n32253 , n32154 , n32251 );
or ( n32254 , n32249 , n32252 , n32253 );
xor ( n32255 , n31702 , n31704 );
xor ( n32256 , n32255 , n31707 );
and ( n32257 , n32254 , n32256 );
xor ( n32258 , n31946 , n31988 );
xor ( n32259 , n32258 , n31991 );
and ( n32260 , n32256 , n32259 );
and ( n32261 , n32254 , n32259 );
or ( n32262 , n32257 , n32260 , n32261 );
and ( n32263 , n32006 , n32262 );
xor ( n32264 , n32006 , n32262 );
xor ( n32265 , n32254 , n32256 );
xor ( n32266 , n32265 , n32259 );
xor ( n32267 , n31776 , n31792 );
xor ( n32268 , n32267 , n31797 );
xor ( n32269 , n31815 , n31831 );
xor ( n32270 , n32269 , n31836 );
and ( n32271 , n32268 , n32270 );
xor ( n32272 , n31859 , n31863 );
xor ( n32273 , n32272 , n31868 );
and ( n32274 , n32270 , n32273 );
and ( n32275 , n32268 , n32273 );
or ( n32276 , n32271 , n32274 , n32275 );
and ( n32277 , n22756 , n23230 );
and ( n32278 , n22425 , n23228 );
nor ( n32279 , n32277 , n32278 );
xnor ( n32280 , n32279 , n22842 );
and ( n32281 , n23381 , n22381 );
and ( n32282 , n23271 , n22379 );
nor ( n32283 , n32281 , n32282 );
xnor ( n32284 , n32283 , n22228 );
and ( n32285 , n32280 , n32284 );
and ( n32286 , n22235 , n23641 );
and ( n32287 , n21955 , n23639 );
nor ( n32288 , n32286 , n32287 );
xnor ( n32289 , n32288 , n23213 );
and ( n32290 , n32285 , n32289 );
and ( n32291 , n29318 , n19688 );
and ( n32292 , n29078 , n19686 );
nor ( n32293 , n32291 , n32292 );
xnor ( n32294 , n32293 , n19655 );
and ( n32295 , n32289 , n32294 );
and ( n32296 , n32285 , n32294 );
or ( n32297 , n32290 , n32295 , n32296 );
and ( n32298 , n19825 , n28628 );
and ( n32299 , n19811 , n28626 );
nor ( n32300 , n32298 , n32299 );
xnor ( n32301 , n32300 , n28096 );
and ( n32302 , n32297 , n32301 );
xor ( n32303 , n31804 , n31808 );
xor ( n32304 , n32303 , n31812 );
and ( n32305 , n32301 , n32304 );
and ( n32306 , n32297 , n32304 );
or ( n32307 , n32302 , n32305 , n32306 );
xor ( n32308 , n31819 , n31823 );
xor ( n32309 , n32308 , n31828 );
xor ( n32310 , n31764 , n31768 );
xor ( n32311 , n32310 , n31773 );
and ( n32312 , n32309 , n32311 );
xor ( n32313 , n31847 , n31851 );
xor ( n32314 , n32313 , n31856 );
and ( n32315 , n32311 , n32314 );
and ( n32316 , n32309 , n32314 );
or ( n32317 , n32312 , n32315 , n32316 );
and ( n32318 , n32307 , n32317 );
xor ( n32319 , n32074 , n32076 );
xor ( n32320 , n32319 , n32079 );
and ( n32321 , n32317 , n32320 );
and ( n32322 , n32307 , n32320 );
or ( n32323 , n32318 , n32321 , n32322 );
and ( n32324 , n32276 , n32323 );
xor ( n32325 , n31871 , n31873 );
xor ( n32326 , n32325 , n31876 );
and ( n32327 , n32323 , n32326 );
and ( n32328 , n32276 , n32326 );
or ( n32329 , n32324 , n32327 , n32328 );
and ( n32330 , n20182 , n27529 );
and ( n32331 , n20080 , n27527 );
nor ( n32332 , n32330 , n32331 );
xnor ( n32333 , n32332 , n27034 );
and ( n32334 , n20618 , n26349 );
and ( n32335 , n20452 , n26347 );
nor ( n32336 , n32334 , n32335 );
xnor ( n32337 , n32336 , n25893 );
and ( n32338 , n32333 , n32337 );
and ( n32339 , n21876 , n23944 );
and ( n32340 , n21704 , n23942 );
nor ( n32341 , n32339 , n32340 );
xnor ( n32342 , n32341 , n23550 );
and ( n32343 , n32337 , n32342 );
and ( n32344 , n32333 , n32342 );
or ( n32345 , n32338 , n32343 , n32344 );
and ( n32346 , n20803 , n26027 );
and ( n32347 , n20666 , n26025 );
nor ( n32348 , n32346 , n32347 );
xnor ( n32349 , n32348 , n25499 );
and ( n32350 , n21072 , n25383 );
and ( n32351 , n20867 , n25381 );
nor ( n32352 , n32350 , n32351 );
xnor ( n32353 , n32352 , n24885 );
and ( n32354 , n32349 , n32353 );
xor ( n32355 , n32043 , n32047 );
xor ( n32356 , n32355 , n32052 );
and ( n32357 , n32353 , n32356 );
and ( n32358 , n32349 , n32356 );
or ( n32359 , n32354 , n32357 , n32358 );
and ( n32360 , n32345 , n32359 );
xor ( n32361 , n31780 , n31784 );
xor ( n32362 , n32361 , n31789 );
and ( n32363 , n32359 , n32362 );
and ( n32364 , n32345 , n32362 );
or ( n32365 , n32360 , n32363 , n32364 );
and ( n32366 , n20360 , n26992 );
and ( n32367 , n20268 , n26990 );
nor ( n32368 , n32366 , n32367 );
xnor ( n32369 , n32368 , n26369 );
and ( n32370 , n21302 , n24902 );
and ( n32371 , n21218 , n24900 );
nor ( n32372 , n32370 , n32371 );
xnor ( n32373 , n32372 , n24397 );
and ( n32374 , n32369 , n32373 );
and ( n32375 , n21612 , n24376 );
and ( n32376 , n21451 , n24374 );
nor ( n32377 , n32375 , n32376 );
xnor ( n32378 , n32377 , n23927 );
and ( n32379 , n32373 , n32378 );
and ( n32380 , n32369 , n32378 );
or ( n32381 , n32374 , n32379 , n32380 );
xor ( n32382 , n32158 , n32162 );
xor ( n32383 , n32382 , n32167 );
and ( n32384 , n32381 , n32383 );
xor ( n32385 , n32055 , n32059 );
xor ( n32386 , n32385 , n32064 );
and ( n32387 , n32383 , n32386 );
and ( n32388 , n32381 , n32386 );
or ( n32389 , n32384 , n32387 , n32388 );
and ( n32390 , n32365 , n32389 );
xor ( n32391 , n31948 , n31950 );
xor ( n32392 , n32391 , n31953 );
and ( n32393 , n32389 , n32392 );
and ( n32394 , n32365 , n32392 );
or ( n32395 , n32390 , n32393 , n32394 );
xor ( n32396 , n31956 , n31958 );
xor ( n32397 , n32396 , n31961 );
and ( n32398 , n32395 , n32397 );
xor ( n32399 , n32070 , n32082 );
xor ( n32400 , n32399 , n32085 );
and ( n32401 , n32397 , n32400 );
and ( n32402 , n32395 , n32400 );
or ( n32403 , n32398 , n32401 , n32402 );
and ( n32404 , n32329 , n32403 );
xor ( n32405 , n32088 , n32090 );
xor ( n32406 , n32405 , n32093 );
and ( n32407 , n32403 , n32406 );
and ( n32408 , n32329 , n32406 );
or ( n32409 , n32404 , n32407 , n32408 );
and ( n32410 , n26851 , n20460 );
and ( n32411 , n26422 , n20458 );
nor ( n32412 , n32410 , n32411 );
xnor ( n32413 , n32412 , n20337 );
and ( n32414 , n27352 , n20276 );
and ( n32415 , n27135 , n20274 );
nor ( n32416 , n32414 , n32415 );
xnor ( n32417 , n32416 , n20175 );
and ( n32418 , n32413 , n32417 );
and ( n32419 , n27757 , n20114 );
and ( n32420 , n27751 , n20112 );
nor ( n32421 , n32419 , n32420 );
xnor ( n32422 , n32421 , n19997 );
and ( n32423 , n32417 , n32422 );
and ( n32424 , n32413 , n32422 );
or ( n32425 , n32418 , n32423 , n32424 );
and ( n32426 , n25284 , n21155 );
and ( n32427 , n24940 , n21153 );
nor ( n32428 , n32426 , n32427 );
xnor ( n32429 , n32428 , n20994 );
and ( n32430 , n25765 , n20955 );
and ( n32431 , n25554 , n20953 );
nor ( n32432 , n32430 , n32431 );
xnor ( n32433 , n32432 , n20780 );
and ( n32434 , n32429 , n32433 );
and ( n32435 , n26319 , n20674 );
and ( n32436 , n25974 , n20672 );
nor ( n32437 , n32435 , n32436 );
xnor ( n32438 , n32437 , n20542 );
and ( n32439 , n32433 , n32438 );
and ( n32440 , n32429 , n32438 );
or ( n32441 , n32434 , n32439 , n32440 );
and ( n32442 , n32425 , n32441 );
xor ( n32443 , n32280 , n32284 );
and ( n32444 , n28810 , n19894 );
and ( n32445 , n28211 , n19892 );
nor ( n32446 , n32444 , n32445 );
xnor ( n32447 , n32446 , n19858 );
and ( n32448 , n32443 , n32447 );
and ( n32449 , n29078 , n19805 );
and ( n32450 , n28700 , n19803 );
nor ( n32451 , n32449 , n32450 );
xnor ( n32452 , n32451 , n19750 );
and ( n32453 , n32447 , n32452 );
and ( n32454 , n32443 , n32452 );
or ( n32455 , n32448 , n32453 , n32454 );
and ( n32456 , n32441 , n32455 );
and ( n32457 , n32425 , n32455 );
or ( n32458 , n32442 , n32456 , n32457 );
xor ( n32459 , n32174 , n32178 );
xor ( n32460 , n32459 , n31810 );
xor ( n32461 , n32186 , n32190 );
xor ( n32462 , n32461 , n32195 );
and ( n32463 , n32460 , n32462 );
xor ( n32464 , n32285 , n32289 );
xor ( n32465 , n32464 , n32294 );
and ( n32466 , n32462 , n32465 );
and ( n32467 , n32460 , n32465 );
or ( n32468 , n32463 , n32466 , n32467 );
and ( n32469 , n32458 , n32468 );
xor ( n32470 , n32026 , n32030 );
xor ( n32471 , n32470 , n32035 );
and ( n32472 , n32468 , n32471 );
and ( n32473 , n32458 , n32471 );
or ( n32474 , n32469 , n32472 , n32473 );
xor ( n32475 , n32124 , n32126 );
xor ( n32476 , n32475 , n32129 );
and ( n32477 , n32474 , n32476 );
xor ( n32478 , n32170 , n32218 );
xor ( n32479 , n32478 , n32221 );
and ( n32480 , n32476 , n32479 );
and ( n32481 , n32474 , n32479 );
or ( n32482 , n32477 , n32480 , n32481 );
xor ( n32483 , n32132 , n32134 );
xor ( n32484 , n32483 , n32137 );
and ( n32485 , n32482 , n32484 );
xor ( n32486 , n32224 , n32226 );
xor ( n32487 , n32486 , n32229 );
and ( n32488 , n32484 , n32487 );
and ( n32489 , n32482 , n32487 );
or ( n32490 , n32485 , n32488 , n32489 );
xor ( n32491 , n32140 , n32142 );
xor ( n32492 , n32491 , n32145 );
and ( n32493 , n32490 , n32492 );
xor ( n32494 , n32232 , n32234 );
xor ( n32495 , n32494 , n32237 );
and ( n32496 , n32492 , n32495 );
and ( n32497 , n32490 , n32495 );
or ( n32498 , n32493 , n32496 , n32497 );
and ( n32499 , n32409 , n32498 );
xor ( n32500 , n32096 , n32148 );
xor ( n32501 , n32500 , n32151 );
and ( n32502 , n32498 , n32501 );
and ( n32503 , n32409 , n32501 );
or ( n32504 , n32499 , n32502 , n32503 );
xor ( n32505 , n31980 , n31982 );
xor ( n32506 , n32505 , n31985 );
and ( n32507 , n32504 , n32506 );
xor ( n32508 , n32154 , n32248 );
xor ( n32509 , n32508 , n32251 );
and ( n32510 , n32506 , n32509 );
and ( n32511 , n32504 , n32509 );
or ( n32512 , n32507 , n32510 , n32511 );
and ( n32513 , n32266 , n32512 );
xor ( n32514 , n32266 , n32512 );
xor ( n32515 , n32504 , n32506 );
xor ( n32516 , n32515 , n32509 );
and ( n32517 , n19637 , n29977 );
and ( n32518 , n19605 , n29974 );
nor ( n32519 , n32517 , n32518 );
xnor ( n32520 , n32519 , n28674 );
and ( n32521 , n19811 , n29276 );
and ( n32522 , n19721 , n29274 );
nor ( n32523 , n32521 , n32522 );
xnor ( n32524 , n32523 , n28677 );
and ( n32525 , n32520 , n32524 );
and ( n32526 , n19881 , n28628 );
and ( n32527 , n19825 , n28626 );
nor ( n32528 , n32526 , n32527 );
xnor ( n32529 , n32528 , n28096 );
and ( n32530 , n32524 , n32529 );
and ( n32531 , n32520 , n32529 );
or ( n32532 , n32525 , n32530 , n32531 );
and ( n32533 , n22198 , n23641 );
and ( n32534 , n22235 , n23639 );
nor ( n32535 , n32533 , n32534 );
xnor ( n32536 , n32535 , n23213 );
and ( n32537 , n23141 , n22859 );
and ( n32538 , n22916 , n22857 );
nor ( n32539 , n32537 , n32538 );
xnor ( n32540 , n32539 , n22418 );
and ( n32541 , n32536 , n32540 );
and ( n32542 , n29623 , n19686 );
not ( n32543 , n32542 );
and ( n32544 , n32543 , n19655 );
and ( n32545 , n32540 , n32544 );
and ( n32546 , n32536 , n32544 );
or ( n32547 , n32541 , n32545 , n32546 );
and ( n32548 , n23968 , n22048 );
and ( n32549 , n23573 , n22046 );
nor ( n32550 , n32548 , n32549 );
xnor ( n32551 , n32550 , n21853 );
and ( n32552 , n24521 , n21741 );
and ( n32553 , n24131 , n21739 );
nor ( n32554 , n32552 , n32553 );
xnor ( n32555 , n32554 , n21605 );
and ( n32556 , n32551 , n32555 );
and ( n32557 , n24621 , n21468 );
and ( n32558 , n24527 , n21466 );
nor ( n32559 , n32557 , n32558 );
xnor ( n32560 , n32559 , n21331 );
and ( n32561 , n32555 , n32560 );
and ( n32562 , n32551 , n32560 );
or ( n32563 , n32556 , n32561 , n32562 );
and ( n32564 , n32547 , n32563 );
and ( n32565 , n20004 , n28062 );
and ( n32566 , n19946 , n28060 );
nor ( n32567 , n32565 , n32566 );
xnor ( n32568 , n32567 , n27549 );
and ( n32569 , n32563 , n32568 );
and ( n32570 , n32547 , n32568 );
or ( n32571 , n32564 , n32569 , n32570 );
and ( n32572 , n32532 , n32571 );
xor ( n32573 , n32010 , n32014 );
xor ( n32574 , n32573 , n32019 );
and ( n32575 , n32571 , n32574 );
and ( n32576 , n32532 , n32574 );
or ( n32577 , n32572 , n32575 , n32576 );
xor ( n32578 , n32112 , n32116 );
xor ( n32579 , n32578 , n32121 );
xor ( n32580 , n32182 , n32198 );
xor ( n32581 , n32580 , n32215 );
and ( n32582 , n32579 , n32581 );
xor ( n32583 , n32297 , n32301 );
xor ( n32584 , n32583 , n32304 );
and ( n32585 , n32581 , n32584 );
and ( n32586 , n32579 , n32584 );
or ( n32587 , n32582 , n32585 , n32586 );
and ( n32588 , n32577 , n32587 );
xor ( n32589 , n32022 , n32038 );
xor ( n32590 , n32589 , n32067 );
and ( n32591 , n32587 , n32590 );
and ( n32592 , n32577 , n32590 );
or ( n32593 , n32588 , n32591 , n32592 );
and ( n32594 , n20080 , n28062 );
and ( n32595 , n20004 , n28060 );
nor ( n32596 , n32594 , n32595 );
xnor ( n32597 , n32596 , n27549 );
and ( n32598 , n20666 , n26349 );
and ( n32599 , n20618 , n26347 );
nor ( n32600 , n32598 , n32599 );
xnor ( n32601 , n32600 , n25893 );
and ( n32602 , n32597 , n32601 );
and ( n32603 , n21955 , n23944 );
and ( n32604 , n21876 , n23942 );
nor ( n32605 , n32603 , n32604 );
xnor ( n32606 , n32605 , n23550 );
and ( n32607 , n32601 , n32606 );
and ( n32608 , n32597 , n32606 );
or ( n32609 , n32602 , n32607 , n32608 );
and ( n32610 , n20452 , n26992 );
and ( n32611 , n20360 , n26990 );
nor ( n32612 , n32610 , n32611 );
xnor ( n32613 , n32612 , n26369 );
and ( n32614 , n21451 , n24902 );
and ( n32615 , n21302 , n24900 );
nor ( n32616 , n32614 , n32615 );
xnor ( n32617 , n32616 , n24397 );
and ( n32618 , n32613 , n32617 );
and ( n32619 , n21704 , n24376 );
and ( n32620 , n21612 , n24374 );
nor ( n32621 , n32619 , n32620 );
xnor ( n32622 , n32621 , n23927 );
and ( n32623 , n32617 , n32622 );
and ( n32624 , n32613 , n32622 );
or ( n32625 , n32618 , n32623 , n32624 );
and ( n32626 , n32609 , n32625 );
and ( n32627 , n22425 , n23641 );
and ( n32628 , n22198 , n23639 );
nor ( n32629 , n32627 , n32628 );
xnor ( n32630 , n32629 , n23213 );
and ( n32631 , n22916 , n23230 );
and ( n32632 , n22756 , n23228 );
nor ( n32633 , n32631 , n32632 );
xnor ( n32634 , n32633 , n22842 );
and ( n32635 , n32630 , n32634 );
and ( n32636 , n23573 , n22381 );
and ( n32637 , n23381 , n22379 );
nor ( n32638 , n32636 , n32637 );
xnor ( n32639 , n32638 , n22228 );
and ( n32640 , n32634 , n32639 );
and ( n32641 , n32630 , n32639 );
or ( n32642 , n32635 , n32640 , n32641 );
and ( n32643 , n29623 , n19688 );
and ( n32644 , n29318 , n19686 );
nor ( n32645 , n32643 , n32644 );
xnor ( n32646 , n32645 , n19655 );
and ( n32647 , n32642 , n32646 );
xor ( n32648 , n32536 , n32540 );
xor ( n32649 , n32648 , n32544 );
and ( n32650 , n32646 , n32649 );
and ( n32651 , n32642 , n32649 );
or ( n32652 , n32647 , n32650 , n32651 );
and ( n32653 , n32625 , n32652 );
and ( n32654 , n32609 , n32652 );
or ( n32655 , n32626 , n32653 , n32654 );
and ( n32656 , n20268 , n27529 );
and ( n32657 , n20182 , n27527 );
nor ( n32658 , n32656 , n32657 );
xnor ( n32659 , n32658 , n27034 );
and ( n32660 , n20867 , n26027 );
and ( n32661 , n20803 , n26025 );
nor ( n32662 , n32660 , n32661 );
xnor ( n32663 , n32662 , n25499 );
and ( n32664 , n32659 , n32663 );
and ( n32665 , n21218 , n25383 );
and ( n32666 , n21072 , n25381 );
nor ( n32667 , n32665 , n32666 );
xnor ( n32668 , n32667 , n24885 );
and ( n32669 , n32663 , n32668 );
and ( n32670 , n32659 , n32668 );
or ( n32671 , n32664 , n32669 , n32670 );
xor ( n32672 , n32203 , n32207 );
xor ( n32673 , n32672 , n32212 );
and ( n32674 , n32671 , n32673 );
xor ( n32675 , n32100 , n32104 );
xor ( n32676 , n32675 , n32109 );
and ( n32677 , n32673 , n32676 );
and ( n32678 , n32671 , n32676 );
or ( n32679 , n32674 , n32677 , n32678 );
and ( n32680 , n32655 , n32679 );
xor ( n32681 , n32309 , n32311 );
xor ( n32682 , n32681 , n32314 );
and ( n32683 , n32679 , n32682 );
and ( n32684 , n32655 , n32682 );
or ( n32685 , n32680 , n32683 , n32684 );
xor ( n32686 , n32268 , n32270 );
xor ( n32687 , n32686 , n32273 );
and ( n32688 , n32685 , n32687 );
xor ( n32689 , n32307 , n32317 );
xor ( n32690 , n32689 , n32320 );
and ( n32691 , n32687 , n32690 );
and ( n32692 , n32685 , n32690 );
or ( n32693 , n32688 , n32691 , n32692 );
and ( n32694 , n32593 , n32693 );
xor ( n32695 , n32276 , n32323 );
xor ( n32696 , n32695 , n32326 );
and ( n32697 , n32693 , n32696 );
and ( n32698 , n32593 , n32696 );
or ( n32699 , n32694 , n32697 , n32698 );
and ( n32700 , n27751 , n20276 );
and ( n32701 , n27352 , n20274 );
nor ( n32702 , n32700 , n32701 );
xnor ( n32703 , n32702 , n20175 );
and ( n32704 , n28211 , n20114 );
and ( n32705 , n27757 , n20112 );
nor ( n32706 , n32704 , n32705 );
xnor ( n32707 , n32706 , n19997 );
and ( n32708 , n32703 , n32707 );
and ( n32709 , n28700 , n19894 );
and ( n32710 , n28810 , n19892 );
nor ( n32711 , n32709 , n32710 );
xnor ( n32712 , n32711 , n19858 );
and ( n32713 , n32707 , n32712 );
and ( n32714 , n32703 , n32712 );
or ( n32715 , n32708 , n32713 , n32714 );
and ( n32716 , n19721 , n29977 );
and ( n32717 , n19637 , n29974 );
nor ( n32718 , n32716 , n32717 );
xnor ( n32719 , n32718 , n28674 );
and ( n32720 , n32715 , n32719 );
and ( n32721 , n19946 , n28628 );
and ( n32722 , n19881 , n28626 );
nor ( n32723 , n32721 , n32722 );
xnor ( n32724 , n32723 , n28096 );
and ( n32725 , n32719 , n32724 );
and ( n32726 , n32715 , n32724 );
or ( n32727 , n32720 , n32725 , n32726 );
and ( n32728 , n24527 , n21741 );
and ( n32729 , n24521 , n21739 );
nor ( n32730 , n32728 , n32729 );
xnor ( n32731 , n32730 , n21605 );
and ( n32732 , n24940 , n21468 );
and ( n32733 , n24621 , n21466 );
nor ( n32734 , n32732 , n32733 );
xnor ( n32735 , n32734 , n21331 );
and ( n32736 , n32731 , n32735 );
and ( n32737 , n25554 , n21155 );
and ( n32738 , n25284 , n21153 );
nor ( n32739 , n32737 , n32738 );
xnor ( n32740 , n32739 , n20994 );
and ( n32741 , n32735 , n32740 );
and ( n32742 , n32731 , n32740 );
or ( n32743 , n32736 , n32741 , n32742 );
and ( n32744 , n25974 , n20955 );
and ( n32745 , n25765 , n20953 );
nor ( n32746 , n32744 , n32745 );
xnor ( n32747 , n32746 , n20780 );
and ( n32748 , n26422 , n20674 );
and ( n32749 , n26319 , n20672 );
nor ( n32750 , n32748 , n32749 );
xnor ( n32751 , n32750 , n20542 );
and ( n32752 , n32747 , n32751 );
and ( n32753 , n27135 , n20460 );
and ( n32754 , n26851 , n20458 );
nor ( n32755 , n32753 , n32754 );
xnor ( n32756 , n32755 , n20337 );
and ( n32757 , n32751 , n32756 );
and ( n32758 , n32747 , n32756 );
or ( n32759 , n32752 , n32757 , n32758 );
and ( n32760 , n32743 , n32759 );
and ( n32761 , n19825 , n29276 );
and ( n32762 , n19811 , n29274 );
nor ( n32763 , n32761 , n32762 );
xnor ( n32764 , n32763 , n28677 );
and ( n32765 , n32759 , n32764 );
and ( n32766 , n32743 , n32764 );
or ( n32767 , n32760 , n32765 , n32766 );
and ( n32768 , n32727 , n32767 );
xor ( n32769 , n32333 , n32337 );
xor ( n32770 , n32769 , n32342 );
and ( n32771 , n32767 , n32770 );
and ( n32772 , n32727 , n32770 );
or ( n32773 , n32768 , n32771 , n32772 );
xor ( n32774 , n32345 , n32359 );
xor ( n32775 , n32774 , n32362 );
and ( n32776 , n32773 , n32775 );
xor ( n32777 , n32381 , n32383 );
xor ( n32778 , n32777 , n32386 );
and ( n32779 , n32775 , n32778 );
and ( n32780 , n32773 , n32778 );
or ( n32781 , n32776 , n32779 , n32780 );
xor ( n32782 , n32577 , n32587 );
xor ( n32783 , n32782 , n32590 );
and ( n32784 , n32781 , n32783 );
xor ( n32785 , n32365 , n32389 );
xor ( n32786 , n32785 , n32392 );
and ( n32787 , n32783 , n32786 );
and ( n32788 , n32781 , n32786 );
or ( n32789 , n32784 , n32787 , n32788 );
and ( n32790 , n23271 , n22859 );
and ( n32791 , n23141 , n22857 );
nor ( n32792 , n32790 , n32791 );
xnor ( n32793 , n32792 , n22418 );
and ( n32794 , n24131 , n22048 );
and ( n32795 , n23968 , n22046 );
nor ( n32796 , n32794 , n32795 );
xnor ( n32797 , n32796 , n21853 );
and ( n32798 , n32793 , n32797 );
and ( n32799 , n32797 , n32542 );
and ( n32800 , n32793 , n32542 );
or ( n32801 , n32798 , n32799 , n32800 );
and ( n32802 , n22756 , n23641 );
and ( n32803 , n22425 , n23639 );
nor ( n32804 , n32802 , n32803 );
xnor ( n32805 , n32804 , n23213 );
and ( n32806 , n23968 , n22381 );
and ( n32807 , n23573 , n22379 );
nor ( n32808 , n32806 , n32807 );
xnor ( n32809 , n32808 , n22228 );
and ( n32810 , n32805 , n32809 );
and ( n32811 , n22235 , n23944 );
and ( n32812 , n21955 , n23942 );
nor ( n32813 , n32811 , n32812 );
xnor ( n32814 , n32813 , n23550 );
and ( n32815 , n32810 , n32814 );
and ( n32816 , n29318 , n19805 );
and ( n32817 , n29078 , n19803 );
nor ( n32818 , n32816 , n32817 );
xnor ( n32819 , n32818 , n19750 );
and ( n32820 , n32814 , n32819 );
and ( n32821 , n32810 , n32819 );
or ( n32822 , n32815 , n32820 , n32821 );
and ( n32823 , n32801 , n32822 );
xor ( n32824 , n32443 , n32447 );
xor ( n32825 , n32824 , n32452 );
and ( n32826 , n32822 , n32825 );
and ( n32827 , n32801 , n32825 );
or ( n32828 , n32823 , n32826 , n32827 );
xor ( n32829 , n32369 , n32373 );
xor ( n32830 , n32829 , n32378 );
and ( n32831 , n32828 , n32830 );
xor ( n32832 , n32349 , n32353 );
xor ( n32833 , n32832 , n32356 );
and ( n32834 , n32830 , n32833 );
and ( n32835 , n32828 , n32833 );
or ( n32836 , n32831 , n32834 , n32835 );
xor ( n32837 , n32532 , n32571 );
xor ( n32838 , n32837 , n32574 );
and ( n32839 , n32836 , n32838 );
xor ( n32840 , n32458 , n32468 );
xor ( n32841 , n32840 , n32471 );
and ( n32842 , n32838 , n32841 );
and ( n32843 , n32836 , n32841 );
or ( n32844 , n32839 , n32842 , n32843 );
xor ( n32845 , n32520 , n32524 );
xor ( n32846 , n32845 , n32529 );
xor ( n32847 , n32547 , n32563 );
xor ( n32848 , n32847 , n32568 );
and ( n32849 , n32846 , n32848 );
xor ( n32850 , n32425 , n32441 );
xor ( n32851 , n32850 , n32455 );
and ( n32852 , n32848 , n32851 );
and ( n32853 , n32846 , n32851 );
or ( n32854 , n32849 , n32852 , n32853 );
and ( n32855 , n21302 , n25383 );
and ( n32856 , n21218 , n25381 );
nor ( n32857 , n32855 , n32856 );
xnor ( n32858 , n32857 , n24885 );
and ( n32859 , n21612 , n24902 );
and ( n32860 , n21451 , n24900 );
nor ( n32861 , n32859 , n32860 );
xnor ( n32862 , n32861 , n24397 );
and ( n32863 , n32858 , n32862 );
and ( n32864 , n21876 , n24376 );
and ( n32865 , n21704 , n24374 );
nor ( n32866 , n32864 , n32865 );
xnor ( n32867 , n32866 , n23927 );
and ( n32868 , n32862 , n32867 );
and ( n32869 , n32858 , n32867 );
or ( n32870 , n32863 , n32868 , n32869 );
and ( n32871 , n23141 , n23230 );
and ( n32872 , n22916 , n23228 );
nor ( n32873 , n32871 , n32872 );
xnor ( n32874 , n32873 , n22842 );
and ( n32875 , n23381 , n22859 );
and ( n32876 , n23271 , n22857 );
nor ( n32877 , n32875 , n32876 );
xnor ( n32878 , n32877 , n22418 );
and ( n32879 , n32874 , n32878 );
and ( n32880 , n29623 , n19803 );
not ( n32881 , n32880 );
and ( n32882 , n32881 , n19750 );
and ( n32883 , n32878 , n32882 );
and ( n32884 , n32874 , n32882 );
or ( n32885 , n32879 , n32883 , n32884 );
and ( n32886 , n20360 , n27529 );
and ( n32887 , n20268 , n27527 );
nor ( n32888 , n32886 , n32887 );
xnor ( n32889 , n32888 , n27034 );
and ( n32890 , n32885 , n32889 );
and ( n32891 , n21072 , n26027 );
and ( n32892 , n20867 , n26025 );
nor ( n32893 , n32891 , n32892 );
xnor ( n32894 , n32893 , n25499 );
and ( n32895 , n32889 , n32894 );
and ( n32896 , n32885 , n32894 );
or ( n32897 , n32890 , n32895 , n32896 );
and ( n32898 , n32870 , n32897 );
and ( n32899 , n20182 , n28062 );
and ( n32900 , n20080 , n28060 );
nor ( n32901 , n32899 , n32900 );
xnor ( n32902 , n32901 , n27549 );
and ( n32903 , n20618 , n26992 );
and ( n32904 , n20452 , n26990 );
nor ( n32905 , n32903 , n32904 );
xnor ( n32906 , n32905 , n26369 );
and ( n32907 , n32902 , n32906 );
xor ( n32908 , n32630 , n32634 );
xor ( n32909 , n32908 , n32639 );
and ( n32910 , n32906 , n32909 );
and ( n32911 , n32902 , n32909 );
or ( n32912 , n32907 , n32910 , n32911 );
and ( n32913 , n32897 , n32912 );
and ( n32914 , n32870 , n32912 );
or ( n32915 , n32898 , n32913 , n32914 );
xor ( n32916 , n32551 , n32555 );
xor ( n32917 , n32916 , n32560 );
xor ( n32918 , n32413 , n32417 );
xor ( n32919 , n32918 , n32422 );
and ( n32920 , n32917 , n32919 );
xor ( n32921 , n32429 , n32433 );
xor ( n32922 , n32921 , n32438 );
and ( n32923 , n32919 , n32922 );
and ( n32924 , n32917 , n32922 );
or ( n32925 , n32920 , n32923 , n32924 );
and ( n32926 , n32915 , n32925 );
xor ( n32927 , n32671 , n32673 );
xor ( n32928 , n32927 , n32676 );
and ( n32929 , n32925 , n32928 );
and ( n32930 , n32915 , n32928 );
or ( n32931 , n32926 , n32929 , n32930 );
and ( n32932 , n32854 , n32931 );
xor ( n32933 , n32579 , n32581 );
xor ( n32934 , n32933 , n32584 );
and ( n32935 , n32931 , n32934 );
and ( n32936 , n32854 , n32934 );
or ( n32937 , n32932 , n32935 , n32936 );
and ( n32938 , n32844 , n32937 );
xor ( n32939 , n32474 , n32476 );
xor ( n32940 , n32939 , n32479 );
and ( n32941 , n32937 , n32940 );
and ( n32942 , n32844 , n32940 );
or ( n32943 , n32938 , n32941 , n32942 );
and ( n32944 , n32789 , n32943 );
xor ( n32945 , n32395 , n32397 );
xor ( n32946 , n32945 , n32400 );
and ( n32947 , n32943 , n32946 );
and ( n32948 , n32789 , n32946 );
or ( n32949 , n32944 , n32947 , n32948 );
and ( n32950 , n32699 , n32949 );
xor ( n32951 , n32329 , n32403 );
xor ( n32952 , n32951 , n32406 );
and ( n32953 , n32949 , n32952 );
and ( n32954 , n32699 , n32952 );
or ( n32955 , n32950 , n32953 , n32954 );
xor ( n32956 , n32240 , n32242 );
xor ( n32957 , n32956 , n32245 );
and ( n32958 , n32955 , n32957 );
xor ( n32959 , n32409 , n32498 );
xor ( n32960 , n32959 , n32501 );
and ( n32961 , n32957 , n32960 );
and ( n32962 , n32955 , n32960 );
or ( n32963 , n32958 , n32961 , n32962 );
and ( n32964 , n32516 , n32963 );
xor ( n32965 , n32516 , n32963 );
xor ( n32966 , n32955 , n32957 );
xor ( n32967 , n32966 , n32960 );
and ( n32968 , n25284 , n21468 );
and ( n32969 , n24940 , n21466 );
nor ( n32970 , n32968 , n32969 );
xnor ( n32971 , n32970 , n21331 );
and ( n32972 , n25765 , n21155 );
and ( n32973 , n25554 , n21153 );
nor ( n32974 , n32972 , n32973 );
xnor ( n32975 , n32974 , n20994 );
and ( n32976 , n32971 , n32975 );
and ( n32977 , n26319 , n20955 );
and ( n32978 , n25974 , n20953 );
nor ( n32979 , n32977 , n32978 );
xnor ( n32980 , n32979 , n20780 );
and ( n32981 , n32975 , n32980 );
and ( n32982 , n32971 , n32980 );
or ( n32983 , n32976 , n32981 , n32982 );
and ( n32984 , n19881 , n29276 );
and ( n32985 , n19825 , n29274 );
nor ( n32986 , n32984 , n32985 );
xnor ( n32987 , n32986 , n28677 );
and ( n32988 , n32983 , n32987 );
and ( n32989 , n20803 , n26349 );
and ( n32990 , n20666 , n26347 );
nor ( n32991 , n32989 , n32990 );
xnor ( n32992 , n32991 , n25893 );
and ( n32993 , n32987 , n32992 );
and ( n32994 , n32983 , n32992 );
or ( n32995 , n32988 , n32993 , n32994 );
and ( n32996 , n26851 , n20674 );
and ( n32997 , n26422 , n20672 );
nor ( n32998 , n32996 , n32997 );
xnor ( n32999 , n32998 , n20542 );
and ( n33000 , n27352 , n20460 );
and ( n33001 , n27135 , n20458 );
nor ( n33002 , n33000 , n33001 );
xnor ( n33003 , n33002 , n20337 );
and ( n33004 , n32999 , n33003 );
and ( n33005 , n27757 , n20276 );
and ( n33006 , n27751 , n20274 );
nor ( n33007 , n33005 , n33006 );
xnor ( n33008 , n33007 , n20175 );
and ( n33009 , n33003 , n33008 );
and ( n33010 , n32999 , n33008 );
or ( n33011 , n33004 , n33009 , n33010 );
xor ( n33012 , n32805 , n32809 );
and ( n33013 , n28810 , n20114 );
and ( n33014 , n28211 , n20112 );
nor ( n33015 , n33013 , n33014 );
xnor ( n33016 , n33015 , n19997 );
and ( n33017 , n33012 , n33016 );
and ( n33018 , n29078 , n19894 );
and ( n33019 , n28700 , n19892 );
nor ( n33020 , n33018 , n33019 );
xnor ( n33021 , n33020 , n19858 );
and ( n33022 , n33016 , n33021 );
and ( n33023 , n33012 , n33021 );
or ( n33024 , n33017 , n33022 , n33023 );
and ( n33025 , n33011 , n33024 );
and ( n33026 , n19811 , n29977 );
and ( n33027 , n19721 , n29974 );
nor ( n33028 , n33026 , n33027 );
xnor ( n33029 , n33028 , n28674 );
and ( n33030 , n33024 , n33029 );
and ( n33031 , n33011 , n33029 );
or ( n33032 , n33025 , n33030 , n33031 );
and ( n33033 , n32995 , n33032 );
and ( n33034 , n22198 , n23944 );
and ( n33035 , n22235 , n23942 );
nor ( n33036 , n33034 , n33035 );
xnor ( n33037 , n33036 , n23550 );
and ( n33038 , n24521 , n22048 );
and ( n33039 , n24131 , n22046 );
nor ( n33040 , n33038 , n33039 );
xnor ( n33041 , n33040 , n21853 );
and ( n33042 , n33037 , n33041 );
and ( n33043 , n24621 , n21741 );
and ( n33044 , n24527 , n21739 );
nor ( n33045 , n33043 , n33044 );
xnor ( n33046 , n33045 , n21605 );
and ( n33047 , n33041 , n33046 );
and ( n33048 , n33037 , n33046 );
or ( n33049 , n33042 , n33047 , n33048 );
and ( n33050 , n20004 , n28628 );
and ( n33051 , n19946 , n28626 );
nor ( n33052 , n33050 , n33051 );
xnor ( n33053 , n33052 , n28096 );
and ( n33054 , n33049 , n33053 );
xor ( n33055 , n32793 , n32797 );
xor ( n33056 , n33055 , n32542 );
and ( n33057 , n33053 , n33056 );
and ( n33058 , n33049 , n33056 );
or ( n33059 , n33054 , n33057 , n33058 );
and ( n33060 , n33032 , n33059 );
and ( n33061 , n32995 , n33059 );
or ( n33062 , n33033 , n33060 , n33061 );
xor ( n33063 , n32609 , n32625 );
xor ( n33064 , n33063 , n32652 );
and ( n33065 , n33062 , n33064 );
xor ( n33066 , n32460 , n32462 );
xor ( n33067 , n33066 , n32465 );
and ( n33068 , n33064 , n33067 );
and ( n33069 , n33062 , n33067 );
or ( n33070 , n33065 , n33068 , n33069 );
xor ( n33071 , n32655 , n32679 );
xor ( n33072 , n33071 , n32682 );
and ( n33073 , n33070 , n33072 );
xor ( n33074 , n32773 , n32775 );
xor ( n33075 , n33074 , n32778 );
and ( n33076 , n33072 , n33075 );
and ( n33077 , n33070 , n33075 );
or ( n33078 , n33073 , n33076 , n33077 );
xor ( n33079 , n32685 , n32687 );
xor ( n33080 , n33079 , n32690 );
and ( n33081 , n33078 , n33080 );
xor ( n33082 , n32781 , n32783 );
xor ( n33083 , n33082 , n32786 );
and ( n33084 , n33080 , n33083 );
and ( n33085 , n33078 , n33083 );
or ( n33086 , n33081 , n33084 , n33085 );
xor ( n33087 , n32482 , n32484 );
xor ( n33088 , n33087 , n32487 );
and ( n33089 , n33086 , n33088 );
xor ( n33090 , n32593 , n32693 );
xor ( n33091 , n33090 , n32696 );
and ( n33092 , n33088 , n33091 );
and ( n33093 , n33086 , n33091 );
or ( n33094 , n33089 , n33092 , n33093 );
xor ( n33095 , n32490 , n32492 );
xor ( n33096 , n33095 , n32495 );
and ( n33097 , n33094 , n33096 );
xor ( n33098 , n32699 , n32949 );
xor ( n33099 , n33098 , n32952 );
and ( n33100 , n33096 , n33099 );
and ( n33101 , n33094 , n33099 );
or ( n33102 , n33097 , n33100 , n33101 );
and ( n33103 , n32967 , n33102 );
xor ( n33104 , n32967 , n33102 );
xor ( n33105 , n33094 , n33096 );
xor ( n33106 , n33105 , n33099 );
and ( n33107 , n20268 , n28062 );
and ( n33108 , n20182 , n28060 );
nor ( n33109 , n33107 , n33108 );
xnor ( n33110 , n33109 , n27549 );
and ( n33111 , n21218 , n26027 );
and ( n33112 , n21072 , n26025 );
nor ( n33113 , n33111 , n33112 );
xnor ( n33114 , n33113 , n25499 );
and ( n33115 , n33110 , n33114 );
and ( n33116 , n21451 , n25383 );
and ( n33117 , n21302 , n25381 );
nor ( n33118 , n33116 , n33117 );
xnor ( n33119 , n33118 , n24885 );
and ( n33120 , n33114 , n33119 );
and ( n33121 , n33110 , n33119 );
or ( n33122 , n33115 , n33120 , n33121 );
xor ( n33123 , n32703 , n32707 );
xor ( n33124 , n33123 , n32712 );
and ( n33125 , n33122 , n33124 );
xor ( n33126 , n32747 , n32751 );
xor ( n33127 , n33126 , n32756 );
and ( n33128 , n33124 , n33127 );
and ( n33129 , n33122 , n33127 );
or ( n33130 , n33125 , n33128 , n33129 );
xor ( n33131 , n32715 , n32719 );
xor ( n33132 , n33131 , n32724 );
and ( n33133 , n33130 , n33132 );
xor ( n33134 , n32917 , n32919 );
xor ( n33135 , n33134 , n32922 );
and ( n33136 , n33132 , n33135 );
and ( n33137 , n33130 , n33135 );
or ( n33138 , n33133 , n33136 , n33137 );
xor ( n33139 , n32727 , n32767 );
xor ( n33140 , n33139 , n32770 );
and ( n33141 , n33138 , n33140 );
xor ( n33142 , n32846 , n32848 );
xor ( n33143 , n33142 , n32851 );
and ( n33144 , n33140 , n33143 );
and ( n33145 , n33138 , n33143 );
or ( n33146 , n33141 , n33144 , n33145 );
and ( n33147 , n22425 , n23944 );
and ( n33148 , n22198 , n23942 );
nor ( n33149 , n33147 , n33148 );
xnor ( n33150 , n33149 , n23550 );
and ( n33151 , n23573 , n22859 );
and ( n33152 , n23381 , n22857 );
nor ( n33153 , n33151 , n33152 );
xnor ( n33154 , n33153 , n22418 );
and ( n33155 , n33150 , n33154 );
and ( n33156 , n24131 , n22381 );
and ( n33157 , n23968 , n22379 );
nor ( n33158 , n33156 , n33157 );
xnor ( n33159 , n33158 , n22228 );
and ( n33160 , n33154 , n33159 );
and ( n33161 , n33150 , n33159 );
or ( n33162 , n33155 , n33160 , n33161 );
and ( n33163 , n23968 , n22859 );
and ( n33164 , n23573 , n22857 );
nor ( n33165 , n33163 , n33164 );
xnor ( n33166 , n33165 , n22418 );
and ( n33167 , n24521 , n22381 );
and ( n33168 , n24131 , n22379 );
nor ( n33169 , n33167 , n33168 );
xnor ( n33170 , n33169 , n22228 );
and ( n33171 , n33166 , n33170 );
and ( n33172 , n22916 , n23641 );
and ( n33173 , n22756 , n23639 );
nor ( n33174 , n33172 , n33173 );
xnor ( n33175 , n33174 , n23213 );
and ( n33176 , n33171 , n33175 );
and ( n33177 , n33175 , n32880 );
and ( n33178 , n33171 , n32880 );
or ( n33179 , n33176 , n33177 , n33178 );
and ( n33180 , n33162 , n33179 );
and ( n33181 , n29623 , n19805 );
and ( n33182 , n29318 , n19803 );
nor ( n33183 , n33181 , n33182 );
xnor ( n33184 , n33183 , n19750 );
and ( n33185 , n33179 , n33184 );
and ( n33186 , n33162 , n33184 );
or ( n33187 , n33180 , n33185 , n33186 );
xor ( n33188 , n32731 , n32735 );
xor ( n33189 , n33188 , n32740 );
and ( n33190 , n33187 , n33189 );
xor ( n33191 , n32810 , n32814 );
xor ( n33192 , n33191 , n32819 );
and ( n33193 , n33189 , n33192 );
and ( n33194 , n33187 , n33192 );
or ( n33195 , n33190 , n33193 , n33194 );
xor ( n33196 , n32613 , n32617 );
xor ( n33197 , n33196 , n32622 );
and ( n33198 , n33195 , n33197 );
xor ( n33199 , n32743 , n32759 );
xor ( n33200 , n33199 , n32764 );
and ( n33201 , n33197 , n33200 );
and ( n33202 , n33195 , n33200 );
or ( n33203 , n33198 , n33201 , n33202 );
xor ( n33204 , n32659 , n32663 );
xor ( n33205 , n33204 , n32668 );
xor ( n33206 , n32597 , n32601 );
xor ( n33207 , n33206 , n32606 );
and ( n33208 , n33205 , n33207 );
xor ( n33209 , n32642 , n32646 );
xor ( n33210 , n33209 , n32649 );
and ( n33211 , n33207 , n33210 );
and ( n33212 , n33205 , n33210 );
or ( n33213 , n33208 , n33211 , n33212 );
and ( n33214 , n33203 , n33213 );
xor ( n33215 , n32828 , n32830 );
xor ( n33216 , n33215 , n32833 );
and ( n33217 , n33213 , n33216 );
and ( n33218 , n33203 , n33216 );
or ( n33219 , n33214 , n33217 , n33218 );
and ( n33220 , n33146 , n33219 );
xor ( n33221 , n32836 , n32838 );
xor ( n33222 , n33221 , n32841 );
and ( n33223 , n33219 , n33222 );
and ( n33224 , n33146 , n33222 );
or ( n33225 , n33220 , n33223 , n33224 );
and ( n33226 , n27135 , n20674 );
and ( n33227 , n26851 , n20672 );
nor ( n33228 , n33226 , n33227 );
xnor ( n33229 , n33228 , n20542 );
and ( n33230 , n27751 , n20460 );
and ( n33231 , n27352 , n20458 );
nor ( n33232 , n33230 , n33231 );
xnor ( n33233 , n33232 , n20337 );
and ( n33234 , n33229 , n33233 );
and ( n33235 , n28700 , n20114 );
and ( n33236 , n28810 , n20112 );
nor ( n33237 , n33235 , n33236 );
xnor ( n33238 , n33237 , n19997 );
and ( n33239 , n33233 , n33238 );
and ( n33240 , n33229 , n33238 );
or ( n33241 , n33234 , n33239 , n33240 );
and ( n33242 , n23271 , n23230 );
and ( n33243 , n23141 , n23228 );
nor ( n33244 , n33242 , n33243 );
xnor ( n33245 , n33244 , n22842 );
and ( n33246 , n24527 , n22048 );
and ( n33247 , n24521 , n22046 );
nor ( n33248 , n33246 , n33247 );
xnor ( n33249 , n33248 , n21853 );
and ( n33250 , n33245 , n33249 );
and ( n33251 , n24940 , n21741 );
and ( n33252 , n24621 , n21739 );
nor ( n33253 , n33251 , n33252 );
xnor ( n33254 , n33253 , n21605 );
and ( n33255 , n33249 , n33254 );
and ( n33256 , n33245 , n33254 );
or ( n33257 , n33250 , n33255 , n33256 );
and ( n33258 , n33241 , n33257 );
and ( n33259 , n19825 , n29977 );
and ( n33260 , n19811 , n29974 );
nor ( n33261 , n33259 , n33260 );
xnor ( n33262 , n33261 , n28674 );
and ( n33263 , n33257 , n33262 );
and ( n33264 , n33241 , n33262 );
or ( n33265 , n33258 , n33263 , n33264 );
xor ( n33266 , n32885 , n32889 );
xor ( n33267 , n33266 , n32894 );
and ( n33268 , n33265 , n33267 );
xor ( n33269 , n32902 , n32906 );
xor ( n33270 , n33269 , n32909 );
and ( n33271 , n33267 , n33270 );
and ( n33272 , n33265 , n33270 );
or ( n33273 , n33268 , n33271 , n33272 );
xor ( n33274 , n32870 , n32897 );
xor ( n33275 , n33274 , n32912 );
and ( n33276 , n33273 , n33275 );
xor ( n33277 , n32801 , n32822 );
xor ( n33278 , n33277 , n32825 );
and ( n33279 , n33275 , n33278 );
and ( n33280 , n33273 , n33278 );
or ( n33281 , n33276 , n33279 , n33280 );
and ( n33282 , n20452 , n27529 );
and ( n33283 , n20360 , n27527 );
nor ( n33284 , n33282 , n33283 );
xnor ( n33285 , n33284 , n27034 );
and ( n33286 , n21704 , n24902 );
and ( n33287 , n21612 , n24900 );
nor ( n33288 , n33286 , n33287 );
xnor ( n33289 , n33288 , n24397 );
and ( n33290 , n33285 , n33289 );
and ( n33291 , n21955 , n24376 );
and ( n33292 , n21876 , n24374 );
nor ( n33293 , n33291 , n33292 );
xnor ( n33294 , n33293 , n23927 );
and ( n33295 , n33289 , n33294 );
and ( n33296 , n33285 , n33294 );
or ( n33297 , n33290 , n33295 , n33296 );
and ( n33298 , n25554 , n21468 );
and ( n33299 , n25284 , n21466 );
nor ( n33300 , n33298 , n33299 );
xnor ( n33301 , n33300 , n21331 );
and ( n33302 , n25974 , n21155 );
and ( n33303 , n25765 , n21153 );
nor ( n33304 , n33302 , n33303 );
xnor ( n33305 , n33304 , n20994 );
and ( n33306 , n33301 , n33305 );
and ( n33307 , n26422 , n20955 );
and ( n33308 , n26319 , n20953 );
nor ( n33309 , n33307 , n33308 );
xnor ( n33310 , n33309 , n20780 );
and ( n33311 , n33305 , n33310 );
and ( n33312 , n33301 , n33310 );
or ( n33313 , n33306 , n33311 , n33312 );
and ( n33314 , n19946 , n29276 );
and ( n33315 , n19881 , n29274 );
nor ( n33316 , n33314 , n33315 );
xnor ( n33317 , n33316 , n28677 );
and ( n33318 , n33313 , n33317 );
and ( n33319 , n20666 , n26992 );
and ( n33320 , n20618 , n26990 );
nor ( n33321 , n33319 , n33320 );
xnor ( n33322 , n33321 , n26369 );
and ( n33323 , n33317 , n33322 );
and ( n33324 , n33313 , n33322 );
or ( n33325 , n33318 , n33323 , n33324 );
and ( n33326 , n33297 , n33325 );
and ( n33327 , n20080 , n28628 );
and ( n33328 , n20004 , n28626 );
nor ( n33329 , n33327 , n33328 );
xnor ( n33330 , n33329 , n28096 );
and ( n33331 , n20867 , n26349 );
and ( n33332 , n20803 , n26347 );
nor ( n33333 , n33331 , n33332 );
xnor ( n33334 , n33333 , n25893 );
and ( n33335 , n33330 , n33334 );
xor ( n33336 , n32874 , n32878 );
xor ( n33337 , n33336 , n32882 );
and ( n33338 , n33334 , n33337 );
and ( n33339 , n33330 , n33337 );
or ( n33340 , n33335 , n33338 , n33339 );
and ( n33341 , n33325 , n33340 );
and ( n33342 , n33297 , n33340 );
or ( n33343 , n33326 , n33341 , n33342 );
and ( n33344 , n22235 , n24376 );
and ( n33345 , n21955 , n24374 );
nor ( n33346 , n33344 , n33345 );
xnor ( n33347 , n33346 , n23927 );
and ( n33348 , n28211 , n20276 );
and ( n33349 , n27757 , n20274 );
nor ( n33350 , n33348 , n33349 );
xnor ( n33351 , n33350 , n20175 );
and ( n33352 , n33347 , n33351 );
and ( n33353 , n29318 , n19894 );
and ( n33354 , n29078 , n19892 );
nor ( n33355 , n33353 , n33354 );
xnor ( n33356 , n33355 , n19858 );
and ( n33357 , n33351 , n33356 );
and ( n33358 , n33347 , n33356 );
or ( n33359 , n33352 , n33357 , n33358 );
xor ( n33360 , n32971 , n32975 );
xor ( n33361 , n33360 , n32980 );
and ( n33362 , n33359 , n33361 );
xor ( n33363 , n33012 , n33016 );
xor ( n33364 , n33363 , n33021 );
and ( n33365 , n33361 , n33364 );
and ( n33366 , n33359 , n33364 );
or ( n33367 , n33362 , n33365 , n33366 );
xor ( n33368 , n32858 , n32862 );
xor ( n33369 , n33368 , n32867 );
and ( n33370 , n33367 , n33369 );
xor ( n33371 , n32983 , n32987 );
xor ( n33372 , n33371 , n32992 );
and ( n33373 , n33369 , n33372 );
and ( n33374 , n33367 , n33372 );
or ( n33375 , n33370 , n33373 , n33374 );
and ( n33376 , n33343 , n33375 );
xor ( n33377 , n33205 , n33207 );
xor ( n33378 , n33377 , n33210 );
and ( n33379 , n33375 , n33378 );
and ( n33380 , n33343 , n33378 );
or ( n33381 , n33376 , n33379 , n33380 );
and ( n33382 , n33281 , n33381 );
xor ( n33383 , n32915 , n32925 );
xor ( n33384 , n33383 , n32928 );
and ( n33385 , n33381 , n33384 );
and ( n33386 , n33281 , n33384 );
or ( n33387 , n33382 , n33385 , n33386 );
xor ( n33388 , n32854 , n32931 );
xor ( n33389 , n33388 , n32934 );
and ( n33390 , n33387 , n33389 );
xor ( n33391 , n33070 , n33072 );
xor ( n33392 , n33391 , n33075 );
and ( n33393 , n33389 , n33392 );
and ( n33394 , n33387 , n33392 );
or ( n33395 , n33390 , n33393 , n33394 );
and ( n33396 , n33225 , n33395 );
xor ( n33397 , n32844 , n32937 );
xor ( n33398 , n33397 , n32940 );
and ( n33399 , n33395 , n33398 );
and ( n33400 , n33225 , n33398 );
or ( n33401 , n33396 , n33399 , n33400 );
xor ( n33402 , n32789 , n32943 );
xor ( n33403 , n33402 , n32946 );
and ( n33404 , n33401 , n33403 );
xor ( n33405 , n33086 , n33088 );
xor ( n33406 , n33405 , n33091 );
and ( n33407 , n33403 , n33406 );
and ( n33408 , n33401 , n33406 );
or ( n33409 , n33404 , n33407 , n33408 );
and ( n33410 , n33106 , n33409 );
xor ( n33411 , n33106 , n33409 );
xor ( n33412 , n33401 , n33403 );
xor ( n33413 , n33412 , n33406 );
xor ( n33414 , n33011 , n33024 );
xor ( n33415 , n33414 , n33029 );
xor ( n33416 , n33049 , n33053 );
xor ( n33417 , n33416 , n33056 );
and ( n33418 , n33415 , n33417 );
xor ( n33419 , n33187 , n33189 );
xor ( n33420 , n33419 , n33192 );
and ( n33421 , n33417 , n33420 );
and ( n33422 , n33415 , n33420 );
or ( n33423 , n33418 , n33421 , n33422 );
xor ( n33424 , n32995 , n33032 );
xor ( n33425 , n33424 , n33059 );
and ( n33426 , n33423 , n33425 );
xor ( n33427 , n33195 , n33197 );
xor ( n33428 , n33427 , n33200 );
and ( n33429 , n33425 , n33428 );
and ( n33430 , n33423 , n33428 );
or ( n33431 , n33426 , n33429 , n33430 );
xor ( n33432 , n33062 , n33064 );
xor ( n33433 , n33432 , n33067 );
and ( n33434 , n33431 , n33433 );
xor ( n33435 , n33203 , n33213 );
xor ( n33436 , n33435 , n33216 );
and ( n33437 , n33433 , n33436 );
and ( n33438 , n33431 , n33436 );
or ( n33439 , n33434 , n33437 , n33438 );
and ( n33440 , n21302 , n26027 );
and ( n33441 , n21218 , n26025 );
nor ( n33442 , n33440 , n33441 );
xnor ( n33443 , n33442 , n25499 );
and ( n33444 , n21612 , n25383 );
and ( n33445 , n21451 , n25381 );
nor ( n33446 , n33444 , n33445 );
xnor ( n33447 , n33446 , n24885 );
and ( n33448 , n33443 , n33447 );
and ( n33449 , n21876 , n24902 );
and ( n33450 , n21704 , n24900 );
nor ( n33451 , n33449 , n33450 );
xnor ( n33452 , n33451 , n24397 );
and ( n33453 , n33447 , n33452 );
and ( n33454 , n33443 , n33452 );
or ( n33455 , n33448 , n33453 , n33454 );
xor ( n33456 , n33037 , n33041 );
xor ( n33457 , n33456 , n33046 );
and ( n33458 , n33455 , n33457 );
xor ( n33459 , n32999 , n33003 );
xor ( n33460 , n33459 , n33008 );
and ( n33461 , n33457 , n33460 );
and ( n33462 , n33455 , n33460 );
or ( n33463 , n33458 , n33461 , n33462 );
and ( n33464 , n22198 , n24376 );
and ( n33465 , n22235 , n24374 );
nor ( n33466 , n33464 , n33465 );
xnor ( n33467 , n33466 , n23927 );
and ( n33468 , n23141 , n23641 );
and ( n33469 , n22916 , n23639 );
nor ( n33470 , n33468 , n33469 );
xnor ( n33471 , n33470 , n23213 );
and ( n33472 , n33467 , n33471 );
and ( n33473 , n23381 , n23230 );
and ( n33474 , n23271 , n23228 );
nor ( n33475 , n33473 , n33474 );
xnor ( n33476 , n33475 , n22842 );
and ( n33477 , n33471 , n33476 );
and ( n33478 , n33467 , n33476 );
or ( n33479 , n33472 , n33477 , n33478 );
and ( n33480 , n20803 , n26992 );
and ( n33481 , n20666 , n26990 );
nor ( n33482 , n33480 , n33481 );
xnor ( n33483 , n33482 , n26369 );
and ( n33484 , n33479 , n33483 );
and ( n33485 , n21072 , n26349 );
and ( n33486 , n20867 , n26347 );
nor ( n33487 , n33485 , n33486 );
xnor ( n33488 , n33487 , n25893 );
and ( n33489 , n33483 , n33488 );
and ( n33490 , n33479 , n33488 );
or ( n33491 , n33484 , n33489 , n33490 );
and ( n33492 , n20360 , n28062 );
and ( n33493 , n20268 , n28060 );
nor ( n33494 , n33492 , n33493 );
xnor ( n33495 , n33494 , n27549 );
and ( n33496 , n20618 , n27529 );
and ( n33497 , n20452 , n27527 );
nor ( n33498 , n33496 , n33497 );
xnor ( n33499 , n33498 , n27034 );
and ( n33500 , n33495 , n33499 );
xor ( n33501 , n33171 , n33175 );
xor ( n33502 , n33501 , n32880 );
and ( n33503 , n33499 , n33502 );
and ( n33504 , n33495 , n33502 );
or ( n33505 , n33500 , n33503 , n33504 );
and ( n33506 , n33491 , n33505 );
xor ( n33507 , n33162 , n33179 );
xor ( n33508 , n33507 , n33184 );
and ( n33509 , n33505 , n33508 );
and ( n33510 , n33491 , n33508 );
or ( n33511 , n33506 , n33509 , n33510 );
and ( n33512 , n33463 , n33511 );
xor ( n33513 , n33122 , n33124 );
xor ( n33514 , n33513 , n33127 );
and ( n33515 , n33511 , n33514 );
and ( n33516 , n33463 , n33514 );
or ( n33517 , n33512 , n33515 , n33516 );
xor ( n33518 , n33130 , n33132 );
xor ( n33519 , n33518 , n33135 );
and ( n33520 , n33517 , n33519 );
xor ( n33521 , n33273 , n33275 );
xor ( n33522 , n33521 , n33278 );
and ( n33523 , n33519 , n33522 );
and ( n33524 , n33517 , n33522 );
or ( n33525 , n33520 , n33523 , n33524 );
xor ( n33526 , n33138 , n33140 );
xor ( n33527 , n33526 , n33143 );
and ( n33528 , n33525 , n33527 );
xor ( n33529 , n33281 , n33381 );
xor ( n33530 , n33529 , n33384 );
and ( n33531 , n33527 , n33530 );
and ( n33532 , n33525 , n33530 );
or ( n33533 , n33528 , n33531 , n33532 );
and ( n33534 , n33439 , n33533 );
xor ( n33535 , n33146 , n33219 );
xor ( n33536 , n33535 , n33222 );
and ( n33537 , n33533 , n33536 );
and ( n33538 , n33439 , n33536 );
or ( n33539 , n33534 , n33537 , n33538 );
xor ( n33540 , n33078 , n33080 );
xor ( n33541 , n33540 , n33083 );
and ( n33542 , n33539 , n33541 );
xor ( n33543 , n33225 , n33395 );
xor ( n33544 , n33543 , n33398 );
and ( n33545 , n33541 , n33544 );
and ( n33546 , n33539 , n33544 );
or ( n33547 , n33542 , n33545 , n33546 );
and ( n33548 , n33413 , n33547 );
xor ( n33549 , n33413 , n33547 );
xor ( n33550 , n33539 , n33541 );
xor ( n33551 , n33550 , n33544 );
and ( n33552 , n27757 , n20460 );
and ( n33553 , n27751 , n20458 );
nor ( n33554 , n33552 , n33553 );
xnor ( n33555 , n33554 , n20337 );
and ( n33556 , n28810 , n20276 );
and ( n33557 , n28211 , n20274 );
nor ( n33558 , n33556 , n33557 );
xnor ( n33559 , n33558 , n20175 );
and ( n33560 , n33555 , n33559 );
and ( n33561 , n29078 , n20114 );
and ( n33562 , n28700 , n20112 );
nor ( n33563 , n33561 , n33562 );
xnor ( n33564 , n33563 , n19997 );
and ( n33565 , n33559 , n33564 );
and ( n33566 , n33555 , n33564 );
or ( n33567 , n33560 , n33565 , n33566 );
and ( n33568 , n26319 , n21155 );
and ( n33569 , n25974 , n21153 );
nor ( n33570 , n33568 , n33569 );
xnor ( n33571 , n33570 , n20994 );
and ( n33572 , n26851 , n20955 );
and ( n33573 , n26422 , n20953 );
nor ( n33574 , n33572 , n33573 );
xnor ( n33575 , n33574 , n20780 );
and ( n33576 , n33571 , n33575 );
and ( n33577 , n27352 , n20674 );
and ( n33578 , n27135 , n20672 );
nor ( n33579 , n33577 , n33578 );
xnor ( n33580 , n33579 , n20542 );
and ( n33581 , n33575 , n33580 );
and ( n33582 , n33571 , n33580 );
or ( n33583 , n33576 , n33581 , n33582 );
and ( n33584 , n33567 , n33583 );
and ( n33585 , n20004 , n29276 );
and ( n33586 , n19946 , n29274 );
nor ( n33587 , n33585 , n33586 );
xnor ( n33588 , n33587 , n28677 );
and ( n33589 , n33583 , n33588 );
and ( n33590 , n33567 , n33588 );
or ( n33591 , n33584 , n33589 , n33590 );
xor ( n33592 , n33285 , n33289 );
xor ( n33593 , n33592 , n33294 );
and ( n33594 , n33591 , n33593 );
xor ( n33595 , n33313 , n33317 );
xor ( n33596 , n33595 , n33322 );
and ( n33597 , n33593 , n33596 );
and ( n33598 , n33591 , n33596 );
or ( n33599 , n33594 , n33597 , n33598 );
xor ( n33600 , n33166 , n33170 );
and ( n33601 , n22756 , n23944 );
and ( n33602 , n22425 , n23942 );
nor ( n33603 , n33601 , n33602 );
xnor ( n33604 , n33603 , n23550 );
and ( n33605 , n33600 , n33604 );
and ( n33606 , n29623 , n19892 );
not ( n33607 , n33606 );
and ( n33608 , n33607 , n19858 );
and ( n33609 , n33604 , n33608 );
and ( n33610 , n33600 , n33608 );
or ( n33611 , n33605 , n33609 , n33610 );
and ( n33612 , n20182 , n28628 );
and ( n33613 , n20080 , n28626 );
nor ( n33614 , n33612 , n33613 );
xnor ( n33615 , n33614 , n28096 );
and ( n33616 , n33611 , n33615 );
xor ( n33617 , n33150 , n33154 );
xor ( n33618 , n33617 , n33159 );
and ( n33619 , n33615 , n33618 );
and ( n33620 , n33611 , n33618 );
or ( n33621 , n33616 , n33619 , n33620 );
xor ( n33622 , n33110 , n33114 );
xor ( n33623 , n33622 , n33119 );
and ( n33624 , n33621 , n33623 );
xor ( n33625 , n33330 , n33334 );
xor ( n33626 , n33625 , n33337 );
and ( n33627 , n33623 , n33626 );
and ( n33628 , n33621 , n33626 );
or ( n33629 , n33624 , n33627 , n33628 );
and ( n33630 , n33599 , n33629 );
xor ( n33631 , n33297 , n33325 );
xor ( n33632 , n33631 , n33340 );
and ( n33633 , n33629 , n33632 );
and ( n33634 , n33599 , n33632 );
or ( n33635 , n33630 , n33633 , n33634 );
and ( n33636 , n24621 , n22048 );
and ( n33637 , n24527 , n22046 );
nor ( n33638 , n33636 , n33637 );
xnor ( n33639 , n33638 , n21853 );
and ( n33640 , n25284 , n21741 );
and ( n33641 , n24940 , n21739 );
nor ( n33642 , n33640 , n33641 );
xnor ( n33643 , n33642 , n21605 );
and ( n33644 , n33639 , n33643 );
and ( n33645 , n25765 , n21468 );
and ( n33646 , n25554 , n21466 );
nor ( n33647 , n33645 , n33646 );
xnor ( n33648 , n33647 , n21331 );
and ( n33649 , n33643 , n33648 );
and ( n33650 , n33639 , n33648 );
or ( n33651 , n33644 , n33649 , n33650 );
and ( n33652 , n23573 , n23230 );
and ( n33653 , n23381 , n23228 );
nor ( n33654 , n33652 , n33653 );
xnor ( n33655 , n33654 , n22842 );
and ( n33656 , n24131 , n22859 );
and ( n33657 , n23968 , n22857 );
nor ( n33658 , n33656 , n33657 );
xnor ( n33659 , n33658 , n22418 );
and ( n33660 , n33655 , n33659 );
and ( n33661 , n24527 , n22381 );
and ( n33662 , n24521 , n22379 );
nor ( n33663 , n33661 , n33662 );
xnor ( n33664 , n33663 , n22228 );
and ( n33665 , n33659 , n33664 );
and ( n33666 , n33655 , n33664 );
or ( n33667 , n33660 , n33665 , n33666 );
and ( n33668 , n23968 , n23230 );
and ( n33669 , n23573 , n23228 );
nor ( n33670 , n33668 , n33669 );
xnor ( n33671 , n33670 , n22842 );
and ( n33672 , n24521 , n22859 );
and ( n33673 , n24131 , n22857 );
nor ( n33674 , n33672 , n33673 );
xnor ( n33675 , n33674 , n22418 );
and ( n33676 , n33671 , n33675 );
and ( n33677 , n23271 , n23641 );
and ( n33678 , n23141 , n23639 );
nor ( n33679 , n33677 , n33678 );
xnor ( n33680 , n33679 , n23213 );
and ( n33681 , n33676 , n33680 );
and ( n33682 , n33680 , n33606 );
and ( n33683 , n33676 , n33606 );
or ( n33684 , n33681 , n33682 , n33683 );
and ( n33685 , n33667 , n33684 );
and ( n33686 , n29623 , n19894 );
and ( n33687 , n29318 , n19892 );
nor ( n33688 , n33686 , n33687 );
xnor ( n33689 , n33688 , n19858 );
and ( n33690 , n33684 , n33689 );
and ( n33691 , n33667 , n33689 );
or ( n33692 , n33685 , n33690 , n33691 );
and ( n33693 , n33651 , n33692 );
and ( n33694 , n19881 , n29977 );
and ( n33695 , n19825 , n29974 );
nor ( n33696 , n33694 , n33695 );
xnor ( n33697 , n33696 , n28674 );
and ( n33698 , n33692 , n33697 );
and ( n33699 , n33651 , n33697 );
or ( n33700 , n33693 , n33698 , n33699 );
xor ( n33701 , n33347 , n33351 );
xor ( n33702 , n33701 , n33356 );
xor ( n33703 , n33229 , n33233 );
xor ( n33704 , n33703 , n33238 );
and ( n33705 , n33702 , n33704 );
xor ( n33706 , n33301 , n33305 );
xor ( n33707 , n33706 , n33310 );
and ( n33708 , n33704 , n33707 );
and ( n33709 , n33702 , n33707 );
or ( n33710 , n33705 , n33708 , n33709 );
and ( n33711 , n33700 , n33710 );
xor ( n33712 , n33241 , n33257 );
xor ( n33713 , n33712 , n33262 );
and ( n33714 , n33710 , n33713 );
and ( n33715 , n33700 , n33713 );
or ( n33716 , n33711 , n33714 , n33715 );
and ( n33717 , n20452 , n28062 );
and ( n33718 , n20360 , n28060 );
nor ( n33719 , n33717 , n33718 );
xnor ( n33720 , n33719 , n27549 );
and ( n33721 , n21704 , n25383 );
and ( n33722 , n21612 , n25381 );
nor ( n33723 , n33721 , n33722 );
xnor ( n33724 , n33723 , n24885 );
and ( n33725 , n33720 , n33724 );
and ( n33726 , n21955 , n24902 );
and ( n33727 , n21876 , n24900 );
nor ( n33728 , n33726 , n33727 );
xnor ( n33729 , n33728 , n24397 );
and ( n33730 , n33724 , n33729 );
and ( n33731 , n33720 , n33729 );
or ( n33732 , n33725 , n33730 , n33731 );
xor ( n33733 , n33245 , n33249 );
xor ( n33734 , n33733 , n33254 );
and ( n33735 , n33732 , n33734 );
xor ( n33736 , n33611 , n33615 );
xor ( n33737 , n33736 , n33618 );
and ( n33738 , n33734 , n33737 );
and ( n33739 , n33732 , n33737 );
or ( n33740 , n33735 , n33738 , n33739 );
xor ( n33741 , n33455 , n33457 );
xor ( n33742 , n33741 , n33460 );
and ( n33743 , n33740 , n33742 );
xor ( n33744 , n33359 , n33361 );
xor ( n33745 , n33744 , n33364 );
and ( n33746 , n33742 , n33745 );
and ( n33747 , n33740 , n33745 );
or ( n33748 , n33743 , n33746 , n33747 );
and ( n33749 , n33716 , n33748 );
xor ( n33750 , n33265 , n33267 );
xor ( n33751 , n33750 , n33270 );
and ( n33752 , n33748 , n33751 );
and ( n33753 , n33716 , n33751 );
or ( n33754 , n33749 , n33752 , n33753 );
and ( n33755 , n33635 , n33754 );
xor ( n33756 , n33343 , n33375 );
xor ( n33757 , n33756 , n33378 );
and ( n33758 , n33754 , n33757 );
and ( n33759 , n33635 , n33757 );
or ( n33760 , n33755 , n33758 , n33759 );
xor ( n33761 , n33367 , n33369 );
xor ( n33762 , n33761 , n33372 );
xor ( n33763 , n33415 , n33417 );
xor ( n33764 , n33763 , n33420 );
and ( n33765 , n33762 , n33764 );
xor ( n33766 , n33463 , n33511 );
xor ( n33767 , n33766 , n33514 );
and ( n33768 , n33764 , n33767 );
and ( n33769 , n33762 , n33767 );
or ( n33770 , n33765 , n33768 , n33769 );
xor ( n33771 , n33423 , n33425 );
xor ( n33772 , n33771 , n33428 );
and ( n33773 , n33770 , n33772 );
xor ( n33774 , n33517 , n33519 );
xor ( n33775 , n33774 , n33522 );
and ( n33776 , n33772 , n33775 );
and ( n33777 , n33770 , n33775 );
or ( n33778 , n33773 , n33776 , n33777 );
and ( n33779 , n33760 , n33778 );
xor ( n33780 , n33431 , n33433 );
xor ( n33781 , n33780 , n33436 );
and ( n33782 , n33778 , n33781 );
and ( n33783 , n33760 , n33781 );
or ( n33784 , n33779 , n33782 , n33783 );
xor ( n33785 , n33387 , n33389 );
xor ( n33786 , n33785 , n33392 );
and ( n33787 , n33784 , n33786 );
xor ( n33788 , n33439 , n33533 );
xor ( n33789 , n33788 , n33536 );
and ( n33790 , n33786 , n33789 );
and ( n33791 , n33784 , n33789 );
or ( n33792 , n33787 , n33790 , n33791 );
and ( n33793 , n33551 , n33792 );
xor ( n33794 , n33551 , n33792 );
xor ( n33795 , n33784 , n33786 );
xor ( n33796 , n33795 , n33789 );
and ( n33797 , n20080 , n29276 );
and ( n33798 , n20004 , n29274 );
nor ( n33799 , n33797 , n33798 );
xnor ( n33800 , n33799 , n28677 );
and ( n33801 , n21451 , n26027 );
and ( n33802 , n21302 , n26025 );
nor ( n33803 , n33801 , n33802 );
xnor ( n33804 , n33803 , n25499 );
and ( n33805 , n33800 , n33804 );
xor ( n33806 , n33467 , n33471 );
xor ( n33807 , n33806 , n33476 );
and ( n33808 , n33804 , n33807 );
and ( n33809 , n33800 , n33807 );
or ( n33810 , n33805 , n33808 , n33809 );
and ( n33811 , n20666 , n27529 );
and ( n33812 , n20618 , n27527 );
nor ( n33813 , n33811 , n33812 );
xnor ( n33814 , n33813 , n27034 );
and ( n33815 , n20867 , n26992 );
and ( n33816 , n20803 , n26990 );
nor ( n33817 , n33815 , n33816 );
xnor ( n33818 , n33817 , n26369 );
and ( n33819 , n33814 , n33818 );
xor ( n33820 , n33600 , n33604 );
xor ( n33821 , n33820 , n33608 );
and ( n33822 , n33818 , n33821 );
and ( n33823 , n33814 , n33821 );
or ( n33824 , n33819 , n33822 , n33823 );
and ( n33825 , n33810 , n33824 );
xor ( n33826 , n33443 , n33447 );
xor ( n33827 , n33826 , n33452 );
and ( n33828 , n33824 , n33827 );
and ( n33829 , n33810 , n33827 );
or ( n33830 , n33825 , n33828 , n33829 );
and ( n33831 , n19946 , n29977 );
and ( n33832 , n19881 , n29974 );
nor ( n33833 , n33831 , n33832 );
xnor ( n33834 , n33833 , n28674 );
and ( n33835 , n20268 , n28628 );
and ( n33836 , n20182 , n28626 );
nor ( n33837 , n33835 , n33836 );
xnor ( n33838 , n33837 , n28096 );
and ( n33839 , n33834 , n33838 );
and ( n33840 , n21218 , n26349 );
and ( n33841 , n21072 , n26347 );
nor ( n33842 , n33840 , n33841 );
xnor ( n33843 , n33842 , n25893 );
and ( n33844 , n33838 , n33843 );
and ( n33845 , n33834 , n33843 );
or ( n33846 , n33839 , n33844 , n33845 );
and ( n33847 , n22425 , n24376 );
and ( n33848 , n22198 , n24374 );
nor ( n33849 , n33847 , n33848 );
xnor ( n33850 , n33849 , n23927 );
and ( n33851 , n22916 , n23944 );
and ( n33852 , n22756 , n23942 );
nor ( n33853 , n33851 , n33852 );
xnor ( n33854 , n33853 , n23550 );
and ( n33855 , n33850 , n33854 );
and ( n33856 , n24940 , n22048 );
and ( n33857 , n24621 , n22046 );
nor ( n33858 , n33856 , n33857 );
xnor ( n33859 , n33858 , n21853 );
and ( n33860 , n33854 , n33859 );
and ( n33861 , n33850 , n33859 );
or ( n33862 , n33855 , n33860 , n33861 );
and ( n33863 , n27135 , n20955 );
and ( n33864 , n26851 , n20953 );
nor ( n33865 , n33863 , n33864 );
xnor ( n33866 , n33865 , n20780 );
and ( n33867 , n27751 , n20674 );
and ( n33868 , n27352 , n20672 );
nor ( n33869 , n33867 , n33868 );
xnor ( n33870 , n33869 , n20542 );
and ( n33871 , n33866 , n33870 );
and ( n33872 , n28211 , n20460 );
and ( n33873 , n27757 , n20458 );
nor ( n33874 , n33872 , n33873 );
xnor ( n33875 , n33874 , n20337 );
and ( n33876 , n33870 , n33875 );
and ( n33877 , n33866 , n33875 );
or ( n33878 , n33871 , n33876 , n33877 );
and ( n33879 , n33862 , n33878 );
and ( n33880 , n28700 , n20276 );
and ( n33881 , n28810 , n20274 );
nor ( n33882 , n33880 , n33881 );
xnor ( n33883 , n33882 , n20175 );
and ( n33884 , n29318 , n20114 );
and ( n33885 , n29078 , n20112 );
nor ( n33886 , n33884 , n33885 );
xnor ( n33887 , n33886 , n19997 );
and ( n33888 , n33883 , n33887 );
xor ( n33889 , n33655 , n33659 );
xor ( n33890 , n33889 , n33664 );
and ( n33891 , n33887 , n33890 );
and ( n33892 , n33883 , n33890 );
or ( n33893 , n33888 , n33891 , n33892 );
and ( n33894 , n33878 , n33893 );
and ( n33895 , n33862 , n33893 );
or ( n33896 , n33879 , n33894 , n33895 );
and ( n33897 , n33846 , n33896 );
xor ( n33898 , n33479 , n33483 );
xor ( n33899 , n33898 , n33488 );
and ( n33900 , n33896 , n33899 );
and ( n33901 , n33846 , n33899 );
or ( n33902 , n33897 , n33900 , n33901 );
and ( n33903 , n33830 , n33902 );
xor ( n33904 , n33491 , n33505 );
xor ( n33905 , n33904 , n33508 );
and ( n33906 , n33902 , n33905 );
and ( n33907 , n33830 , n33905 );
or ( n33908 , n33903 , n33906 , n33907 );
xor ( n33909 , n33555 , n33559 );
xor ( n33910 , n33909 , n33564 );
xor ( n33911 , n33571 , n33575 );
xor ( n33912 , n33911 , n33580 );
and ( n33913 , n33910 , n33912 );
xor ( n33914 , n33639 , n33643 );
xor ( n33915 , n33914 , n33648 );
and ( n33916 , n33912 , n33915 );
and ( n33917 , n33910 , n33915 );
or ( n33918 , n33913 , n33916 , n33917 );
and ( n33919 , n25554 , n21741 );
and ( n33920 , n25284 , n21739 );
nor ( n33921 , n33919 , n33920 );
xnor ( n33922 , n33921 , n21605 );
and ( n33923 , n25974 , n21468 );
and ( n33924 , n25765 , n21466 );
nor ( n33925 , n33923 , n33924 );
xnor ( n33926 , n33925 , n21331 );
and ( n33927 , n33922 , n33926 );
and ( n33928 , n26422 , n21155 );
and ( n33929 , n26319 , n21153 );
nor ( n33930 , n33928 , n33929 );
xnor ( n33931 , n33930 , n20994 );
and ( n33932 , n33926 , n33931 );
and ( n33933 , n33922 , n33931 );
or ( n33934 , n33927 , n33932 , n33933 );
and ( n33935 , n22756 , n24376 );
and ( n33936 , n22425 , n24374 );
nor ( n33937 , n33935 , n33936 );
xnor ( n33938 , n33937 , n23927 );
and ( n33939 , n23141 , n23944 );
and ( n33940 , n22916 , n23942 );
nor ( n33941 , n33939 , n33940 );
xnor ( n33942 , n33941 , n23550 );
and ( n33943 , n33938 , n33942 );
and ( n33944 , n29623 , n20112 );
not ( n33945 , n33944 );
and ( n33946 , n33945 , n19997 );
and ( n33947 , n33942 , n33946 );
and ( n33948 , n33938 , n33946 );
or ( n33949 , n33943 , n33947 , n33948 );
xor ( n33950 , n33671 , n33675 );
and ( n33951 , n23381 , n23641 );
and ( n33952 , n23271 , n23639 );
nor ( n33953 , n33951 , n33952 );
xnor ( n33954 , n33953 , n23213 );
and ( n33955 , n33950 , n33954 );
and ( n33956 , n24621 , n22381 );
and ( n33957 , n24527 , n22379 );
nor ( n33958 , n33956 , n33957 );
xnor ( n33959 , n33958 , n22228 );
and ( n33960 , n33954 , n33959 );
and ( n33961 , n33950 , n33959 );
or ( n33962 , n33955 , n33960 , n33961 );
and ( n33963 , n33949 , n33962 );
and ( n33964 , n22235 , n24902 );
and ( n33965 , n21955 , n24900 );
nor ( n33966 , n33964 , n33965 );
xnor ( n33967 , n33966 , n24397 );
and ( n33968 , n33962 , n33967 );
and ( n33969 , n33949 , n33967 );
or ( n33970 , n33963 , n33968 , n33969 );
and ( n33971 , n33934 , n33970 );
xor ( n33972 , n33667 , n33684 );
xor ( n33973 , n33972 , n33689 );
and ( n33974 , n33970 , n33973 );
and ( n33975 , n33934 , n33973 );
or ( n33976 , n33971 , n33974 , n33975 );
and ( n33977 , n33918 , n33976 );
xor ( n33978 , n33495 , n33499 );
xor ( n33979 , n33978 , n33502 );
and ( n33980 , n33976 , n33979 );
and ( n33981 , n33918 , n33979 );
or ( n33982 , n33977 , n33980 , n33981 );
xor ( n33983 , n33591 , n33593 );
xor ( n33984 , n33983 , n33596 );
and ( n33985 , n33982 , n33984 );
xor ( n33986 , n33621 , n33623 );
xor ( n33987 , n33986 , n33626 );
and ( n33988 , n33984 , n33987 );
and ( n33989 , n33982 , n33987 );
or ( n33990 , n33985 , n33988 , n33989 );
and ( n33991 , n33908 , n33990 );
xor ( n33992 , n33599 , n33629 );
xor ( n33993 , n33992 , n33632 );
and ( n33994 , n33990 , n33993 );
and ( n33995 , n33908 , n33993 );
or ( n33996 , n33991 , n33994 , n33995 );
xor ( n33997 , n33567 , n33583 );
xor ( n33998 , n33997 , n33588 );
xor ( n33999 , n33651 , n33692 );
xor ( n34000 , n33999 , n33697 );
and ( n34001 , n33998 , n34000 );
xor ( n34002 , n33702 , n33704 );
xor ( n34003 , n34002 , n33707 );
and ( n34004 , n34000 , n34003 );
and ( n34005 , n33998 , n34003 );
or ( n34006 , n34001 , n34004 , n34005 );
xor ( n34007 , n33700 , n33710 );
xor ( n34008 , n34007 , n33713 );
and ( n34009 , n34006 , n34008 );
xor ( n34010 , n33740 , n33742 );
xor ( n34011 , n34010 , n33745 );
and ( n34012 , n34008 , n34011 );
and ( n34013 , n34006 , n34011 );
or ( n34014 , n34009 , n34012 , n34013 );
xor ( n34015 , n33716 , n33748 );
xor ( n34016 , n34015 , n33751 );
and ( n34017 , n34014 , n34016 );
xor ( n34018 , n33762 , n33764 );
xor ( n34019 , n34018 , n33767 );
and ( n34020 , n34016 , n34019 );
and ( n34021 , n34014 , n34019 );
or ( n34022 , n34017 , n34020 , n34021 );
and ( n34023 , n33996 , n34022 );
xor ( n34024 , n33635 , n33754 );
xor ( n34025 , n34024 , n33757 );
and ( n34026 , n34022 , n34025 );
and ( n34027 , n33996 , n34025 );
or ( n34028 , n34023 , n34026 , n34027 );
xor ( n34029 , n33525 , n33527 );
xor ( n34030 , n34029 , n33530 );
and ( n34031 , n34028 , n34030 );
xor ( n34032 , n33760 , n33778 );
xor ( n34033 , n34032 , n33781 );
and ( n34034 , n34030 , n34033 );
and ( n34035 , n34028 , n34033 );
or ( n34036 , n34031 , n34034 , n34035 );
and ( n34037 , n33796 , n34036 );
xor ( n34038 , n33796 , n34036 );
xor ( n34039 , n34028 , n34030 );
xor ( n34040 , n34039 , n34033 );
and ( n34041 , n20803 , n27529 );
and ( n34042 , n20666 , n27527 );
nor ( n34043 , n34041 , n34042 );
xnor ( n34044 , n34043 , n27034 );
and ( n34045 , n21612 , n26027 );
and ( n34046 , n21451 , n26025 );
nor ( n34047 , n34045 , n34046 );
xnor ( n34048 , n34047 , n25499 );
and ( n34049 , n34044 , n34048 );
and ( n34050 , n21876 , n25383 );
and ( n34051 , n21704 , n25381 );
nor ( n34052 , n34050 , n34051 );
xnor ( n34053 , n34052 , n24885 );
and ( n34054 , n34048 , n34053 );
and ( n34055 , n34044 , n34053 );
or ( n34056 , n34049 , n34054 , n34055 );
and ( n34057 , n20182 , n29276 );
and ( n34058 , n20080 , n29274 );
nor ( n34059 , n34057 , n34058 );
xnor ( n34060 , n34059 , n28677 );
and ( n34061 , n20618 , n28062 );
and ( n34062 , n20452 , n28060 );
nor ( n34063 , n34061 , n34062 );
xnor ( n34064 , n34063 , n27549 );
and ( n34065 , n34060 , n34064 );
and ( n34066 , n21072 , n26992 );
and ( n34067 , n20867 , n26990 );
nor ( n34068 , n34066 , n34067 );
xnor ( n34069 , n34068 , n26369 );
and ( n34070 , n34064 , n34069 );
and ( n34071 , n34060 , n34069 );
or ( n34072 , n34065 , n34070 , n34071 );
and ( n34073 , n34056 , n34072 );
and ( n34074 , n20360 , n28628 );
and ( n34075 , n20268 , n28626 );
nor ( n34076 , n34074 , n34075 );
xnor ( n34077 , n34076 , n28096 );
and ( n34078 , n21302 , n26349 );
and ( n34079 , n21218 , n26347 );
nor ( n34080 , n34078 , n34079 );
xnor ( n34081 , n34080 , n25893 );
and ( n34082 , n34077 , n34081 );
xor ( n34083 , n33676 , n33680 );
xor ( n34084 , n34083 , n33606 );
and ( n34085 , n34081 , n34084 );
and ( n34086 , n34077 , n34084 );
or ( n34087 , n34082 , n34085 , n34086 );
and ( n34088 , n34072 , n34087 );
and ( n34089 , n34056 , n34087 );
or ( n34090 , n34073 , n34088 , n34089 );
and ( n34091 , n27352 , n20955 );
and ( n34092 , n27135 , n20953 );
nor ( n34093 , n34091 , n34092 );
xnor ( n34094 , n34093 , n20780 );
and ( n34095 , n27757 , n20674 );
and ( n34096 , n27751 , n20672 );
nor ( n34097 , n34095 , n34096 );
xnor ( n34098 , n34097 , n20542 );
and ( n34099 , n34094 , n34098 );
and ( n34100 , n28810 , n20460 );
and ( n34101 , n28211 , n20458 );
nor ( n34102 , n34100 , n34101 );
xnor ( n34103 , n34102 , n20337 );
and ( n34104 , n34098 , n34103 );
and ( n34105 , n34094 , n34103 );
or ( n34106 , n34099 , n34104 , n34105 );
and ( n34107 , n20004 , n29977 );
and ( n34108 , n19946 , n29974 );
nor ( n34109 , n34107 , n34108 );
xnor ( n34110 , n34109 , n28674 );
and ( n34111 , n34106 , n34110 );
xor ( n34112 , n33850 , n33854 );
xor ( n34113 , n34112 , n33859 );
and ( n34114 , n34110 , n34113 );
and ( n34115 , n34106 , n34113 );
or ( n34116 , n34111 , n34114 , n34115 );
xor ( n34117 , n33834 , n33838 );
xor ( n34118 , n34117 , n33843 );
and ( n34119 , n34116 , n34118 );
xor ( n34120 , n33800 , n33804 );
xor ( n34121 , n34120 , n33807 );
and ( n34122 , n34118 , n34121 );
and ( n34123 , n34116 , n34121 );
or ( n34124 , n34119 , n34122 , n34123 );
and ( n34125 , n34090 , n34124 );
xor ( n34126 , n33810 , n33824 );
xor ( n34127 , n34126 , n33827 );
and ( n34128 , n34124 , n34127 );
and ( n34129 , n34090 , n34127 );
or ( n34130 , n34125 , n34128 , n34129 );
xor ( n34131 , n33720 , n33724 );
xor ( n34132 , n34131 , n33729 );
xor ( n34133 , n33862 , n33878 );
xor ( n34134 , n34133 , n33893 );
and ( n34135 , n34132 , n34134 );
xor ( n34136 , n33814 , n33818 );
xor ( n34137 , n34136 , n33821 );
and ( n34138 , n34134 , n34137 );
and ( n34139 , n34132 , n34137 );
or ( n34140 , n34135 , n34138 , n34139 );
xor ( n34141 , n33846 , n33896 );
xor ( n34142 , n34141 , n33899 );
and ( n34143 , n34140 , n34142 );
xor ( n34144 , n33732 , n33734 );
xor ( n34145 , n34144 , n33737 );
and ( n34146 , n34142 , n34145 );
and ( n34147 , n34140 , n34145 );
or ( n34148 , n34143 , n34146 , n34147 );
and ( n34149 , n34130 , n34148 );
xor ( n34150 , n33830 , n33902 );
xor ( n34151 , n34150 , n33905 );
and ( n34152 , n34148 , n34151 );
and ( n34153 , n34130 , n34151 );
or ( n34154 , n34149 , n34152 , n34153 );
and ( n34155 , n25765 , n21741 );
and ( n34156 , n25554 , n21739 );
nor ( n34157 , n34155 , n34156 );
xnor ( n34158 , n34157 , n21605 );
and ( n34159 , n26319 , n21468 );
and ( n34160 , n25974 , n21466 );
nor ( n34161 , n34159 , n34160 );
xnor ( n34162 , n34161 , n21331 );
and ( n34163 , n34158 , n34162 );
and ( n34164 , n26851 , n21155 );
and ( n34165 , n26422 , n21153 );
nor ( n34166 , n34164 , n34165 );
xnor ( n34167 , n34166 , n20994 );
and ( n34168 , n34162 , n34167 );
and ( n34169 , n34158 , n34167 );
or ( n34170 , n34163 , n34168 , n34169 );
and ( n34171 , n24131 , n23230 );
and ( n34172 , n23968 , n23228 );
nor ( n34173 , n34171 , n34172 );
xnor ( n34174 , n34173 , n22842 );
and ( n34175 , n24527 , n22859 );
and ( n34176 , n24521 , n22857 );
nor ( n34177 , n34175 , n34176 );
xnor ( n34178 , n34177 , n22418 );
and ( n34179 , n34174 , n34178 );
and ( n34180 , n24940 , n22381 );
and ( n34181 , n24621 , n22379 );
nor ( n34182 , n34180 , n34181 );
xnor ( n34183 , n34182 , n22228 );
and ( n34184 , n34178 , n34183 );
and ( n34185 , n34174 , n34183 );
or ( n34186 , n34179 , n34184 , n34185 );
and ( n34187 , n22198 , n24902 );
and ( n34188 , n22235 , n24900 );
nor ( n34189 , n34187 , n34188 );
xnor ( n34190 , n34189 , n24397 );
and ( n34191 , n34186 , n34190 );
and ( n34192 , n25284 , n22048 );
and ( n34193 , n24940 , n22046 );
nor ( n34194 , n34192 , n34193 );
xnor ( n34195 , n34194 , n21853 );
and ( n34196 , n34190 , n34195 );
and ( n34197 , n34186 , n34195 );
or ( n34198 , n34191 , n34196 , n34197 );
and ( n34199 , n34170 , n34198 );
and ( n34200 , n29078 , n20276 );
and ( n34201 , n28700 , n20274 );
nor ( n34202 , n34200 , n34201 );
xnor ( n34203 , n34202 , n20175 );
and ( n34204 , n29623 , n20114 );
and ( n34205 , n29318 , n20112 );
nor ( n34206 , n34204 , n34205 );
xnor ( n34207 , n34206 , n19997 );
and ( n34208 , n34203 , n34207 );
xor ( n34209 , n33950 , n33954 );
xor ( n34210 , n34209 , n33959 );
and ( n34211 , n34207 , n34210 );
and ( n34212 , n34203 , n34210 );
or ( n34213 , n34208 , n34211 , n34212 );
and ( n34214 , n34198 , n34213 );
and ( n34215 , n34170 , n34213 );
or ( n34216 , n34199 , n34214 , n34215 );
xor ( n34217 , n33922 , n33926 );
xor ( n34218 , n34217 , n33931 );
xor ( n34219 , n33866 , n33870 );
xor ( n34220 , n34219 , n33875 );
and ( n34221 , n34218 , n34220 );
xor ( n34222 , n33883 , n33887 );
xor ( n34223 , n34222 , n33890 );
and ( n34224 , n34220 , n34223 );
and ( n34225 , n34218 , n34223 );
or ( n34226 , n34221 , n34224 , n34225 );
and ( n34227 , n34216 , n34226 );
xor ( n34228 , n33910 , n33912 );
xor ( n34229 , n34228 , n33915 );
and ( n34230 , n34226 , n34229 );
and ( n34231 , n34216 , n34229 );
or ( n34232 , n34227 , n34230 , n34231 );
xor ( n34233 , n33918 , n33976 );
xor ( n34234 , n34233 , n33979 );
and ( n34235 , n34232 , n34234 );
xor ( n34236 , n33998 , n34000 );
xor ( n34237 , n34236 , n34003 );
and ( n34238 , n34234 , n34237 );
and ( n34239 , n34232 , n34237 );
or ( n34240 , n34235 , n34238 , n34239 );
xor ( n34241 , n33982 , n33984 );
xor ( n34242 , n34241 , n33987 );
and ( n34243 , n34240 , n34242 );
xor ( n34244 , n34006 , n34008 );
xor ( n34245 , n34244 , n34011 );
and ( n34246 , n34242 , n34245 );
and ( n34247 , n34240 , n34245 );
or ( n34248 , n34243 , n34246 , n34247 );
and ( n34249 , n34154 , n34248 );
xor ( n34250 , n33908 , n33990 );
xor ( n34251 , n34250 , n33993 );
and ( n34252 , n34248 , n34251 );
and ( n34253 , n34154 , n34251 );
or ( n34254 , n34249 , n34252 , n34253 );
xor ( n34255 , n33770 , n33772 );
xor ( n34256 , n34255 , n33775 );
and ( n34257 , n34254 , n34256 );
xor ( n34258 , n33996 , n34022 );
xor ( n34259 , n34258 , n34025 );
and ( n34260 , n34256 , n34259 );
and ( n34261 , n34254 , n34259 );
or ( n34262 , n34257 , n34260 , n34261 );
and ( n34263 , n34040 , n34262 );
xor ( n34264 , n34040 , n34262 );
xor ( n34265 , n34254 , n34256 );
xor ( n34266 , n34265 , n34259 );
and ( n34267 , n20666 , n28062 );
and ( n34268 , n20618 , n28060 );
nor ( n34269 , n34267 , n34268 );
xnor ( n34270 , n34269 , n27549 );
and ( n34271 , n20867 , n27529 );
and ( n34272 , n20803 , n27527 );
nor ( n34273 , n34271 , n34272 );
xnor ( n34274 , n34273 , n27034 );
and ( n34275 , n34270 , n34274 );
and ( n34276 , n21955 , n25383 );
and ( n34277 , n21876 , n25381 );
nor ( n34278 , n34276 , n34277 );
xnor ( n34279 , n34278 , n24885 );
and ( n34280 , n34274 , n34279 );
and ( n34281 , n34270 , n34279 );
or ( n34282 , n34275 , n34280 , n34281 );
xor ( n34283 , n34044 , n34048 );
xor ( n34284 , n34283 , n34053 );
and ( n34285 , n34282 , n34284 );
xor ( n34286 , n33949 , n33962 );
xor ( n34287 , n34286 , n33967 );
and ( n34288 , n34284 , n34287 );
and ( n34289 , n34282 , n34287 );
or ( n34290 , n34285 , n34288 , n34289 );
and ( n34291 , n25554 , n22048 );
and ( n34292 , n25284 , n22046 );
nor ( n34293 , n34291 , n34292 );
xnor ( n34294 , n34293 , n21853 );
and ( n34295 , n25974 , n21741 );
and ( n34296 , n25765 , n21739 );
nor ( n34297 , n34295 , n34296 );
xnor ( n34298 , n34297 , n21605 );
and ( n34299 , n34294 , n34298 );
xor ( n34300 , n34174 , n34178 );
xor ( n34301 , n34300 , n34183 );
and ( n34302 , n34298 , n34301 );
and ( n34303 , n34294 , n34301 );
or ( n34304 , n34299 , n34302 , n34303 );
and ( n34305 , n23968 , n23641 );
and ( n34306 , n23573 , n23639 );
nor ( n34307 , n34305 , n34306 );
xnor ( n34308 , n34307 , n23213 );
and ( n34309 , n24521 , n23230 );
and ( n34310 , n24131 , n23228 );
nor ( n34311 , n34309 , n34310 );
xnor ( n34312 , n34311 , n22842 );
xor ( n34313 , n34308 , n34312 );
and ( n34314 , n24621 , n22859 );
and ( n34315 , n24527 , n22857 );
nor ( n34316 , n34314 , n34315 );
xnor ( n34317 , n34316 , n22418 );
and ( n34318 , n34313 , n34317 );
and ( n34319 , n25284 , n22381 );
and ( n34320 , n24940 , n22379 );
nor ( n34321 , n34319 , n34320 );
xnor ( n34322 , n34321 , n22228 );
and ( n34323 , n34317 , n34322 );
and ( n34324 , n34313 , n34322 );
or ( n34325 , n34318 , n34323 , n34324 );
and ( n34326 , n22235 , n25383 );
and ( n34327 , n21955 , n25381 );
nor ( n34328 , n34326 , n34327 );
xnor ( n34329 , n34328 , n24885 );
and ( n34330 , n34325 , n34329 );
and ( n34331 , n34308 , n34312 );
and ( n34332 , n22916 , n24376 );
and ( n34333 , n22756 , n24374 );
nor ( n34334 , n34332 , n34333 );
xnor ( n34335 , n34334 , n23927 );
xor ( n34336 , n34331 , n34335 );
and ( n34337 , n23573 , n23641 );
and ( n34338 , n23381 , n23639 );
nor ( n34339 , n34337 , n34338 );
xnor ( n34340 , n34339 , n23213 );
xor ( n34341 , n34336 , n34340 );
and ( n34342 , n34329 , n34341 );
and ( n34343 , n34325 , n34341 );
or ( n34344 , n34330 , n34342 , n34343 );
and ( n34345 , n34304 , n34344 );
xor ( n34346 , n34203 , n34207 );
xor ( n34347 , n34346 , n34210 );
and ( n34348 , n34344 , n34347 );
and ( n34349 , n34304 , n34347 );
or ( n34350 , n34345 , n34348 , n34349 );
xor ( n34351 , n34170 , n34198 );
xor ( n34352 , n34351 , n34213 );
and ( n34353 , n34350 , n34352 );
xor ( n34354 , n34106 , n34110 );
xor ( n34355 , n34354 , n34113 );
and ( n34356 , n34352 , n34355 );
and ( n34357 , n34350 , n34355 );
or ( n34358 , n34353 , n34356 , n34357 );
and ( n34359 , n34290 , n34358 );
xor ( n34360 , n34056 , n34072 );
xor ( n34361 , n34360 , n34087 );
and ( n34362 , n34358 , n34361 );
and ( n34363 , n34290 , n34361 );
or ( n34364 , n34359 , n34362 , n34363 );
and ( n34365 , n20452 , n28628 );
and ( n34366 , n20360 , n28626 );
nor ( n34367 , n34365 , n34366 );
xnor ( n34368 , n34367 , n28096 );
and ( n34369 , n21218 , n26992 );
and ( n34370 , n21072 , n26990 );
nor ( n34371 , n34369 , n34370 );
xnor ( n34372 , n34371 , n26369 );
and ( n34373 , n34368 , n34372 );
and ( n34374 , n21451 , n26349 );
and ( n34375 , n21302 , n26347 );
nor ( n34376 , n34374 , n34375 );
xnor ( n34377 , n34376 , n25893 );
and ( n34378 , n34372 , n34377 );
and ( n34379 , n34368 , n34377 );
or ( n34380 , n34373 , n34378 , n34379 );
and ( n34381 , n22425 , n24902 );
and ( n34382 , n22198 , n24900 );
nor ( n34383 , n34381 , n34382 );
xnor ( n34384 , n34383 , n24397 );
and ( n34385 , n23271 , n23944 );
and ( n34386 , n23141 , n23942 );
nor ( n34387 , n34385 , n34386 );
xnor ( n34388 , n34387 , n23550 );
and ( n34389 , n34384 , n34388 );
and ( n34390 , n34388 , n33944 );
and ( n34391 , n34384 , n33944 );
or ( n34392 , n34389 , n34390 , n34391 );
and ( n34393 , n34331 , n34335 );
and ( n34394 , n34335 , n34340 );
and ( n34395 , n34331 , n34340 );
or ( n34396 , n34393 , n34394 , n34395 );
and ( n34397 , n34392 , n34396 );
and ( n34398 , n21704 , n26027 );
and ( n34399 , n21612 , n26025 );
nor ( n34400 , n34398 , n34399 );
xnor ( n34401 , n34400 , n25499 );
and ( n34402 , n34396 , n34401 );
and ( n34403 , n34392 , n34401 );
or ( n34404 , n34397 , n34402 , n34403 );
and ( n34405 , n34380 , n34404 );
and ( n34406 , n20080 , n29977 );
and ( n34407 , n20004 , n29974 );
nor ( n34408 , n34406 , n34407 );
xnor ( n34409 , n34408 , n28674 );
and ( n34410 , n20268 , n29276 );
and ( n34411 , n20182 , n29274 );
nor ( n34412 , n34410 , n34411 );
xnor ( n34413 , n34412 , n28677 );
and ( n34414 , n34409 , n34413 );
xor ( n34415 , n33938 , n33942 );
xor ( n34416 , n34415 , n33946 );
and ( n34417 , n34413 , n34416 );
and ( n34418 , n34409 , n34416 );
or ( n34419 , n34414 , n34417 , n34418 );
and ( n34420 , n34404 , n34419 );
and ( n34421 , n34380 , n34419 );
or ( n34422 , n34405 , n34420 , n34421 );
and ( n34423 , n28211 , n20674 );
and ( n34424 , n27757 , n20672 );
nor ( n34425 , n34423 , n34424 );
xnor ( n34426 , n34425 , n20542 );
and ( n34427 , n28700 , n20460 );
and ( n34428 , n28810 , n20458 );
nor ( n34429 , n34427 , n34428 );
xnor ( n34430 , n34429 , n20337 );
and ( n34431 , n34426 , n34430 );
and ( n34432 , n29318 , n20276 );
and ( n34433 , n29078 , n20274 );
nor ( n34434 , n34432 , n34433 );
xnor ( n34435 , n34434 , n20175 );
and ( n34436 , n34430 , n34435 );
and ( n34437 , n34426 , n34435 );
or ( n34438 , n34431 , n34436 , n34437 );
and ( n34439 , n26422 , n21468 );
and ( n34440 , n26319 , n21466 );
nor ( n34441 , n34439 , n34440 );
xnor ( n34442 , n34441 , n21331 );
and ( n34443 , n27135 , n21155 );
and ( n34444 , n26851 , n21153 );
nor ( n34445 , n34443 , n34444 );
xnor ( n34446 , n34445 , n20994 );
and ( n34447 , n34442 , n34446 );
and ( n34448 , n27751 , n20955 );
and ( n34449 , n27352 , n20953 );
nor ( n34450 , n34448 , n34449 );
xnor ( n34451 , n34450 , n20780 );
and ( n34452 , n34446 , n34451 );
and ( n34453 , n34442 , n34451 );
or ( n34454 , n34447 , n34452 , n34453 );
and ( n34455 , n34438 , n34454 );
xor ( n34456 , n34186 , n34190 );
xor ( n34457 , n34456 , n34195 );
and ( n34458 , n34454 , n34457 );
and ( n34459 , n34438 , n34457 );
or ( n34460 , n34455 , n34458 , n34459 );
xor ( n34461 , n34060 , n34064 );
xor ( n34462 , n34461 , n34069 );
and ( n34463 , n34460 , n34462 );
xor ( n34464 , n34077 , n34081 );
xor ( n34465 , n34464 , n34084 );
and ( n34466 , n34462 , n34465 );
and ( n34467 , n34460 , n34465 );
or ( n34468 , n34463 , n34466 , n34467 );
and ( n34469 , n34422 , n34468 );
xor ( n34470 , n33934 , n33970 );
xor ( n34471 , n34470 , n33973 );
and ( n34472 , n34468 , n34471 );
and ( n34473 , n34422 , n34471 );
or ( n34474 , n34469 , n34472 , n34473 );
and ( n34475 , n34364 , n34474 );
xor ( n34476 , n34090 , n34124 );
xor ( n34477 , n34476 , n34127 );
and ( n34478 , n34474 , n34477 );
and ( n34479 , n34364 , n34477 );
or ( n34480 , n34475 , n34478 , n34479 );
xor ( n34481 , n34116 , n34118 );
xor ( n34482 , n34481 , n34121 );
xor ( n34483 , n34132 , n34134 );
xor ( n34484 , n34483 , n34137 );
and ( n34485 , n34482 , n34484 );
xor ( n34486 , n34216 , n34226 );
xor ( n34487 , n34486 , n34229 );
and ( n34488 , n34484 , n34487 );
and ( n34489 , n34482 , n34487 );
or ( n34490 , n34485 , n34488 , n34489 );
and ( n34491 , n27352 , n21155 );
and ( n34492 , n27135 , n21153 );
nor ( n34493 , n34491 , n34492 );
xnor ( n34494 , n34493 , n20994 );
and ( n34495 , n27757 , n20955 );
and ( n34496 , n27751 , n20953 );
nor ( n34497 , n34495 , n34496 );
xnor ( n34498 , n34497 , n20780 );
and ( n34499 , n34494 , n34498 );
and ( n34500 , n29078 , n20460 );
and ( n34501 , n28700 , n20458 );
nor ( n34502 , n34500 , n34501 );
xnor ( n34503 , n34502 , n20337 );
and ( n34504 , n34498 , n34503 );
and ( n34505 , n34494 , n34503 );
or ( n34506 , n34499 , n34504 , n34505 );
and ( n34507 , n24131 , n23641 );
and ( n34508 , n23968 , n23639 );
nor ( n34509 , n34507 , n34508 );
xnor ( n34510 , n34509 , n23213 );
and ( n34511 , n24527 , n23230 );
and ( n34512 , n24521 , n23228 );
nor ( n34513 , n34511 , n34512 );
xnor ( n34514 , n34513 , n22842 );
and ( n34515 , n34510 , n34514 );
and ( n34516 , n24940 , n22859 );
and ( n34517 , n24621 , n22857 );
nor ( n34518 , n34516 , n34517 );
xnor ( n34519 , n34518 , n22418 );
and ( n34520 , n34514 , n34519 );
and ( n34521 , n34510 , n34519 );
or ( n34522 , n34515 , n34520 , n34521 );
and ( n34523 , n22198 , n25383 );
and ( n34524 , n22235 , n25381 );
nor ( n34525 , n34523 , n34524 );
xnor ( n34526 , n34525 , n24885 );
and ( n34527 , n34522 , n34526 );
and ( n34528 , n22756 , n24902 );
and ( n34529 , n22425 , n24900 );
nor ( n34530 , n34528 , n34529 );
xnor ( n34531 , n34530 , n24397 );
and ( n34532 , n34526 , n34531 );
and ( n34533 , n34522 , n34531 );
or ( n34534 , n34527 , n34532 , n34533 );
and ( n34535 , n34506 , n34534 );
and ( n34536 , n21612 , n26349 );
and ( n34537 , n21451 , n26347 );
nor ( n34538 , n34536 , n34537 );
xnor ( n34539 , n34538 , n25893 );
and ( n34540 , n34534 , n34539 );
and ( n34541 , n34506 , n34539 );
or ( n34542 , n34535 , n34540 , n34541 );
xor ( n34543 , n34270 , n34274 );
xor ( n34544 , n34543 , n34279 );
and ( n34545 , n34542 , n34544 );
xor ( n34546 , n34368 , n34372 );
xor ( n34547 , n34546 , n34377 );
and ( n34548 , n34544 , n34547 );
and ( n34549 , n34542 , n34547 );
or ( n34550 , n34545 , n34548 , n34549 );
xor ( n34551 , n34380 , n34404 );
xor ( n34552 , n34551 , n34419 );
and ( n34553 , n34550 , n34552 );
xor ( n34554 , n34282 , n34284 );
xor ( n34555 , n34554 , n34287 );
and ( n34556 , n34552 , n34555 );
and ( n34557 , n34550 , n34555 );
or ( n34558 , n34553 , n34556 , n34557 );
and ( n34559 , n23141 , n24376 );
and ( n34560 , n22916 , n24374 );
nor ( n34561 , n34559 , n34560 );
xnor ( n34562 , n34561 , n23927 );
and ( n34563 , n23381 , n23944 );
and ( n34564 , n23271 , n23942 );
nor ( n34565 , n34563 , n34564 );
xnor ( n34566 , n34565 , n23550 );
and ( n34567 , n34562 , n34566 );
and ( n34568 , n29623 , n20274 );
not ( n34569 , n34568 );
and ( n34570 , n34569 , n20175 );
and ( n34571 , n34566 , n34570 );
and ( n34572 , n34562 , n34570 );
or ( n34573 , n34567 , n34571 , n34572 );
and ( n34574 , n20360 , n29276 );
and ( n34575 , n20268 , n29274 );
nor ( n34576 , n34574 , n34575 );
xnor ( n34577 , n34576 , n28677 );
and ( n34578 , n34573 , n34577 );
and ( n34579 , n21876 , n26027 );
and ( n34580 , n21704 , n26025 );
nor ( n34581 , n34579 , n34580 );
xnor ( n34582 , n34581 , n25499 );
and ( n34583 , n34577 , n34582 );
and ( n34584 , n34573 , n34582 );
or ( n34585 , n34578 , n34583 , n34584 );
xor ( n34586 , n34094 , n34098 );
xor ( n34587 , n34586 , n34103 );
and ( n34588 , n34585 , n34587 );
xor ( n34589 , n34158 , n34162 );
xor ( n34590 , n34589 , n34167 );
and ( n34591 , n34587 , n34590 );
and ( n34592 , n34585 , n34590 );
or ( n34593 , n34588 , n34591 , n34592 );
and ( n34594 , n20182 , n29977 );
and ( n34595 , n20080 , n29974 );
nor ( n34596 , n34594 , n34595 );
xnor ( n34597 , n34596 , n28674 );
and ( n34598 , n20618 , n28628 );
and ( n34599 , n20452 , n28626 );
nor ( n34600 , n34598 , n34599 );
xnor ( n34601 , n34600 , n28096 );
and ( n34602 , n34597 , n34601 );
and ( n34603 , n21302 , n26992 );
and ( n34604 , n21218 , n26990 );
nor ( n34605 , n34603 , n34604 );
xnor ( n34606 , n34605 , n26369 );
and ( n34607 , n34601 , n34606 );
and ( n34608 , n34597 , n34606 );
or ( n34609 , n34602 , n34607 , n34608 );
and ( n34610 , n20803 , n28062 );
and ( n34611 , n20666 , n28060 );
nor ( n34612 , n34610 , n34611 );
xnor ( n34613 , n34612 , n27549 );
and ( n34614 , n21072 , n27529 );
and ( n34615 , n20867 , n27527 );
nor ( n34616 , n34614 , n34615 );
xnor ( n34617 , n34616 , n27034 );
and ( n34618 , n34613 , n34617 );
xor ( n34619 , n34384 , n34388 );
xor ( n34620 , n34619 , n33944 );
and ( n34621 , n34617 , n34620 );
and ( n34622 , n34613 , n34620 );
or ( n34623 , n34618 , n34621 , n34622 );
and ( n34624 , n34609 , n34623 );
xor ( n34625 , n34392 , n34396 );
xor ( n34626 , n34625 , n34401 );
and ( n34627 , n34623 , n34626 );
and ( n34628 , n34609 , n34626 );
or ( n34629 , n34624 , n34627 , n34628 );
and ( n34630 , n34593 , n34629 );
xor ( n34631 , n34218 , n34220 );
xor ( n34632 , n34631 , n34223 );
and ( n34633 , n34629 , n34632 );
and ( n34634 , n34593 , n34632 );
or ( n34635 , n34630 , n34633 , n34634 );
and ( n34636 , n34558 , n34635 );
xor ( n34637 , n34422 , n34468 );
xor ( n34638 , n34637 , n34471 );
and ( n34639 , n34635 , n34638 );
and ( n34640 , n34558 , n34638 );
or ( n34641 , n34636 , n34639 , n34640 );
and ( n34642 , n34490 , n34641 );
xor ( n34643 , n34140 , n34142 );
xor ( n34644 , n34643 , n34145 );
and ( n34645 , n34641 , n34644 );
and ( n34646 , n34490 , n34644 );
or ( n34647 , n34642 , n34645 , n34646 );
and ( n34648 , n34480 , n34647 );
xor ( n34649 , n34130 , n34148 );
xor ( n34650 , n34649 , n34151 );
and ( n34651 , n34647 , n34650 );
and ( n34652 , n34480 , n34650 );
or ( n34653 , n34648 , n34651 , n34652 );
xor ( n34654 , n34154 , n34248 );
xor ( n34655 , n34654 , n34251 );
and ( n34656 , n34653 , n34655 );
xor ( n34657 , n34014 , n34016 );
xor ( n34658 , n34657 , n34019 );
and ( n34659 , n34655 , n34658 );
and ( n34660 , n34653 , n34658 );
or ( n34661 , n34656 , n34659 , n34660 );
and ( n34662 , n34266 , n34661 );
xor ( n34663 , n34266 , n34661 );
xor ( n34664 , n34653 , n34655 );
xor ( n34665 , n34664 , n34658 );
and ( n34666 , n25765 , n22048 );
and ( n34667 , n25554 , n22046 );
nor ( n34668 , n34666 , n34667 );
xnor ( n34669 , n34668 , n21853 );
and ( n34670 , n26319 , n21741 );
and ( n34671 , n25974 , n21739 );
nor ( n34672 , n34670 , n34671 );
xnor ( n34673 , n34672 , n21605 );
and ( n34674 , n34669 , n34673 );
and ( n34675 , n26851 , n21468 );
and ( n34676 , n26422 , n21466 );
nor ( n34677 , n34675 , n34676 );
xnor ( n34678 , n34677 , n21331 );
and ( n34679 , n34673 , n34678 );
and ( n34680 , n34669 , n34678 );
or ( n34681 , n34674 , n34679 , n34680 );
and ( n34682 , n28810 , n20674 );
and ( n34683 , n28211 , n20672 );
nor ( n34684 , n34682 , n34683 );
xnor ( n34685 , n34684 , n20542 );
and ( n34686 , n29623 , n20276 );
and ( n34687 , n29318 , n20274 );
nor ( n34688 , n34686 , n34687 );
xnor ( n34689 , n34688 , n20175 );
and ( n34690 , n34685 , n34689 );
xor ( n34691 , n34313 , n34317 );
xor ( n34692 , n34691 , n34322 );
and ( n34693 , n34689 , n34692 );
and ( n34694 , n34685 , n34692 );
or ( n34695 , n34690 , n34693 , n34694 );
and ( n34696 , n34681 , n34695 );
xor ( n34697 , n34426 , n34430 );
xor ( n34698 , n34697 , n34435 );
and ( n34699 , n34695 , n34698 );
and ( n34700 , n34681 , n34698 );
or ( n34701 , n34696 , n34699 , n34700 );
xor ( n34702 , n34409 , n34413 );
xor ( n34703 , n34702 , n34416 );
and ( n34704 , n34701 , n34703 );
xor ( n34705 , n34438 , n34454 );
xor ( n34706 , n34705 , n34457 );
and ( n34707 , n34703 , n34706 );
and ( n34708 , n34701 , n34706 );
or ( n34709 , n34704 , n34707 , n34708 );
xor ( n34710 , n34460 , n34462 );
xor ( n34711 , n34710 , n34465 );
and ( n34712 , n34709 , n34711 );
xor ( n34713 , n34350 , n34352 );
xor ( n34714 , n34713 , n34355 );
and ( n34715 , n34711 , n34714 );
and ( n34716 , n34709 , n34714 );
or ( n34717 , n34712 , n34715 , n34716 );
xor ( n34718 , n34290 , n34358 );
xor ( n34719 , n34718 , n34361 );
and ( n34720 , n34717 , n34719 );
xor ( n34721 , n34482 , n34484 );
xor ( n34722 , n34721 , n34487 );
and ( n34723 , n34719 , n34722 );
and ( n34724 , n34717 , n34722 );
or ( n34725 , n34720 , n34723 , n34724 );
xor ( n34726 , n34232 , n34234 );
xor ( n34727 , n34726 , n34237 );
and ( n34728 , n34725 , n34727 );
xor ( n34729 , n34364 , n34474 );
xor ( n34730 , n34729 , n34477 );
and ( n34731 , n34727 , n34730 );
and ( n34732 , n34725 , n34730 );
or ( n34733 , n34728 , n34731 , n34732 );
xor ( n34734 , n34240 , n34242 );
xor ( n34735 , n34734 , n34245 );
and ( n34736 , n34733 , n34735 );
xor ( n34737 , n34480 , n34647 );
xor ( n34738 , n34737 , n34650 );
and ( n34739 , n34735 , n34738 );
and ( n34740 , n34733 , n34738 );
or ( n34741 , n34736 , n34739 , n34740 );
and ( n34742 , n34665 , n34741 );
xor ( n34743 , n34665 , n34741 );
xor ( n34744 , n34733 , n34735 );
xor ( n34745 , n34744 , n34738 );
and ( n34746 , n22425 , n25383 );
and ( n34747 , n22198 , n25381 );
nor ( n34748 , n34746 , n34747 );
xnor ( n34749 , n34748 , n24885 );
and ( n34750 , n22916 , n24902 );
and ( n34751 , n22756 , n24900 );
nor ( n34752 , n34750 , n34751 );
xnor ( n34753 , n34752 , n24397 );
and ( n34754 , n34749 , n34753 );
and ( n34755 , n23271 , n24376 );
and ( n34756 , n23141 , n24374 );
nor ( n34757 , n34755 , n34756 );
xnor ( n34758 , n34757 , n23927 );
and ( n34759 , n34753 , n34758 );
and ( n34760 , n34749 , n34758 );
or ( n34761 , n34754 , n34759 , n34760 );
and ( n34762 , n23968 , n23944 );
and ( n34763 , n23573 , n23942 );
nor ( n34764 , n34762 , n34763 );
xnor ( n34765 , n34764 , n23550 );
and ( n34766 , n24521 , n23641 );
and ( n34767 , n24131 , n23639 );
nor ( n34768 , n34766 , n34767 );
xnor ( n34769 , n34768 , n23213 );
and ( n34770 , n34765 , n34769 );
and ( n34771 , n23573 , n23944 );
and ( n34772 , n23381 , n23942 );
nor ( n34773 , n34771 , n34772 );
xnor ( n34774 , n34773 , n23550 );
and ( n34775 , n34770 , n34774 );
and ( n34776 , n25554 , n22381 );
and ( n34777 , n25284 , n22379 );
nor ( n34778 , n34776 , n34777 );
xnor ( n34779 , n34778 , n22228 );
and ( n34780 , n34774 , n34779 );
and ( n34781 , n34770 , n34779 );
or ( n34782 , n34775 , n34780 , n34781 );
and ( n34783 , n34761 , n34782 );
xor ( n34784 , n34522 , n34526 );
xor ( n34785 , n34784 , n34531 );
and ( n34786 , n34782 , n34785 );
and ( n34787 , n34761 , n34785 );
or ( n34788 , n34783 , n34786 , n34787 );
xor ( n34789 , n34442 , n34446 );
xor ( n34790 , n34789 , n34451 );
and ( n34791 , n34788 , n34790 );
xor ( n34792 , n34294 , n34298 );
xor ( n34793 , n34792 , n34301 );
and ( n34794 , n34790 , n34793 );
and ( n34795 , n34788 , n34793 );
or ( n34796 , n34791 , n34794 , n34795 );
and ( n34797 , n20452 , n29276 );
and ( n34798 , n20360 , n29274 );
nor ( n34799 , n34797 , n34798 );
xnor ( n34800 , n34799 , n28677 );
and ( n34801 , n20867 , n28062 );
and ( n34802 , n20803 , n28060 );
nor ( n34803 , n34801 , n34802 );
xnor ( n34804 , n34803 , n27549 );
and ( n34805 , n34800 , n34804 );
and ( n34806 , n21955 , n26027 );
and ( n34807 , n21876 , n26025 );
nor ( n34808 , n34806 , n34807 );
xnor ( n34809 , n34808 , n25499 );
and ( n34810 , n34804 , n34809 );
and ( n34811 , n34800 , n34809 );
or ( n34812 , n34805 , n34810 , n34811 );
and ( n34813 , n21218 , n27529 );
and ( n34814 , n21072 , n27527 );
nor ( n34815 , n34813 , n34814 );
xnor ( n34816 , n34815 , n27034 );
and ( n34817 , n21451 , n26992 );
and ( n34818 , n21302 , n26990 );
nor ( n34819 , n34817 , n34818 );
xnor ( n34820 , n34819 , n26369 );
and ( n34821 , n34816 , n34820 );
xor ( n34822 , n34562 , n34566 );
xor ( n34823 , n34822 , n34570 );
and ( n34824 , n34820 , n34823 );
and ( n34825 , n34816 , n34823 );
or ( n34826 , n34821 , n34824 , n34825 );
and ( n34827 , n34812 , n34826 );
xor ( n34828 , n34325 , n34329 );
xor ( n34829 , n34828 , n34341 );
and ( n34830 , n34826 , n34829 );
and ( n34831 , n34812 , n34829 );
or ( n34832 , n34827 , n34830 , n34831 );
and ( n34833 , n34796 , n34832 );
xor ( n34834 , n34585 , n34587 );
xor ( n34835 , n34834 , n34590 );
and ( n34836 , n34832 , n34835 );
and ( n34837 , n34796 , n34835 );
or ( n34838 , n34833 , n34836 , n34837 );
and ( n34839 , n20268 , n29977 );
and ( n34840 , n20182 , n29974 );
nor ( n34841 , n34839 , n34840 );
xnor ( n34842 , n34841 , n28674 );
and ( n34843 , n20666 , n28628 );
and ( n34844 , n20618 , n28626 );
nor ( n34845 , n34843 , n34844 );
xnor ( n34846 , n34845 , n28096 );
and ( n34847 , n34842 , n34846 );
and ( n34848 , n21704 , n26349 );
and ( n34849 , n21612 , n26347 );
nor ( n34850 , n34848 , n34849 );
xnor ( n34851 , n34850 , n25893 );
and ( n34852 , n34846 , n34851 );
and ( n34853 , n34842 , n34851 );
or ( n34854 , n34847 , n34852 , n34853 );
and ( n34855 , n27751 , n21155 );
and ( n34856 , n27352 , n21153 );
nor ( n34857 , n34855 , n34856 );
xnor ( n34858 , n34857 , n20994 );
and ( n34859 , n28211 , n20955 );
and ( n34860 , n27757 , n20953 );
nor ( n34861 , n34859 , n34860 );
xnor ( n34862 , n34861 , n20780 );
and ( n34863 , n34858 , n34862 );
and ( n34864 , n28700 , n20674 );
and ( n34865 , n28810 , n20672 );
nor ( n34866 , n34864 , n34865 );
xnor ( n34867 , n34866 , n20542 );
and ( n34868 , n34862 , n34867 );
and ( n34869 , n34858 , n34867 );
or ( n34870 , n34863 , n34868 , n34869 );
and ( n34871 , n25974 , n22048 );
and ( n34872 , n25765 , n22046 );
nor ( n34873 , n34871 , n34872 );
xnor ( n34874 , n34873 , n21853 );
and ( n34875 , n26422 , n21741 );
and ( n34876 , n26319 , n21739 );
nor ( n34877 , n34875 , n34876 );
xnor ( n34878 , n34877 , n21605 );
and ( n34879 , n34874 , n34878 );
and ( n34880 , n27135 , n21468 );
and ( n34881 , n26851 , n21466 );
nor ( n34882 , n34880 , n34881 );
xnor ( n34883 , n34882 , n21331 );
and ( n34884 , n34878 , n34883 );
and ( n34885 , n34874 , n34883 );
or ( n34886 , n34879 , n34884 , n34885 );
and ( n34887 , n34870 , n34886 );
and ( n34888 , n24621 , n23230 );
and ( n34889 , n24527 , n23228 );
nor ( n34890 , n34888 , n34889 );
xnor ( n34891 , n34890 , n22842 );
and ( n34892 , n25284 , n22859 );
and ( n34893 , n24940 , n22857 );
nor ( n34894 , n34892 , n34893 );
xnor ( n34895 , n34894 , n22418 );
and ( n34896 , n34891 , n34895 );
and ( n34897 , n25765 , n22381 );
and ( n34898 , n25554 , n22379 );
nor ( n34899 , n34897 , n34898 );
xnor ( n34900 , n34899 , n22228 );
and ( n34901 , n34895 , n34900 );
and ( n34902 , n34891 , n34900 );
or ( n34903 , n34896 , n34901 , n34902 );
and ( n34904 , n34903 , n34568 );
xor ( n34905 , n34510 , n34514 );
xor ( n34906 , n34905 , n34519 );
and ( n34907 , n34568 , n34906 );
and ( n34908 , n34903 , n34906 );
or ( n34909 , n34904 , n34907 , n34908 );
and ( n34910 , n34886 , n34909 );
and ( n34911 , n34870 , n34909 );
or ( n34912 , n34887 , n34910 , n34911 );
and ( n34913 , n34854 , n34912 );
xor ( n34914 , n34573 , n34577 );
xor ( n34915 , n34914 , n34582 );
and ( n34916 , n34912 , n34915 );
and ( n34917 , n34854 , n34915 );
or ( n34918 , n34913 , n34916 , n34917 );
xor ( n34919 , n34597 , n34601 );
xor ( n34920 , n34919 , n34606 );
xor ( n34921 , n34506 , n34534 );
xor ( n34922 , n34921 , n34539 );
and ( n34923 , n34920 , n34922 );
xor ( n34924 , n34613 , n34617 );
xor ( n34925 , n34924 , n34620 );
and ( n34926 , n34922 , n34925 );
and ( n34927 , n34920 , n34925 );
or ( n34928 , n34923 , n34926 , n34927 );
and ( n34929 , n34918 , n34928 );
xor ( n34930 , n34304 , n34344 );
xor ( n34931 , n34930 , n34347 );
and ( n34932 , n34928 , n34931 );
and ( n34933 , n34918 , n34931 );
or ( n34934 , n34929 , n34932 , n34933 );
and ( n34935 , n34838 , n34934 );
xor ( n34936 , n34593 , n34629 );
xor ( n34937 , n34936 , n34632 );
and ( n34938 , n34934 , n34937 );
and ( n34939 , n34838 , n34937 );
or ( n34940 , n34935 , n34938 , n34939 );
xor ( n34941 , n34765 , n34769 );
and ( n34942 , n23141 , n24902 );
and ( n34943 , n22916 , n24900 );
nor ( n34944 , n34942 , n34943 );
xnor ( n34945 , n34944 , n24397 );
and ( n34946 , n34941 , n34945 );
and ( n34947 , n23381 , n24376 );
and ( n34948 , n23271 , n24374 );
nor ( n34949 , n34947 , n34948 );
xnor ( n34950 , n34949 , n23927 );
and ( n34951 , n34945 , n34950 );
and ( n34952 , n34941 , n34950 );
or ( n34953 , n34946 , n34951 , n34952 );
and ( n34954 , n29318 , n20460 );
and ( n34955 , n29078 , n20458 );
nor ( n34956 , n34954 , n34955 );
xnor ( n34957 , n34956 , n20337 );
and ( n34958 , n34953 , n34957 );
xor ( n34959 , n34770 , n34774 );
xor ( n34960 , n34959 , n34779 );
and ( n34961 , n34957 , n34960 );
and ( n34962 , n34953 , n34960 );
or ( n34963 , n34958 , n34961 , n34962 );
xor ( n34964 , n34494 , n34498 );
xor ( n34965 , n34964 , n34503 );
and ( n34966 , n34963 , n34965 );
xor ( n34967 , n34685 , n34689 );
xor ( n34968 , n34967 , n34692 );
and ( n34969 , n34965 , n34968 );
and ( n34970 , n34963 , n34968 );
or ( n34971 , n34966 , n34969 , n34970 );
xor ( n34972 , n34681 , n34695 );
xor ( n34973 , n34972 , n34698 );
and ( n34974 , n34971 , n34973 );
xor ( n34975 , n34788 , n34790 );
xor ( n34976 , n34975 , n34793 );
and ( n34977 , n34973 , n34976 );
and ( n34978 , n34971 , n34976 );
or ( n34979 , n34974 , n34977 , n34978 );
xor ( n34980 , n34609 , n34623 );
xor ( n34981 , n34980 , n34626 );
and ( n34982 , n34979 , n34981 );
xor ( n34983 , n34542 , n34544 );
xor ( n34984 , n34983 , n34547 );
and ( n34985 , n34981 , n34984 );
and ( n34986 , n34979 , n34984 );
or ( n34987 , n34982 , n34985 , n34986 );
xor ( n34988 , n34550 , n34552 );
xor ( n34989 , n34988 , n34555 );
and ( n34990 , n34987 , n34989 );
xor ( n34991 , n34709 , n34711 );
xor ( n34992 , n34991 , n34714 );
and ( n34993 , n34989 , n34992 );
and ( n34994 , n34987 , n34992 );
or ( n34995 , n34990 , n34993 , n34994 );
and ( n34996 , n34940 , n34995 );
xor ( n34997 , n34558 , n34635 );
xor ( n34998 , n34997 , n34638 );
and ( n34999 , n34995 , n34998 );
and ( n35000 , n34940 , n34998 );
or ( n35001 , n34996 , n34999 , n35000 );
xor ( n35002 , n34490 , n34641 );
xor ( n35003 , n35002 , n34644 );
and ( n35004 , n35001 , n35003 );
xor ( n35005 , n34725 , n34727 );
xor ( n35006 , n35005 , n34730 );
and ( n35007 , n35003 , n35006 );
and ( n35008 , n35001 , n35006 );
or ( n35009 , n35004 , n35007 , n35008 );
and ( n35010 , n34745 , n35009 );
xor ( n35011 , n34745 , n35009 );
xor ( n35012 , n35001 , n35003 );
xor ( n35013 , n35012 , n35006 );
and ( n35014 , n20803 , n28628 );
and ( n35015 , n20666 , n28626 );
nor ( n35016 , n35014 , n35015 );
xnor ( n35017 , n35016 , n28096 );
and ( n35018 , n21302 , n27529 );
and ( n35019 , n21218 , n27527 );
nor ( n35020 , n35018 , n35019 );
xnor ( n35021 , n35020 , n27034 );
and ( n35022 , n35017 , n35021 );
and ( n35023 , n21612 , n26992 );
and ( n35024 , n21451 , n26990 );
nor ( n35025 , n35023 , n35024 );
xnor ( n35026 , n35025 , n26369 );
and ( n35027 , n35021 , n35026 );
and ( n35028 , n35017 , n35026 );
or ( n35029 , n35022 , n35027 , n35028 );
and ( n35030 , n20360 , n29977 );
and ( n35031 , n20268 , n29974 );
nor ( n35032 , n35030 , n35031 );
xnor ( n35033 , n35032 , n28674 );
and ( n35034 , n20618 , n29276 );
and ( n35035 , n20452 , n29274 );
nor ( n35036 , n35034 , n35035 );
xnor ( n35037 , n35036 , n28677 );
and ( n35038 , n35033 , n35037 );
xor ( n35039 , n34749 , n34753 );
xor ( n35040 , n35039 , n34758 );
and ( n35041 , n35037 , n35040 );
and ( n35042 , n35033 , n35040 );
or ( n35043 , n35038 , n35041 , n35042 );
and ( n35044 , n35029 , n35043 );
xor ( n35045 , n34842 , n34846 );
xor ( n35046 , n35045 , n34851 );
and ( n35047 , n35043 , n35046 );
and ( n35048 , n35029 , n35046 );
or ( n35049 , n35044 , n35047 , n35048 );
and ( n35050 , n24131 , n23944 );
and ( n35051 , n23968 , n23942 );
nor ( n35052 , n35050 , n35051 );
xnor ( n35053 , n35052 , n23550 );
and ( n35054 , n24527 , n23641 );
and ( n35055 , n24521 , n23639 );
nor ( n35056 , n35054 , n35055 );
xnor ( n35057 , n35056 , n23213 );
and ( n35058 , n35053 , n35057 );
and ( n35059 , n24940 , n23230 );
and ( n35060 , n24621 , n23228 );
nor ( n35061 , n35059 , n35060 );
xnor ( n35062 , n35061 , n22842 );
and ( n35063 , n35057 , n35062 );
and ( n35064 , n35053 , n35062 );
or ( n35065 , n35058 , n35063 , n35064 );
and ( n35066 , n22756 , n25383 );
and ( n35067 , n22425 , n25381 );
nor ( n35068 , n35066 , n35067 );
xnor ( n35069 , n35068 , n24885 );
and ( n35070 , n35065 , n35069 );
and ( n35071 , n29623 , n20458 );
not ( n35072 , n35071 );
and ( n35073 , n35072 , n20337 );
and ( n35074 , n35069 , n35073 );
and ( n35075 , n35065 , n35073 );
or ( n35076 , n35070 , n35074 , n35075 );
and ( n35077 , n21072 , n28062 );
and ( n35078 , n20867 , n28060 );
nor ( n35079 , n35077 , n35078 );
xnor ( n35080 , n35079 , n27549 );
and ( n35081 , n35076 , n35080 );
and ( n35082 , n22235 , n26027 );
and ( n35083 , n21955 , n26025 );
nor ( n35084 , n35082 , n35083 );
xnor ( n35085 , n35084 , n25499 );
and ( n35086 , n35080 , n35085 );
and ( n35087 , n35076 , n35085 );
or ( n35088 , n35081 , n35086 , n35087 );
xor ( n35089 , n34669 , n34673 );
xor ( n35090 , n35089 , n34678 );
and ( n35091 , n35088 , n35090 );
xor ( n35092 , n34761 , n34782 );
xor ( n35093 , n35092 , n34785 );
and ( n35094 , n35090 , n35093 );
and ( n35095 , n35088 , n35093 );
or ( n35096 , n35091 , n35094 , n35095 );
and ( n35097 , n35049 , n35096 );
and ( n35098 , n27757 , n21155 );
and ( n35099 , n27751 , n21153 );
nor ( n35100 , n35098 , n35099 );
xnor ( n35101 , n35100 , n20994 );
and ( n35102 , n29078 , n20674 );
and ( n35103 , n28700 , n20672 );
nor ( n35104 , n35102 , n35103 );
xnor ( n35105 , n35104 , n20542 );
and ( n35106 , n35101 , n35105 );
and ( n35107 , n29623 , n20460 );
and ( n35108 , n29318 , n20458 );
nor ( n35109 , n35107 , n35108 );
xnor ( n35110 , n35109 , n20337 );
and ( n35111 , n35105 , n35110 );
and ( n35112 , n35101 , n35110 );
or ( n35113 , n35106 , n35111 , n35112 );
and ( n35114 , n21876 , n26349 );
and ( n35115 , n21704 , n26347 );
nor ( n35116 , n35114 , n35115 );
xnor ( n35117 , n35116 , n25893 );
and ( n35118 , n35113 , n35117 );
xor ( n35119 , n34903 , n34568 );
xor ( n35120 , n35119 , n34906 );
and ( n35121 , n35117 , n35120 );
and ( n35122 , n35113 , n35120 );
or ( n35123 , n35118 , n35121 , n35122 );
xor ( n35124 , n34800 , n34804 );
xor ( n35125 , n35124 , n34809 );
and ( n35126 , n35123 , n35125 );
xor ( n35127 , n34816 , n34820 );
xor ( n35128 , n35127 , n34823 );
and ( n35129 , n35125 , n35128 );
and ( n35130 , n35123 , n35128 );
or ( n35131 , n35126 , n35129 , n35130 );
and ( n35132 , n35096 , n35131 );
and ( n35133 , n35049 , n35131 );
or ( n35134 , n35097 , n35132 , n35133 );
xor ( n35135 , n34701 , n34703 );
xor ( n35136 , n35135 , n34706 );
and ( n35137 , n35134 , n35136 );
xor ( n35138 , n34796 , n34832 );
xor ( n35139 , n35138 , n34835 );
and ( n35140 , n35136 , n35139 );
and ( n35141 , n35134 , n35139 );
or ( n35142 , n35137 , n35140 , n35141 );
xor ( n35143 , n34854 , n34912 );
xor ( n35144 , n35143 , n34915 );
xor ( n35145 , n34812 , n34826 );
xor ( n35146 , n35145 , n34829 );
and ( n35147 , n35144 , n35146 );
xor ( n35148 , n34920 , n34922 );
xor ( n35149 , n35148 , n34925 );
and ( n35150 , n35146 , n35149 );
and ( n35151 , n35144 , n35149 );
or ( n35152 , n35147 , n35150 , n35151 );
xor ( n35153 , n34979 , n34981 );
xor ( n35154 , n35153 , n34984 );
and ( n35155 , n35152 , n35154 );
xor ( n35156 , n34918 , n34928 );
xor ( n35157 , n35156 , n34931 );
and ( n35158 , n35154 , n35157 );
and ( n35159 , n35152 , n35157 );
or ( n35160 , n35155 , n35158 , n35159 );
and ( n35161 , n35142 , n35160 );
xor ( n35162 , n34838 , n34934 );
xor ( n35163 , n35162 , n34937 );
and ( n35164 , n35160 , n35163 );
and ( n35165 , n35142 , n35163 );
or ( n35166 , n35161 , n35164 , n35165 );
xor ( n35167 , n34717 , n34719 );
xor ( n35168 , n35167 , n34722 );
and ( n35169 , n35166 , n35168 );
xor ( n35170 , n34940 , n34995 );
xor ( n35171 , n35170 , n34998 );
and ( n35172 , n35168 , n35171 );
and ( n35173 , n35166 , n35171 );
or ( n35174 , n35169 , n35172 , n35173 );
and ( n35175 , n35013 , n35174 );
xor ( n35176 , n35013 , n35174 );
xor ( n35177 , n35166 , n35168 );
xor ( n35178 , n35177 , n35171 );
and ( n35179 , n27135 , n21741 );
and ( n35180 , n26851 , n21739 );
nor ( n35181 , n35179 , n35180 );
xnor ( n35182 , n35181 , n21605 );
and ( n35183 , n27751 , n21468 );
and ( n35184 , n27352 , n21466 );
nor ( n35185 , n35183 , n35184 );
xnor ( n35186 , n35185 , n21331 );
and ( n35187 , n35182 , n35186 );
and ( n35188 , n23573 , n24376 );
and ( n35189 , n23381 , n24374 );
nor ( n35190 , n35188 , n35189 );
xnor ( n35191 , n35190 , n23927 );
and ( n35192 , n25554 , n22859 );
and ( n35193 , n25284 , n22857 );
nor ( n35194 , n35192 , n35193 );
xnor ( n35195 , n35194 , n22418 );
xor ( n35196 , n35191 , n35195 );
and ( n35197 , n25974 , n22381 );
and ( n35198 , n25765 , n22379 );
nor ( n35199 , n35197 , n35198 );
xnor ( n35200 , n35199 , n22228 );
xor ( n35201 , n35196 , n35200 );
and ( n35202 , n35186 , n35201 );
and ( n35203 , n35182 , n35201 );
or ( n35204 , n35187 , n35202 , n35203 );
and ( n35205 , n26422 , n22048 );
and ( n35206 , n26319 , n22046 );
nor ( n35207 , n35205 , n35206 );
xnor ( n35208 , n35207 , n21853 );
and ( n35209 , n28700 , n20955 );
and ( n35210 , n28810 , n20953 );
nor ( n35211 , n35209 , n35210 );
xnor ( n35212 , n35211 , n20780 );
and ( n35213 , n35208 , n35212 );
xor ( n35214 , n35053 , n35057 );
xor ( n35215 , n35214 , n35062 );
and ( n35216 , n35212 , n35215 );
and ( n35217 , n35208 , n35215 );
or ( n35218 , n35213 , n35216 , n35217 );
and ( n35219 , n35204 , n35218 );
and ( n35220 , n22198 , n26027 );
and ( n35221 , n22235 , n26025 );
nor ( n35222 , n35220 , n35221 );
xnor ( n35223 , n35222 , n25499 );
and ( n35224 , n26319 , n22048 );
and ( n35225 , n25974 , n22046 );
nor ( n35226 , n35224 , n35225 );
xnor ( n35227 , n35226 , n21853 );
xor ( n35228 , n35223 , n35227 );
xor ( n35229 , n34891 , n34895 );
xor ( n35230 , n35229 , n34900 );
xor ( n35231 , n35228 , n35230 );
and ( n35232 , n35218 , n35231 );
and ( n35233 , n35204 , n35231 );
or ( n35234 , n35219 , n35232 , n35233 );
xor ( n35235 , n35017 , n35021 );
xor ( n35236 , n35235 , n35026 );
and ( n35237 , n35234 , n35236 );
xor ( n35238 , n34953 , n34957 );
xor ( n35239 , n35238 , n34960 );
and ( n35240 , n35236 , n35239 );
and ( n35241 , n35234 , n35239 );
or ( n35242 , n35237 , n35240 , n35241 );
and ( n35243 , n22235 , n26349 );
and ( n35244 , n21955 , n26347 );
nor ( n35245 , n35243 , n35244 );
xnor ( n35246 , n35245 , n25893 );
and ( n35247 , n28211 , n21155 );
and ( n35248 , n27757 , n21153 );
nor ( n35249 , n35247 , n35248 );
xnor ( n35250 , n35249 , n20994 );
and ( n35251 , n35246 , n35250 );
and ( n35252 , n29318 , n20674 );
and ( n35253 , n29078 , n20672 );
nor ( n35254 , n35252 , n35253 );
xnor ( n35255 , n35254 , n20542 );
and ( n35256 , n35250 , n35255 );
and ( n35257 , n35246 , n35255 );
or ( n35258 , n35251 , n35256 , n35257 );
and ( n35259 , n26851 , n21741 );
and ( n35260 , n26422 , n21739 );
nor ( n35261 , n35259 , n35260 );
xnor ( n35262 , n35261 , n21605 );
and ( n35263 , n27352 , n21468 );
and ( n35264 , n27135 , n21466 );
nor ( n35265 , n35263 , n35264 );
xnor ( n35266 , n35265 , n21331 );
xor ( n35267 , n35262 , n35266 );
and ( n35268 , n28810 , n20955 );
and ( n35269 , n28211 , n20953 );
nor ( n35270 , n35268 , n35269 );
xnor ( n35271 , n35270 , n20780 );
xor ( n35272 , n35267 , n35271 );
and ( n35273 , n35258 , n35272 );
xor ( n35274 , n35101 , n35105 );
xor ( n35275 , n35274 , n35110 );
and ( n35276 , n35272 , n35275 );
and ( n35277 , n35258 , n35275 );
or ( n35278 , n35273 , n35276 , n35277 );
and ( n35279 , n35262 , n35266 );
and ( n35280 , n35266 , n35271 );
and ( n35281 , n35262 , n35271 );
or ( n35282 , n35279 , n35280 , n35281 );
and ( n35283 , n35191 , n35195 );
and ( n35284 , n35195 , n35200 );
and ( n35285 , n35191 , n35200 );
or ( n35286 , n35283 , n35284 , n35285 );
and ( n35287 , n24621 , n23641 );
and ( n35288 , n24527 , n23639 );
nor ( n35289 , n35287 , n35288 );
xnor ( n35290 , n35289 , n23213 );
and ( n35291 , n25284 , n23230 );
and ( n35292 , n24940 , n23228 );
nor ( n35293 , n35291 , n35292 );
xnor ( n35294 , n35293 , n22842 );
and ( n35295 , n35290 , n35294 );
and ( n35296 , n25765 , n22859 );
and ( n35297 , n25554 , n22857 );
nor ( n35298 , n35296 , n35297 );
xnor ( n35299 , n35298 , n22418 );
and ( n35300 , n35294 , n35299 );
and ( n35301 , n35290 , n35299 );
or ( n35302 , n35295 , n35300 , n35301 );
and ( n35303 , n23271 , n24902 );
and ( n35304 , n23141 , n24900 );
nor ( n35305 , n35303 , n35304 );
xnor ( n35306 , n35305 , n24397 );
and ( n35307 , n35302 , n35306 );
and ( n35308 , n35306 , n35071 );
and ( n35309 , n35302 , n35071 );
or ( n35310 , n35307 , n35308 , n35309 );
and ( n35311 , n35286 , n35310 );
and ( n35312 , n23968 , n24376 );
and ( n35313 , n23573 , n24374 );
nor ( n35314 , n35312 , n35313 );
xnor ( n35315 , n35314 , n23927 );
and ( n35316 , n24521 , n23944 );
and ( n35317 , n24131 , n23942 );
nor ( n35318 , n35316 , n35317 );
xnor ( n35319 , n35318 , n23550 );
and ( n35320 , n35315 , n35319 );
and ( n35321 , n22425 , n26027 );
and ( n35322 , n22198 , n26025 );
nor ( n35323 , n35321 , n35322 );
xnor ( n35324 , n35323 , n25499 );
and ( n35325 , n35320 , n35324 );
and ( n35326 , n22916 , n25383 );
and ( n35327 , n22756 , n25381 );
nor ( n35328 , n35326 , n35327 );
xnor ( n35329 , n35328 , n24885 );
and ( n35330 , n35324 , n35329 );
and ( n35331 , n35320 , n35329 );
or ( n35332 , n35325 , n35330 , n35331 );
and ( n35333 , n35310 , n35332 );
and ( n35334 , n35286 , n35332 );
or ( n35335 , n35311 , n35333 , n35334 );
xor ( n35336 , n35282 , n35335 );
and ( n35337 , n35223 , n35227 );
and ( n35338 , n35227 , n35230 );
and ( n35339 , n35223 , n35230 );
or ( n35340 , n35337 , n35338 , n35339 );
xor ( n35341 , n35336 , n35340 );
and ( n35342 , n35278 , n35341 );
xor ( n35343 , n35033 , n35037 );
xor ( n35344 , n35343 , n35040 );
and ( n35345 , n35341 , n35344 );
and ( n35346 , n35278 , n35344 );
or ( n35347 , n35342 , n35345 , n35346 );
and ( n35348 , n35242 , n35347 );
xor ( n35349 , n35088 , n35090 );
xor ( n35350 , n35349 , n35093 );
and ( n35351 , n35347 , n35350 );
and ( n35352 , n35242 , n35350 );
or ( n35353 , n35348 , n35351 , n35352 );
and ( n35354 , n20618 , n29977 );
and ( n35355 , n20452 , n29974 );
nor ( n35356 , n35354 , n35355 );
xnor ( n35357 , n35356 , n28674 );
and ( n35358 , n21612 , n27529 );
and ( n35359 , n21451 , n27527 );
nor ( n35360 , n35358 , n35359 );
xnor ( n35361 , n35360 , n27034 );
and ( n35362 , n35357 , n35361 );
and ( n35363 , n21876 , n26992 );
and ( n35364 , n21704 , n26990 );
nor ( n35365 , n35363 , n35364 );
xnor ( n35366 , n35365 , n26369 );
and ( n35367 , n35361 , n35366 );
and ( n35368 , n35357 , n35366 );
or ( n35369 , n35362 , n35367 , n35368 );
and ( n35370 , n23141 , n25383 );
and ( n35371 , n22916 , n25381 );
nor ( n35372 , n35370 , n35371 );
xnor ( n35373 , n35372 , n24885 );
and ( n35374 , n23381 , n24902 );
and ( n35375 , n23271 , n24900 );
nor ( n35376 , n35374 , n35375 );
xnor ( n35377 , n35376 , n24397 );
and ( n35378 , n35373 , n35377 );
and ( n35379 , n29623 , n20672 );
not ( n35380 , n35379 );
and ( n35381 , n35380 , n20542 );
and ( n35382 , n35377 , n35381 );
and ( n35383 , n35373 , n35381 );
or ( n35384 , n35378 , n35382 , n35383 );
xor ( n35385 , n35315 , n35319 );
and ( n35386 , n22756 , n26027 );
and ( n35387 , n22425 , n26025 );
nor ( n35388 , n35386 , n35387 );
xnor ( n35389 , n35388 , n25499 );
and ( n35390 , n35385 , n35389 );
and ( n35391 , n26319 , n22381 );
and ( n35392 , n25974 , n22379 );
nor ( n35393 , n35391 , n35392 );
xnor ( n35394 , n35393 , n22228 );
and ( n35395 , n35389 , n35394 );
and ( n35396 , n35385 , n35394 );
or ( n35397 , n35390 , n35395 , n35396 );
and ( n35398 , n35384 , n35397 );
and ( n35399 , n21302 , n28062 );
and ( n35400 , n21218 , n28060 );
nor ( n35401 , n35399 , n35400 );
xnor ( n35402 , n35401 , n27549 );
and ( n35403 , n35397 , n35402 );
and ( n35404 , n35384 , n35402 );
or ( n35405 , n35398 , n35403 , n35404 );
and ( n35406 , n35369 , n35405 );
xor ( n35407 , n35286 , n35310 );
xor ( n35408 , n35407 , n35332 );
and ( n35409 , n35405 , n35408 );
and ( n35410 , n35369 , n35408 );
or ( n35411 , n35406 , n35409 , n35410 );
xor ( n35412 , n34858 , n34862 );
xor ( n35413 , n35412 , n34867 );
xor ( n35414 , n34874 , n34878 );
xor ( n35415 , n35414 , n34883 );
xor ( n35416 , n35413 , n35415 );
xor ( n35417 , n35076 , n35080 );
xor ( n35418 , n35417 , n35085 );
xor ( n35419 , n35416 , n35418 );
and ( n35420 , n35411 , n35419 );
xor ( n35421 , n35113 , n35117 );
xor ( n35422 , n35421 , n35120 );
and ( n35423 , n35419 , n35422 );
and ( n35424 , n35411 , n35422 );
or ( n35425 , n35420 , n35423 , n35424 );
xor ( n35426 , n35123 , n35125 );
xor ( n35427 , n35426 , n35128 );
and ( n35428 , n35425 , n35427 );
and ( n35429 , n35282 , n35335 );
and ( n35430 , n35335 , n35340 );
and ( n35431 , n35282 , n35340 );
or ( n35432 , n35429 , n35430 , n35431 );
xor ( n35433 , n34870 , n34886 );
xor ( n35434 , n35433 , n34909 );
xor ( n35435 , n35432 , n35434 );
xor ( n35436 , n34963 , n34965 );
xor ( n35437 , n35436 , n34968 );
xor ( n35438 , n35435 , n35437 );
and ( n35439 , n35427 , n35438 );
and ( n35440 , n35425 , n35438 );
or ( n35441 , n35428 , n35439 , n35440 );
and ( n35442 , n35353 , n35441 );
xor ( n35443 , n35049 , n35096 );
xor ( n35444 , n35443 , n35131 );
and ( n35445 , n35441 , n35444 );
and ( n35446 , n35353 , n35444 );
or ( n35447 , n35442 , n35445 , n35446 );
and ( n35448 , n20452 , n29977 );
and ( n35449 , n20360 , n29974 );
nor ( n35450 , n35448 , n35449 );
xnor ( n35451 , n35450 , n28674 );
and ( n35452 , n20666 , n29276 );
and ( n35453 , n20618 , n29274 );
nor ( n35454 , n35452 , n35453 );
xnor ( n35455 , n35454 , n28677 );
and ( n35456 , n35451 , n35455 );
and ( n35457 , n21218 , n28062 );
and ( n35458 , n21072 , n28060 );
nor ( n35459 , n35457 , n35458 );
xnor ( n35460 , n35459 , n27549 );
and ( n35461 , n35455 , n35460 );
and ( n35462 , n35451 , n35460 );
or ( n35463 , n35456 , n35461 , n35462 );
and ( n35464 , n20867 , n28628 );
and ( n35465 , n20803 , n28626 );
nor ( n35466 , n35464 , n35465 );
xnor ( n35467 , n35466 , n28096 );
and ( n35468 , n21704 , n26992 );
and ( n35469 , n21612 , n26990 );
nor ( n35470 , n35468 , n35469 );
xnor ( n35471 , n35470 , n26369 );
and ( n35472 , n35467 , n35471 );
and ( n35473 , n21955 , n26349 );
and ( n35474 , n21876 , n26347 );
nor ( n35475 , n35473 , n35474 );
xnor ( n35476 , n35475 , n25893 );
and ( n35477 , n35471 , n35476 );
and ( n35478 , n35467 , n35476 );
or ( n35479 , n35472 , n35477 , n35478 );
and ( n35480 , n35463 , n35479 );
and ( n35481 , n21451 , n27529 );
and ( n35482 , n21302 , n27527 );
nor ( n35483 , n35481 , n35482 );
xnor ( n35484 , n35483 , n27034 );
xor ( n35485 , n35065 , n35069 );
xor ( n35486 , n35485 , n35073 );
and ( n35487 , n35484 , n35486 );
xor ( n35488 , n34941 , n34945 );
xor ( n35489 , n35488 , n34950 );
and ( n35490 , n35486 , n35489 );
and ( n35491 , n35484 , n35489 );
or ( n35492 , n35487 , n35490 , n35491 );
and ( n35493 , n35479 , n35492 );
and ( n35494 , n35463 , n35492 );
or ( n35495 , n35480 , n35493 , n35494 );
and ( n35496 , n35413 , n35415 );
and ( n35497 , n35415 , n35418 );
and ( n35498 , n35413 , n35418 );
or ( n35499 , n35496 , n35497 , n35498 );
and ( n35500 , n35495 , n35499 );
xor ( n35501 , n35029 , n35043 );
xor ( n35502 , n35501 , n35046 );
and ( n35503 , n35499 , n35502 );
and ( n35504 , n35495 , n35502 );
or ( n35505 , n35500 , n35503 , n35504 );
and ( n35506 , n35432 , n35434 );
and ( n35507 , n35434 , n35437 );
and ( n35508 , n35432 , n35437 );
or ( n35509 , n35506 , n35507 , n35508 );
and ( n35510 , n35505 , n35509 );
xor ( n35511 , n34971 , n34973 );
xor ( n35512 , n35511 , n34976 );
and ( n35513 , n35509 , n35512 );
and ( n35514 , n35505 , n35512 );
or ( n35515 , n35510 , n35513 , n35514 );
and ( n35516 , n35447 , n35515 );
xor ( n35517 , n35134 , n35136 );
xor ( n35518 , n35517 , n35139 );
and ( n35519 , n35515 , n35518 );
and ( n35520 , n35447 , n35518 );
or ( n35521 , n35516 , n35519 , n35520 );
xor ( n35522 , n34987 , n34989 );
xor ( n35523 , n35522 , n34992 );
and ( n35524 , n35521 , n35523 );
xor ( n35525 , n35142 , n35160 );
xor ( n35526 , n35525 , n35163 );
and ( n35527 , n35523 , n35526 );
and ( n35528 , n35521 , n35526 );
or ( n35529 , n35524 , n35527 , n35528 );
and ( n35530 , n35178 , n35529 );
xor ( n35531 , n35178 , n35529 );
xor ( n35532 , n35521 , n35523 );
xor ( n35533 , n35532 , n35526 );
and ( n35534 , n24527 , n23944 );
and ( n35535 , n24521 , n23942 );
nor ( n35536 , n35534 , n35535 );
xnor ( n35537 , n35536 , n23550 );
and ( n35538 , n25974 , n22859 );
and ( n35539 , n25765 , n22857 );
nor ( n35540 , n35538 , n35539 );
xnor ( n35541 , n35540 , n22418 );
and ( n35542 , n35537 , n35541 );
and ( n35543 , n26422 , n22381 );
and ( n35544 , n26319 , n22379 );
nor ( n35545 , n35543 , n35544 );
xnor ( n35546 , n35545 , n22228 );
and ( n35547 , n35541 , n35546 );
and ( n35548 , n35537 , n35546 );
or ( n35549 , n35542 , n35547 , n35548 );
and ( n35550 , n26851 , n22048 );
and ( n35551 , n26422 , n22046 );
nor ( n35552 , n35550 , n35551 );
xnor ( n35553 , n35552 , n21853 );
and ( n35554 , n35549 , n35553 );
and ( n35555 , n27352 , n21741 );
and ( n35556 , n27135 , n21739 );
nor ( n35557 , n35555 , n35556 );
xnor ( n35558 , n35557 , n21605 );
and ( n35559 , n35553 , n35558 );
and ( n35560 , n35549 , n35558 );
or ( n35561 , n35554 , n35559 , n35560 );
and ( n35562 , n24131 , n24376 );
and ( n35563 , n23968 , n24374 );
nor ( n35564 , n35562 , n35563 );
xnor ( n35565 , n35564 , n23927 );
and ( n35566 , n24940 , n23641 );
and ( n35567 , n24621 , n23639 );
nor ( n35568 , n35566 , n35567 );
xnor ( n35569 , n35568 , n23213 );
and ( n35570 , n35565 , n35569 );
and ( n35571 , n25554 , n23230 );
and ( n35572 , n25284 , n23228 );
nor ( n35573 , n35571 , n35572 );
xnor ( n35574 , n35573 , n22842 );
and ( n35575 , n35569 , n35574 );
and ( n35576 , n35565 , n35574 );
or ( n35577 , n35570 , n35575 , n35576 );
and ( n35578 , n22198 , n26349 );
and ( n35579 , n22235 , n26347 );
nor ( n35580 , n35578 , n35579 );
xnor ( n35581 , n35580 , n25893 );
and ( n35582 , n35577 , n35581 );
xor ( n35583 , n35290 , n35294 );
xor ( n35584 , n35583 , n35299 );
and ( n35585 , n35581 , n35584 );
and ( n35586 , n35577 , n35584 );
or ( n35587 , n35582 , n35585 , n35586 );
and ( n35588 , n35561 , n35587 );
and ( n35589 , n21072 , n28628 );
and ( n35590 , n20867 , n28626 );
nor ( n35591 , n35589 , n35590 );
xnor ( n35592 , n35591 , n28096 );
and ( n35593 , n35587 , n35592 );
and ( n35594 , n35561 , n35592 );
or ( n35595 , n35588 , n35593 , n35594 );
and ( n35596 , n20803 , n29276 );
and ( n35597 , n20666 , n29274 );
nor ( n35598 , n35596 , n35597 );
xnor ( n35599 , n35598 , n28677 );
xor ( n35600 , n35302 , n35306 );
xor ( n35601 , n35600 , n35071 );
and ( n35602 , n35599 , n35601 );
xor ( n35603 , n35320 , n35324 );
xor ( n35604 , n35603 , n35329 );
and ( n35605 , n35601 , n35604 );
and ( n35606 , n35599 , n35604 );
or ( n35607 , n35602 , n35605 , n35606 );
and ( n35608 , n35595 , n35607 );
xor ( n35609 , n35451 , n35455 );
xor ( n35610 , n35609 , n35460 );
and ( n35611 , n35607 , n35610 );
and ( n35612 , n35595 , n35610 );
or ( n35613 , n35608 , n35611 , n35612 );
xor ( n35614 , n35463 , n35479 );
xor ( n35615 , n35614 , n35492 );
and ( n35616 , n35613 , n35615 );
xor ( n35617 , n35234 , n35236 );
xor ( n35618 , n35617 , n35239 );
and ( n35619 , n35615 , n35618 );
and ( n35620 , n35613 , n35618 );
or ( n35621 , n35616 , n35619 , n35620 );
xor ( n35622 , n35495 , n35499 );
xor ( n35623 , n35622 , n35502 );
and ( n35624 , n35621 , n35623 );
xor ( n35625 , n35242 , n35347 );
xor ( n35626 , n35625 , n35350 );
and ( n35627 , n35623 , n35626 );
and ( n35628 , n35621 , n35626 );
or ( n35629 , n35624 , n35627 , n35628 );
xor ( n35630 , n35144 , n35146 );
xor ( n35631 , n35630 , n35149 );
and ( n35632 , n35629 , n35631 );
xor ( n35633 , n35505 , n35509 );
xor ( n35634 , n35633 , n35512 );
and ( n35635 , n35631 , n35634 );
and ( n35636 , n35629 , n35634 );
or ( n35637 , n35632 , n35635 , n35636 );
xor ( n35638 , n35152 , n35154 );
xor ( n35639 , n35638 , n35157 );
and ( n35640 , n35637 , n35639 );
xor ( n35641 , n35447 , n35515 );
xor ( n35642 , n35641 , n35518 );
and ( n35643 , n35639 , n35642 );
and ( n35644 , n35637 , n35642 );
or ( n35645 , n35640 , n35643 , n35644 );
and ( n35646 , n35533 , n35645 );
xor ( n35647 , n35533 , n35645 );
xor ( n35648 , n35637 , n35639 );
xor ( n35649 , n35648 , n35642 );
and ( n35650 , n27757 , n21468 );
and ( n35651 , n27751 , n21466 );
nor ( n35652 , n35650 , n35651 );
xnor ( n35653 , n35652 , n21331 );
and ( n35654 , n28810 , n21155 );
and ( n35655 , n28211 , n21153 );
nor ( n35656 , n35654 , n35655 );
xnor ( n35657 , n35656 , n20994 );
and ( n35658 , n35653 , n35657 );
and ( n35659 , n29623 , n20674 );
and ( n35660 , n29318 , n20672 );
nor ( n35661 , n35659 , n35660 );
xnor ( n35662 , n35661 , n20542 );
and ( n35663 , n35657 , n35662 );
and ( n35664 , n35653 , n35662 );
or ( n35665 , n35658 , n35663 , n35664 );
xor ( n35666 , n35182 , n35186 );
xor ( n35667 , n35666 , n35201 );
and ( n35668 , n35665 , n35667 );
xor ( n35669 , n35208 , n35212 );
xor ( n35670 , n35669 , n35215 );
and ( n35671 , n35667 , n35670 );
and ( n35672 , n35665 , n35670 );
or ( n35673 , n35668 , n35671 , n35672 );
xor ( n35674 , n35467 , n35471 );
xor ( n35675 , n35674 , n35476 );
and ( n35676 , n35673 , n35675 );
xor ( n35677 , n35484 , n35486 );
xor ( n35678 , n35677 , n35489 );
and ( n35679 , n35675 , n35678 );
and ( n35680 , n35673 , n35678 );
or ( n35681 , n35676 , n35679 , n35680 );
and ( n35682 , n20867 , n29276 );
and ( n35683 , n20803 , n29274 );
nor ( n35684 , n35682 , n35683 );
xnor ( n35685 , n35684 , n28677 );
and ( n35686 , n21955 , n26992 );
and ( n35687 , n21876 , n26990 );
nor ( n35688 , n35686 , n35687 );
xnor ( n35689 , n35688 , n26369 );
and ( n35690 , n35685 , n35689 );
xor ( n35691 , n35373 , n35377 );
xor ( n35692 , n35691 , n35381 );
and ( n35693 , n35689 , n35692 );
and ( n35694 , n35685 , n35692 );
or ( n35695 , n35690 , n35693 , n35694 );
and ( n35696 , n24521 , n24376 );
and ( n35697 , n24131 , n24374 );
nor ( n35698 , n35696 , n35697 );
xnor ( n35699 , n35698 , n23927 );
and ( n35700 , n25765 , n23230 );
and ( n35701 , n25554 , n23228 );
nor ( n35702 , n35700 , n35701 );
xnor ( n35703 , n35702 , n22842 );
and ( n35704 , n35699 , n35703 );
and ( n35705 , n23271 , n25383 );
and ( n35706 , n23141 , n25381 );
nor ( n35707 , n35705 , n35706 );
xnor ( n35708 , n35707 , n24885 );
and ( n35709 , n35704 , n35708 );
and ( n35710 , n23573 , n24902 );
and ( n35711 , n23381 , n24900 );
nor ( n35712 , n35710 , n35711 );
xnor ( n35713 , n35712 , n24397 );
and ( n35714 , n35708 , n35713 );
and ( n35715 , n35704 , n35713 );
or ( n35716 , n35709 , n35714 , n35715 );
and ( n35717 , n29078 , n20955 );
and ( n35718 , n28700 , n20953 );
nor ( n35719 , n35717 , n35718 );
xnor ( n35720 , n35719 , n20780 );
and ( n35721 , n35716 , n35720 );
xor ( n35722 , n35385 , n35389 );
xor ( n35723 , n35722 , n35394 );
and ( n35724 , n35720 , n35723 );
and ( n35725 , n35716 , n35723 );
or ( n35726 , n35721 , n35724 , n35725 );
and ( n35727 , n35695 , n35726 );
xor ( n35728 , n35246 , n35250 );
xor ( n35729 , n35728 , n35255 );
and ( n35730 , n35726 , n35729 );
and ( n35731 , n35695 , n35729 );
or ( n35732 , n35727 , n35730 , n35731 );
xor ( n35733 , n35258 , n35272 );
xor ( n35734 , n35733 , n35275 );
and ( n35735 , n35732 , n35734 );
xor ( n35736 , n35204 , n35218 );
xor ( n35737 , n35736 , n35231 );
and ( n35738 , n35734 , n35737 );
and ( n35739 , n35732 , n35737 );
or ( n35740 , n35735 , n35738 , n35739 );
and ( n35741 , n35681 , n35740 );
xor ( n35742 , n35278 , n35341 );
xor ( n35743 , n35742 , n35344 );
and ( n35744 , n35740 , n35743 );
and ( n35745 , n35681 , n35743 );
or ( n35746 , n35741 , n35744 , n35745 );
and ( n35747 , n22425 , n26349 );
and ( n35748 , n22198 , n26347 );
nor ( n35749 , n35747 , n35748 );
xnor ( n35750 , n35749 , n25893 );
and ( n35751 , n22916 , n26027 );
and ( n35752 , n22756 , n26025 );
nor ( n35753 , n35751 , n35752 );
xnor ( n35754 , n35753 , n25499 );
and ( n35755 , n35750 , n35754 );
and ( n35756 , n35754 , n35379 );
and ( n35757 , n35750 , n35379 );
or ( n35758 , n35755 , n35756 , n35757 );
and ( n35759 , n21451 , n28062 );
and ( n35760 , n21302 , n28060 );
nor ( n35761 , n35759 , n35760 );
xnor ( n35762 , n35761 , n27549 );
and ( n35763 , n35758 , n35762 );
and ( n35764 , n21704 , n27529 );
and ( n35765 , n21612 , n27527 );
nor ( n35766 , n35764 , n35765 );
xnor ( n35767 , n35766 , n27034 );
and ( n35768 , n35762 , n35767 );
and ( n35769 , n35758 , n35767 );
or ( n35770 , n35763 , n35768 , n35769 );
and ( n35771 , n23968 , n24902 );
and ( n35772 , n23573 , n24900 );
nor ( n35773 , n35771 , n35772 );
xnor ( n35774 , n35773 , n24397 );
and ( n35775 , n24621 , n23944 );
and ( n35776 , n24527 , n23942 );
nor ( n35777 , n35775 , n35776 );
xnor ( n35778 , n35777 , n23550 );
and ( n35779 , n35774 , n35778 );
and ( n35780 , n25284 , n23641 );
and ( n35781 , n24940 , n23639 );
nor ( n35782 , n35780 , n35781 );
xnor ( n35783 , n35782 , n23213 );
and ( n35784 , n35778 , n35783 );
and ( n35785 , n35774 , n35783 );
or ( n35786 , n35779 , n35784 , n35785 );
xor ( n35787 , n35565 , n35569 );
xor ( n35788 , n35787 , n35574 );
and ( n35789 , n35786 , n35788 );
xor ( n35790 , n35537 , n35541 );
xor ( n35791 , n35790 , n35546 );
and ( n35792 , n35788 , n35791 );
and ( n35793 , n35786 , n35791 );
or ( n35794 , n35789 , n35792 , n35793 );
and ( n35795 , n20666 , n29977 );
and ( n35796 , n20618 , n29974 );
nor ( n35797 , n35795 , n35796 );
xnor ( n35798 , n35797 , n28674 );
and ( n35799 , n35794 , n35798 );
and ( n35800 , n21218 , n28628 );
and ( n35801 , n21072 , n28626 );
nor ( n35802 , n35800 , n35801 );
xnor ( n35803 , n35802 , n28096 );
and ( n35804 , n35798 , n35803 );
and ( n35805 , n35794 , n35803 );
or ( n35806 , n35799 , n35804 , n35805 );
and ( n35807 , n35770 , n35806 );
xor ( n35808 , n35384 , n35397 );
xor ( n35809 , n35808 , n35402 );
and ( n35810 , n35806 , n35809 );
and ( n35811 , n35770 , n35809 );
or ( n35812 , n35807 , n35810 , n35811 );
and ( n35813 , n27135 , n22048 );
and ( n35814 , n26851 , n22046 );
nor ( n35815 , n35813 , n35814 );
xnor ( n35816 , n35815 , n21853 );
and ( n35817 , n27751 , n21741 );
and ( n35818 , n27352 , n21739 );
nor ( n35819 , n35817 , n35818 );
xnor ( n35820 , n35819 , n21605 );
and ( n35821 , n35816 , n35820 );
and ( n35822 , n28211 , n21468 );
and ( n35823 , n27757 , n21466 );
nor ( n35824 , n35822 , n35823 );
xnor ( n35825 , n35824 , n21331 );
and ( n35826 , n35820 , n35825 );
and ( n35827 , n35816 , n35825 );
or ( n35828 , n35821 , n35826 , n35827 );
xor ( n35829 , n35699 , n35703 );
and ( n35830 , n26319 , n22859 );
and ( n35831 , n25974 , n22857 );
nor ( n35832 , n35830 , n35831 );
xnor ( n35833 , n35832 , n22418 );
and ( n35834 , n35829 , n35833 );
and ( n35835 , n26851 , n22381 );
and ( n35836 , n26422 , n22379 );
nor ( n35837 , n35835 , n35836 );
xnor ( n35838 , n35837 , n22228 );
and ( n35839 , n35833 , n35838 );
and ( n35840 , n35829 , n35838 );
or ( n35841 , n35834 , n35839 , n35840 );
and ( n35842 , n28700 , n21155 );
and ( n35843 , n28810 , n21153 );
nor ( n35844 , n35842 , n35843 );
xnor ( n35845 , n35844 , n20994 );
and ( n35846 , n35841 , n35845 );
and ( n35847 , n29318 , n20955 );
and ( n35848 , n29078 , n20953 );
nor ( n35849 , n35847 , n35848 );
xnor ( n35850 , n35849 , n20780 );
and ( n35851 , n35845 , n35850 );
and ( n35852 , n35841 , n35850 );
or ( n35853 , n35846 , n35851 , n35852 );
and ( n35854 , n35828 , n35853 );
xor ( n35855 , n35577 , n35581 );
xor ( n35856 , n35855 , n35584 );
and ( n35857 , n35853 , n35856 );
and ( n35858 , n35828 , n35856 );
or ( n35859 , n35854 , n35857 , n35858 );
xor ( n35860 , n35357 , n35361 );
xor ( n35861 , n35860 , n35366 );
and ( n35862 , n35859 , n35861 );
xor ( n35863 , n35561 , n35587 );
xor ( n35864 , n35863 , n35592 );
and ( n35865 , n35861 , n35864 );
and ( n35866 , n35859 , n35864 );
or ( n35867 , n35862 , n35865 , n35866 );
and ( n35868 , n35812 , n35867 );
xor ( n35869 , n35369 , n35405 );
xor ( n35870 , n35869 , n35408 );
and ( n35871 , n35867 , n35870 );
and ( n35872 , n35812 , n35870 );
or ( n35873 , n35868 , n35871 , n35872 );
xor ( n35874 , n35411 , n35419 );
xor ( n35875 , n35874 , n35422 );
and ( n35876 , n35873 , n35875 );
xor ( n35877 , n35613 , n35615 );
xor ( n35878 , n35877 , n35618 );
and ( n35879 , n35875 , n35878 );
and ( n35880 , n35873 , n35878 );
or ( n35881 , n35876 , n35879 , n35880 );
and ( n35882 , n35746 , n35881 );
xor ( n35883 , n35425 , n35427 );
xor ( n35884 , n35883 , n35438 );
and ( n35885 , n35881 , n35884 );
and ( n35886 , n35746 , n35884 );
or ( n35887 , n35882 , n35885 , n35886 );
xor ( n35888 , n35353 , n35441 );
xor ( n35889 , n35888 , n35444 );
and ( n35890 , n35887 , n35889 );
xor ( n35891 , n35629 , n35631 );
xor ( n35892 , n35891 , n35634 );
and ( n35893 , n35889 , n35892 );
and ( n35894 , n35887 , n35892 );
or ( n35895 , n35890 , n35893 , n35894 );
and ( n35896 , n35649 , n35895 );
xor ( n35897 , n35649 , n35895 );
xor ( n35898 , n35887 , n35889 );
xor ( n35899 , n35898 , n35892 );
and ( n35900 , n22756 , n26349 );
and ( n35901 , n22425 , n26347 );
nor ( n35902 , n35900 , n35901 );
xnor ( n35903 , n35902 , n25893 );
and ( n35904 , n23141 , n26027 );
and ( n35905 , n22916 , n26025 );
nor ( n35906 , n35904 , n35905 );
xnor ( n35907 , n35906 , n25499 );
and ( n35908 , n35903 , n35907 );
and ( n35909 , n23381 , n25383 );
and ( n35910 , n23271 , n25381 );
nor ( n35911 , n35909 , n35910 );
xnor ( n35912 , n35911 , n24885 );
and ( n35913 , n35907 , n35912 );
and ( n35914 , n35903 , n35912 );
or ( n35915 , n35908 , n35913 , n35914 );
and ( n35916 , n22235 , n26992 );
and ( n35917 , n21955 , n26990 );
nor ( n35918 , n35916 , n35917 );
xnor ( n35919 , n35918 , n26369 );
and ( n35920 , n35915 , n35919 );
xor ( n35921 , n35704 , n35708 );
xor ( n35922 , n35921 , n35713 );
and ( n35923 , n35919 , n35922 );
and ( n35924 , n35915 , n35922 );
or ( n35925 , n35920 , n35923 , n35924 );
xor ( n35926 , n35653 , n35657 );
xor ( n35927 , n35926 , n35662 );
and ( n35928 , n35925 , n35927 );
xor ( n35929 , n35549 , n35553 );
xor ( n35930 , n35929 , n35558 );
and ( n35931 , n35927 , n35930 );
and ( n35932 , n35925 , n35930 );
or ( n35933 , n35928 , n35931 , n35932 );
and ( n35934 , n21072 , n29276 );
and ( n35935 , n20867 , n29274 );
nor ( n35936 , n35934 , n35935 );
xnor ( n35937 , n35936 , n28677 );
and ( n35938 , n21302 , n28628 );
and ( n35939 , n21218 , n28626 );
nor ( n35940 , n35938 , n35939 );
xnor ( n35941 , n35940 , n28096 );
and ( n35942 , n35937 , n35941 );
and ( n35943 , n21876 , n27529 );
and ( n35944 , n21704 , n27527 );
nor ( n35945 , n35943 , n35944 );
xnor ( n35946 , n35945 , n27034 );
and ( n35947 , n35941 , n35946 );
and ( n35948 , n35937 , n35946 );
or ( n35949 , n35942 , n35947 , n35948 );
and ( n35950 , n24131 , n24902 );
and ( n35951 , n23968 , n24900 );
nor ( n35952 , n35950 , n35951 );
xnor ( n35953 , n35952 , n24397 );
and ( n35954 , n24527 , n24376 );
and ( n35955 , n24521 , n24374 );
nor ( n35956 , n35954 , n35955 );
xnor ( n35957 , n35956 , n23927 );
and ( n35958 , n35953 , n35957 );
and ( n35959 , n25974 , n23230 );
and ( n35960 , n25765 , n23228 );
nor ( n35961 , n35959 , n35960 );
xnor ( n35962 , n35961 , n22842 );
and ( n35963 , n35957 , n35962 );
and ( n35964 , n35953 , n35962 );
or ( n35965 , n35958 , n35963 , n35964 );
and ( n35966 , n24940 , n23944 );
and ( n35967 , n24621 , n23942 );
nor ( n35968 , n35966 , n35967 );
xnor ( n35969 , n35968 , n23550 );
and ( n35970 , n25554 , n23641 );
and ( n35971 , n25284 , n23639 );
nor ( n35972 , n35970 , n35971 );
xnor ( n35973 , n35972 , n23213 );
and ( n35974 , n35969 , n35973 );
and ( n35975 , n26422 , n22859 );
and ( n35976 , n26319 , n22857 );
nor ( n35977 , n35975 , n35976 );
xnor ( n35978 , n35977 , n22418 );
and ( n35979 , n35973 , n35978 );
and ( n35980 , n35969 , n35978 );
or ( n35981 , n35974 , n35979 , n35980 );
and ( n35982 , n35965 , n35981 );
and ( n35983 , n29623 , n20953 );
not ( n35984 , n35983 );
and ( n35985 , n35984 , n20780 );
and ( n35986 , n35981 , n35985 );
and ( n35987 , n35965 , n35985 );
or ( n35988 , n35982 , n35986 , n35987 );
and ( n35989 , n21612 , n28062 );
and ( n35990 , n21451 , n28060 );
nor ( n35991 , n35989 , n35990 );
xnor ( n35992 , n35991 , n27549 );
and ( n35993 , n35988 , n35992 );
xor ( n35994 , n35750 , n35754 );
xor ( n35995 , n35994 , n35379 );
and ( n35996 , n35992 , n35995 );
and ( n35997 , n35988 , n35995 );
or ( n35998 , n35993 , n35996 , n35997 );
and ( n35999 , n35949 , n35998 );
xor ( n36000 , n35716 , n35720 );
xor ( n36001 , n36000 , n35723 );
and ( n36002 , n35998 , n36001 );
and ( n36003 , n35949 , n36001 );
or ( n36004 , n35999 , n36002 , n36003 );
and ( n36005 , n35933 , n36004 );
xor ( n36006 , n35599 , n35601 );
xor ( n36007 , n36006 , n35604 );
and ( n36008 , n36004 , n36007 );
and ( n36009 , n35933 , n36007 );
or ( n36010 , n36005 , n36008 , n36009 );
xor ( n36011 , n35595 , n35607 );
xor ( n36012 , n36011 , n35610 );
and ( n36013 , n36010 , n36012 );
xor ( n36014 , n35673 , n35675 );
xor ( n36015 , n36014 , n35678 );
and ( n36016 , n36012 , n36015 );
and ( n36017 , n36010 , n36015 );
or ( n36018 , n36013 , n36016 , n36017 );
xor ( n36019 , n35695 , n35726 );
xor ( n36020 , n36019 , n35729 );
xor ( n36021 , n35770 , n35806 );
xor ( n36022 , n36021 , n35809 );
and ( n36023 , n36020 , n36022 );
xor ( n36024 , n35665 , n35667 );
xor ( n36025 , n36024 , n35670 );
and ( n36026 , n36022 , n36025 );
and ( n36027 , n36020 , n36025 );
or ( n36028 , n36023 , n36026 , n36027 );
xor ( n36029 , n35812 , n35867 );
xor ( n36030 , n36029 , n35870 );
and ( n36031 , n36028 , n36030 );
xor ( n36032 , n35732 , n35734 );
xor ( n36033 , n36032 , n35737 );
and ( n36034 , n36030 , n36033 );
and ( n36035 , n36028 , n36033 );
or ( n36036 , n36031 , n36034 , n36035 );
and ( n36037 , n36018 , n36036 );
xor ( n36038 , n35681 , n35740 );
xor ( n36039 , n36038 , n35743 );
and ( n36040 , n36036 , n36039 );
and ( n36041 , n36018 , n36039 );
or ( n36042 , n36037 , n36040 , n36041 );
xor ( n36043 , n35621 , n35623 );
xor ( n36044 , n36043 , n35626 );
and ( n36045 , n36042 , n36044 );
xor ( n36046 , n35746 , n35881 );
xor ( n36047 , n36046 , n35884 );
and ( n36048 , n36044 , n36047 );
and ( n36049 , n36042 , n36047 );
or ( n36050 , n36045 , n36048 , n36049 );
and ( n36051 , n35899 , n36050 );
xor ( n36052 , n35899 , n36050 );
xor ( n36053 , n36042 , n36044 );
xor ( n36054 , n36053 , n36047 );
xor ( n36055 , n35758 , n35762 );
xor ( n36056 , n36055 , n35767 );
xor ( n36057 , n35794 , n35798 );
xor ( n36058 , n36057 , n35803 );
and ( n36059 , n36056 , n36058 );
xor ( n36060 , n35685 , n35689 );
xor ( n36061 , n36060 , n35692 );
and ( n36062 , n36058 , n36061 );
and ( n36063 , n36056 , n36061 );
or ( n36064 , n36059 , n36062 , n36063 );
and ( n36065 , n24521 , n24902 );
and ( n36066 , n24131 , n24900 );
nor ( n36067 , n36065 , n36066 );
xnor ( n36068 , n36067 , n24397 );
and ( n36069 , n26319 , n23230 );
and ( n36070 , n25974 , n23228 );
nor ( n36071 , n36069 , n36070 );
xnor ( n36072 , n36071 , n22842 );
and ( n36073 , n36068 , n36072 );
and ( n36074 , n23573 , n25383 );
and ( n36075 , n23381 , n25381 );
nor ( n36076 , n36074 , n36075 );
xnor ( n36077 , n36076 , n24885 );
and ( n36078 , n36073 , n36077 );
and ( n36079 , n27135 , n22381 );
and ( n36080 , n26851 , n22379 );
nor ( n36081 , n36079 , n36080 );
xnor ( n36082 , n36081 , n22228 );
and ( n36083 , n36077 , n36082 );
and ( n36084 , n36073 , n36082 );
or ( n36085 , n36078 , n36083 , n36084 );
and ( n36086 , n29078 , n21155 );
and ( n36087 , n28700 , n21153 );
nor ( n36088 , n36086 , n36087 );
xnor ( n36089 , n36088 , n20994 );
and ( n36090 , n36085 , n36089 );
and ( n36091 , n29623 , n20955 );
and ( n36092 , n29318 , n20953 );
nor ( n36093 , n36091 , n36092 );
xnor ( n36094 , n36093 , n20780 );
and ( n36095 , n36089 , n36094 );
and ( n36096 , n36085 , n36094 );
or ( n36097 , n36090 , n36095 , n36096 );
and ( n36098 , n22198 , n26992 );
and ( n36099 , n22235 , n26990 );
nor ( n36100 , n36098 , n36099 );
xnor ( n36101 , n36100 , n26369 );
and ( n36102 , n27352 , n22048 );
and ( n36103 , n27135 , n22046 );
nor ( n36104 , n36102 , n36103 );
xnor ( n36105 , n36104 , n21853 );
and ( n36106 , n36101 , n36105 );
xor ( n36107 , n35774 , n35778 );
xor ( n36108 , n36107 , n35783 );
and ( n36109 , n36105 , n36108 );
and ( n36110 , n36101 , n36108 );
or ( n36111 , n36106 , n36109 , n36110 );
and ( n36112 , n36097 , n36111 );
xor ( n36113 , n35816 , n35820 );
xor ( n36114 , n36113 , n35825 );
and ( n36115 , n36111 , n36114 );
and ( n36116 , n36097 , n36114 );
or ( n36117 , n36112 , n36115 , n36116 );
and ( n36118 , n27757 , n21741 );
and ( n36119 , n27751 , n21739 );
nor ( n36120 , n36118 , n36119 );
xnor ( n36121 , n36120 , n21605 );
and ( n36122 , n28810 , n21468 );
and ( n36123 , n28211 , n21466 );
nor ( n36124 , n36122 , n36123 );
xnor ( n36125 , n36124 , n21331 );
and ( n36126 , n36121 , n36125 );
xor ( n36127 , n35829 , n35833 );
xor ( n36128 , n36127 , n35838 );
and ( n36129 , n36125 , n36128 );
and ( n36130 , n36121 , n36128 );
or ( n36131 , n36126 , n36129 , n36130 );
and ( n36132 , n20803 , n29977 );
and ( n36133 , n20666 , n29974 );
nor ( n36134 , n36132 , n36133 );
xnor ( n36135 , n36134 , n28674 );
and ( n36136 , n36131 , n36135 );
xor ( n36137 , n35786 , n35788 );
xor ( n36138 , n36137 , n35791 );
and ( n36139 , n36135 , n36138 );
and ( n36140 , n36131 , n36138 );
or ( n36141 , n36136 , n36139 , n36140 );
and ( n36142 , n36117 , n36141 );
xor ( n36143 , n35828 , n35853 );
xor ( n36144 , n36143 , n35856 );
and ( n36145 , n36141 , n36144 );
and ( n36146 , n36117 , n36144 );
or ( n36147 , n36142 , n36145 , n36146 );
and ( n36148 , n36064 , n36147 );
xor ( n36149 , n35859 , n35861 );
xor ( n36150 , n36149 , n35864 );
and ( n36151 , n36147 , n36150 );
and ( n36152 , n36064 , n36150 );
or ( n36153 , n36148 , n36151 , n36152 );
and ( n36154 , n23968 , n25383 );
and ( n36155 , n23573 , n25381 );
nor ( n36156 , n36154 , n36155 );
xnor ( n36157 , n36156 , n24885 );
and ( n36158 , n24621 , n24376 );
and ( n36159 , n24527 , n24374 );
nor ( n36160 , n36158 , n36159 );
xnor ( n36161 , n36160 , n23927 );
and ( n36162 , n36157 , n36161 );
and ( n36163 , n25765 , n23641 );
and ( n36164 , n25554 , n23639 );
nor ( n36165 , n36163 , n36164 );
xnor ( n36166 , n36165 , n23213 );
and ( n36167 , n36161 , n36166 );
and ( n36168 , n36157 , n36166 );
or ( n36169 , n36162 , n36167 , n36168 );
and ( n36170 , n22916 , n26349 );
and ( n36171 , n22756 , n26347 );
nor ( n36172 , n36170 , n36171 );
xnor ( n36173 , n36172 , n25893 );
and ( n36174 , n36169 , n36173 );
xor ( n36175 , n35953 , n35957 );
xor ( n36176 , n36175 , n35962 );
and ( n36177 , n36173 , n36176 );
and ( n36178 , n36169 , n36176 );
or ( n36179 , n36174 , n36177 , n36178 );
and ( n36180 , n20867 , n29977 );
and ( n36181 , n20803 , n29974 );
nor ( n36182 , n36180 , n36181 );
xnor ( n36183 , n36182 , n28674 );
and ( n36184 , n36179 , n36183 );
and ( n36185 , n21955 , n27529 );
and ( n36186 , n21876 , n27527 );
nor ( n36187 , n36185 , n36186 );
xnor ( n36188 , n36187 , n27034 );
and ( n36189 , n36183 , n36188 );
and ( n36190 , n36179 , n36188 );
or ( n36191 , n36184 , n36189 , n36190 );
xor ( n36192 , n35841 , n35845 );
xor ( n36193 , n36192 , n35850 );
and ( n36194 , n36191 , n36193 );
xor ( n36195 , n35915 , n35919 );
xor ( n36196 , n36195 , n35922 );
and ( n36197 , n36193 , n36196 );
and ( n36198 , n36191 , n36196 );
or ( n36199 , n36194 , n36197 , n36198 );
xor ( n36200 , n35925 , n35927 );
xor ( n36201 , n36200 , n35930 );
and ( n36202 , n36199 , n36201 );
xor ( n36203 , n35949 , n35998 );
xor ( n36204 , n36203 , n36001 );
and ( n36205 , n36201 , n36204 );
and ( n36206 , n36199 , n36204 );
or ( n36207 , n36202 , n36205 , n36206 );
xor ( n36208 , n35933 , n36004 );
xor ( n36209 , n36208 , n36007 );
and ( n36210 , n36207 , n36209 );
xor ( n36211 , n36020 , n36022 );
xor ( n36212 , n36211 , n36025 );
and ( n36213 , n36209 , n36212 );
and ( n36214 , n36207 , n36212 );
or ( n36215 , n36210 , n36213 , n36214 );
and ( n36216 , n36153 , n36215 );
xor ( n36217 , n36010 , n36012 );
xor ( n36218 , n36217 , n36015 );
and ( n36219 , n36215 , n36218 );
and ( n36220 , n36153 , n36218 );
or ( n36221 , n36216 , n36219 , n36220 );
xor ( n36222 , n35873 , n35875 );
xor ( n36223 , n36222 , n35878 );
and ( n36224 , n36221 , n36223 );
xor ( n36225 , n36018 , n36036 );
xor ( n36226 , n36225 , n36039 );
and ( n36227 , n36223 , n36226 );
and ( n36228 , n36221 , n36226 );
or ( n36229 , n36224 , n36227 , n36228 );
and ( n36230 , n36054 , n36229 );
xor ( n36231 , n36054 , n36229 );
and ( n36232 , n21218 , n29276 );
and ( n36233 , n21072 , n29274 );
nor ( n36234 , n36232 , n36233 );
xnor ( n36235 , n36234 , n28677 );
and ( n36236 , n21451 , n28628 );
and ( n36237 , n21302 , n28626 );
nor ( n36238 , n36236 , n36237 );
xnor ( n36239 , n36238 , n28096 );
and ( n36240 , n36235 , n36239 );
xor ( n36241 , n35903 , n35907 );
xor ( n36242 , n36241 , n35912 );
and ( n36243 , n36239 , n36242 );
and ( n36244 , n36235 , n36242 );
or ( n36245 , n36240 , n36243 , n36244 );
and ( n36246 , n22425 , n26992 );
and ( n36247 , n22198 , n26990 );
nor ( n36248 , n36246 , n36247 );
xnor ( n36249 , n36248 , n26369 );
and ( n36250 , n23271 , n26027 );
and ( n36251 , n23141 , n26025 );
nor ( n36252 , n36250 , n36251 );
xnor ( n36253 , n36252 , n25499 );
and ( n36254 , n36249 , n36253 );
and ( n36255 , n36253 , n35983 );
and ( n36256 , n36249 , n35983 );
or ( n36257 , n36254 , n36255 , n36256 );
and ( n36258 , n21704 , n28062 );
and ( n36259 , n21612 , n28060 );
nor ( n36260 , n36258 , n36259 );
xnor ( n36261 , n36260 , n27549 );
and ( n36262 , n36257 , n36261 );
xor ( n36263 , n35965 , n35981 );
xor ( n36264 , n36263 , n35985 );
and ( n36265 , n36261 , n36264 );
and ( n36266 , n36257 , n36264 );
or ( n36267 , n36262 , n36265 , n36266 );
and ( n36268 , n36245 , n36267 );
and ( n36269 , n28211 , n21741 );
and ( n36270 , n27757 , n21739 );
nor ( n36271 , n36269 , n36270 );
xnor ( n36272 , n36271 , n21605 );
and ( n36273 , n28700 , n21468 );
and ( n36274 , n28810 , n21466 );
nor ( n36275 , n36273 , n36274 );
xnor ( n36276 , n36275 , n21331 );
and ( n36277 , n36272 , n36276 );
and ( n36278 , n29318 , n21155 );
and ( n36279 , n29078 , n21153 );
nor ( n36280 , n36278 , n36279 );
xnor ( n36281 , n36280 , n20994 );
and ( n36282 , n36276 , n36281 );
and ( n36283 , n36272 , n36281 );
or ( n36284 , n36277 , n36282 , n36283 );
and ( n36285 , n25284 , n23944 );
and ( n36286 , n24940 , n23942 );
nor ( n36287 , n36285 , n36286 );
xnor ( n36288 , n36287 , n23550 );
and ( n36289 , n26851 , n22859 );
and ( n36290 , n26422 , n22857 );
nor ( n36291 , n36289 , n36290 );
xnor ( n36292 , n36291 , n22418 );
and ( n36293 , n36288 , n36292 );
and ( n36294 , n27352 , n22381 );
and ( n36295 , n27135 , n22379 );
nor ( n36296 , n36294 , n36295 );
xnor ( n36297 , n36296 , n22228 );
and ( n36298 , n36292 , n36297 );
and ( n36299 , n36288 , n36297 );
or ( n36300 , n36293 , n36298 , n36299 );
and ( n36301 , n27751 , n22048 );
and ( n36302 , n27352 , n22046 );
nor ( n36303 , n36301 , n36302 );
xnor ( n36304 , n36303 , n21853 );
and ( n36305 , n36300 , n36304 );
xor ( n36306 , n35969 , n35973 );
xor ( n36307 , n36306 , n35978 );
and ( n36308 , n36304 , n36307 );
and ( n36309 , n36300 , n36307 );
or ( n36310 , n36305 , n36308 , n36309 );
and ( n36311 , n36284 , n36310 );
xor ( n36312 , n36101 , n36105 );
xor ( n36313 , n36312 , n36108 );
and ( n36314 , n36310 , n36313 );
and ( n36315 , n36284 , n36313 );
or ( n36316 , n36311 , n36314 , n36315 );
and ( n36317 , n36267 , n36316 );
and ( n36318 , n36245 , n36316 );
or ( n36319 , n36268 , n36317 , n36318 );
xor ( n36320 , n35937 , n35941 );
xor ( n36321 , n36320 , n35946 );
xor ( n36322 , n35988 , n35992 );
xor ( n36323 , n36322 , n35995 );
and ( n36324 , n36321 , n36323 );
xor ( n36325 , n36097 , n36111 );
xor ( n36326 , n36325 , n36114 );
and ( n36327 , n36323 , n36326 );
and ( n36328 , n36321 , n36326 );
or ( n36329 , n36324 , n36327 , n36328 );
and ( n36330 , n36319 , n36329 );
xor ( n36331 , n36056 , n36058 );
xor ( n36332 , n36331 , n36061 );
and ( n36333 , n36329 , n36332 );
and ( n36334 , n36319 , n36332 );
or ( n36335 , n36330 , n36333 , n36334 );
and ( n36336 , n24527 , n24902 );
and ( n36337 , n24521 , n24900 );
nor ( n36338 , n36336 , n36337 );
xnor ( n36339 , n36338 , n24397 );
and ( n36340 , n25554 , n23944 );
and ( n36341 , n25284 , n23942 );
nor ( n36342 , n36340 , n36341 );
xnor ( n36343 , n36342 , n23550 );
and ( n36344 , n36339 , n36343 );
and ( n36345 , n26422 , n23230 );
and ( n36346 , n26319 , n23228 );
nor ( n36347 , n36345 , n36346 );
xnor ( n36348 , n36347 , n22842 );
and ( n36349 , n36343 , n36348 );
and ( n36350 , n36339 , n36348 );
or ( n36351 , n36344 , n36349 , n36350 );
and ( n36352 , n24131 , n25383 );
and ( n36353 , n23968 , n25381 );
nor ( n36354 , n36352 , n36353 );
xnor ( n36355 , n36354 , n24885 );
and ( n36356 , n24940 , n24376 );
and ( n36357 , n24621 , n24374 );
nor ( n36358 , n36356 , n36357 );
xnor ( n36359 , n36358 , n23927 );
and ( n36360 , n36355 , n36359 );
and ( n36361 , n25974 , n23641 );
and ( n36362 , n25765 , n23639 );
nor ( n36363 , n36361 , n36362 );
xnor ( n36364 , n36363 , n23213 );
and ( n36365 , n36359 , n36364 );
and ( n36366 , n36355 , n36364 );
or ( n36367 , n36360 , n36365 , n36366 );
and ( n36368 , n36351 , n36367 );
and ( n36369 , n22756 , n26992 );
and ( n36370 , n22425 , n26990 );
nor ( n36371 , n36369 , n36370 );
xnor ( n36372 , n36371 , n26369 );
and ( n36373 , n36367 , n36372 );
and ( n36374 , n36351 , n36372 );
or ( n36375 , n36368 , n36373 , n36374 );
xor ( n36376 , n36068 , n36072 );
and ( n36377 , n23381 , n26027 );
and ( n36378 , n23271 , n26025 );
nor ( n36379 , n36377 , n36378 );
xnor ( n36380 , n36379 , n25499 );
and ( n36381 , n36376 , n36380 );
and ( n36382 , n29623 , n21153 );
not ( n36383 , n36382 );
and ( n36384 , n36383 , n20994 );
and ( n36385 , n36380 , n36384 );
and ( n36386 , n36376 , n36384 );
or ( n36387 , n36381 , n36385 , n36386 );
and ( n36388 , n36375 , n36387 );
xor ( n36389 , n36073 , n36077 );
xor ( n36390 , n36389 , n36082 );
and ( n36391 , n36387 , n36390 );
and ( n36392 , n36375 , n36390 );
or ( n36393 , n36388 , n36391 , n36392 );
xor ( n36394 , n36085 , n36089 );
xor ( n36395 , n36394 , n36094 );
and ( n36396 , n36393 , n36395 );
xor ( n36397 , n36121 , n36125 );
xor ( n36398 , n36397 , n36128 );
and ( n36399 , n36395 , n36398 );
and ( n36400 , n36393 , n36398 );
or ( n36401 , n36396 , n36399 , n36400 );
xor ( n36402 , n36245 , n36267 );
xor ( n36403 , n36402 , n36316 );
and ( n36404 , n36401 , n36403 );
xor ( n36405 , n36131 , n36135 );
xor ( n36406 , n36405 , n36138 );
and ( n36407 , n36403 , n36406 );
and ( n36408 , n36401 , n36406 );
or ( n36409 , n36404 , n36407 , n36408 );
and ( n36410 , n21302 , n29276 );
and ( n36411 , n21218 , n29274 );
nor ( n36412 , n36410 , n36411 );
xnor ( n36413 , n36412 , n28677 );
and ( n36414 , n21876 , n28062 );
and ( n36415 , n21704 , n28060 );
nor ( n36416 , n36414 , n36415 );
xnor ( n36417 , n36416 , n27549 );
and ( n36418 , n36413 , n36417 );
and ( n36419 , n22235 , n27529 );
and ( n36420 , n21955 , n27527 );
nor ( n36421 , n36419 , n36420 );
xnor ( n36422 , n36421 , n27034 );
and ( n36423 , n36417 , n36422 );
and ( n36424 , n36413 , n36422 );
or ( n36425 , n36418 , n36423 , n36424 );
and ( n36426 , n21072 , n29977 );
and ( n36427 , n20867 , n29974 );
nor ( n36428 , n36426 , n36427 );
xnor ( n36429 , n36428 , n28674 );
and ( n36430 , n21612 , n28628 );
and ( n36431 , n21451 , n28626 );
nor ( n36432 , n36430 , n36431 );
xnor ( n36433 , n36432 , n28096 );
and ( n36434 , n36429 , n36433 );
xor ( n36435 , n36249 , n36253 );
xor ( n36436 , n36435 , n35983 );
and ( n36437 , n36433 , n36436 );
and ( n36438 , n36429 , n36436 );
or ( n36439 , n36434 , n36437 , n36438 );
and ( n36440 , n36425 , n36439 );
xor ( n36441 , n36257 , n36261 );
xor ( n36442 , n36441 , n36264 );
and ( n36443 , n36439 , n36442 );
and ( n36444 , n36425 , n36442 );
or ( n36445 , n36440 , n36443 , n36444 );
and ( n36446 , n23141 , n26349 );
and ( n36447 , n22916 , n26347 );
nor ( n36448 , n36446 , n36447 );
xnor ( n36449 , n36448 , n25893 );
xor ( n36450 , n36157 , n36161 );
xor ( n36451 , n36450 , n36166 );
and ( n36452 , n36449 , n36451 );
xor ( n36453 , n36288 , n36292 );
xor ( n36454 , n36453 , n36297 );
and ( n36455 , n36451 , n36454 );
and ( n36456 , n36449 , n36454 );
or ( n36457 , n36452 , n36455 , n36456 );
xor ( n36458 , n36169 , n36173 );
xor ( n36459 , n36458 , n36176 );
and ( n36460 , n36457 , n36459 );
xor ( n36461 , n36300 , n36304 );
xor ( n36462 , n36461 , n36307 );
and ( n36463 , n36459 , n36462 );
and ( n36464 , n36457 , n36462 );
or ( n36465 , n36460 , n36463 , n36464 );
xor ( n36466 , n36179 , n36183 );
xor ( n36467 , n36466 , n36188 );
and ( n36468 , n36465 , n36467 );
xor ( n36469 , n36235 , n36239 );
xor ( n36470 , n36469 , n36242 );
and ( n36471 , n36467 , n36470 );
and ( n36472 , n36465 , n36470 );
or ( n36473 , n36468 , n36471 , n36472 );
and ( n36474 , n36445 , n36473 );
xor ( n36475 , n36191 , n36193 );
xor ( n36476 , n36475 , n36196 );
and ( n36477 , n36473 , n36476 );
and ( n36478 , n36445 , n36476 );
or ( n36479 , n36474 , n36477 , n36478 );
and ( n36480 , n36409 , n36479 );
xor ( n36481 , n36117 , n36141 );
xor ( n36482 , n36481 , n36144 );
and ( n36483 , n36479 , n36482 );
and ( n36484 , n36409 , n36482 );
or ( n36485 , n36480 , n36483 , n36484 );
and ( n36486 , n36335 , n36485 );
xor ( n36487 , n36064 , n36147 );
xor ( n36488 , n36487 , n36150 );
and ( n36489 , n36485 , n36488 );
and ( n36490 , n36335 , n36488 );
or ( n36491 , n36486 , n36489 , n36490 );
xor ( n36492 , n36028 , n36030 );
xor ( n36493 , n36492 , n36033 );
and ( n36494 , n36491 , n36493 );
xor ( n36495 , n36153 , n36215 );
xor ( n36496 , n36495 , n36218 );
and ( n36497 , n36493 , n36496 );
and ( n36498 , n36491 , n36496 );
or ( n36499 , n36494 , n36497 , n36498 );
xor ( n36500 , n36221 , n36223 );
xor ( n36501 , n36500 , n36226 );
and ( n36502 , n36499 , n36501 );
xor ( n36503 , n36499 , n36501 );
xor ( n36504 , n36491 , n36493 );
xor ( n36505 , n36504 , n36496 );
and ( n36506 , n28810 , n21741 );
and ( n36507 , n28211 , n21739 );
nor ( n36508 , n36506 , n36507 );
xnor ( n36509 , n36508 , n21605 );
and ( n36510 , n29078 , n21468 );
and ( n36511 , n28700 , n21466 );
nor ( n36512 , n36510 , n36511 );
xnor ( n36513 , n36512 , n21331 );
and ( n36514 , n36509 , n36513 );
and ( n36515 , n29623 , n21155 );
and ( n36516 , n29318 , n21153 );
nor ( n36517 , n36515 , n36516 );
xnor ( n36518 , n36517 , n20994 );
and ( n36519 , n36513 , n36518 );
and ( n36520 , n36509 , n36518 );
or ( n36521 , n36514 , n36519 , n36520 );
and ( n36522 , n25765 , n23944 );
and ( n36523 , n25554 , n23942 );
nor ( n36524 , n36522 , n36523 );
xnor ( n36525 , n36524 , n23550 );
and ( n36526 , n26851 , n23230 );
and ( n36527 , n26422 , n23228 );
nor ( n36528 , n36526 , n36527 );
xnor ( n36529 , n36528 , n22842 );
and ( n36530 , n36525 , n36529 );
and ( n36531 , n27135 , n22859 );
and ( n36532 , n26851 , n22857 );
nor ( n36533 , n36531 , n36532 );
xnor ( n36534 , n36533 , n22418 );
and ( n36535 , n36530 , n36534 );
and ( n36536 , n27751 , n22381 );
and ( n36537 , n27352 , n22379 );
nor ( n36538 , n36536 , n36537 );
xnor ( n36539 , n36538 , n22228 );
and ( n36540 , n36534 , n36539 );
and ( n36541 , n36530 , n36539 );
or ( n36542 , n36535 , n36540 , n36541 );
and ( n36543 , n22198 , n27529 );
and ( n36544 , n22235 , n27527 );
nor ( n36545 , n36543 , n36544 );
xnor ( n36546 , n36545 , n27034 );
and ( n36547 , n36542 , n36546 );
and ( n36548 , n27757 , n22048 );
and ( n36549 , n27751 , n22046 );
nor ( n36550 , n36548 , n36549 );
xnor ( n36551 , n36550 , n21853 );
and ( n36552 , n36546 , n36551 );
and ( n36553 , n36542 , n36551 );
or ( n36554 , n36547 , n36552 , n36553 );
and ( n36555 , n36521 , n36554 );
xor ( n36556 , n36272 , n36276 );
xor ( n36557 , n36556 , n36281 );
and ( n36558 , n36554 , n36557 );
and ( n36559 , n36521 , n36557 );
or ( n36560 , n36555 , n36558 , n36559 );
xor ( n36561 , n36284 , n36310 );
xor ( n36562 , n36561 , n36313 );
and ( n36563 , n36560 , n36562 );
xor ( n36564 , n36393 , n36395 );
xor ( n36565 , n36564 , n36398 );
and ( n36566 , n36562 , n36565 );
and ( n36567 , n36560 , n36565 );
or ( n36568 , n36563 , n36566 , n36567 );
and ( n36569 , n21218 , n29977 );
and ( n36570 , n21072 , n29974 );
nor ( n36571 , n36569 , n36570 );
xnor ( n36572 , n36571 , n28674 );
and ( n36573 , n21704 , n28628 );
and ( n36574 , n21612 , n28626 );
nor ( n36575 , n36573 , n36574 );
xnor ( n36576 , n36575 , n28096 );
and ( n36577 , n36572 , n36576 );
xor ( n36578 , n36351 , n36367 );
xor ( n36579 , n36578 , n36372 );
and ( n36580 , n36576 , n36579 );
and ( n36581 , n36572 , n36579 );
or ( n36582 , n36577 , n36580 , n36581 );
and ( n36583 , n21451 , n29276 );
and ( n36584 , n21302 , n29274 );
nor ( n36585 , n36583 , n36584 );
xnor ( n36586 , n36585 , n28677 );
and ( n36587 , n21955 , n28062 );
and ( n36588 , n21876 , n28060 );
nor ( n36589 , n36587 , n36588 );
xnor ( n36590 , n36589 , n27549 );
and ( n36591 , n36586 , n36590 );
xor ( n36592 , n36376 , n36380 );
xor ( n36593 , n36592 , n36384 );
and ( n36594 , n36590 , n36593 );
and ( n36595 , n36586 , n36593 );
or ( n36596 , n36591 , n36594 , n36595 );
and ( n36597 , n36582 , n36596 );
xor ( n36598 , n36375 , n36387 );
xor ( n36599 , n36598 , n36390 );
and ( n36600 , n36596 , n36599 );
and ( n36601 , n36582 , n36599 );
or ( n36602 , n36597 , n36600 , n36601 );
and ( n36603 , n24521 , n25383 );
and ( n36604 , n24131 , n25381 );
nor ( n36605 , n36603 , n36604 );
xnor ( n36606 , n36605 , n24885 );
and ( n36607 , n24621 , n24902 );
and ( n36608 , n24527 , n24900 );
nor ( n36609 , n36607 , n36608 );
xnor ( n36610 , n36609 , n24397 );
and ( n36611 , n36606 , n36610 );
and ( n36612 , n25284 , n24376 );
and ( n36613 , n24940 , n24374 );
nor ( n36614 , n36612 , n36613 );
xnor ( n36615 , n36614 , n23927 );
and ( n36616 , n36610 , n36615 );
and ( n36617 , n36606 , n36615 );
or ( n36618 , n36611 , n36616 , n36617 );
and ( n36619 , n23968 , n26027 );
and ( n36620 , n23573 , n26025 );
nor ( n36621 , n36619 , n36620 );
xnor ( n36622 , n36621 , n25499 );
and ( n36623 , n26319 , n23641 );
and ( n36624 , n25974 , n23639 );
nor ( n36625 , n36623 , n36624 );
xnor ( n36626 , n36625 , n23213 );
and ( n36627 , n36622 , n36626 );
and ( n36628 , n27352 , n22859 );
and ( n36629 , n27135 , n22857 );
nor ( n36630 , n36628 , n36629 );
xnor ( n36631 , n36630 , n22418 );
and ( n36632 , n36626 , n36631 );
and ( n36633 , n36622 , n36631 );
or ( n36634 , n36627 , n36632 , n36633 );
and ( n36635 , n36618 , n36634 );
and ( n36636 , n36634 , n36382 );
and ( n36637 , n36618 , n36382 );
or ( n36638 , n36635 , n36636 , n36637 );
and ( n36639 , n22916 , n26992 );
and ( n36640 , n22756 , n26990 );
nor ( n36641 , n36639 , n36640 );
xnor ( n36642 , n36641 , n26369 );
and ( n36643 , n23271 , n26349 );
and ( n36644 , n23141 , n26347 );
nor ( n36645 , n36643 , n36644 );
xnor ( n36646 , n36645 , n25893 );
and ( n36647 , n36642 , n36646 );
xor ( n36648 , n36355 , n36359 );
xor ( n36649 , n36648 , n36364 );
and ( n36650 , n36646 , n36649 );
and ( n36651 , n36642 , n36649 );
or ( n36652 , n36647 , n36650 , n36651 );
and ( n36653 , n36638 , n36652 );
and ( n36654 , n22425 , n27529 );
and ( n36655 , n22198 , n27527 );
nor ( n36656 , n36654 , n36655 );
xnor ( n36657 , n36656 , n27034 );
and ( n36658 , n23573 , n26027 );
and ( n36659 , n23381 , n26025 );
nor ( n36660 , n36658 , n36659 );
xnor ( n36661 , n36660 , n25499 );
and ( n36662 , n36657 , n36661 );
xor ( n36663 , n36339 , n36343 );
xor ( n36664 , n36663 , n36348 );
and ( n36665 , n36661 , n36664 );
and ( n36666 , n36657 , n36664 );
or ( n36667 , n36662 , n36665 , n36666 );
and ( n36668 , n36652 , n36667 );
and ( n36669 , n36638 , n36667 );
or ( n36670 , n36653 , n36668 , n36669 );
xor ( n36671 , n36413 , n36417 );
xor ( n36672 , n36671 , n36422 );
and ( n36673 , n36670 , n36672 );
xor ( n36674 , n36457 , n36459 );
xor ( n36675 , n36674 , n36462 );
and ( n36676 , n36672 , n36675 );
and ( n36677 , n36670 , n36675 );
or ( n36678 , n36673 , n36676 , n36677 );
and ( n36679 , n36602 , n36678 );
xor ( n36680 , n36425 , n36439 );
xor ( n36681 , n36680 , n36442 );
and ( n36682 , n36678 , n36681 );
and ( n36683 , n36602 , n36681 );
or ( n36684 , n36679 , n36682 , n36683 );
and ( n36685 , n36568 , n36684 );
xor ( n36686 , n36321 , n36323 );
xor ( n36687 , n36686 , n36326 );
and ( n36688 , n36684 , n36687 );
and ( n36689 , n36568 , n36687 );
or ( n36690 , n36685 , n36688 , n36689 );
xor ( n36691 , n36199 , n36201 );
xor ( n36692 , n36691 , n36204 );
and ( n36693 , n36690 , n36692 );
xor ( n36694 , n36319 , n36329 );
xor ( n36695 , n36694 , n36332 );
and ( n36696 , n36692 , n36695 );
and ( n36697 , n36690 , n36695 );
or ( n36698 , n36693 , n36696 , n36697 );
xor ( n36699 , n36335 , n36485 );
xor ( n36700 , n36699 , n36488 );
and ( n36701 , n36698 , n36700 );
xor ( n36702 , n36207 , n36209 );
xor ( n36703 , n36702 , n36212 );
and ( n36704 , n36700 , n36703 );
and ( n36705 , n36698 , n36703 );
or ( n36706 , n36701 , n36704 , n36705 );
and ( n36707 , n36505 , n36706 );
xor ( n36708 , n36505 , n36706 );
xor ( n36709 , n36698 , n36700 );
xor ( n36710 , n36709 , n36703 );
and ( n36711 , n28211 , n22048 );
and ( n36712 , n27757 , n22046 );
nor ( n36713 , n36711 , n36712 );
xnor ( n36714 , n36713 , n21853 );
and ( n36715 , n28700 , n21741 );
and ( n36716 , n28810 , n21739 );
nor ( n36717 , n36715 , n36716 );
xnor ( n36718 , n36717 , n21605 );
and ( n36719 , n36714 , n36718 );
xor ( n36720 , n36530 , n36534 );
xor ( n36721 , n36720 , n36539 );
and ( n36722 , n36718 , n36721 );
and ( n36723 , n36714 , n36721 );
or ( n36724 , n36719 , n36722 , n36723 );
xor ( n36725 , n36542 , n36546 );
xor ( n36726 , n36725 , n36551 );
and ( n36727 , n36724 , n36726 );
xor ( n36728 , n36449 , n36451 );
xor ( n36729 , n36728 , n36454 );
and ( n36730 , n36726 , n36729 );
and ( n36731 , n36724 , n36729 );
or ( n36732 , n36727 , n36730 , n36731 );
xor ( n36733 , n36429 , n36433 );
xor ( n36734 , n36733 , n36436 );
and ( n36735 , n36732 , n36734 );
xor ( n36736 , n36521 , n36554 );
xor ( n36737 , n36736 , n36557 );
and ( n36738 , n36734 , n36737 );
and ( n36739 , n36732 , n36737 );
or ( n36740 , n36735 , n36738 , n36739 );
xor ( n36741 , n36465 , n36467 );
xor ( n36742 , n36741 , n36470 );
and ( n36743 , n36740 , n36742 );
xor ( n36744 , n36560 , n36562 );
xor ( n36745 , n36744 , n36565 );
and ( n36746 , n36742 , n36745 );
and ( n36747 , n36740 , n36745 );
or ( n36748 , n36743 , n36746 , n36747 );
xor ( n36749 , n36401 , n36403 );
xor ( n36750 , n36749 , n36406 );
and ( n36751 , n36748 , n36750 );
xor ( n36752 , n36445 , n36473 );
xor ( n36753 , n36752 , n36476 );
and ( n36754 , n36750 , n36753 );
and ( n36755 , n36748 , n36753 );
or ( n36756 , n36751 , n36754 , n36755 );
xor ( n36757 , n36409 , n36479 );
xor ( n36758 , n36757 , n36482 );
and ( n36759 , n36756 , n36758 );
xor ( n36760 , n36690 , n36692 );
xor ( n36761 , n36760 , n36695 );
and ( n36762 , n36758 , n36761 );
and ( n36763 , n36756 , n36761 );
or ( n36764 , n36759 , n36762 , n36763 );
and ( n36765 , n36710 , n36764 );
xor ( n36766 , n36710 , n36764 );
xor ( n36767 , n36756 , n36758 );
xor ( n36768 , n36767 , n36761 );
and ( n36769 , n21302 , n29977 );
and ( n36770 , n21218 , n29974 );
nor ( n36771 , n36769 , n36770 );
xnor ( n36772 , n36771 , n28674 );
and ( n36773 , n21876 , n28628 );
and ( n36774 , n21704 , n28626 );
nor ( n36775 , n36773 , n36774 );
xnor ( n36776 , n36775 , n28096 );
and ( n36777 , n36772 , n36776 );
xor ( n36778 , n36618 , n36634 );
xor ( n36779 , n36778 , n36382 );
and ( n36780 , n36776 , n36779 );
and ( n36781 , n36772 , n36779 );
or ( n36782 , n36777 , n36780 , n36781 );
and ( n36783 , n21612 , n29276 );
and ( n36784 , n21451 , n29274 );
nor ( n36785 , n36783 , n36784 );
xnor ( n36786 , n36785 , n28677 );
xor ( n36787 , n36642 , n36646 );
xor ( n36788 , n36787 , n36649 );
and ( n36789 , n36786 , n36788 );
xor ( n36790 , n36657 , n36661 );
xor ( n36791 , n36790 , n36664 );
and ( n36792 , n36788 , n36791 );
and ( n36793 , n36786 , n36791 );
or ( n36794 , n36789 , n36792 , n36793 );
and ( n36795 , n36782 , n36794 );
xor ( n36796 , n36638 , n36652 );
xor ( n36797 , n36796 , n36667 );
and ( n36798 , n36794 , n36797 );
and ( n36799 , n36782 , n36797 );
or ( n36800 , n36795 , n36798 , n36799 );
and ( n36801 , n24940 , n24902 );
and ( n36802 , n24621 , n24900 );
nor ( n36803 , n36801 , n36802 );
xnor ( n36804 , n36803 , n24397 );
and ( n36805 , n26422 , n23641 );
and ( n36806 , n26319 , n23639 );
nor ( n36807 , n36805 , n36806 );
xnor ( n36808 , n36807 , n23213 );
and ( n36809 , n36804 , n36808 );
and ( n36810 , n27751 , n22859 );
and ( n36811 , n27352 , n22857 );
nor ( n36812 , n36810 , n36811 );
xnor ( n36813 , n36812 , n22418 );
and ( n36814 , n36808 , n36813 );
and ( n36815 , n36804 , n36813 );
or ( n36816 , n36809 , n36814 , n36815 );
and ( n36817 , n23141 , n26992 );
and ( n36818 , n22916 , n26990 );
nor ( n36819 , n36817 , n36818 );
xnor ( n36820 , n36819 , n26369 );
and ( n36821 , n36816 , n36820 );
and ( n36822 , n23381 , n26349 );
and ( n36823 , n23271 , n26347 );
nor ( n36824 , n36822 , n36823 );
xnor ( n36825 , n36824 , n25893 );
and ( n36826 , n36820 , n36825 );
and ( n36827 , n36816 , n36825 );
or ( n36828 , n36821 , n36826 , n36827 );
and ( n36829 , n22198 , n28062 );
and ( n36830 , n22235 , n28060 );
nor ( n36831 , n36829 , n36830 );
xnor ( n36832 , n36831 , n27549 );
xor ( n36833 , n36606 , n36610 );
xor ( n36834 , n36833 , n36615 );
and ( n36835 , n36832 , n36834 );
xor ( n36836 , n36622 , n36626 );
xor ( n36837 , n36836 , n36631 );
and ( n36838 , n36834 , n36837 );
and ( n36839 , n36832 , n36837 );
or ( n36840 , n36835 , n36838 , n36839 );
and ( n36841 , n36828 , n36840 );
and ( n36842 , n22235 , n28062 );
and ( n36843 , n21955 , n28060 );
nor ( n36844 , n36842 , n36843 );
xnor ( n36845 , n36844 , n27549 );
and ( n36846 , n36840 , n36845 );
and ( n36847 , n36828 , n36845 );
or ( n36848 , n36841 , n36846 , n36847 );
and ( n36849 , n25765 , n24376 );
and ( n36850 , n25554 , n24374 );
nor ( n36851 , n36849 , n36850 );
xnor ( n36852 , n36851 , n23927 );
and ( n36853 , n26319 , n23944 );
and ( n36854 , n25974 , n23942 );
nor ( n36855 , n36853 , n36854 );
xnor ( n36856 , n36855 , n23550 );
and ( n36857 , n36852 , n36856 );
and ( n36858 , n24131 , n26027 );
and ( n36859 , n23968 , n26025 );
nor ( n36860 , n36858 , n36859 );
xnor ( n36861 , n36860 , n25499 );
and ( n36862 , n36857 , n36861 );
and ( n36863 , n24527 , n25383 );
and ( n36864 , n24521 , n25381 );
nor ( n36865 , n36863 , n36864 );
xnor ( n36866 , n36865 , n24885 );
and ( n36867 , n36861 , n36866 );
and ( n36868 , n36857 , n36866 );
or ( n36869 , n36862 , n36867 , n36868 );
and ( n36870 , n22756 , n27529 );
and ( n36871 , n22425 , n27527 );
nor ( n36872 , n36870 , n36871 );
xnor ( n36873 , n36872 , n27034 );
and ( n36874 , n36869 , n36873 );
and ( n36875 , n29623 , n21466 );
not ( n36876 , n36875 );
and ( n36877 , n36876 , n21331 );
and ( n36878 , n36873 , n36877 );
and ( n36879 , n36869 , n36877 );
or ( n36880 , n36874 , n36878 , n36879 );
xor ( n36881 , n36525 , n36529 );
and ( n36882 , n25554 , n24376 );
and ( n36883 , n25284 , n24374 );
nor ( n36884 , n36882 , n36883 );
xnor ( n36885 , n36884 , n23927 );
and ( n36886 , n25974 , n23944 );
and ( n36887 , n25765 , n23942 );
nor ( n36888 , n36886 , n36887 );
xnor ( n36889 , n36888 , n23550 );
and ( n36890 , n36885 , n36889 );
and ( n36891 , n27135 , n23230 );
and ( n36892 , n26851 , n23228 );
nor ( n36893 , n36891 , n36892 );
xnor ( n36894 , n36893 , n22842 );
and ( n36895 , n36889 , n36894 );
and ( n36896 , n36885 , n36894 );
or ( n36897 , n36890 , n36895 , n36896 );
and ( n36898 , n36881 , n36897 );
and ( n36899 , n27757 , n22381 );
and ( n36900 , n27751 , n22379 );
nor ( n36901 , n36899 , n36900 );
xnor ( n36902 , n36901 , n22228 );
and ( n36903 , n36897 , n36902 );
and ( n36904 , n36881 , n36902 );
or ( n36905 , n36898 , n36903 , n36904 );
and ( n36906 , n36880 , n36905 );
and ( n36907 , n29318 , n21468 );
and ( n36908 , n29078 , n21466 );
nor ( n36909 , n36907 , n36908 );
xnor ( n36910 , n36909 , n21331 );
and ( n36911 , n36905 , n36910 );
and ( n36912 , n36880 , n36910 );
or ( n36913 , n36906 , n36911 , n36912 );
and ( n36914 , n36848 , n36913 );
xor ( n36915 , n36509 , n36513 );
xor ( n36916 , n36915 , n36518 );
and ( n36917 , n36913 , n36916 );
and ( n36918 , n36848 , n36916 );
or ( n36919 , n36914 , n36917 , n36918 );
and ( n36920 , n36800 , n36919 );
xor ( n36921 , n36582 , n36596 );
xor ( n36922 , n36921 , n36599 );
and ( n36923 , n36919 , n36922 );
and ( n36924 , n36800 , n36922 );
or ( n36925 , n36920 , n36923 , n36924 );
and ( n36926 , n28810 , n22048 );
and ( n36927 , n28211 , n22046 );
nor ( n36928 , n36926 , n36927 );
xnor ( n36929 , n36928 , n21853 );
and ( n36930 , n29078 , n21741 );
and ( n36931 , n28700 , n21739 );
nor ( n36932 , n36930 , n36931 );
xnor ( n36933 , n36932 , n21605 );
and ( n36934 , n36929 , n36933 );
and ( n36935 , n29623 , n21468 );
and ( n36936 , n29318 , n21466 );
nor ( n36937 , n36935 , n36936 );
xnor ( n36938 , n36937 , n21331 );
and ( n36939 , n36933 , n36938 );
and ( n36940 , n36929 , n36938 );
or ( n36941 , n36934 , n36939 , n36940 );
and ( n36942 , n23968 , n26349 );
and ( n36943 , n23573 , n26347 );
nor ( n36944 , n36942 , n36943 );
xnor ( n36945 , n36944 , n25893 );
and ( n36946 , n24621 , n25383 );
and ( n36947 , n24527 , n25381 );
nor ( n36948 , n36946 , n36947 );
xnor ( n36949 , n36948 , n24885 );
and ( n36950 , n36945 , n36949 );
and ( n36951 , n27352 , n23230 );
and ( n36952 , n27135 , n23228 );
nor ( n36953 , n36951 , n36952 );
xnor ( n36954 , n36953 , n22842 );
and ( n36955 , n36949 , n36954 );
and ( n36956 , n36945 , n36954 );
or ( n36957 , n36950 , n36955 , n36956 );
and ( n36958 , n22916 , n27529 );
and ( n36959 , n22756 , n27527 );
nor ( n36960 , n36958 , n36959 );
xnor ( n36961 , n36960 , n27034 );
and ( n36962 , n36957 , n36961 );
and ( n36963 , n36961 , n36875 );
and ( n36964 , n36957 , n36875 );
or ( n36965 , n36962 , n36963 , n36964 );
and ( n36966 , n23573 , n26349 );
and ( n36967 , n23381 , n26347 );
nor ( n36968 , n36966 , n36967 );
xnor ( n36969 , n36968 , n25893 );
and ( n36970 , n28211 , n22381 );
and ( n36971 , n27757 , n22379 );
nor ( n36972 , n36970 , n36971 );
xnor ( n36973 , n36972 , n22228 );
and ( n36974 , n36969 , n36973 );
xor ( n36975 , n36885 , n36889 );
xor ( n36976 , n36975 , n36894 );
and ( n36977 , n36973 , n36976 );
and ( n36978 , n36969 , n36976 );
or ( n36979 , n36974 , n36977 , n36978 );
and ( n36980 , n36965 , n36979 );
xor ( n36981 , n36881 , n36897 );
xor ( n36982 , n36981 , n36902 );
and ( n36983 , n36979 , n36982 );
and ( n36984 , n36965 , n36982 );
or ( n36985 , n36980 , n36983 , n36984 );
and ( n36986 , n36941 , n36985 );
xor ( n36987 , n36880 , n36905 );
xor ( n36988 , n36987 , n36910 );
and ( n36989 , n36985 , n36988 );
and ( n36990 , n36941 , n36988 );
or ( n36991 , n36986 , n36989 , n36990 );
xor ( n36992 , n36572 , n36576 );
xor ( n36993 , n36992 , n36579 );
and ( n36994 , n36991 , n36993 );
xor ( n36995 , n36586 , n36590 );
xor ( n36996 , n36995 , n36593 );
and ( n36997 , n36993 , n36996 );
and ( n36998 , n36991 , n36996 );
or ( n36999 , n36994 , n36997 , n36998 );
xor ( n37000 , n36732 , n36734 );
xor ( n37001 , n37000 , n36737 );
and ( n37002 , n36999 , n37001 );
xor ( n37003 , n36670 , n36672 );
xor ( n37004 , n37003 , n36675 );
and ( n37005 , n37001 , n37004 );
and ( n37006 , n36999 , n37004 );
or ( n37007 , n37002 , n37005 , n37006 );
and ( n37008 , n36925 , n37007 );
xor ( n37009 , n36602 , n36678 );
xor ( n37010 , n37009 , n36681 );
and ( n37011 , n37007 , n37010 );
and ( n37012 , n36925 , n37010 );
or ( n37013 , n37008 , n37011 , n37012 );
xor ( n37014 , n36568 , n36684 );
xor ( n37015 , n37014 , n36687 );
and ( n37016 , n37013 , n37015 );
xor ( n37017 , n36748 , n36750 );
xor ( n37018 , n37017 , n36753 );
and ( n37019 , n37015 , n37018 );
and ( n37020 , n37013 , n37018 );
or ( n37021 , n37016 , n37019 , n37020 );
and ( n37022 , n36768 , n37021 );
xor ( n37023 , n36768 , n37021 );
xor ( n37024 , n37013 , n37015 );
xor ( n37025 , n37024 , n37018 );
and ( n37026 , n21451 , n29977 );
and ( n37027 , n21302 , n29974 );
nor ( n37028 , n37026 , n37027 );
xnor ( n37029 , n37028 , n28674 );
and ( n37030 , n21704 , n29276 );
and ( n37031 , n21612 , n29274 );
nor ( n37032 , n37030 , n37031 );
xnor ( n37033 , n37032 , n28677 );
and ( n37034 , n37029 , n37033 );
xor ( n37035 , n36869 , n36873 );
xor ( n37036 , n37035 , n36877 );
and ( n37037 , n37033 , n37036 );
and ( n37038 , n37029 , n37036 );
or ( n37039 , n37034 , n37037 , n37038 );
xor ( n37040 , n36828 , n36840 );
xor ( n37041 , n37040 , n36845 );
and ( n37042 , n37039 , n37041 );
xor ( n37043 , n36714 , n36718 );
xor ( n37044 , n37043 , n36721 );
and ( n37045 , n37041 , n37044 );
and ( n37046 , n37039 , n37044 );
or ( n37047 , n37042 , n37045 , n37046 );
xor ( n37048 , n36848 , n36913 );
xor ( n37049 , n37048 , n36916 );
and ( n37050 , n37047 , n37049 );
xor ( n37051 , n36724 , n36726 );
xor ( n37052 , n37051 , n36729 );
and ( n37053 , n37049 , n37052 );
and ( n37054 , n37047 , n37052 );
or ( n37055 , n37050 , n37053 , n37054 );
xor ( n37056 , n36852 , n36856 );
and ( n37057 , n24521 , n26027 );
and ( n37058 , n24131 , n26025 );
nor ( n37059 , n37057 , n37058 );
xnor ( n37060 , n37059 , n25499 );
and ( n37061 , n37056 , n37060 );
and ( n37062 , n25284 , n24902 );
and ( n37063 , n24940 , n24900 );
nor ( n37064 , n37062 , n37063 );
xnor ( n37065 , n37064 , n24397 );
and ( n37066 , n37060 , n37065 );
and ( n37067 , n37056 , n37065 );
or ( n37068 , n37061 , n37066 , n37067 );
and ( n37069 , n22425 , n28062 );
and ( n37070 , n22198 , n28060 );
nor ( n37071 , n37069 , n37070 );
xnor ( n37072 , n37071 , n27549 );
and ( n37073 , n37068 , n37072 );
and ( n37074 , n23271 , n26992 );
and ( n37075 , n23141 , n26990 );
nor ( n37076 , n37074 , n37075 );
xnor ( n37077 , n37076 , n26369 );
and ( n37078 , n37072 , n37077 );
and ( n37079 , n37068 , n37077 );
or ( n37080 , n37073 , n37078 , n37079 );
and ( n37081 , n21955 , n28628 );
and ( n37082 , n21876 , n28626 );
nor ( n37083 , n37081 , n37082 );
xnor ( n37084 , n37083 , n28096 );
and ( n37085 , n37080 , n37084 );
xor ( n37086 , n36816 , n36820 );
xor ( n37087 , n37086 , n36825 );
and ( n37088 , n37084 , n37087 );
and ( n37089 , n37080 , n37087 );
or ( n37090 , n37085 , n37088 , n37089 );
xor ( n37091 , n36772 , n36776 );
xor ( n37092 , n37091 , n36779 );
and ( n37093 , n37090 , n37092 );
xor ( n37094 , n36786 , n36788 );
xor ( n37095 , n37094 , n36791 );
and ( n37096 , n37092 , n37095 );
and ( n37097 , n37090 , n37095 );
or ( n37098 , n37093 , n37096 , n37097 );
xor ( n37099 , n36782 , n36794 );
xor ( n37100 , n37099 , n36797 );
and ( n37101 , n37098 , n37100 );
xor ( n37102 , n36991 , n36993 );
xor ( n37103 , n37102 , n36996 );
and ( n37104 , n37100 , n37103 );
and ( n37105 , n37098 , n37103 );
or ( n37106 , n37101 , n37104 , n37105 );
and ( n37107 , n37055 , n37106 );
xor ( n37108 , n36800 , n36919 );
xor ( n37109 , n37108 , n36922 );
and ( n37110 , n37106 , n37109 );
and ( n37111 , n37055 , n37109 );
or ( n37112 , n37107 , n37110 , n37111 );
xor ( n37113 , n36740 , n36742 );
xor ( n37114 , n37113 , n36745 );
and ( n37115 , n37112 , n37114 );
xor ( n37116 , n36925 , n37007 );
xor ( n37117 , n37116 , n37010 );
and ( n37118 , n37114 , n37117 );
and ( n37119 , n37112 , n37117 );
or ( n37120 , n37115 , n37118 , n37119 );
and ( n37121 , n37025 , n37120 );
xor ( n37122 , n37025 , n37120 );
xor ( n37123 , n37112 , n37114 );
xor ( n37124 , n37123 , n37117 );
and ( n37125 , n22235 , n28628 );
and ( n37126 , n21955 , n28626 );
nor ( n37127 , n37125 , n37126 );
xnor ( n37128 , n37127 , n28096 );
and ( n37129 , n28700 , n22048 );
and ( n37130 , n28810 , n22046 );
nor ( n37131 , n37129 , n37130 );
xnor ( n37132 , n37131 , n21853 );
and ( n37133 , n37128 , n37132 );
and ( n37134 , n29318 , n21741 );
and ( n37135 , n29078 , n21739 );
nor ( n37136 , n37134 , n37135 );
xnor ( n37137 , n37136 , n21605 );
and ( n37138 , n37132 , n37137 );
and ( n37139 , n37128 , n37137 );
or ( n37140 , n37133 , n37138 , n37139 );
and ( n37141 , n26851 , n23641 );
and ( n37142 , n26422 , n23639 );
nor ( n37143 , n37141 , n37142 );
xnor ( n37144 , n37143 , n23213 );
and ( n37145 , n27757 , n22859 );
and ( n37146 , n27751 , n22857 );
nor ( n37147 , n37145 , n37146 );
xnor ( n37148 , n37147 , n22418 );
and ( n37149 , n37144 , n37148 );
and ( n37150 , n28810 , n22381 );
and ( n37151 , n28211 , n22379 );
nor ( n37152 , n37150 , n37151 );
xnor ( n37153 , n37152 , n22228 );
and ( n37154 , n37148 , n37153 );
and ( n37155 , n37144 , n37153 );
or ( n37156 , n37149 , n37154 , n37155 );
xor ( n37157 , n36804 , n36808 );
xor ( n37158 , n37157 , n36813 );
and ( n37159 , n37156 , n37158 );
xor ( n37160 , n36857 , n36861 );
xor ( n37161 , n37160 , n36866 );
and ( n37162 , n37158 , n37161 );
and ( n37163 , n37156 , n37161 );
or ( n37164 , n37159 , n37162 , n37163 );
and ( n37165 , n37140 , n37164 );
xor ( n37166 , n36832 , n36834 );
xor ( n37167 , n37166 , n36837 );
and ( n37168 , n37164 , n37167 );
and ( n37169 , n37140 , n37167 );
or ( n37170 , n37165 , n37168 , n37169 );
and ( n37171 , n25554 , n24902 );
and ( n37172 , n25284 , n24900 );
nor ( n37173 , n37171 , n37172 );
xnor ( n37174 , n37173 , n24397 );
and ( n37175 , n25974 , n24376 );
and ( n37176 , n25765 , n24374 );
nor ( n37177 , n37175 , n37176 );
xnor ( n37178 , n37177 , n23927 );
and ( n37179 , n37174 , n37178 );
and ( n37180 , n26422 , n23944 );
and ( n37181 , n26319 , n23942 );
nor ( n37182 , n37180 , n37181 );
xnor ( n37183 , n37182 , n23550 );
and ( n37184 , n37178 , n37183 );
and ( n37185 , n37174 , n37183 );
or ( n37186 , n37179 , n37184 , n37185 );
and ( n37187 , n23141 , n27529 );
and ( n37188 , n22916 , n27527 );
nor ( n37189 , n37187 , n37188 );
xnor ( n37190 , n37189 , n27034 );
and ( n37191 , n37186 , n37190 );
and ( n37192 , n29623 , n21739 );
not ( n37193 , n37192 );
and ( n37194 , n37193 , n21605 );
and ( n37195 , n37190 , n37194 );
and ( n37196 , n37186 , n37194 );
or ( n37197 , n37191 , n37195 , n37196 );
and ( n37198 , n24131 , n26349 );
and ( n37199 , n23968 , n26347 );
nor ( n37200 , n37198 , n37199 );
xnor ( n37201 , n37200 , n25893 );
and ( n37202 , n24527 , n26027 );
and ( n37203 , n24521 , n26025 );
nor ( n37204 , n37202 , n37203 );
xnor ( n37205 , n37204 , n25499 );
and ( n37206 , n37201 , n37205 );
and ( n37207 , n27135 , n23641 );
and ( n37208 , n26851 , n23639 );
nor ( n37209 , n37207 , n37208 );
xnor ( n37210 , n37209 , n23213 );
and ( n37211 , n37205 , n37210 );
and ( n37212 , n37201 , n37210 );
or ( n37213 , n37206 , n37211 , n37212 );
and ( n37214 , n25765 , n24902 );
and ( n37215 , n25554 , n24900 );
nor ( n37216 , n37214 , n37215 );
xnor ( n37217 , n37216 , n24397 );
and ( n37218 , n26319 , n24376 );
and ( n37219 , n25974 , n24374 );
nor ( n37220 , n37218 , n37219 );
xnor ( n37221 , n37220 , n23927 );
and ( n37222 , n37217 , n37221 );
and ( n37223 , n24940 , n25383 );
and ( n37224 , n24621 , n25381 );
nor ( n37225 , n37223 , n37224 );
xnor ( n37226 , n37225 , n24885 );
and ( n37227 , n37222 , n37226 );
and ( n37228 , n27751 , n23230 );
and ( n37229 , n27352 , n23228 );
nor ( n37230 , n37228 , n37229 );
xnor ( n37231 , n37230 , n22842 );
and ( n37232 , n37226 , n37231 );
and ( n37233 , n37222 , n37231 );
or ( n37234 , n37227 , n37232 , n37233 );
and ( n37235 , n37213 , n37234 );
and ( n37236 , n22756 , n28062 );
and ( n37237 , n22425 , n28060 );
nor ( n37238 , n37236 , n37237 );
xnor ( n37239 , n37238 , n27549 );
and ( n37240 , n37234 , n37239 );
and ( n37241 , n37213 , n37239 );
or ( n37242 , n37235 , n37240 , n37241 );
and ( n37243 , n37197 , n37242 );
xor ( n37244 , n36969 , n36973 );
xor ( n37245 , n37244 , n36976 );
and ( n37246 , n37242 , n37245 );
and ( n37247 , n37197 , n37245 );
or ( n37248 , n37243 , n37246 , n37247 );
xor ( n37249 , n36929 , n36933 );
xor ( n37250 , n37249 , n36938 );
and ( n37251 , n37248 , n37250 );
xor ( n37252 , n36965 , n36979 );
xor ( n37253 , n37252 , n36982 );
and ( n37254 , n37250 , n37253 );
and ( n37255 , n37248 , n37253 );
or ( n37256 , n37251 , n37254 , n37255 );
and ( n37257 , n37170 , n37256 );
xor ( n37258 , n36941 , n36985 );
xor ( n37259 , n37258 , n36988 );
and ( n37260 , n37256 , n37259 );
and ( n37261 , n37170 , n37259 );
or ( n37262 , n37257 , n37260 , n37261 );
and ( n37263 , n22198 , n28628 );
and ( n37264 , n22235 , n28626 );
nor ( n37265 , n37263 , n37264 );
xnor ( n37266 , n37265 , n28096 );
and ( n37267 , n23381 , n26992 );
and ( n37268 , n23271 , n26990 );
nor ( n37269 , n37267 , n37268 );
xnor ( n37270 , n37269 , n26369 );
and ( n37271 , n37266 , n37270 );
xor ( n37272 , n36945 , n36949 );
xor ( n37273 , n37272 , n36954 );
and ( n37274 , n37270 , n37273 );
and ( n37275 , n37266 , n37273 );
or ( n37276 , n37271 , n37274 , n37275 );
and ( n37277 , n29078 , n22048 );
and ( n37278 , n28700 , n22046 );
nor ( n37279 , n37277 , n37278 );
xnor ( n37280 , n37279 , n21853 );
xor ( n37281 , n37144 , n37148 );
xor ( n37282 , n37281 , n37153 );
and ( n37283 , n37280 , n37282 );
xor ( n37284 , n37056 , n37060 );
xor ( n37285 , n37284 , n37065 );
and ( n37286 , n37282 , n37285 );
and ( n37287 , n37280 , n37285 );
or ( n37288 , n37283 , n37286 , n37287 );
and ( n37289 , n37276 , n37288 );
xor ( n37290 , n36957 , n36961 );
xor ( n37291 , n37290 , n36875 );
and ( n37292 , n37288 , n37291 );
and ( n37293 , n37276 , n37291 );
or ( n37294 , n37289 , n37292 , n37293 );
and ( n37295 , n21612 , n29977 );
and ( n37296 , n21451 , n29974 );
nor ( n37297 , n37295 , n37296 );
xnor ( n37298 , n37297 , n28674 );
and ( n37299 , n21876 , n29276 );
and ( n37300 , n21704 , n29274 );
nor ( n37301 , n37299 , n37300 );
xnor ( n37302 , n37301 , n28677 );
and ( n37303 , n37298 , n37302 );
xor ( n37304 , n37068 , n37072 );
xor ( n37305 , n37304 , n37077 );
and ( n37306 , n37302 , n37305 );
and ( n37307 , n37298 , n37305 );
or ( n37308 , n37303 , n37306 , n37307 );
and ( n37309 , n37294 , n37308 );
xor ( n37310 , n37029 , n37033 );
xor ( n37311 , n37310 , n37036 );
and ( n37312 , n37308 , n37311 );
and ( n37313 , n37294 , n37311 );
or ( n37314 , n37309 , n37312 , n37313 );
xor ( n37315 , n37039 , n37041 );
xor ( n37316 , n37315 , n37044 );
and ( n37317 , n37314 , n37316 );
xor ( n37318 , n37090 , n37092 );
xor ( n37319 , n37318 , n37095 );
and ( n37320 , n37316 , n37319 );
and ( n37321 , n37314 , n37319 );
or ( n37322 , n37317 , n37320 , n37321 );
and ( n37323 , n37262 , n37322 );
xor ( n37324 , n37047 , n37049 );
xor ( n37325 , n37324 , n37052 );
and ( n37326 , n37322 , n37325 );
and ( n37327 , n37262 , n37325 );
or ( n37328 , n37323 , n37326 , n37327 );
xor ( n37329 , n36999 , n37001 );
xor ( n37330 , n37329 , n37004 );
and ( n37331 , n37328 , n37330 );
xor ( n37332 , n37055 , n37106 );
xor ( n37333 , n37332 , n37109 );
and ( n37334 , n37330 , n37333 );
and ( n37335 , n37328 , n37333 );
or ( n37336 , n37331 , n37334 , n37335 );
and ( n37337 , n37124 , n37336 );
xor ( n37338 , n37124 , n37336 );
and ( n37339 , n22916 , n28062 );
and ( n37340 , n22756 , n28060 );
nor ( n37341 , n37339 , n37340 );
xnor ( n37342 , n37341 , n27549 );
and ( n37343 , n23573 , n26992 );
and ( n37344 , n23381 , n26990 );
nor ( n37345 , n37343 , n37344 );
xnor ( n37346 , n37345 , n26369 );
and ( n37347 , n37342 , n37346 );
and ( n37348 , n37346 , n37192 );
and ( n37349 , n37342 , n37192 );
or ( n37350 , n37347 , n37348 , n37349 );
and ( n37351 , n28211 , n22859 );
and ( n37352 , n27757 , n22857 );
nor ( n37353 , n37351 , n37352 );
xnor ( n37354 , n37353 , n22418 );
and ( n37355 , n28700 , n22381 );
and ( n37356 , n28810 , n22379 );
nor ( n37357 , n37355 , n37356 );
xnor ( n37358 , n37357 , n22228 );
and ( n37359 , n37354 , n37358 );
xor ( n37360 , n37174 , n37178 );
xor ( n37361 , n37360 , n37183 );
and ( n37362 , n37358 , n37361 );
and ( n37363 , n37354 , n37361 );
or ( n37364 , n37359 , n37362 , n37363 );
and ( n37365 , n37350 , n37364 );
and ( n37366 , n29623 , n21741 );
and ( n37367 , n29318 , n21739 );
nor ( n37368 , n37366 , n37367 );
xnor ( n37369 , n37368 , n21605 );
and ( n37370 , n37364 , n37369 );
and ( n37371 , n37350 , n37369 );
or ( n37372 , n37365 , n37370 , n37371 );
xor ( n37373 , n37128 , n37132 );
xor ( n37374 , n37373 , n37137 );
and ( n37375 , n37372 , n37374 );
xor ( n37376 , n37156 , n37158 );
xor ( n37377 , n37376 , n37161 );
and ( n37378 , n37374 , n37377 );
and ( n37379 , n37372 , n37377 );
or ( n37380 , n37375 , n37378 , n37379 );
xor ( n37381 , n37080 , n37084 );
xor ( n37382 , n37381 , n37087 );
and ( n37383 , n37380 , n37382 );
xor ( n37384 , n37140 , n37164 );
xor ( n37385 , n37384 , n37167 );
and ( n37386 , n37382 , n37385 );
and ( n37387 , n37380 , n37385 );
or ( n37388 , n37383 , n37386 , n37387 );
and ( n37389 , n29318 , n22048 );
and ( n37390 , n29078 , n22046 );
nor ( n37391 , n37389 , n37390 );
xnor ( n37392 , n37391 , n21853 );
xor ( n37393 , n37201 , n37205 );
xor ( n37394 , n37393 , n37210 );
and ( n37395 , n37392 , n37394 );
xor ( n37396 , n37222 , n37226 );
xor ( n37397 , n37396 , n37231 );
and ( n37398 , n37394 , n37397 );
and ( n37399 , n37392 , n37397 );
or ( n37400 , n37395 , n37398 , n37399 );
xor ( n37401 , n37266 , n37270 );
xor ( n37402 , n37401 , n37273 );
and ( n37403 , n37400 , n37402 );
xor ( n37404 , n37280 , n37282 );
xor ( n37405 , n37404 , n37285 );
and ( n37406 , n37402 , n37405 );
and ( n37407 , n37400 , n37405 );
or ( n37408 , n37403 , n37406 , n37407 );
xor ( n37409 , n37276 , n37288 );
xor ( n37410 , n37409 , n37291 );
and ( n37411 , n37408 , n37410 );
xor ( n37412 , n37298 , n37302 );
xor ( n37413 , n37412 , n37305 );
and ( n37414 , n37410 , n37413 );
and ( n37415 , n37408 , n37413 );
or ( n37416 , n37411 , n37414 , n37415 );
and ( n37417 , n25284 , n25383 );
and ( n37418 , n24940 , n25381 );
nor ( n37419 , n37417 , n37418 );
xnor ( n37420 , n37419 , n24885 );
and ( n37421 , n26851 , n23944 );
and ( n37422 , n26422 , n23942 );
nor ( n37423 , n37421 , n37422 );
xnor ( n37424 , n37423 , n23550 );
and ( n37425 , n37420 , n37424 );
and ( n37426 , n27757 , n23230 );
and ( n37427 , n27751 , n23228 );
nor ( n37428 , n37426 , n37427 );
xnor ( n37429 , n37428 , n22842 );
and ( n37430 , n37424 , n37429 );
and ( n37431 , n37420 , n37429 );
or ( n37432 , n37425 , n37430 , n37431 );
xor ( n37433 , n37217 , n37221 );
and ( n37434 , n23968 , n26992 );
and ( n37435 , n23573 , n26990 );
nor ( n37436 , n37434 , n37435 );
xnor ( n37437 , n37436 , n26369 );
and ( n37438 , n37433 , n37437 );
and ( n37439 , n24621 , n26027 );
and ( n37440 , n24527 , n26025 );
nor ( n37441 , n37439 , n37440 );
xnor ( n37442 , n37441 , n25499 );
and ( n37443 , n37437 , n37442 );
and ( n37444 , n37433 , n37442 );
or ( n37445 , n37438 , n37443 , n37444 );
and ( n37446 , n37432 , n37445 );
and ( n37447 , n23271 , n27529 );
and ( n37448 , n23141 , n27527 );
nor ( n37449 , n37447 , n37448 );
xnor ( n37450 , n37449 , n27034 );
and ( n37451 , n37445 , n37450 );
and ( n37452 , n37432 , n37450 );
or ( n37453 , n37446 , n37451 , n37452 );
and ( n37454 , n21955 , n29276 );
and ( n37455 , n21876 , n29274 );
nor ( n37456 , n37454 , n37455 );
xnor ( n37457 , n37456 , n28677 );
and ( n37458 , n37453 , n37457 );
xor ( n37459 , n37186 , n37190 );
xor ( n37460 , n37459 , n37194 );
and ( n37461 , n37457 , n37460 );
and ( n37462 , n37453 , n37460 );
or ( n37463 , n37458 , n37461 , n37462 );
and ( n37464 , n24521 , n26349 );
and ( n37465 , n24131 , n26347 );
nor ( n37466 , n37464 , n37465 );
xnor ( n37467 , n37466 , n25893 );
and ( n37468 , n27352 , n23641 );
and ( n37469 , n27135 , n23639 );
nor ( n37470 , n37468 , n37469 );
xnor ( n37471 , n37470 , n23213 );
and ( n37472 , n37467 , n37471 );
and ( n37473 , n28810 , n22859 );
and ( n37474 , n28211 , n22857 );
nor ( n37475 , n37473 , n37474 );
xnor ( n37476 , n37475 , n22418 );
and ( n37477 , n37471 , n37476 );
and ( n37478 , n37467 , n37476 );
or ( n37479 , n37472 , n37477 , n37478 );
and ( n37480 , n25974 , n24902 );
and ( n37481 , n25765 , n24900 );
nor ( n37482 , n37480 , n37481 );
xnor ( n37483 , n37482 , n24397 );
and ( n37484 , n26422 , n24376 );
and ( n37485 , n26319 , n24374 );
nor ( n37486 , n37484 , n37485 );
xnor ( n37487 , n37486 , n23927 );
and ( n37488 , n37483 , n37487 );
and ( n37489 , n27135 , n23944 );
and ( n37490 , n26851 , n23942 );
nor ( n37491 , n37489 , n37490 );
xnor ( n37492 , n37491 , n23550 );
and ( n37493 , n37487 , n37492 );
and ( n37494 , n37483 , n37492 );
or ( n37495 , n37488 , n37493 , n37494 );
and ( n37496 , n29078 , n22381 );
and ( n37497 , n28700 , n22379 );
nor ( n37498 , n37496 , n37497 );
xnor ( n37499 , n37498 , n22228 );
and ( n37500 , n37495 , n37499 );
and ( n37501 , n29623 , n22046 );
not ( n37502 , n37501 );
and ( n37503 , n37502 , n21853 );
and ( n37504 , n37499 , n37503 );
and ( n37505 , n37495 , n37503 );
or ( n37506 , n37500 , n37504 , n37505 );
and ( n37507 , n37479 , n37506 );
and ( n37508 , n22425 , n28628 );
and ( n37509 , n22198 , n28626 );
nor ( n37510 , n37508 , n37509 );
xnor ( n37511 , n37510 , n28096 );
and ( n37512 , n37506 , n37511 );
and ( n37513 , n37479 , n37511 );
or ( n37514 , n37507 , n37512 , n37513 );
and ( n37515 , n21704 , n29977 );
and ( n37516 , n21612 , n29974 );
nor ( n37517 , n37515 , n37516 );
xnor ( n37518 , n37517 , n28674 );
and ( n37519 , n37514 , n37518 );
xor ( n37520 , n37213 , n37234 );
xor ( n37521 , n37520 , n37239 );
and ( n37522 , n37518 , n37521 );
and ( n37523 , n37514 , n37521 );
or ( n37524 , n37519 , n37522 , n37523 );
and ( n37525 , n37463 , n37524 );
xor ( n37526 , n37197 , n37242 );
xor ( n37527 , n37526 , n37245 );
and ( n37528 , n37524 , n37527 );
and ( n37529 , n37463 , n37527 );
or ( n37530 , n37525 , n37528 , n37529 );
and ( n37531 , n37416 , n37530 );
xor ( n37532 , n37248 , n37250 );
xor ( n37533 , n37532 , n37253 );
and ( n37534 , n37530 , n37533 );
and ( n37535 , n37416 , n37533 );
or ( n37536 , n37531 , n37534 , n37535 );
and ( n37537 , n37388 , n37536 );
xor ( n37538 , n37170 , n37256 );
xor ( n37539 , n37538 , n37259 );
and ( n37540 , n37536 , n37539 );
and ( n37541 , n37388 , n37539 );
or ( n37542 , n37537 , n37540 , n37541 );
xor ( n37543 , n37098 , n37100 );
xor ( n37544 , n37543 , n37103 );
and ( n37545 , n37542 , n37544 );
xor ( n37546 , n37262 , n37322 );
xor ( n37547 , n37546 , n37325 );
and ( n37548 , n37544 , n37547 );
and ( n37549 , n37542 , n37547 );
or ( n37550 , n37545 , n37548 , n37549 );
xor ( n37551 , n37328 , n37330 );
xor ( n37552 , n37551 , n37333 );
and ( n37553 , n37550 , n37552 );
xor ( n37554 , n37550 , n37552 );
xor ( n37555 , n37542 , n37544 );
xor ( n37556 , n37555 , n37547 );
and ( n37557 , n27751 , n23641 );
and ( n37558 , n27352 , n23639 );
nor ( n37559 , n37557 , n37558 );
xnor ( n37560 , n37559 , n23213 );
and ( n37561 , n28700 , n22859 );
and ( n37562 , n28810 , n22857 );
nor ( n37563 , n37561 , n37562 );
xnor ( n37564 , n37563 , n22418 );
and ( n37565 , n37560 , n37564 );
and ( n37566 , n29318 , n22381 );
and ( n37567 , n29078 , n22379 );
nor ( n37568 , n37566 , n37567 );
xnor ( n37569 , n37568 , n22228 );
and ( n37570 , n37564 , n37569 );
and ( n37571 , n37560 , n37569 );
or ( n37572 , n37565 , n37570 , n37571 );
and ( n37573 , n22198 , n29276 );
and ( n37574 , n22235 , n29274 );
nor ( n37575 , n37573 , n37574 );
xnor ( n37576 , n37575 , n28677 );
and ( n37577 , n37572 , n37576 );
xor ( n37578 , n37467 , n37471 );
xor ( n37579 , n37578 , n37476 );
and ( n37580 , n37576 , n37579 );
and ( n37581 , n37572 , n37579 );
or ( n37582 , n37577 , n37580 , n37581 );
and ( n37583 , n21876 , n29977 );
and ( n37584 , n21704 , n29974 );
nor ( n37585 , n37583 , n37584 );
xnor ( n37586 , n37585 , n28674 );
and ( n37587 , n37582 , n37586 );
and ( n37588 , n22235 , n29276 );
and ( n37589 , n21955 , n29274 );
nor ( n37590 , n37588 , n37589 );
xnor ( n37591 , n37590 , n28677 );
and ( n37592 , n37586 , n37591 );
and ( n37593 , n37582 , n37591 );
or ( n37594 , n37587 , n37592 , n37593 );
and ( n37595 , n24940 , n26027 );
and ( n37596 , n24621 , n26025 );
nor ( n37597 , n37595 , n37596 );
xnor ( n37598 , n37597 , n25499 );
and ( n37599 , n25554 , n25383 );
and ( n37600 , n25284 , n25381 );
nor ( n37601 , n37599 , n37600 );
xnor ( n37602 , n37601 , n24885 );
and ( n37603 , n37598 , n37602 );
and ( n37604 , n28211 , n23230 );
and ( n37605 , n27757 , n23228 );
nor ( n37606 , n37604 , n37605 );
xnor ( n37607 , n37606 , n22842 );
and ( n37608 , n37602 , n37607 );
and ( n37609 , n37598 , n37607 );
or ( n37610 , n37603 , n37608 , n37609 );
and ( n37611 , n23141 , n28062 );
and ( n37612 , n22916 , n28060 );
nor ( n37613 , n37611 , n37612 );
xnor ( n37614 , n37613 , n27549 );
and ( n37615 , n37610 , n37614 );
and ( n37616 , n23381 , n27529 );
and ( n37617 , n23271 , n27527 );
nor ( n37618 , n37616 , n37617 );
xnor ( n37619 , n37618 , n27034 );
and ( n37620 , n37614 , n37619 );
and ( n37621 , n37610 , n37619 );
or ( n37622 , n37615 , n37620 , n37621 );
and ( n37623 , n25765 , n25383 );
and ( n37624 , n25554 , n25381 );
nor ( n37625 , n37623 , n37624 );
xnor ( n37626 , n37625 , n24885 );
and ( n37627 , n26319 , n24902 );
and ( n37628 , n25974 , n24900 );
nor ( n37629 , n37627 , n37628 );
xnor ( n37630 , n37629 , n24397 );
and ( n37631 , n37626 , n37630 );
and ( n37632 , n24131 , n26992 );
and ( n37633 , n23968 , n26990 );
nor ( n37634 , n37632 , n37633 );
xnor ( n37635 , n37634 , n26369 );
and ( n37636 , n37631 , n37635 );
and ( n37637 , n24527 , n26349 );
and ( n37638 , n24521 , n26347 );
nor ( n37639 , n37637 , n37638 );
xnor ( n37640 , n37639 , n25893 );
and ( n37641 , n37635 , n37640 );
and ( n37642 , n37631 , n37640 );
or ( n37643 , n37636 , n37641 , n37642 );
and ( n37644 , n22756 , n28628 );
and ( n37645 , n22425 , n28626 );
nor ( n37646 , n37644 , n37645 );
xnor ( n37647 , n37646 , n28096 );
and ( n37648 , n37643 , n37647 );
xor ( n37649 , n37420 , n37424 );
xor ( n37650 , n37649 , n37429 );
and ( n37651 , n37647 , n37650 );
and ( n37652 , n37643 , n37650 );
or ( n37653 , n37648 , n37651 , n37652 );
and ( n37654 , n37622 , n37653 );
xor ( n37655 , n37354 , n37358 );
xor ( n37656 , n37655 , n37361 );
and ( n37657 , n37653 , n37656 );
and ( n37658 , n37622 , n37656 );
or ( n37659 , n37654 , n37657 , n37658 );
and ( n37660 , n37594 , n37659 );
xor ( n37661 , n37350 , n37364 );
xor ( n37662 , n37661 , n37369 );
and ( n37663 , n37659 , n37662 );
and ( n37664 , n37594 , n37662 );
or ( n37665 , n37660 , n37663 , n37664 );
xor ( n37666 , n37342 , n37346 );
xor ( n37667 , n37666 , n37192 );
xor ( n37668 , n37479 , n37506 );
xor ( n37669 , n37668 , n37511 );
and ( n37670 , n37667 , n37669 );
xor ( n37671 , n37432 , n37445 );
xor ( n37672 , n37671 , n37450 );
and ( n37673 , n37669 , n37672 );
and ( n37674 , n37667 , n37672 );
or ( n37675 , n37670 , n37673 , n37674 );
xor ( n37676 , n37453 , n37457 );
xor ( n37677 , n37676 , n37460 );
and ( n37678 , n37675 , n37677 );
xor ( n37679 , n37514 , n37518 );
xor ( n37680 , n37679 , n37521 );
and ( n37681 , n37677 , n37680 );
and ( n37682 , n37675 , n37680 );
or ( n37683 , n37678 , n37681 , n37682 );
and ( n37684 , n37665 , n37683 );
xor ( n37685 , n37372 , n37374 );
xor ( n37686 , n37685 , n37377 );
and ( n37687 , n37683 , n37686 );
and ( n37688 , n37665 , n37686 );
or ( n37689 , n37684 , n37687 , n37688 );
xor ( n37690 , n37294 , n37308 );
xor ( n37691 , n37690 , n37311 );
and ( n37692 , n37689 , n37691 );
xor ( n37693 , n37380 , n37382 );
xor ( n37694 , n37693 , n37385 );
and ( n37695 , n37691 , n37694 );
and ( n37696 , n37689 , n37694 );
or ( n37697 , n37692 , n37695 , n37696 );
xor ( n37698 , n37388 , n37536 );
xor ( n37699 , n37698 , n37539 );
and ( n37700 , n37697 , n37699 );
xor ( n37701 , n37314 , n37316 );
xor ( n37702 , n37701 , n37319 );
and ( n37703 , n37699 , n37702 );
and ( n37704 , n37697 , n37702 );
or ( n37705 , n37700 , n37703 , n37704 );
and ( n37706 , n37556 , n37705 );
xor ( n37707 , n37556 , n37705 );
xor ( n37708 , n37697 , n37699 );
xor ( n37709 , n37708 , n37702 );
and ( n37710 , n26851 , n24376 );
and ( n37711 , n26422 , n24374 );
nor ( n37712 , n37710 , n37711 );
xnor ( n37713 , n37712 , n23927 );
and ( n37714 , n27352 , n23944 );
and ( n37715 , n27135 , n23942 );
nor ( n37716 , n37714 , n37715 );
xnor ( n37717 , n37716 , n23550 );
and ( n37718 , n37713 , n37717 );
and ( n37719 , n29623 , n22379 );
not ( n37720 , n37719 );
and ( n37721 , n37720 , n22228 );
and ( n37722 , n37717 , n37721 );
and ( n37723 , n37713 , n37721 );
or ( n37724 , n37718 , n37722 , n37723 );
and ( n37725 , n23573 , n27529 );
and ( n37726 , n23381 , n27527 );
nor ( n37727 , n37725 , n37726 );
xnor ( n37728 , n37727 , n27034 );
and ( n37729 , n37724 , n37728 );
and ( n37730 , n37728 , n37501 );
and ( n37731 , n37724 , n37501 );
or ( n37732 , n37729 , n37730 , n37731 );
and ( n37733 , n29623 , n22048 );
and ( n37734 , n29318 , n22046 );
nor ( n37735 , n37733 , n37734 );
xnor ( n37736 , n37735 , n21853 );
and ( n37737 , n37732 , n37736 );
xor ( n37738 , n37433 , n37437 );
xor ( n37739 , n37738 , n37442 );
and ( n37740 , n37736 , n37739 );
and ( n37741 , n37732 , n37739 );
or ( n37742 , n37737 , n37740 , n37741 );
xor ( n37743 , n37626 , n37630 );
and ( n37744 , n25284 , n26027 );
and ( n37745 , n24940 , n26025 );
nor ( n37746 , n37744 , n37745 );
xnor ( n37747 , n37746 , n25499 );
and ( n37748 , n37743 , n37747 );
and ( n37749 , n28810 , n23230 );
and ( n37750 , n28211 , n23228 );
nor ( n37751 , n37749 , n37750 );
xnor ( n37752 , n37751 , n22842 );
and ( n37753 , n37747 , n37752 );
and ( n37754 , n37743 , n37752 );
or ( n37755 , n37748 , n37753 , n37754 );
and ( n37756 , n22425 , n29276 );
and ( n37757 , n22198 , n29274 );
nor ( n37758 , n37756 , n37757 );
xnor ( n37759 , n37758 , n28677 );
and ( n37760 , n37755 , n37759 );
and ( n37761 , n23271 , n28062 );
and ( n37762 , n23141 , n28060 );
nor ( n37763 , n37761 , n37762 );
xnor ( n37764 , n37763 , n27549 );
and ( n37765 , n37759 , n37764 );
and ( n37766 , n37755 , n37764 );
or ( n37767 , n37760 , n37765 , n37766 );
and ( n37768 , n23968 , n27529 );
and ( n37769 , n23573 , n27527 );
nor ( n37770 , n37768 , n37769 );
xnor ( n37771 , n37770 , n27034 );
and ( n37772 , n24521 , n26992 );
and ( n37773 , n24131 , n26990 );
nor ( n37774 , n37772 , n37773 );
xnor ( n37775 , n37774 , n26369 );
and ( n37776 , n37771 , n37775 );
and ( n37777 , n27757 , n23641 );
and ( n37778 , n27751 , n23639 );
nor ( n37779 , n37777 , n37778 );
xnor ( n37780 , n37779 , n23213 );
and ( n37781 , n37775 , n37780 );
and ( n37782 , n37771 , n37780 );
or ( n37783 , n37776 , n37781 , n37782 );
xor ( n37784 , n37483 , n37487 );
xor ( n37785 , n37784 , n37492 );
and ( n37786 , n37783 , n37785 );
xor ( n37787 , n37598 , n37602 );
xor ( n37788 , n37787 , n37607 );
and ( n37789 , n37785 , n37788 );
and ( n37790 , n37783 , n37788 );
or ( n37791 , n37786 , n37789 , n37790 );
and ( n37792 , n37767 , n37791 );
xor ( n37793 , n37495 , n37499 );
xor ( n37794 , n37793 , n37503 );
and ( n37795 , n37791 , n37794 );
and ( n37796 , n37767 , n37794 );
or ( n37797 , n37792 , n37795 , n37796 );
and ( n37798 , n37742 , n37797 );
xor ( n37799 , n37392 , n37394 );
xor ( n37800 , n37799 , n37397 );
and ( n37801 , n37797 , n37800 );
and ( n37802 , n37742 , n37800 );
or ( n37803 , n37798 , n37801 , n37802 );
xor ( n37804 , n37594 , n37659 );
xor ( n37805 , n37804 , n37662 );
and ( n37806 , n37803 , n37805 );
xor ( n37807 , n37400 , n37402 );
xor ( n37808 , n37807 , n37405 );
and ( n37809 , n37805 , n37808 );
and ( n37810 , n37803 , n37808 );
or ( n37811 , n37806 , n37809 , n37810 );
xor ( n37812 , n37408 , n37410 );
xor ( n37813 , n37812 , n37413 );
and ( n37814 , n37811 , n37813 );
xor ( n37815 , n37463 , n37524 );
xor ( n37816 , n37815 , n37527 );
and ( n37817 , n37813 , n37816 );
and ( n37818 , n37811 , n37816 );
or ( n37819 , n37814 , n37817 , n37818 );
xor ( n37820 , n37416 , n37530 );
xor ( n37821 , n37820 , n37533 );
and ( n37822 , n37819 , n37821 );
xor ( n37823 , n37689 , n37691 );
xor ( n37824 , n37823 , n37694 );
and ( n37825 , n37821 , n37824 );
and ( n37826 , n37819 , n37824 );
or ( n37827 , n37822 , n37825 , n37826 );
and ( n37828 , n37709 , n37827 );
xor ( n37829 , n37709 , n37827 );
xor ( n37830 , n37819 , n37821 );
xor ( n37831 , n37830 , n37824 );
and ( n37832 , n24621 , n26349 );
and ( n37833 , n24527 , n26347 );
nor ( n37834 , n37832 , n37833 );
xnor ( n37835 , n37834 , n25893 );
and ( n37836 , n29078 , n22859 );
and ( n37837 , n28700 , n22857 );
nor ( n37838 , n37836 , n37837 );
xnor ( n37839 , n37838 , n22418 );
and ( n37840 , n37835 , n37839 );
and ( n37841 , n29623 , n22381 );
and ( n37842 , n29318 , n22379 );
nor ( n37843 , n37841 , n37842 );
xnor ( n37844 , n37843 , n22228 );
and ( n37845 , n37839 , n37844 );
and ( n37846 , n37835 , n37844 );
or ( n37847 , n37840 , n37845 , n37846 );
and ( n37848 , n22916 , n28628 );
and ( n37849 , n22756 , n28626 );
nor ( n37850 , n37848 , n37849 );
xnor ( n37851 , n37850 , n28096 );
and ( n37852 , n37847 , n37851 );
xor ( n37853 , n37560 , n37564 );
xor ( n37854 , n37853 , n37569 );
and ( n37855 , n37851 , n37854 );
and ( n37856 , n37847 , n37854 );
or ( n37857 , n37852 , n37855 , n37856 );
and ( n37858 , n21955 , n29977 );
and ( n37859 , n21876 , n29974 );
nor ( n37860 , n37858 , n37859 );
xnor ( n37861 , n37860 , n28674 );
and ( n37862 , n37857 , n37861 );
xor ( n37863 , n37610 , n37614 );
xor ( n37864 , n37863 , n37619 );
and ( n37865 , n37861 , n37864 );
and ( n37866 , n37857 , n37864 );
or ( n37867 , n37862 , n37865 , n37866 );
xor ( n37868 , n37667 , n37669 );
xor ( n37869 , n37868 , n37672 );
and ( n37870 , n37867 , n37869 );
xor ( n37871 , n37622 , n37653 );
xor ( n37872 , n37871 , n37656 );
and ( n37873 , n37869 , n37872 );
and ( n37874 , n37867 , n37872 );
or ( n37875 , n37870 , n37873 , n37874 );
and ( n37876 , n25974 , n25383 );
and ( n37877 , n25765 , n25381 );
nor ( n37878 , n37876 , n37877 );
xnor ( n37879 , n37878 , n24885 );
and ( n37880 , n26422 , n24902 );
and ( n37881 , n26319 , n24900 );
nor ( n37882 , n37880 , n37881 );
xnor ( n37883 , n37882 , n24397 );
and ( n37884 , n37879 , n37883 );
and ( n37885 , n37883 , n37719 );
and ( n37886 , n37879 , n37719 );
or ( n37887 , n37884 , n37885 , n37886 );
and ( n37888 , n25765 , n26027 );
and ( n37889 , n25554 , n26025 );
nor ( n37890 , n37888 , n37889 );
xnor ( n37891 , n37890 , n25499 );
and ( n37892 , n26319 , n25383 );
and ( n37893 , n25974 , n25381 );
nor ( n37894 , n37892 , n37893 );
xnor ( n37895 , n37894 , n24885 );
and ( n37896 , n37891 , n37895 );
and ( n37897 , n27135 , n24376 );
and ( n37898 , n26851 , n24374 );
nor ( n37899 , n37897 , n37898 );
xnor ( n37900 , n37899 , n23927 );
and ( n37901 , n37896 , n37900 );
and ( n37902 , n27751 , n23944 );
and ( n37903 , n27352 , n23942 );
nor ( n37904 , n37902 , n37903 );
xnor ( n37905 , n37904 , n23550 );
and ( n37906 , n37900 , n37905 );
and ( n37907 , n37896 , n37905 );
or ( n37908 , n37901 , n37906 , n37907 );
and ( n37909 , n37887 , n37908 );
xor ( n37910 , n37713 , n37717 );
xor ( n37911 , n37910 , n37721 );
and ( n37912 , n37908 , n37911 );
and ( n37913 , n37887 , n37911 );
or ( n37914 , n37909 , n37912 , n37913 );
xor ( n37915 , n37631 , n37635 );
xor ( n37916 , n37915 , n37640 );
and ( n37917 , n37914 , n37916 );
xor ( n37918 , n37724 , n37728 );
xor ( n37919 , n37918 , n37501 );
and ( n37920 , n37916 , n37919 );
and ( n37921 , n37914 , n37919 );
or ( n37922 , n37917 , n37920 , n37921 );
xor ( n37923 , n37572 , n37576 );
xor ( n37924 , n37923 , n37579 );
and ( n37925 , n37922 , n37924 );
xor ( n37926 , n37643 , n37647 );
xor ( n37927 , n37926 , n37650 );
and ( n37928 , n37924 , n37927 );
and ( n37929 , n37922 , n37927 );
or ( n37930 , n37925 , n37928 , n37929 );
xor ( n37931 , n37582 , n37586 );
xor ( n37932 , n37931 , n37591 );
and ( n37933 , n37930 , n37932 );
xor ( n37934 , n37742 , n37797 );
xor ( n37935 , n37934 , n37800 );
and ( n37936 , n37932 , n37935 );
and ( n37937 , n37930 , n37935 );
or ( n37938 , n37933 , n37936 , n37937 );
and ( n37939 , n37875 , n37938 );
xor ( n37940 , n37675 , n37677 );
xor ( n37941 , n37940 , n37680 );
and ( n37942 , n37938 , n37941 );
and ( n37943 , n37875 , n37941 );
or ( n37944 , n37939 , n37942 , n37943 );
xor ( n37945 , n37665 , n37683 );
xor ( n37946 , n37945 , n37686 );
and ( n37947 , n37944 , n37946 );
xor ( n37948 , n37811 , n37813 );
xor ( n37949 , n37948 , n37816 );
and ( n37950 , n37946 , n37949 );
and ( n37951 , n37944 , n37949 );
or ( n37952 , n37947 , n37950 , n37951 );
and ( n37953 , n37831 , n37952 );
xor ( n37954 , n37831 , n37952 );
xor ( n37955 , n37944 , n37946 );
xor ( n37956 , n37955 , n37949 );
and ( n37957 , n24527 , n26992 );
and ( n37958 , n24521 , n26990 );
nor ( n37959 , n37957 , n37958 );
xnor ( n37960 , n37959 , n26369 );
and ( n37961 , n24940 , n26349 );
and ( n37962 , n24621 , n26347 );
nor ( n37963 , n37961 , n37962 );
xnor ( n37964 , n37963 , n25893 );
and ( n37965 , n37960 , n37964 );
and ( n37966 , n28211 , n23641 );
and ( n37967 , n27757 , n23639 );
nor ( n37968 , n37966 , n37967 );
xnor ( n37969 , n37968 , n23213 );
and ( n37970 , n37964 , n37969 );
and ( n37971 , n37960 , n37969 );
or ( n37972 , n37965 , n37970 , n37971 );
and ( n37973 , n22198 , n29977 );
and ( n37974 , n22235 , n29974 );
nor ( n37975 , n37973 , n37974 );
xnor ( n37976 , n37975 , n28674 );
and ( n37977 , n37972 , n37976 );
and ( n37978 , n23141 , n28628 );
and ( n37979 , n22916 , n28626 );
nor ( n37980 , n37978 , n37979 );
xnor ( n37981 , n37980 , n28096 );
and ( n37982 , n37976 , n37981 );
and ( n37983 , n37972 , n37981 );
or ( n37984 , n37977 , n37982 , n37983 );
xor ( n37985 , n37835 , n37839 );
xor ( n37986 , n37985 , n37844 );
xor ( n37987 , n37771 , n37775 );
xor ( n37988 , n37987 , n37780 );
and ( n37989 , n37986 , n37988 );
xor ( n37990 , n37743 , n37747 );
xor ( n37991 , n37990 , n37752 );
and ( n37992 , n37988 , n37991 );
and ( n37993 , n37986 , n37991 );
or ( n37994 , n37989 , n37992 , n37993 );
and ( n37995 , n37984 , n37994 );
xor ( n37996 , n37783 , n37785 );
xor ( n37997 , n37996 , n37788 );
and ( n37998 , n37994 , n37997 );
and ( n37999 , n37984 , n37997 );
or ( n38000 , n37995 , n37998 , n37999 );
xor ( n38001 , n37732 , n37736 );
xor ( n38002 , n38001 , n37739 );
and ( n38003 , n38000 , n38002 );
xor ( n38004 , n37767 , n37791 );
xor ( n38005 , n38004 , n37794 );
and ( n38006 , n38002 , n38005 );
and ( n38007 , n38000 , n38005 );
or ( n38008 , n38003 , n38006 , n38007 );
and ( n38009 , n24131 , n27529 );
and ( n38010 , n23968 , n27527 );
nor ( n38011 , n38009 , n38010 );
xnor ( n38012 , n38011 , n27034 );
and ( n38013 , n25554 , n26027 );
and ( n38014 , n25284 , n26025 );
nor ( n38015 , n38013 , n38014 );
xnor ( n38016 , n38015 , n25499 );
and ( n38017 , n38012 , n38016 );
and ( n38018 , n28700 , n23230 );
and ( n38019 , n28810 , n23228 );
nor ( n38020 , n38018 , n38019 );
xnor ( n38021 , n38020 , n22842 );
and ( n38022 , n38016 , n38021 );
and ( n38023 , n38012 , n38021 );
or ( n38024 , n38017 , n38022 , n38023 );
and ( n38025 , n22756 , n29276 );
and ( n38026 , n22425 , n29274 );
nor ( n38027 , n38025 , n38026 );
xnor ( n38028 , n38027 , n28677 );
and ( n38029 , n38024 , n38028 );
and ( n38030 , n23381 , n28062 );
and ( n38031 , n23271 , n28060 );
nor ( n38032 , n38030 , n38031 );
xnor ( n38033 , n38032 , n27549 );
and ( n38034 , n38028 , n38033 );
and ( n38035 , n38024 , n38033 );
or ( n38036 , n38029 , n38034 , n38035 );
and ( n38037 , n22235 , n29977 );
and ( n38038 , n21955 , n29974 );
nor ( n38039 , n38037 , n38038 );
xnor ( n38040 , n38039 , n28674 );
and ( n38041 , n38036 , n38040 );
xor ( n38042 , n37755 , n37759 );
xor ( n38043 , n38042 , n37764 );
and ( n38044 , n38040 , n38043 );
and ( n38045 , n38036 , n38043 );
or ( n38046 , n38041 , n38044 , n38045 );
xor ( n38047 , n37857 , n37861 );
xor ( n38048 , n38047 , n37864 );
and ( n38049 , n38046 , n38048 );
xor ( n38050 , n37922 , n37924 );
xor ( n38051 , n38050 , n37927 );
and ( n38052 , n38048 , n38051 );
and ( n38053 , n38046 , n38051 );
or ( n38054 , n38049 , n38052 , n38053 );
and ( n38055 , n38008 , n38054 );
xor ( n38056 , n37867 , n37869 );
xor ( n38057 , n38056 , n37872 );
and ( n38058 , n38054 , n38057 );
and ( n38059 , n38008 , n38057 );
or ( n38060 , n38055 , n38058 , n38059 );
xor ( n38061 , n37803 , n37805 );
xor ( n38062 , n38061 , n37808 );
and ( n38063 , n38060 , n38062 );
xor ( n38064 , n37875 , n37938 );
xor ( n38065 , n38064 , n37941 );
and ( n38066 , n38062 , n38065 );
and ( n38067 , n38060 , n38065 );
or ( n38068 , n38063 , n38066 , n38067 );
and ( n38069 , n37956 , n38068 );
xor ( n38070 , n37956 , n38068 );
xor ( n38071 , n38060 , n38062 );
xor ( n38072 , n38071 , n38065 );
and ( n38073 , n26851 , n24902 );
and ( n38074 , n26422 , n24900 );
nor ( n38075 , n38073 , n38074 );
xnor ( n38076 , n38075 , n24397 );
and ( n38077 , n27352 , n24376 );
and ( n38078 , n27135 , n24374 );
nor ( n38079 , n38077 , n38078 );
xnor ( n38080 , n38079 , n23927 );
and ( n38081 , n38076 , n38080 );
and ( n38082 , n29623 , n22857 );
not ( n38083 , n38082 );
and ( n38084 , n38083 , n22418 );
and ( n38085 , n38080 , n38084 );
and ( n38086 , n38076 , n38084 );
or ( n38087 , n38081 , n38085 , n38086 );
and ( n38088 , n23573 , n28062 );
and ( n38089 , n23381 , n28060 );
nor ( n38090 , n38088 , n38089 );
xnor ( n38091 , n38090 , n27549 );
and ( n38092 , n38087 , n38091 );
and ( n38093 , n29318 , n22859 );
and ( n38094 , n29078 , n22857 );
nor ( n38095 , n38093 , n38094 );
xnor ( n38096 , n38095 , n22418 );
and ( n38097 , n38091 , n38096 );
and ( n38098 , n38087 , n38096 );
or ( n38099 , n38092 , n38097 , n38098 );
xor ( n38100 , n37891 , n37895 );
and ( n38101 , n27757 , n23944 );
and ( n38102 , n27751 , n23942 );
nor ( n38103 , n38101 , n38102 );
xnor ( n38104 , n38103 , n23550 );
and ( n38105 , n38100 , n38104 );
and ( n38106 , n29078 , n23230 );
and ( n38107 , n28700 , n23228 );
nor ( n38108 , n38106 , n38107 );
xnor ( n38109 , n38108 , n22842 );
and ( n38110 , n38104 , n38109 );
and ( n38111 , n38100 , n38109 );
or ( n38112 , n38105 , n38110 , n38111 );
xor ( n38113 , n37879 , n37883 );
xor ( n38114 , n38113 , n37719 );
and ( n38115 , n38112 , n38114 );
xor ( n38116 , n37896 , n37900 );
xor ( n38117 , n38116 , n37905 );
and ( n38118 , n38114 , n38117 );
and ( n38119 , n38112 , n38117 );
or ( n38120 , n38115 , n38118 , n38119 );
and ( n38121 , n38099 , n38120 );
xor ( n38122 , n37887 , n37908 );
xor ( n38123 , n38122 , n37911 );
and ( n38124 , n38120 , n38123 );
and ( n38125 , n38099 , n38123 );
or ( n38126 , n38121 , n38124 , n38125 );
xor ( n38127 , n37847 , n37851 );
xor ( n38128 , n38127 , n37854 );
and ( n38129 , n38126 , n38128 );
xor ( n38130 , n37914 , n37916 );
xor ( n38131 , n38130 , n37919 );
and ( n38132 , n38128 , n38131 );
and ( n38133 , n38126 , n38131 );
or ( n38134 , n38129 , n38132 , n38133 );
and ( n38135 , n24621 , n26992 );
and ( n38136 , n24527 , n26990 );
nor ( n38137 , n38135 , n38136 );
xnor ( n38138 , n38137 , n26369 );
and ( n38139 , n25284 , n26349 );
and ( n38140 , n24940 , n26347 );
nor ( n38141 , n38139 , n38140 );
xnor ( n38142 , n38141 , n25893 );
and ( n38143 , n38138 , n38142 );
and ( n38144 , n28810 , n23641 );
and ( n38145 , n28211 , n23639 );
nor ( n38146 , n38144 , n38145 );
xnor ( n38147 , n38146 , n23213 );
and ( n38148 , n38142 , n38147 );
and ( n38149 , n38138 , n38147 );
or ( n38150 , n38143 , n38148 , n38149 );
and ( n38151 , n22425 , n29977 );
and ( n38152 , n22198 , n29974 );
nor ( n38153 , n38151 , n38152 );
xnor ( n38154 , n38153 , n28674 );
and ( n38155 , n38150 , n38154 );
and ( n38156 , n22916 , n29276 );
and ( n38157 , n22756 , n29274 );
nor ( n38158 , n38156 , n38157 );
xnor ( n38159 , n38158 , n28677 );
and ( n38160 , n38154 , n38159 );
and ( n38161 , n38150 , n38159 );
or ( n38162 , n38155 , n38160 , n38161 );
and ( n38163 , n25974 , n26027 );
and ( n38164 , n25765 , n26025 );
nor ( n38165 , n38163 , n38164 );
xnor ( n38166 , n38165 , n25499 );
and ( n38167 , n26422 , n25383 );
and ( n38168 , n26319 , n25381 );
nor ( n38169 , n38167 , n38168 );
xnor ( n38170 , n38169 , n24885 );
and ( n38171 , n38166 , n38170 );
and ( n38172 , n38170 , n38082 );
and ( n38173 , n38166 , n38082 );
or ( n38174 , n38171 , n38172 , n38173 );
and ( n38175 , n23968 , n28062 );
and ( n38176 , n23573 , n28060 );
nor ( n38177 , n38175 , n38176 );
xnor ( n38178 , n38177 , n27549 );
and ( n38179 , n38174 , n38178 );
and ( n38180 , n24521 , n27529 );
and ( n38181 , n24131 , n27527 );
nor ( n38182 , n38180 , n38181 );
xnor ( n38183 , n38182 , n27034 );
and ( n38184 , n38178 , n38183 );
and ( n38185 , n38174 , n38183 );
or ( n38186 , n38179 , n38184 , n38185 );
and ( n38187 , n23271 , n28628 );
and ( n38188 , n23141 , n28626 );
nor ( n38189 , n38187 , n38188 );
xnor ( n38190 , n38189 , n28096 );
and ( n38191 , n38186 , n38190 );
xor ( n38192 , n38012 , n38016 );
xor ( n38193 , n38192 , n38021 );
and ( n38194 , n38190 , n38193 );
and ( n38195 , n38186 , n38193 );
or ( n38196 , n38191 , n38194 , n38195 );
and ( n38197 , n38162 , n38196 );
xor ( n38198 , n37972 , n37976 );
xor ( n38199 , n38198 , n37981 );
and ( n38200 , n38196 , n38199 );
and ( n38201 , n38162 , n38199 );
or ( n38202 , n38197 , n38200 , n38201 );
xor ( n38203 , n38036 , n38040 );
xor ( n38204 , n38203 , n38043 );
and ( n38205 , n38202 , n38204 );
xor ( n38206 , n37984 , n37994 );
xor ( n38207 , n38206 , n37997 );
and ( n38208 , n38204 , n38207 );
and ( n38209 , n38202 , n38207 );
or ( n38210 , n38205 , n38208 , n38209 );
and ( n38211 , n38134 , n38210 );
xor ( n38212 , n38000 , n38002 );
xor ( n38213 , n38212 , n38005 );
and ( n38214 , n38210 , n38213 );
and ( n38215 , n38134 , n38213 );
or ( n38216 , n38211 , n38214 , n38215 );
xor ( n38217 , n37930 , n37932 );
xor ( n38218 , n38217 , n37935 );
and ( n38219 , n38216 , n38218 );
xor ( n38220 , n38008 , n38054 );
xor ( n38221 , n38220 , n38057 );
and ( n38222 , n38218 , n38221 );
and ( n38223 , n38216 , n38221 );
or ( n38224 , n38219 , n38222 , n38223 );
and ( n38225 , n38072 , n38224 );
xor ( n38226 , n38072 , n38224 );
and ( n38227 , n27135 , n24902 );
and ( n38228 , n26851 , n24900 );
nor ( n38229 , n38227 , n38228 );
xnor ( n38230 , n38229 , n24397 );
and ( n38231 , n27751 , n24376 );
and ( n38232 , n27352 , n24374 );
nor ( n38233 , n38231 , n38232 );
xnor ( n38234 , n38233 , n23927 );
and ( n38235 , n38230 , n38234 );
and ( n38236 , n28211 , n23944 );
and ( n38237 , n27757 , n23942 );
nor ( n38238 , n38236 , n38237 );
xnor ( n38239 , n38238 , n23550 );
and ( n38240 , n38234 , n38239 );
and ( n38241 , n38230 , n38239 );
or ( n38242 , n38235 , n38240 , n38241 );
and ( n38243 , n25765 , n26349 );
and ( n38244 , n25554 , n26347 );
nor ( n38245 , n38243 , n38244 );
xnor ( n38246 , n38245 , n25893 );
and ( n38247 , n26319 , n26027 );
and ( n38248 , n25974 , n26025 );
nor ( n38249 , n38247 , n38248 );
xnor ( n38250 , n38249 , n25499 );
and ( n38251 , n38246 , n38250 );
and ( n38252 , n25554 , n26349 );
and ( n38253 , n25284 , n26347 );
nor ( n38254 , n38252 , n38253 );
xnor ( n38255 , n38254 , n25893 );
and ( n38256 , n38251 , n38255 );
and ( n38257 , n29318 , n23230 );
and ( n38258 , n29078 , n23228 );
nor ( n38259 , n38257 , n38258 );
xnor ( n38260 , n38259 , n22842 );
and ( n38261 , n38255 , n38260 );
and ( n38262 , n38251 , n38260 );
or ( n38263 , n38256 , n38261 , n38262 );
and ( n38264 , n38242 , n38263 );
and ( n38265 , n29623 , n22859 );
and ( n38266 , n29318 , n22857 );
nor ( n38267 , n38265 , n38266 );
xnor ( n38268 , n38267 , n22418 );
and ( n38269 , n38263 , n38268 );
and ( n38270 , n38242 , n38268 );
or ( n38271 , n38264 , n38269 , n38270 );
xor ( n38272 , n37960 , n37964 );
xor ( n38273 , n38272 , n37969 );
and ( n38274 , n38271 , n38273 );
xor ( n38275 , n38087 , n38091 );
xor ( n38276 , n38275 , n38096 );
and ( n38277 , n38273 , n38276 );
and ( n38278 , n38271 , n38276 );
or ( n38279 , n38274 , n38277 , n38278 );
xor ( n38280 , n38024 , n38028 );
xor ( n38281 , n38280 , n38033 );
and ( n38282 , n38279 , n38281 );
xor ( n38283 , n37986 , n37988 );
xor ( n38284 , n38283 , n37991 );
and ( n38285 , n38281 , n38284 );
and ( n38286 , n38279 , n38284 );
or ( n38287 , n38282 , n38285 , n38286 );
and ( n38288 , n26851 , n25383 );
and ( n38289 , n26422 , n25381 );
nor ( n38290 , n38288 , n38289 );
xnor ( n38291 , n38290 , n24885 );
and ( n38292 , n27352 , n24902 );
and ( n38293 , n27135 , n24900 );
nor ( n38294 , n38292 , n38293 );
xnor ( n38295 , n38294 , n24397 );
and ( n38296 , n38291 , n38295 );
and ( n38297 , n29623 , n23228 );
not ( n38298 , n38297 );
and ( n38299 , n38298 , n22842 );
and ( n38300 , n38295 , n38299 );
and ( n38301 , n38291 , n38299 );
or ( n38302 , n38296 , n38300 , n38301 );
and ( n38303 , n24940 , n26992 );
and ( n38304 , n24621 , n26990 );
nor ( n38305 , n38303 , n38304 );
xnor ( n38306 , n38305 , n26369 );
and ( n38307 , n38302 , n38306 );
xor ( n38308 , n38166 , n38170 );
xor ( n38309 , n38308 , n38082 );
and ( n38310 , n38306 , n38309 );
and ( n38311 , n38302 , n38309 );
or ( n38312 , n38307 , n38310 , n38311 );
xor ( n38313 , n38138 , n38142 );
xor ( n38314 , n38313 , n38147 );
and ( n38315 , n38312 , n38314 );
xor ( n38316 , n38174 , n38178 );
xor ( n38317 , n38316 , n38183 );
and ( n38318 , n38314 , n38317 );
and ( n38319 , n38312 , n38317 );
or ( n38320 , n38315 , n38318 , n38319 );
xor ( n38321 , n38150 , n38154 );
xor ( n38322 , n38321 , n38159 );
and ( n38323 , n38320 , n38322 );
xor ( n38324 , n38186 , n38190 );
xor ( n38325 , n38324 , n38193 );
and ( n38326 , n38322 , n38325 );
and ( n38327 , n38320 , n38325 );
or ( n38328 , n38323 , n38326 , n38327 );
and ( n38329 , n24131 , n28062 );
and ( n38330 , n23968 , n28060 );
nor ( n38331 , n38329 , n38330 );
xnor ( n38332 , n38331 , n27549 );
and ( n38333 , n24527 , n27529 );
and ( n38334 , n24521 , n27527 );
nor ( n38335 , n38333 , n38334 );
xnor ( n38336 , n38335 , n27034 );
and ( n38337 , n38332 , n38336 );
and ( n38338 , n28700 , n23641 );
and ( n38339 , n28810 , n23639 );
nor ( n38340 , n38338 , n38339 );
xnor ( n38341 , n38340 , n23213 );
and ( n38342 , n38336 , n38341 );
and ( n38343 , n38332 , n38341 );
or ( n38344 , n38337 , n38342 , n38343 );
and ( n38345 , n22756 , n29977 );
and ( n38346 , n22425 , n29974 );
nor ( n38347 , n38345 , n38346 );
xnor ( n38348 , n38347 , n28674 );
and ( n38349 , n38344 , n38348 );
and ( n38350 , n23381 , n28628 );
and ( n38351 , n23271 , n28626 );
nor ( n38352 , n38350 , n38351 );
xnor ( n38353 , n38352 , n28096 );
and ( n38354 , n38348 , n38353 );
and ( n38355 , n38344 , n38353 );
or ( n38356 , n38349 , n38354 , n38355 );
and ( n38357 , n23141 , n29276 );
and ( n38358 , n22916 , n29274 );
nor ( n38359 , n38357 , n38358 );
xnor ( n38360 , n38359 , n28677 );
xor ( n38361 , n38076 , n38080 );
xor ( n38362 , n38361 , n38084 );
and ( n38363 , n38360 , n38362 );
xor ( n38364 , n38100 , n38104 );
xor ( n38365 , n38364 , n38109 );
and ( n38366 , n38362 , n38365 );
and ( n38367 , n38360 , n38365 );
or ( n38368 , n38363 , n38366 , n38367 );
and ( n38369 , n38356 , n38368 );
xor ( n38370 , n38112 , n38114 );
xor ( n38371 , n38370 , n38117 );
and ( n38372 , n38368 , n38371 );
and ( n38373 , n38356 , n38371 );
or ( n38374 , n38369 , n38372 , n38373 );
and ( n38375 , n38328 , n38374 );
xor ( n38376 , n38099 , n38120 );
xor ( n38377 , n38376 , n38123 );
and ( n38378 , n38374 , n38377 );
and ( n38379 , n38328 , n38377 );
or ( n38380 , n38375 , n38378 , n38379 );
and ( n38381 , n38287 , n38380 );
xor ( n38382 , n38126 , n38128 );
xor ( n38383 , n38382 , n38131 );
and ( n38384 , n38380 , n38383 );
and ( n38385 , n38287 , n38383 );
or ( n38386 , n38381 , n38384 , n38385 );
xor ( n38387 , n38046 , n38048 );
xor ( n38388 , n38387 , n38051 );
and ( n38389 , n38386 , n38388 );
xor ( n38390 , n38134 , n38210 );
xor ( n38391 , n38390 , n38213 );
and ( n38392 , n38388 , n38391 );
and ( n38393 , n38386 , n38391 );
or ( n38394 , n38389 , n38392 , n38393 );
xor ( n38395 , n38216 , n38218 );
xor ( n38396 , n38395 , n38221 );
and ( n38397 , n38394 , n38396 );
xor ( n38398 , n38394 , n38396 );
xor ( n38399 , n38386 , n38388 );
xor ( n38400 , n38399 , n38391 );
xor ( n38401 , n38162 , n38196 );
xor ( n38402 , n38401 , n38199 );
xor ( n38403 , n38279 , n38281 );
xor ( n38404 , n38403 , n38284 );
and ( n38405 , n38402 , n38404 );
xor ( n38406 , n38328 , n38374 );
xor ( n38407 , n38406 , n38377 );
and ( n38408 , n38404 , n38407 );
and ( n38409 , n38402 , n38407 );
or ( n38410 , n38405 , n38408 , n38409 );
xor ( n38411 , n38202 , n38204 );
xor ( n38412 , n38411 , n38207 );
and ( n38413 , n38410 , n38412 );
xor ( n38414 , n38287 , n38380 );
xor ( n38415 , n38414 , n38383 );
and ( n38416 , n38412 , n38415 );
and ( n38417 , n38410 , n38415 );
or ( n38418 , n38413 , n38416 , n38417 );
and ( n38419 , n38400 , n38418 );
xor ( n38420 , n38400 , n38418 );
xor ( n38421 , n38410 , n38412 );
xor ( n38422 , n38421 , n38415 );
and ( n38423 , n25974 , n26349 );
and ( n38424 , n25765 , n26347 );
nor ( n38425 , n38423 , n38424 );
xnor ( n38426 , n38425 , n25893 );
and ( n38427 , n26422 , n26027 );
and ( n38428 , n26319 , n26025 );
nor ( n38429 , n38427 , n38428 );
xnor ( n38430 , n38429 , n25499 );
and ( n38431 , n38426 , n38430 );
and ( n38432 , n27135 , n25383 );
and ( n38433 , n26851 , n25381 );
nor ( n38434 , n38432 , n38433 );
xnor ( n38435 , n38434 , n24885 );
and ( n38436 , n38430 , n38435 );
and ( n38437 , n38426 , n38435 );
or ( n38438 , n38431 , n38436 , n38437 );
and ( n38439 , n24521 , n28062 );
and ( n38440 , n24131 , n28060 );
nor ( n38441 , n38439 , n38440 );
xnor ( n38442 , n38441 , n27549 );
and ( n38443 , n38438 , n38442 );
and ( n38444 , n29623 , n23230 );
and ( n38445 , n29318 , n23228 );
nor ( n38446 , n38444 , n38445 );
xnor ( n38447 , n38446 , n22842 );
and ( n38448 , n38442 , n38447 );
and ( n38449 , n38438 , n38447 );
or ( n38450 , n38443 , n38448 , n38449 );
and ( n38451 , n22916 , n29977 );
and ( n38452 , n22756 , n29974 );
nor ( n38453 , n38451 , n38452 );
xnor ( n38454 , n38453 , n28674 );
and ( n38455 , n38450 , n38454 );
and ( n38456 , n23271 , n29276 );
and ( n38457 , n23141 , n29274 );
nor ( n38458 , n38456 , n38457 );
xnor ( n38459 , n38458 , n28677 );
and ( n38460 , n38454 , n38459 );
and ( n38461 , n38450 , n38459 );
or ( n38462 , n38455 , n38460 , n38461 );
xor ( n38463 , n38246 , n38250 );
and ( n38464 , n27757 , n24376 );
and ( n38465 , n27751 , n24374 );
nor ( n38466 , n38464 , n38465 );
xnor ( n38467 , n38466 , n23927 );
and ( n38468 , n38463 , n38467 );
and ( n38469 , n28810 , n23944 );
and ( n38470 , n28211 , n23942 );
nor ( n38471 , n38469 , n38470 );
xnor ( n38472 , n38471 , n23550 );
and ( n38473 , n38467 , n38472 );
and ( n38474 , n38463 , n38472 );
or ( n38475 , n38468 , n38473 , n38474 );
and ( n38476 , n23573 , n28628 );
and ( n38477 , n23381 , n28626 );
nor ( n38478 , n38476 , n38477 );
xnor ( n38479 , n38478 , n28096 );
and ( n38480 , n38475 , n38479 );
xor ( n38481 , n38230 , n38234 );
xor ( n38482 , n38481 , n38239 );
and ( n38483 , n38479 , n38482 );
and ( n38484 , n38475 , n38482 );
or ( n38485 , n38480 , n38483 , n38484 );
and ( n38486 , n38462 , n38485 );
xor ( n38487 , n38242 , n38263 );
xor ( n38488 , n38487 , n38268 );
and ( n38489 , n38485 , n38488 );
and ( n38490 , n38462 , n38488 );
or ( n38491 , n38486 , n38489 , n38490 );
and ( n38492 , n23968 , n28628 );
and ( n38493 , n23573 , n28626 );
nor ( n38494 , n38492 , n38493 );
xnor ( n38495 , n38494 , n28096 );
and ( n38496 , n24621 , n27529 );
and ( n38497 , n24527 , n27527 );
nor ( n38498 , n38496 , n38497 );
xnor ( n38499 , n38498 , n27034 );
and ( n38500 , n38495 , n38499 );
and ( n38501 , n25284 , n26992 );
and ( n38502 , n24940 , n26990 );
nor ( n38503 , n38501 , n38502 );
xnor ( n38504 , n38503 , n26369 );
and ( n38505 , n38499 , n38504 );
and ( n38506 , n38495 , n38504 );
or ( n38507 , n38500 , n38505 , n38506 );
xor ( n38508 , n38332 , n38336 );
xor ( n38509 , n38508 , n38341 );
and ( n38510 , n38507 , n38509 );
xor ( n38511 , n38251 , n38255 );
xor ( n38512 , n38511 , n38260 );
and ( n38513 , n38509 , n38512 );
and ( n38514 , n38507 , n38512 );
or ( n38515 , n38510 , n38513 , n38514 );
xor ( n38516 , n38344 , n38348 );
xor ( n38517 , n38516 , n38353 );
and ( n38518 , n38515 , n38517 );
xor ( n38519 , n38360 , n38362 );
xor ( n38520 , n38519 , n38365 );
and ( n38521 , n38517 , n38520 );
and ( n38522 , n38515 , n38520 );
or ( n38523 , n38518 , n38521 , n38522 );
and ( n38524 , n38491 , n38523 );
xor ( n38525 , n38271 , n38273 );
xor ( n38526 , n38525 , n38276 );
and ( n38527 , n38523 , n38526 );
and ( n38528 , n38491 , n38526 );
or ( n38529 , n38524 , n38527 , n38528 );
and ( n38530 , n27751 , n24902 );
and ( n38531 , n27352 , n24900 );
nor ( n38532 , n38530 , n38531 );
xnor ( n38533 , n38532 , n24397 );
and ( n38534 , n28211 , n24376 );
and ( n38535 , n27757 , n24374 );
nor ( n38536 , n38534 , n38535 );
xnor ( n38537 , n38536 , n23927 );
and ( n38538 , n38533 , n38537 );
and ( n38539 , n38537 , n38297 );
and ( n38540 , n38533 , n38297 );
or ( n38541 , n38538 , n38539 , n38540 );
and ( n38542 , n29078 , n23641 );
and ( n38543 , n28700 , n23639 );
nor ( n38544 , n38542 , n38543 );
xnor ( n38545 , n38544 , n23213 );
and ( n38546 , n38541 , n38545 );
xor ( n38547 , n38291 , n38295 );
xor ( n38548 , n38547 , n38299 );
and ( n38549 , n38545 , n38548 );
and ( n38550 , n38541 , n38548 );
or ( n38551 , n38546 , n38549 , n38550 );
xor ( n38552 , n38302 , n38306 );
xor ( n38553 , n38552 , n38309 );
and ( n38554 , n38551 , n38553 );
xor ( n38555 , n38475 , n38479 );
xor ( n38556 , n38555 , n38482 );
and ( n38557 , n38553 , n38556 );
and ( n38558 , n38551 , n38556 );
or ( n38559 , n38554 , n38557 , n38558 );
xor ( n38560 , n38312 , n38314 );
xor ( n38561 , n38560 , n38317 );
and ( n38562 , n38559 , n38561 );
xor ( n38563 , n38462 , n38485 );
xor ( n38564 , n38563 , n38488 );
and ( n38565 , n38561 , n38564 );
and ( n38566 , n38559 , n38564 );
or ( n38567 , n38562 , n38565 , n38566 );
xor ( n38568 , n38320 , n38322 );
xor ( n38569 , n38568 , n38325 );
and ( n38570 , n38567 , n38569 );
xor ( n38571 , n38356 , n38368 );
xor ( n38572 , n38571 , n38371 );
and ( n38573 , n38569 , n38572 );
and ( n38574 , n38567 , n38572 );
or ( n38575 , n38570 , n38573 , n38574 );
and ( n38576 , n38529 , n38575 );
xor ( n38577 , n38402 , n38404 );
xor ( n38578 , n38577 , n38407 );
and ( n38579 , n38575 , n38578 );
and ( n38580 , n38529 , n38578 );
or ( n38581 , n38576 , n38579 , n38580 );
and ( n38582 , n38422 , n38581 );
xor ( n38583 , n38422 , n38581 );
xor ( n38584 , n38529 , n38575 );
xor ( n38585 , n38584 , n38578 );
and ( n38586 , n26319 , n26349 );
and ( n38587 , n25974 , n26347 );
nor ( n38588 , n38586 , n38587 );
xnor ( n38589 , n38588 , n25893 );
and ( n38590 , n26851 , n26027 );
and ( n38591 , n26422 , n26025 );
nor ( n38592 , n38590 , n38591 );
xnor ( n38593 , n38592 , n25499 );
and ( n38594 , n38589 , n38593 );
and ( n38595 , n25554 , n26992 );
and ( n38596 , n25284 , n26990 );
nor ( n38597 , n38595 , n38596 );
xnor ( n38598 , n38597 , n26369 );
and ( n38599 , n38594 , n38598 );
and ( n38600 , n28700 , n23944 );
and ( n38601 , n28810 , n23942 );
nor ( n38602 , n38600 , n38601 );
xnor ( n38603 , n38602 , n23550 );
and ( n38604 , n38598 , n38603 );
and ( n38605 , n38594 , n38603 );
or ( n38606 , n38599 , n38604 , n38605 );
and ( n38607 , n23381 , n29276 );
and ( n38608 , n23271 , n29274 );
nor ( n38609 , n38607 , n38608 );
xnor ( n38610 , n38609 , n28677 );
and ( n38611 , n38606 , n38610 );
xor ( n38612 , n38463 , n38467 );
xor ( n38613 , n38612 , n38472 );
and ( n38614 , n38610 , n38613 );
and ( n38615 , n38606 , n38613 );
or ( n38616 , n38611 , n38614 , n38615 );
and ( n38617 , n24527 , n28062 );
and ( n38618 , n24521 , n28060 );
nor ( n38619 , n38617 , n38618 );
xnor ( n38620 , n38619 , n27549 );
and ( n38621 , n24940 , n27529 );
and ( n38622 , n24621 , n27527 );
nor ( n38623 , n38621 , n38622 );
xnor ( n38624 , n38623 , n27034 );
and ( n38625 , n38620 , n38624 );
xor ( n38626 , n38426 , n38430 );
xor ( n38627 , n38626 , n38435 );
and ( n38628 , n38624 , n38627 );
and ( n38629 , n38620 , n38627 );
or ( n38630 , n38625 , n38628 , n38629 );
and ( n38631 , n23141 , n29977 );
and ( n38632 , n22916 , n29974 );
nor ( n38633 , n38631 , n38632 );
xnor ( n38634 , n38633 , n28674 );
and ( n38635 , n38630 , n38634 );
xor ( n38636 , n38495 , n38499 );
xor ( n38637 , n38636 , n38504 );
and ( n38638 , n38634 , n38637 );
and ( n38639 , n38630 , n38637 );
or ( n38640 , n38635 , n38638 , n38639 );
and ( n38641 , n38616 , n38640 );
xor ( n38642 , n38450 , n38454 );
xor ( n38643 , n38642 , n38459 );
and ( n38644 , n38640 , n38643 );
and ( n38645 , n38616 , n38643 );
or ( n38646 , n38641 , n38644 , n38645 );
and ( n38647 , n25765 , n26992 );
and ( n38648 , n25554 , n26990 );
nor ( n38649 , n38647 , n38648 );
xnor ( n38650 , n38649 , n26369 );
and ( n38651 , n27352 , n25383 );
and ( n38652 , n27135 , n25381 );
nor ( n38653 , n38651 , n38652 );
xnor ( n38654 , n38653 , n24885 );
and ( n38655 , n38650 , n38654 );
and ( n38656 , n27757 , n24902 );
and ( n38657 , n27751 , n24900 );
nor ( n38658 , n38656 , n38657 );
xnor ( n38659 , n38658 , n24397 );
and ( n38660 , n38654 , n38659 );
and ( n38661 , n38650 , n38659 );
or ( n38662 , n38655 , n38660 , n38661 );
and ( n38663 , n24131 , n28628 );
and ( n38664 , n23968 , n28626 );
nor ( n38665 , n38663 , n38664 );
xnor ( n38666 , n38665 , n28096 );
and ( n38667 , n38662 , n38666 );
and ( n38668 , n29318 , n23641 );
and ( n38669 , n29078 , n23639 );
nor ( n38670 , n38668 , n38669 );
xnor ( n38671 , n38670 , n23213 );
and ( n38672 , n38666 , n38671 );
and ( n38673 , n38662 , n38671 );
or ( n38674 , n38667 , n38672 , n38673 );
xor ( n38675 , n38438 , n38442 );
xor ( n38676 , n38675 , n38447 );
and ( n38677 , n38674 , n38676 );
xor ( n38678 , n38541 , n38545 );
xor ( n38679 , n38678 , n38548 );
and ( n38680 , n38676 , n38679 );
and ( n38681 , n38674 , n38679 );
or ( n38682 , n38677 , n38680 , n38681 );
xor ( n38683 , n38507 , n38509 );
xor ( n38684 , n38683 , n38512 );
and ( n38685 , n38682 , n38684 );
xor ( n38686 , n38551 , n38553 );
xor ( n38687 , n38686 , n38556 );
and ( n38688 , n38684 , n38687 );
and ( n38689 , n38682 , n38687 );
or ( n38690 , n38685 , n38688 , n38689 );
and ( n38691 , n38646 , n38690 );
xor ( n38692 , n38515 , n38517 );
xor ( n38693 , n38692 , n38520 );
and ( n38694 , n38690 , n38693 );
and ( n38695 , n38646 , n38693 );
or ( n38696 , n38691 , n38694 , n38695 );
xor ( n38697 , n38491 , n38523 );
xor ( n38698 , n38697 , n38526 );
and ( n38699 , n38696 , n38698 );
xor ( n38700 , n38567 , n38569 );
xor ( n38701 , n38700 , n38572 );
and ( n38702 , n38698 , n38701 );
and ( n38703 , n38696 , n38701 );
or ( n38704 , n38699 , n38702 , n38703 );
and ( n38705 , n38585 , n38704 );
xor ( n38706 , n38585 , n38704 );
xor ( n38707 , n38696 , n38698 );
xor ( n38708 , n38707 , n38701 );
xor ( n38709 , n38589 , n38593 );
and ( n38710 , n28810 , n24376 );
and ( n38711 , n28211 , n24374 );
nor ( n38712 , n38710 , n38711 );
xnor ( n38713 , n38712 , n23927 );
and ( n38714 , n38709 , n38713 );
and ( n38715 , n29078 , n23944 );
and ( n38716 , n28700 , n23942 );
nor ( n38717 , n38715 , n38716 );
xnor ( n38718 , n38717 , n23550 );
and ( n38719 , n38713 , n38718 );
and ( n38720 , n38709 , n38718 );
or ( n38721 , n38714 , n38719 , n38720 );
and ( n38722 , n23573 , n29276 );
and ( n38723 , n23381 , n29274 );
nor ( n38724 , n38722 , n38723 );
xnor ( n38725 , n38724 , n28677 );
and ( n38726 , n38721 , n38725 );
xor ( n38727 , n38594 , n38598 );
xor ( n38728 , n38727 , n38603 );
and ( n38729 , n38725 , n38728 );
and ( n38730 , n38721 , n38728 );
or ( n38731 , n38726 , n38729 , n38730 );
and ( n38732 , n25974 , n26992 );
and ( n38733 , n25765 , n26990 );
nor ( n38734 , n38732 , n38733 );
xnor ( n38735 , n38734 , n26369 );
and ( n38736 , n26422 , n26349 );
and ( n38737 , n26319 , n26347 );
nor ( n38738 , n38736 , n38737 );
xnor ( n38739 , n38738 , n25893 );
and ( n38740 , n38735 , n38739 );
and ( n38741 , n27135 , n26027 );
and ( n38742 , n26851 , n26025 );
nor ( n38743 , n38741 , n38742 );
xnor ( n38744 , n38743 , n25499 );
and ( n38745 , n38739 , n38744 );
and ( n38746 , n38735 , n38744 );
or ( n38747 , n38740 , n38745 , n38746 );
and ( n38748 , n24621 , n28062 );
and ( n38749 , n24527 , n28060 );
nor ( n38750 , n38748 , n38749 );
xnor ( n38751 , n38750 , n27549 );
and ( n38752 , n38747 , n38751 );
and ( n38753 , n29623 , n23639 );
not ( n38754 , n38753 );
and ( n38755 , n38754 , n23213 );
and ( n38756 , n38751 , n38755 );
and ( n38757 , n38747 , n38755 );
or ( n38758 , n38752 , n38756 , n38757 );
and ( n38759 , n23271 , n29977 );
and ( n38760 , n23141 , n29974 );
nor ( n38761 , n38759 , n38760 );
xnor ( n38762 , n38761 , n28674 );
and ( n38763 , n38758 , n38762 );
xor ( n38764 , n38533 , n38537 );
xor ( n38765 , n38764 , n38297 );
and ( n38766 , n38762 , n38765 );
and ( n38767 , n38758 , n38765 );
or ( n38768 , n38763 , n38766 , n38767 );
and ( n38769 , n38731 , n38768 );
xor ( n38770 , n38606 , n38610 );
xor ( n38771 , n38770 , n38613 );
and ( n38772 , n38768 , n38771 );
and ( n38773 , n38731 , n38771 );
or ( n38774 , n38769 , n38772 , n38773 );
and ( n38775 , n24521 , n28628 );
and ( n38776 , n24131 , n28626 );
nor ( n38777 , n38775 , n38776 );
xnor ( n38778 , n38777 , n28096 );
and ( n38779 , n25284 , n27529 );
and ( n38780 , n24940 , n27527 );
nor ( n38781 , n38779 , n38780 );
xnor ( n38782 , n38781 , n27034 );
and ( n38783 , n38778 , n38782 );
and ( n38784 , n29623 , n23641 );
and ( n38785 , n29318 , n23639 );
nor ( n38786 , n38784 , n38785 );
xnor ( n38787 , n38786 , n23213 );
and ( n38788 , n38782 , n38787 );
and ( n38789 , n38778 , n38787 );
or ( n38790 , n38783 , n38788 , n38789 );
and ( n38791 , n28700 , n24376 );
and ( n38792 , n28810 , n24374 );
nor ( n38793 , n38791 , n38792 );
xnor ( n38794 , n38793 , n23927 );
and ( n38795 , n29318 , n23944 );
and ( n38796 , n29078 , n23942 );
nor ( n38797 , n38795 , n38796 );
xnor ( n38798 , n38797 , n23550 );
and ( n38799 , n38794 , n38798 );
and ( n38800 , n38798 , n38753 );
and ( n38801 , n38794 , n38753 );
or ( n38802 , n38799 , n38800 , n38801 );
and ( n38803 , n26851 , n26349 );
and ( n38804 , n26422 , n26347 );
nor ( n38805 , n38803 , n38804 );
xnor ( n38806 , n38805 , n25893 );
and ( n38807 , n27352 , n26027 );
and ( n38808 , n27135 , n26025 );
nor ( n38809 , n38807 , n38808 );
xnor ( n38810 , n38809 , n25499 );
and ( n38811 , n38806 , n38810 );
and ( n38812 , n27751 , n25383 );
and ( n38813 , n27352 , n25381 );
nor ( n38814 , n38812 , n38813 );
xnor ( n38815 , n38814 , n24885 );
and ( n38816 , n38811 , n38815 );
and ( n38817 , n28211 , n24902 );
and ( n38818 , n27757 , n24900 );
nor ( n38819 , n38817 , n38818 );
xnor ( n38820 , n38819 , n24397 );
and ( n38821 , n38815 , n38820 );
and ( n38822 , n38811 , n38820 );
or ( n38823 , n38816 , n38821 , n38822 );
and ( n38824 , n38802 , n38823 );
and ( n38825 , n23968 , n29276 );
and ( n38826 , n23573 , n29274 );
nor ( n38827 , n38825 , n38826 );
xnor ( n38828 , n38827 , n28677 );
and ( n38829 , n38823 , n38828 );
and ( n38830 , n38802 , n38828 );
or ( n38831 , n38824 , n38829 , n38830 );
and ( n38832 , n38790 , n38831 );
xor ( n38833 , n38662 , n38666 );
xor ( n38834 , n38833 , n38671 );
and ( n38835 , n38831 , n38834 );
and ( n38836 , n38790 , n38834 );
or ( n38837 , n38832 , n38835 , n38836 );
xor ( n38838 , n38630 , n38634 );
xor ( n38839 , n38838 , n38637 );
and ( n38840 , n38837 , n38839 );
xor ( n38841 , n38674 , n38676 );
xor ( n38842 , n38841 , n38679 );
and ( n38843 , n38839 , n38842 );
and ( n38844 , n38837 , n38842 );
or ( n38845 , n38840 , n38843 , n38844 );
and ( n38846 , n38774 , n38845 );
xor ( n38847 , n38616 , n38640 );
xor ( n38848 , n38847 , n38643 );
and ( n38849 , n38845 , n38848 );
and ( n38850 , n38774 , n38848 );
or ( n38851 , n38846 , n38849 , n38850 );
xor ( n38852 , n38559 , n38561 );
xor ( n38853 , n38852 , n38564 );
and ( n38854 , n38851 , n38853 );
xor ( n38855 , n38646 , n38690 );
xor ( n38856 , n38855 , n38693 );
and ( n38857 , n38853 , n38856 );
and ( n38858 , n38851 , n38856 );
or ( n38859 , n38854 , n38857 , n38858 );
and ( n38860 , n38708 , n38859 );
xor ( n38861 , n38708 , n38859 );
xor ( n38862 , n38851 , n38853 );
xor ( n38863 , n38862 , n38856 );
and ( n38864 , n24131 , n29276 );
and ( n38865 , n23968 , n29274 );
nor ( n38866 , n38864 , n38865 );
xnor ( n38867 , n38866 , n28677 );
and ( n38868 , n24527 , n28628 );
and ( n38869 , n24521 , n28626 );
nor ( n38870 , n38868 , n38869 );
xnor ( n38871 , n38870 , n28096 );
and ( n38872 , n38867 , n38871 );
and ( n38873 , n24940 , n28062 );
and ( n38874 , n24621 , n28060 );
nor ( n38875 , n38873 , n38874 );
xnor ( n38876 , n38875 , n27549 );
and ( n38877 , n38871 , n38876 );
and ( n38878 , n38867 , n38876 );
or ( n38879 , n38872 , n38877 , n38878 );
and ( n38880 , n23381 , n29977 );
and ( n38881 , n23271 , n29974 );
nor ( n38882 , n38880 , n38881 );
xnor ( n38883 , n38882 , n28674 );
and ( n38884 , n38879 , n38883 );
xor ( n38885 , n38747 , n38751 );
xor ( n38886 , n38885 , n38755 );
and ( n38887 , n38883 , n38886 );
and ( n38888 , n38879 , n38886 );
or ( n38889 , n38884 , n38887 , n38888 );
xor ( n38890 , n38806 , n38810 );
and ( n38891 , n26319 , n26992 );
and ( n38892 , n25974 , n26990 );
nor ( n38893 , n38891 , n38892 );
xnor ( n38894 , n38893 , n26369 );
and ( n38895 , n38890 , n38894 );
and ( n38896 , n29623 , n23942 );
not ( n38897 , n38896 );
and ( n38898 , n38897 , n23550 );
and ( n38899 , n38894 , n38898 );
and ( n38900 , n38890 , n38898 );
or ( n38901 , n38895 , n38899 , n38900 );
and ( n38902 , n25554 , n27529 );
and ( n38903 , n25284 , n27527 );
nor ( n38904 , n38902 , n38903 );
xnor ( n38905 , n38904 , n27034 );
and ( n38906 , n38901 , n38905 );
xor ( n38907 , n38735 , n38739 );
xor ( n38908 , n38907 , n38744 );
and ( n38909 , n38905 , n38908 );
and ( n38910 , n38901 , n38908 );
or ( n38911 , n38906 , n38909 , n38910 );
xor ( n38912 , n38650 , n38654 );
xor ( n38913 , n38912 , n38659 );
and ( n38914 , n38911 , n38913 );
xor ( n38915 , n38709 , n38713 );
xor ( n38916 , n38915 , n38718 );
and ( n38917 , n38913 , n38916 );
and ( n38918 , n38911 , n38916 );
or ( n38919 , n38914 , n38917 , n38918 );
and ( n38920 , n38889 , n38919 );
xor ( n38921 , n38620 , n38624 );
xor ( n38922 , n38921 , n38627 );
and ( n38923 , n38919 , n38922 );
and ( n38924 , n38889 , n38922 );
or ( n38925 , n38920 , n38923 , n38924 );
xor ( n38926 , n38721 , n38725 );
xor ( n38927 , n38926 , n38728 );
xor ( n38928 , n38758 , n38762 );
xor ( n38929 , n38928 , n38765 );
and ( n38930 , n38927 , n38929 );
xor ( n38931 , n38790 , n38831 );
xor ( n38932 , n38931 , n38834 );
and ( n38933 , n38929 , n38932 );
and ( n38934 , n38927 , n38932 );
or ( n38935 , n38930 , n38933 , n38934 );
and ( n38936 , n38925 , n38935 );
xor ( n38937 , n38731 , n38768 );
xor ( n38938 , n38937 , n38771 );
and ( n38939 , n38935 , n38938 );
and ( n38940 , n38925 , n38938 );
or ( n38941 , n38936 , n38939 , n38940 );
xor ( n38942 , n38774 , n38845 );
xor ( n38943 , n38942 , n38848 );
and ( n38944 , n38941 , n38943 );
xor ( n38945 , n38682 , n38684 );
xor ( n38946 , n38945 , n38687 );
and ( n38947 , n38943 , n38946 );
and ( n38948 , n38941 , n38946 );
or ( n38949 , n38944 , n38947 , n38948 );
and ( n38950 , n38863 , n38949 );
xor ( n38951 , n38863 , n38949 );
xor ( n38952 , n38941 , n38943 );
xor ( n38953 , n38952 , n38946 );
and ( n38954 , n25765 , n27529 );
and ( n38955 , n25554 , n27527 );
nor ( n38956 , n38954 , n38955 );
xnor ( n38957 , n38956 , n27034 );
and ( n38958 , n27757 , n25383 );
and ( n38959 , n27751 , n25381 );
nor ( n38960 , n38958 , n38959 );
xnor ( n38961 , n38960 , n24885 );
and ( n38962 , n38957 , n38961 );
and ( n38963 , n29078 , n24376 );
and ( n38964 , n28700 , n24374 );
nor ( n38965 , n38963 , n38964 );
xnor ( n38966 , n38965 , n23927 );
and ( n38967 , n38961 , n38966 );
and ( n38968 , n38957 , n38966 );
or ( n38969 , n38962 , n38967 , n38968 );
and ( n38970 , n26422 , n26992 );
and ( n38971 , n26319 , n26990 );
nor ( n38972 , n38970 , n38971 );
xnor ( n38973 , n38972 , n26369 );
and ( n38974 , n27135 , n26349 );
and ( n38975 , n26851 , n26347 );
nor ( n38976 , n38974 , n38975 );
xnor ( n38977 , n38976 , n25893 );
and ( n38978 , n38973 , n38977 );
and ( n38979 , n27751 , n26027 );
and ( n38980 , n27352 , n26025 );
nor ( n38981 , n38979 , n38980 );
xnor ( n38982 , n38981 , n25499 );
and ( n38983 , n38977 , n38982 );
and ( n38984 , n38973 , n38982 );
or ( n38985 , n38978 , n38983 , n38984 );
and ( n38986 , n28810 , n24902 );
and ( n38987 , n28211 , n24900 );
nor ( n38988 , n38986 , n38987 );
xnor ( n38989 , n38988 , n24397 );
and ( n38990 , n38985 , n38989 );
and ( n38991 , n29623 , n23944 );
and ( n38992 , n29318 , n23942 );
nor ( n38993 , n38991 , n38992 );
xnor ( n38994 , n38993 , n23550 );
and ( n38995 , n38989 , n38994 );
and ( n38996 , n38985 , n38994 );
or ( n38997 , n38990 , n38995 , n38996 );
and ( n38998 , n38969 , n38997 );
xor ( n38999 , n38811 , n38815 );
xor ( n39000 , n38999 , n38820 );
and ( n39001 , n38997 , n39000 );
and ( n39002 , n38969 , n39000 );
or ( n39003 , n38998 , n39001 , n39002 );
xor ( n39004 , n38778 , n38782 );
xor ( n39005 , n39004 , n38787 );
and ( n39006 , n39003 , n39005 );
xor ( n39007 , n38802 , n38823 );
xor ( n39008 , n39007 , n38828 );
and ( n39009 , n39005 , n39008 );
and ( n39010 , n39003 , n39008 );
or ( n39011 , n39006 , n39009 , n39010 );
and ( n39012 , n23573 , n29977 );
and ( n39013 , n23381 , n29974 );
nor ( n39014 , n39012 , n39013 );
xnor ( n39015 , n39014 , n28674 );
xor ( n39016 , n38794 , n38798 );
xor ( n39017 , n39016 , n38753 );
and ( n39018 , n39015 , n39017 );
xor ( n39019 , n38901 , n38905 );
xor ( n39020 , n39019 , n38908 );
and ( n39021 , n39017 , n39020 );
and ( n39022 , n39015 , n39020 );
or ( n39023 , n39018 , n39021 , n39022 );
xor ( n39024 , n38879 , n38883 );
xor ( n39025 , n39024 , n38886 );
and ( n39026 , n39023 , n39025 );
xor ( n39027 , n38911 , n38913 );
xor ( n39028 , n39027 , n38916 );
and ( n39029 , n39025 , n39028 );
and ( n39030 , n39023 , n39028 );
or ( n39031 , n39026 , n39029 , n39030 );
and ( n39032 , n39011 , n39031 );
xor ( n39033 , n38889 , n38919 );
xor ( n39034 , n39033 , n38922 );
and ( n39035 , n39031 , n39034 );
and ( n39036 , n39011 , n39034 );
or ( n39037 , n39032 , n39035 , n39036 );
xor ( n39038 , n38837 , n38839 );
xor ( n39039 , n39038 , n38842 );
and ( n39040 , n39037 , n39039 );
xor ( n39041 , n38925 , n38935 );
xor ( n39042 , n39041 , n38938 );
and ( n39043 , n39039 , n39042 );
and ( n39044 , n39037 , n39042 );
or ( n39045 , n39040 , n39043 , n39044 );
and ( n39046 , n38953 , n39045 );
xor ( n39047 , n38953 , n39045 );
xor ( n39048 , n39037 , n39039 );
xor ( n39049 , n39048 , n39042 );
and ( n39050 , n26851 , n26992 );
and ( n39051 , n26422 , n26990 );
nor ( n39052 , n39050 , n39051 );
xnor ( n39053 , n39052 , n26369 );
and ( n39054 , n27352 , n26349 );
and ( n39055 , n27135 , n26347 );
nor ( n39056 , n39054 , n39055 );
xnor ( n39057 , n39056 , n25893 );
and ( n39058 , n39053 , n39057 );
and ( n39059 , n25974 , n27529 );
and ( n39060 , n25765 , n27527 );
nor ( n39061 , n39059 , n39060 );
xnor ( n39062 , n39061 , n27034 );
and ( n39063 , n39058 , n39062 );
and ( n39064 , n39062 , n38896 );
and ( n39065 , n39058 , n38896 );
or ( n39066 , n39063 , n39064 , n39065 );
and ( n39067 , n23968 , n29977 );
and ( n39068 , n23573 , n29974 );
nor ( n39069 , n39067 , n39068 );
xnor ( n39070 , n39069 , n28674 );
and ( n39071 , n39066 , n39070 );
and ( n39072 , n25284 , n28062 );
and ( n39073 , n24940 , n28060 );
nor ( n39074 , n39072 , n39073 );
xnor ( n39075 , n39074 , n27549 );
and ( n39076 , n39070 , n39075 );
and ( n39077 , n39066 , n39075 );
or ( n39078 , n39071 , n39076 , n39077 );
and ( n39079 , n24521 , n29276 );
and ( n39080 , n24131 , n29274 );
nor ( n39081 , n39079 , n39080 );
xnor ( n39082 , n39081 , n28677 );
and ( n39083 , n24621 , n28628 );
and ( n39084 , n24527 , n28626 );
nor ( n39085 , n39083 , n39084 );
xnor ( n39086 , n39085 , n28096 );
and ( n39087 , n39082 , n39086 );
xor ( n39088 , n38890 , n38894 );
xor ( n39089 , n39088 , n38898 );
and ( n39090 , n39086 , n39089 );
and ( n39091 , n39082 , n39089 );
or ( n39092 , n39087 , n39090 , n39091 );
and ( n39093 , n39078 , n39092 );
xor ( n39094 , n38867 , n38871 );
xor ( n39095 , n39094 , n38876 );
and ( n39096 , n39092 , n39095 );
and ( n39097 , n39078 , n39095 );
or ( n39098 , n39093 , n39096 , n39097 );
and ( n39099 , n28211 , n25383 );
and ( n39100 , n27757 , n25381 );
nor ( n39101 , n39099 , n39100 );
xnor ( n39102 , n39101 , n24885 );
and ( n39103 , n28700 , n24902 );
and ( n39104 , n28810 , n24900 );
nor ( n39105 , n39103 , n39104 );
xnor ( n39106 , n39105 , n24397 );
and ( n39107 , n39102 , n39106 );
xor ( n39108 , n38973 , n38977 );
xor ( n39109 , n39108 , n38982 );
and ( n39110 , n39106 , n39109 );
and ( n39111 , n39102 , n39109 );
or ( n39112 , n39107 , n39110 , n39111 );
xor ( n39113 , n38957 , n38961 );
xor ( n39114 , n39113 , n38966 );
and ( n39115 , n39112 , n39114 );
xor ( n39116 , n38985 , n38989 );
xor ( n39117 , n39116 , n38994 );
and ( n39118 , n39114 , n39117 );
and ( n39119 , n39112 , n39117 );
or ( n39120 , n39115 , n39118 , n39119 );
xor ( n39121 , n38969 , n38997 );
xor ( n39122 , n39121 , n39000 );
and ( n39123 , n39120 , n39122 );
xor ( n39124 , n39015 , n39017 );
xor ( n39125 , n39124 , n39020 );
and ( n39126 , n39122 , n39125 );
and ( n39127 , n39120 , n39125 );
or ( n39128 , n39123 , n39126 , n39127 );
and ( n39129 , n39098 , n39128 );
xor ( n39130 , n39003 , n39005 );
xor ( n39131 , n39130 , n39008 );
and ( n39132 , n39128 , n39131 );
and ( n39133 , n39098 , n39131 );
or ( n39134 , n39129 , n39132 , n39133 );
xor ( n39135 , n38927 , n38929 );
xor ( n39136 , n39135 , n38932 );
and ( n39137 , n39134 , n39136 );
xor ( n39138 , n39011 , n39031 );
xor ( n39139 , n39138 , n39034 );
and ( n39140 , n39136 , n39139 );
and ( n39141 , n39134 , n39139 );
or ( n39142 , n39137 , n39140 , n39141 );
and ( n39143 , n39049 , n39142 );
xor ( n39144 , n39049 , n39142 );
xor ( n39145 , n39134 , n39136 );
xor ( n39146 , n39145 , n39139 );
xor ( n39147 , n39053 , n39057 );
and ( n39148 , n27757 , n26027 );
and ( n39149 , n27751 , n26025 );
nor ( n39150 , n39148 , n39149 );
xnor ( n39151 , n39150 , n25499 );
and ( n39152 , n39147 , n39151 );
and ( n39153 , n29623 , n24374 );
not ( n39154 , n39153 );
and ( n39155 , n39154 , n23927 );
and ( n39156 , n39151 , n39155 );
and ( n39157 , n39147 , n39155 );
or ( n39158 , n39152 , n39156 , n39157 );
and ( n39159 , n25554 , n28062 );
and ( n39160 , n25284 , n28060 );
nor ( n39161 , n39159 , n39160 );
xnor ( n39162 , n39161 , n27549 );
and ( n39163 , n39158 , n39162 );
and ( n39164 , n29318 , n24376 );
and ( n39165 , n29078 , n24374 );
nor ( n39166 , n39164 , n39165 );
xnor ( n39167 , n39166 , n23927 );
and ( n39168 , n39162 , n39167 );
and ( n39169 , n39158 , n39167 );
or ( n39170 , n39163 , n39168 , n39169 );
and ( n39171 , n25765 , n28062 );
and ( n39172 , n25554 , n28060 );
nor ( n39173 , n39171 , n39172 );
xnor ( n39174 , n39173 , n27549 );
and ( n39175 , n26319 , n27529 );
and ( n39176 , n25974 , n27527 );
nor ( n39177 , n39175 , n39176 );
xnor ( n39178 , n39177 , n27034 );
and ( n39179 , n39174 , n39178 );
and ( n39180 , n28810 , n25383 );
and ( n39181 , n28211 , n25381 );
nor ( n39182 , n39180 , n39181 );
xnor ( n39183 , n39182 , n24885 );
and ( n39184 , n39178 , n39183 );
and ( n39185 , n39174 , n39183 );
or ( n39186 , n39179 , n39184 , n39185 );
and ( n39187 , n24527 , n29276 );
and ( n39188 , n24521 , n29274 );
nor ( n39189 , n39187 , n39188 );
xnor ( n39190 , n39189 , n28677 );
and ( n39191 , n39186 , n39190 );
xor ( n39192 , n39058 , n39062 );
xor ( n39193 , n39192 , n38896 );
and ( n39194 , n39190 , n39193 );
and ( n39195 , n39186 , n39193 );
or ( n39196 , n39191 , n39194 , n39195 );
and ( n39197 , n39170 , n39196 );
xor ( n39198 , n39082 , n39086 );
xor ( n39199 , n39198 , n39089 );
and ( n39200 , n39196 , n39199 );
and ( n39201 , n39170 , n39199 );
or ( n39202 , n39197 , n39200 , n39201 );
and ( n39203 , n27135 , n26992 );
and ( n39204 , n26851 , n26990 );
nor ( n39205 , n39203 , n39204 );
xnor ( n39206 , n39205 , n26369 );
and ( n39207 , n27751 , n26349 );
and ( n39208 , n27352 , n26347 );
nor ( n39209 , n39207 , n39208 );
xnor ( n39210 , n39209 , n25893 );
and ( n39211 , n39206 , n39210 );
and ( n39212 , n28211 , n26027 );
and ( n39213 , n27757 , n26025 );
nor ( n39214 , n39212 , n39213 );
xnor ( n39215 , n39214 , n25499 );
and ( n39216 , n39210 , n39215 );
and ( n39217 , n39206 , n39215 );
or ( n39218 , n39211 , n39216 , n39217 );
and ( n39219 , n29078 , n24902 );
and ( n39220 , n28700 , n24900 );
nor ( n39221 , n39219 , n39220 );
xnor ( n39222 , n39221 , n24397 );
and ( n39223 , n39218 , n39222 );
and ( n39224 , n29623 , n24376 );
and ( n39225 , n29318 , n24374 );
nor ( n39226 , n39224 , n39225 );
xnor ( n39227 , n39226 , n23927 );
and ( n39228 , n39222 , n39227 );
and ( n39229 , n39218 , n39227 );
or ( n39230 , n39223 , n39228 , n39229 );
and ( n39231 , n24131 , n29977 );
and ( n39232 , n23968 , n29974 );
nor ( n39233 , n39231 , n39232 );
xnor ( n39234 , n39233 , n28674 );
and ( n39235 , n39230 , n39234 );
and ( n39236 , n24940 , n28628 );
and ( n39237 , n24621 , n28626 );
nor ( n39238 , n39236 , n39237 );
xnor ( n39239 , n39238 , n28096 );
and ( n39240 , n39234 , n39239 );
and ( n39241 , n39230 , n39239 );
or ( n39242 , n39235 , n39240 , n39241 );
xor ( n39243 , n39066 , n39070 );
xor ( n39244 , n39243 , n39075 );
and ( n39245 , n39242 , n39244 );
xor ( n39246 , n39112 , n39114 );
xor ( n39247 , n39246 , n39117 );
and ( n39248 , n39244 , n39247 );
and ( n39249 , n39242 , n39247 );
or ( n39250 , n39245 , n39248 , n39249 );
and ( n39251 , n39202 , n39250 );
xor ( n39252 , n39078 , n39092 );
xor ( n39253 , n39252 , n39095 );
and ( n39254 , n39250 , n39253 );
and ( n39255 , n39202 , n39253 );
or ( n39256 , n39251 , n39254 , n39255 );
xor ( n39257 , n39023 , n39025 );
xor ( n39258 , n39257 , n39028 );
and ( n39259 , n39256 , n39258 );
xor ( n39260 , n39098 , n39128 );
xor ( n39261 , n39260 , n39131 );
and ( n39262 , n39258 , n39261 );
and ( n39263 , n39256 , n39261 );
or ( n39264 , n39259 , n39262 , n39263 );
and ( n39265 , n39146 , n39264 );
xor ( n39266 , n39146 , n39264 );
and ( n39267 , n28700 , n25383 );
and ( n39268 , n28810 , n25381 );
nor ( n39269 , n39267 , n39268 );
xnor ( n39270 , n39269 , n24885 );
and ( n39271 , n39270 , n39153 );
xor ( n39272 , n39206 , n39210 );
xor ( n39273 , n39272 , n39215 );
and ( n39274 , n39153 , n39273 );
and ( n39275 , n39270 , n39273 );
or ( n39276 , n39271 , n39274 , n39275 );
and ( n39277 , n24521 , n29977 );
and ( n39278 , n24131 , n29974 );
nor ( n39279 , n39277 , n39278 );
xnor ( n39280 , n39279 , n28674 );
and ( n39281 , n39276 , n39280 );
and ( n39282 , n25284 , n28628 );
and ( n39283 , n24940 , n28626 );
nor ( n39284 , n39282 , n39283 );
xnor ( n39285 , n39284 , n28096 );
and ( n39286 , n39280 , n39285 );
and ( n39287 , n39276 , n39285 );
or ( n39288 , n39281 , n39286 , n39287 );
xor ( n39289 , n39158 , n39162 );
xor ( n39290 , n39289 , n39167 );
and ( n39291 , n39288 , n39290 );
xor ( n39292 , n39102 , n39106 );
xor ( n39293 , n39292 , n39109 );
and ( n39294 , n39290 , n39293 );
and ( n39295 , n39288 , n39293 );
or ( n39296 , n39291 , n39294 , n39295 );
and ( n39297 , n26851 , n27529 );
and ( n39298 , n26422 , n27527 );
nor ( n39299 , n39297 , n39298 );
xnor ( n39300 , n39299 , n27034 );
and ( n39301 , n27352 , n26992 );
and ( n39302 , n27135 , n26990 );
nor ( n39303 , n39301 , n39302 );
xnor ( n39304 , n39303 , n26369 );
and ( n39305 , n39300 , n39304 );
and ( n39306 , n25974 , n28062 );
and ( n39307 , n25765 , n28060 );
nor ( n39308 , n39306 , n39307 );
xnor ( n39309 , n39308 , n27549 );
and ( n39310 , n39305 , n39309 );
and ( n39311 , n26422 , n27529 );
and ( n39312 , n26319 , n27527 );
nor ( n39313 , n39311 , n39312 );
xnor ( n39314 , n39313 , n27034 );
and ( n39315 , n39309 , n39314 );
and ( n39316 , n39305 , n39314 );
or ( n39317 , n39310 , n39315 , n39316 );
and ( n39318 , n24621 , n29276 );
and ( n39319 , n24527 , n29274 );
nor ( n39320 , n39318 , n39319 );
xnor ( n39321 , n39320 , n28677 );
and ( n39322 , n39317 , n39321 );
xor ( n39323 , n39147 , n39151 );
xor ( n39324 , n39323 , n39155 );
and ( n39325 , n39321 , n39324 );
and ( n39326 , n39317 , n39324 );
or ( n39327 , n39322 , n39325 , n39326 );
xor ( n39328 , n39230 , n39234 );
xor ( n39329 , n39328 , n39239 );
and ( n39330 , n39327 , n39329 );
xor ( n39331 , n39186 , n39190 );
xor ( n39332 , n39331 , n39193 );
and ( n39333 , n39329 , n39332 );
and ( n39334 , n39327 , n39332 );
or ( n39335 , n39330 , n39333 , n39334 );
and ( n39336 , n39296 , n39335 );
xor ( n39337 , n39170 , n39196 );
xor ( n39338 , n39337 , n39199 );
and ( n39339 , n39335 , n39338 );
and ( n39340 , n39296 , n39338 );
or ( n39341 , n39336 , n39339 , n39340 );
xor ( n39342 , n39202 , n39250 );
xor ( n39343 , n39342 , n39253 );
and ( n39344 , n39341 , n39343 );
xor ( n39345 , n39120 , n39122 );
xor ( n39346 , n39345 , n39125 );
and ( n39347 , n39343 , n39346 );
and ( n39348 , n39341 , n39346 );
or ( n39349 , n39344 , n39347 , n39348 );
xor ( n39350 , n39256 , n39258 );
xor ( n39351 , n39350 , n39261 );
and ( n39352 , n39349 , n39351 );
xor ( n39353 , n39349 , n39351 );
xor ( n39354 , n39341 , n39343 );
xor ( n39355 , n39354 , n39346 );
xor ( n39356 , n39300 , n39304 );
and ( n39357 , n27757 , n26349 );
and ( n39358 , n27751 , n26347 );
nor ( n39359 , n39357 , n39358 );
xnor ( n39360 , n39359 , n25893 );
and ( n39361 , n39356 , n39360 );
and ( n39362 , n28810 , n26027 );
and ( n39363 , n28211 , n26025 );
nor ( n39364 , n39362 , n39363 );
xnor ( n39365 , n39364 , n25499 );
and ( n39366 , n39360 , n39365 );
and ( n39367 , n39356 , n39365 );
or ( n39368 , n39361 , n39366 , n39367 );
and ( n39369 , n29318 , n24902 );
and ( n39370 , n29078 , n24900 );
nor ( n39371 , n39369 , n39370 );
xnor ( n39372 , n39371 , n24397 );
and ( n39373 , n39368 , n39372 );
xor ( n39374 , n39305 , n39309 );
xor ( n39375 , n39374 , n39314 );
and ( n39376 , n39372 , n39375 );
and ( n39377 , n39368 , n39375 );
or ( n39378 , n39373 , n39376 , n39377 );
xor ( n39379 , n39174 , n39178 );
xor ( n39380 , n39379 , n39183 );
and ( n39381 , n39378 , n39380 );
xor ( n39382 , n39218 , n39222 );
xor ( n39383 , n39382 , n39227 );
and ( n39384 , n39380 , n39383 );
and ( n39385 , n39378 , n39383 );
or ( n39386 , n39381 , n39384 , n39385 );
and ( n39387 , n27135 , n27529 );
and ( n39388 , n26851 , n27527 );
nor ( n39389 , n39387 , n39388 );
xnor ( n39390 , n39389 , n27034 );
and ( n39391 , n27751 , n26992 );
and ( n39392 , n27352 , n26990 );
nor ( n39393 , n39391 , n39392 );
xnor ( n39394 , n39393 , n26369 );
and ( n39395 , n39390 , n39394 );
and ( n39396 , n28211 , n26349 );
and ( n39397 , n27757 , n26347 );
nor ( n39398 , n39396 , n39397 );
xnor ( n39399 , n39398 , n25893 );
and ( n39400 , n39394 , n39399 );
and ( n39401 , n39390 , n39399 );
or ( n39402 , n39395 , n39400 , n39401 );
and ( n39403 , n26319 , n28062 );
and ( n39404 , n25974 , n28060 );
nor ( n39405 , n39403 , n39404 );
xnor ( n39406 , n39405 , n27549 );
and ( n39407 , n39402 , n39406 );
and ( n39408 , n29623 , n24900 );
not ( n39409 , n39408 );
and ( n39410 , n39409 , n24397 );
and ( n39411 , n39406 , n39410 );
and ( n39412 , n39402 , n39410 );
or ( n39413 , n39407 , n39411 , n39412 );
and ( n39414 , n24940 , n29276 );
and ( n39415 , n24621 , n29274 );
nor ( n39416 , n39414 , n39415 );
xnor ( n39417 , n39416 , n28677 );
and ( n39418 , n39413 , n39417 );
and ( n39419 , n25554 , n28628 );
and ( n39420 , n25284 , n28626 );
nor ( n39421 , n39419 , n39420 );
xnor ( n39422 , n39421 , n28096 );
and ( n39423 , n39417 , n39422 );
and ( n39424 , n39413 , n39422 );
or ( n39425 , n39418 , n39423 , n39424 );
and ( n39426 , n25765 , n28628 );
and ( n39427 , n25554 , n28626 );
nor ( n39428 , n39426 , n39427 );
xnor ( n39429 , n39428 , n28096 );
and ( n39430 , n29078 , n25383 );
and ( n39431 , n28700 , n25381 );
nor ( n39432 , n39430 , n39431 );
xnor ( n39433 , n39432 , n24885 );
and ( n39434 , n39429 , n39433 );
xor ( n39435 , n39356 , n39360 );
xor ( n39436 , n39435 , n39365 );
and ( n39437 , n39433 , n39436 );
and ( n39438 , n39429 , n39436 );
or ( n39439 , n39434 , n39437 , n39438 );
and ( n39440 , n24527 , n29977 );
and ( n39441 , n24521 , n29974 );
nor ( n39442 , n39440 , n39441 );
xnor ( n39443 , n39442 , n28674 );
and ( n39444 , n39439 , n39443 );
xor ( n39445 , n39270 , n39153 );
xor ( n39446 , n39445 , n39273 );
and ( n39447 , n39443 , n39446 );
and ( n39448 , n39439 , n39446 );
or ( n39449 , n39444 , n39447 , n39448 );
and ( n39450 , n39425 , n39449 );
xor ( n39451 , n39317 , n39321 );
xor ( n39452 , n39451 , n39324 );
and ( n39453 , n39449 , n39452 );
and ( n39454 , n39425 , n39452 );
or ( n39455 , n39450 , n39453 , n39454 );
and ( n39456 , n39386 , n39455 );
xor ( n39457 , n39288 , n39290 );
xor ( n39458 , n39457 , n39293 );
and ( n39459 , n39455 , n39458 );
and ( n39460 , n39386 , n39458 );
or ( n39461 , n39456 , n39459 , n39460 );
xor ( n39462 , n39242 , n39244 );
xor ( n39463 , n39462 , n39247 );
and ( n39464 , n39461 , n39463 );
xor ( n39465 , n39296 , n39335 );
xor ( n39466 , n39465 , n39338 );
and ( n39467 , n39463 , n39466 );
and ( n39468 , n39461 , n39466 );
or ( n39469 , n39464 , n39467 , n39468 );
and ( n39470 , n39355 , n39469 );
xor ( n39471 , n39355 , n39469 );
xor ( n39472 , n39461 , n39463 );
xor ( n39473 , n39472 , n39466 );
and ( n39474 , n27352 , n27529 );
and ( n39475 , n27135 , n27527 );
nor ( n39476 , n39474 , n39475 );
xnor ( n39477 , n39476 , n27034 );
and ( n39478 , n27757 , n26992 );
and ( n39479 , n27751 , n26990 );
nor ( n39480 , n39478 , n39479 );
xnor ( n39481 , n39480 , n26369 );
and ( n39482 , n39477 , n39481 );
and ( n39483 , n26422 , n28062 );
and ( n39484 , n26319 , n28060 );
nor ( n39485 , n39483 , n39484 );
xnor ( n39486 , n39485 , n27549 );
and ( n39487 , n39482 , n39486 );
and ( n39488 , n28700 , n26027 );
and ( n39489 , n28810 , n26025 );
nor ( n39490 , n39488 , n39489 );
xnor ( n39491 , n39490 , n25499 );
and ( n39492 , n39486 , n39491 );
and ( n39493 , n39482 , n39491 );
or ( n39494 , n39487 , n39492 , n39493 );
and ( n39495 , n25974 , n28628 );
and ( n39496 , n25765 , n28626 );
nor ( n39497 , n39495 , n39496 );
xnor ( n39498 , n39497 , n28096 );
and ( n39499 , n39498 , n39408 );
xor ( n39500 , n39390 , n39394 );
xor ( n39501 , n39500 , n39399 );
and ( n39502 , n39408 , n39501 );
and ( n39503 , n39498 , n39501 );
or ( n39504 , n39499 , n39502 , n39503 );
and ( n39505 , n39494 , n39504 );
and ( n39506 , n29623 , n24902 );
and ( n39507 , n29318 , n24900 );
nor ( n39508 , n39506 , n39507 );
xnor ( n39509 , n39508 , n24397 );
and ( n39510 , n39504 , n39509 );
and ( n39511 , n39494 , n39509 );
or ( n39512 , n39505 , n39510 , n39511 );
xor ( n39513 , n39413 , n39417 );
xor ( n39514 , n39513 , n39422 );
and ( n39515 , n39512 , n39514 );
xor ( n39516 , n39368 , n39372 );
xor ( n39517 , n39516 , n39375 );
and ( n39518 , n39514 , n39517 );
and ( n39519 , n39512 , n39517 );
or ( n39520 , n39515 , n39518 , n39519 );
xor ( n39521 , n39276 , n39280 );
xor ( n39522 , n39521 , n39285 );
and ( n39523 , n39520 , n39522 );
xor ( n39524 , n39378 , n39380 );
xor ( n39525 , n39524 , n39383 );
and ( n39526 , n39522 , n39525 );
and ( n39527 , n39520 , n39525 );
or ( n39528 , n39523 , n39526 , n39527 );
xor ( n39529 , n39327 , n39329 );
xor ( n39530 , n39529 , n39332 );
and ( n39531 , n39528 , n39530 );
xor ( n39532 , n39386 , n39455 );
xor ( n39533 , n39532 , n39458 );
and ( n39534 , n39530 , n39533 );
and ( n39535 , n39528 , n39533 );
or ( n39536 , n39531 , n39534 , n39535 );
and ( n39537 , n39473 , n39536 );
xor ( n39538 , n39473 , n39536 );
and ( n39539 , n24621 , n29977 );
and ( n39540 , n24527 , n29974 );
nor ( n39541 , n39539 , n39540 );
xnor ( n39542 , n39541 , n28674 );
and ( n39543 , n25284 , n29276 );
and ( n39544 , n24940 , n29274 );
nor ( n39545 , n39543 , n39544 );
xnor ( n39546 , n39545 , n28677 );
and ( n39547 , n39542 , n39546 );
xor ( n39548 , n39402 , n39406 );
xor ( n39549 , n39548 , n39410 );
and ( n39550 , n39546 , n39549 );
and ( n39551 , n39542 , n39549 );
or ( n39552 , n39547 , n39550 , n39551 );
and ( n39553 , n26851 , n28062 );
and ( n39554 , n26422 , n28060 );
nor ( n39555 , n39553 , n39554 );
xnor ( n39556 , n39555 , n27549 );
and ( n39557 , n28810 , n26349 );
and ( n39558 , n28211 , n26347 );
nor ( n39559 , n39557 , n39558 );
xnor ( n39560 , n39559 , n25893 );
and ( n39561 , n39556 , n39560 );
and ( n39562 , n29078 , n26027 );
and ( n39563 , n28700 , n26025 );
nor ( n39564 , n39562 , n39563 );
xnor ( n39565 , n39564 , n25499 );
and ( n39566 , n39560 , n39565 );
and ( n39567 , n39556 , n39565 );
or ( n39568 , n39561 , n39566 , n39567 );
xor ( n39569 , n39477 , n39481 );
and ( n39570 , n27135 , n28062 );
and ( n39571 , n26851 , n28060 );
nor ( n39572 , n39570 , n39571 );
xnor ( n39573 , n39572 , n27549 );
and ( n39574 , n27751 , n27529 );
and ( n39575 , n27352 , n27527 );
nor ( n39576 , n39574 , n39575 );
xnor ( n39577 , n39576 , n27034 );
and ( n39578 , n39573 , n39577 );
and ( n39579 , n28211 , n26992 );
and ( n39580 , n27757 , n26990 );
nor ( n39581 , n39579 , n39580 );
xnor ( n39582 , n39581 , n26369 );
and ( n39583 , n39577 , n39582 );
and ( n39584 , n39573 , n39582 );
or ( n39585 , n39578 , n39583 , n39584 );
and ( n39586 , n39569 , n39585 );
and ( n39587 , n29623 , n25381 );
not ( n39588 , n39587 );
and ( n39589 , n39588 , n24885 );
and ( n39590 , n39585 , n39589 );
and ( n39591 , n39569 , n39589 );
or ( n39592 , n39586 , n39590 , n39591 );
and ( n39593 , n39568 , n39592 );
and ( n39594 , n29318 , n25383 );
and ( n39595 , n29078 , n25381 );
nor ( n39596 , n39594 , n39595 );
xnor ( n39597 , n39596 , n24885 );
and ( n39598 , n39592 , n39597 );
and ( n39599 , n39568 , n39597 );
or ( n39600 , n39593 , n39598 , n39599 );
xor ( n39601 , n39494 , n39504 );
xor ( n39602 , n39601 , n39509 );
and ( n39603 , n39600 , n39602 );
xor ( n39604 , n39429 , n39433 );
xor ( n39605 , n39604 , n39436 );
and ( n39606 , n39602 , n39605 );
and ( n39607 , n39600 , n39605 );
or ( n39608 , n39603 , n39606 , n39607 );
and ( n39609 , n39552 , n39608 );
xor ( n39610 , n39439 , n39443 );
xor ( n39611 , n39610 , n39446 );
and ( n39612 , n39608 , n39611 );
and ( n39613 , n39552 , n39611 );
or ( n39614 , n39609 , n39612 , n39613 );
xor ( n39615 , n39425 , n39449 );
xor ( n39616 , n39615 , n39452 );
and ( n39617 , n39614 , n39616 );
xor ( n39618 , n39520 , n39522 );
xor ( n39619 , n39618 , n39525 );
and ( n39620 , n39616 , n39619 );
and ( n39621 , n39614 , n39619 );
or ( n39622 , n39617 , n39620 , n39621 );
xor ( n39623 , n39528 , n39530 );
xor ( n39624 , n39623 , n39533 );
and ( n39625 , n39622 , n39624 );
xor ( n39626 , n39622 , n39624 );
xor ( n39627 , n39614 , n39616 );
xor ( n39628 , n39627 , n39619 );
and ( n39629 , n24940 , n29977 );
and ( n39630 , n24621 , n29974 );
nor ( n39631 , n39629 , n39630 );
xnor ( n39632 , n39631 , n28674 );
and ( n39633 , n25554 , n29276 );
and ( n39634 , n25284 , n29274 );
nor ( n39635 , n39633 , n39634 );
xnor ( n39636 , n39635 , n28677 );
and ( n39637 , n39632 , n39636 );
xor ( n39638 , n39482 , n39486 );
xor ( n39639 , n39638 , n39491 );
and ( n39640 , n39636 , n39639 );
and ( n39641 , n39632 , n39639 );
or ( n39642 , n39637 , n39640 , n39641 );
and ( n39643 , n25765 , n29276 );
and ( n39644 , n25554 , n29274 );
nor ( n39645 , n39643 , n39644 );
xnor ( n39646 , n39645 , n28677 );
and ( n39647 , n26319 , n28628 );
and ( n39648 , n25974 , n28626 );
nor ( n39649 , n39647 , n39648 );
xnor ( n39650 , n39649 , n28096 );
and ( n39651 , n39646 , n39650 );
and ( n39652 , n29623 , n25383 );
and ( n39653 , n29318 , n25381 );
nor ( n39654 , n39652 , n39653 );
xnor ( n39655 , n39654 , n24885 );
and ( n39656 , n39650 , n39655 );
and ( n39657 , n39646 , n39655 );
or ( n39658 , n39651 , n39656 , n39657 );
xor ( n39659 , n39568 , n39592 );
xor ( n39660 , n39659 , n39597 );
and ( n39661 , n39658 , n39660 );
xor ( n39662 , n39498 , n39408 );
xor ( n39663 , n39662 , n39501 );
and ( n39664 , n39660 , n39663 );
and ( n39665 , n39658 , n39663 );
or ( n39666 , n39661 , n39664 , n39665 );
and ( n39667 , n39642 , n39666 );
xor ( n39668 , n39542 , n39546 );
xor ( n39669 , n39668 , n39549 );
and ( n39670 , n39666 , n39669 );
and ( n39671 , n39642 , n39669 );
or ( n39672 , n39667 , n39670 , n39671 );
xor ( n39673 , n39512 , n39514 );
xor ( n39674 , n39673 , n39517 );
and ( n39675 , n39672 , n39674 );
xor ( n39676 , n39552 , n39608 );
xor ( n39677 , n39676 , n39611 );
and ( n39678 , n39674 , n39677 );
and ( n39679 , n39672 , n39677 );
or ( n39680 , n39675 , n39678 , n39679 );
and ( n39681 , n39628 , n39680 );
xor ( n39682 , n39628 , n39680 );
xor ( n39683 , n39672 , n39674 );
xor ( n39684 , n39683 , n39677 );
and ( n39685 , n27757 , n27529 );
and ( n39686 , n27751 , n27527 );
nor ( n39687 , n39685 , n39686 );
xnor ( n39688 , n39687 , n27034 );
and ( n39689 , n28810 , n26992 );
and ( n39690 , n28211 , n26990 );
nor ( n39691 , n39689 , n39690 );
xnor ( n39692 , n39691 , n26369 );
xor ( n39693 , n39688 , n39692 );
and ( n39694 , n27352 , n28062 );
and ( n39695 , n27135 , n28060 );
nor ( n39696 , n39694 , n39695 );
xnor ( n39697 , n39696 , n27549 );
and ( n39698 , n39693 , n39697 );
and ( n39699 , n29623 , n26025 );
not ( n39700 , n39699 );
and ( n39701 , n39700 , n25499 );
and ( n39702 , n39697 , n39701 );
and ( n39703 , n39693 , n39701 );
or ( n39704 , n39698 , n39702 , n39703 );
and ( n39705 , n26422 , n28628 );
and ( n39706 , n26319 , n28626 );
nor ( n39707 , n39705 , n39706 );
xnor ( n39708 , n39707 , n28096 );
and ( n39709 , n39704 , n39708 );
and ( n39710 , n39708 , n39587 );
and ( n39711 , n39704 , n39587 );
or ( n39712 , n39709 , n39710 , n39711 );
and ( n39713 , n26851 , n28628 );
and ( n39714 , n26422 , n28626 );
nor ( n39715 , n39713 , n39714 );
xnor ( n39716 , n39715 , n28096 );
and ( n39717 , n29078 , n26349 );
and ( n39718 , n28700 , n26347 );
nor ( n39719 , n39717 , n39718 );
xnor ( n39720 , n39719 , n25893 );
and ( n39721 , n39716 , n39720 );
and ( n39722 , n29623 , n26027 );
and ( n39723 , n29318 , n26025 );
nor ( n39724 , n39722 , n39723 );
xnor ( n39725 , n39724 , n25499 );
and ( n39726 , n39720 , n39725 );
and ( n39727 , n39716 , n39725 );
or ( n39728 , n39721 , n39726 , n39727 );
and ( n39729 , n25974 , n29276 );
and ( n39730 , n25765 , n29274 );
nor ( n39731 , n39729 , n39730 );
xnor ( n39732 , n39731 , n28677 );
and ( n39733 , n39728 , n39732 );
xor ( n39734 , n39573 , n39577 );
xor ( n39735 , n39734 , n39582 );
and ( n39736 , n39732 , n39735 );
and ( n39737 , n39728 , n39735 );
or ( n39738 , n39733 , n39736 , n39737 );
and ( n39739 , n39712 , n39738 );
and ( n39740 , n25284 , n29977 );
and ( n39741 , n24940 , n29974 );
nor ( n39742 , n39740 , n39741 );
xnor ( n39743 , n39742 , n28674 );
and ( n39744 , n39738 , n39743 );
and ( n39745 , n39712 , n39743 );
or ( n39746 , n39739 , n39744 , n39745 );
and ( n39747 , n39688 , n39692 );
and ( n39748 , n28700 , n26349 );
and ( n39749 , n28810 , n26347 );
nor ( n39750 , n39748 , n39749 );
xnor ( n39751 , n39750 , n25893 );
and ( n39752 , n39747 , n39751 );
and ( n39753 , n29318 , n26027 );
and ( n39754 , n29078 , n26025 );
nor ( n39755 , n39753 , n39754 );
xnor ( n39756 , n39755 , n25499 );
and ( n39757 , n39751 , n39756 );
and ( n39758 , n39747 , n39756 );
or ( n39759 , n39752 , n39757 , n39758 );
xor ( n39760 , n39556 , n39560 );
xor ( n39761 , n39760 , n39565 );
and ( n39762 , n39759 , n39761 );
xor ( n39763 , n39569 , n39585 );
xor ( n39764 , n39763 , n39589 );
and ( n39765 , n39761 , n39764 );
and ( n39766 , n39759 , n39764 );
or ( n39767 , n39762 , n39765 , n39766 );
and ( n39768 , n39746 , n39767 );
xor ( n39769 , n39632 , n39636 );
xor ( n39770 , n39769 , n39639 );
and ( n39771 , n39767 , n39770 );
and ( n39772 , n39746 , n39770 );
or ( n39773 , n39768 , n39771 , n39772 );
xor ( n39774 , n39600 , n39602 );
xor ( n39775 , n39774 , n39605 );
and ( n39776 , n39773 , n39775 );
xor ( n39777 , n39642 , n39666 );
xor ( n39778 , n39777 , n39669 );
and ( n39779 , n39775 , n39778 );
and ( n39780 , n39773 , n39778 );
or ( n39781 , n39776 , n39779 , n39780 );
and ( n39782 , n39684 , n39781 );
xor ( n39783 , n39684 , n39781 );
xor ( n39784 , n39773 , n39775 );
xor ( n39785 , n39784 , n39778 );
and ( n39786 , n27751 , n28062 );
and ( n39787 , n27352 , n28060 );
nor ( n39788 , n39786 , n39787 );
xnor ( n39789 , n39788 , n27549 );
and ( n39790 , n28211 , n27529 );
and ( n39791 , n27757 , n27527 );
nor ( n39792 , n39790 , n39791 );
xnor ( n39793 , n39792 , n27034 );
and ( n39794 , n39789 , n39793 );
and ( n39795 , n28700 , n26992 );
and ( n39796 , n28810 , n26990 );
nor ( n39797 , n39795 , n39796 );
xnor ( n39798 , n39797 , n26369 );
and ( n39799 , n39793 , n39798 );
and ( n39800 , n39789 , n39798 );
or ( n39801 , n39794 , n39799 , n39800 );
and ( n39802 , n27757 , n28062 );
and ( n39803 , n27751 , n28060 );
nor ( n39804 , n39802 , n39803 );
xnor ( n39805 , n39804 , n27549 );
and ( n39806 , n28810 , n27529 );
and ( n39807 , n28211 , n27527 );
nor ( n39808 , n39806 , n39807 );
xnor ( n39809 , n39808 , n27034 );
and ( n39810 , n39805 , n39809 );
and ( n39811 , n27135 , n28628 );
and ( n39812 , n26851 , n28626 );
nor ( n39813 , n39811 , n39812 );
xnor ( n39814 , n39813 , n28096 );
and ( n39815 , n39810 , n39814 );
and ( n39816 , n39814 , n39699 );
and ( n39817 , n39810 , n39699 );
or ( n39818 , n39815 , n39816 , n39817 );
and ( n39819 , n39801 , n39818 );
xor ( n39820 , n39693 , n39697 );
xor ( n39821 , n39820 , n39701 );
and ( n39822 , n39818 , n39821 );
and ( n39823 , n39801 , n39821 );
or ( n39824 , n39819 , n39822 , n39823 );
and ( n39825 , n25554 , n29977 );
and ( n39826 , n25284 , n29974 );
nor ( n39827 , n39825 , n39826 );
xnor ( n39828 , n39827 , n28674 );
and ( n39829 , n39824 , n39828 );
xor ( n39830 , n39747 , n39751 );
xor ( n39831 , n39830 , n39756 );
and ( n39832 , n39828 , n39831 );
and ( n39833 , n39824 , n39831 );
or ( n39834 , n39829 , n39832 , n39833 );
xor ( n39835 , n39646 , n39650 );
xor ( n39836 , n39835 , n39655 );
and ( n39837 , n39834 , n39836 );
xor ( n39838 , n39759 , n39761 );
xor ( n39839 , n39838 , n39764 );
and ( n39840 , n39836 , n39839 );
and ( n39841 , n39834 , n39839 );
or ( n39842 , n39837 , n39840 , n39841 );
xor ( n39843 , n39658 , n39660 );
xor ( n39844 , n39843 , n39663 );
and ( n39845 , n39842 , n39844 );
xor ( n39846 , n39746 , n39767 );
xor ( n39847 , n39846 , n39770 );
and ( n39848 , n39844 , n39847 );
and ( n39849 , n39842 , n39847 );
or ( n39850 , n39845 , n39848 , n39849 );
and ( n39851 , n39785 , n39850 );
xor ( n39852 , n39785 , n39850 );
xor ( n39853 , n39842 , n39844 );
xor ( n39854 , n39853 , n39847 );
and ( n39855 , n25765 , n29977 );
and ( n39856 , n25554 , n29974 );
nor ( n39857 , n39855 , n39856 );
xnor ( n39858 , n39857 , n28674 );
and ( n39859 , n26319 , n29276 );
and ( n39860 , n25974 , n29274 );
nor ( n39861 , n39859 , n39860 );
xnor ( n39862 , n39861 , n28677 );
and ( n39863 , n39858 , n39862 );
xor ( n39864 , n39716 , n39720 );
xor ( n39865 , n39864 , n39725 );
and ( n39866 , n39862 , n39865 );
and ( n39867 , n39858 , n39865 );
or ( n39868 , n39863 , n39866 , n39867 );
xor ( n39869 , n39704 , n39708 );
xor ( n39870 , n39869 , n39587 );
and ( n39871 , n39868 , n39870 );
xor ( n39872 , n39728 , n39732 );
xor ( n39873 , n39872 , n39735 );
and ( n39874 , n39870 , n39873 );
and ( n39875 , n39868 , n39873 );
or ( n39876 , n39871 , n39874 , n39875 );
xor ( n39877 , n39712 , n39738 );
xor ( n39878 , n39877 , n39743 );
and ( n39879 , n39876 , n39878 );
xor ( n39880 , n39834 , n39836 );
xor ( n39881 , n39880 , n39839 );
and ( n39882 , n39878 , n39881 );
and ( n39883 , n39876 , n39881 );
or ( n39884 , n39879 , n39882 , n39883 );
and ( n39885 , n39854 , n39884 );
xor ( n39886 , n39854 , n39884 );
and ( n39887 , n26422 , n29276 );
and ( n39888 , n26319 , n29274 );
nor ( n39889 , n39887 , n39888 );
xnor ( n39890 , n39889 , n28677 );
and ( n39891 , n29318 , n26349 );
and ( n39892 , n29078 , n26347 );
nor ( n39893 , n39891 , n39892 );
xnor ( n39894 , n39893 , n25893 );
and ( n39895 , n39890 , n39894 );
xor ( n39896 , n39789 , n39793 );
xor ( n39897 , n39896 , n39798 );
and ( n39898 , n39894 , n39897 );
and ( n39899 , n39890 , n39897 );
or ( n39900 , n39895 , n39898 , n39899 );
and ( n39901 , n27352 , n28628 );
and ( n39902 , n27135 , n28626 );
nor ( n39903 , n39901 , n39902 );
xnor ( n39904 , n39903 , n28096 );
and ( n39905 , n29078 , n26992 );
and ( n39906 , n28700 , n26990 );
nor ( n39907 , n39905 , n39906 );
xnor ( n39908 , n39907 , n26369 );
and ( n39909 , n39904 , n39908 );
and ( n39910 , n29623 , n26347 );
not ( n39911 , n39910 );
and ( n39912 , n39911 , n25893 );
and ( n39913 , n39908 , n39912 );
and ( n39914 , n39904 , n39912 );
or ( n39915 , n39909 , n39913 , n39914 );
and ( n39916 , n25974 , n29977 );
and ( n39917 , n25765 , n29974 );
nor ( n39918 , n39916 , n39917 );
xnor ( n39919 , n39918 , n28674 );
and ( n39920 , n39915 , n39919 );
xor ( n39921 , n39810 , n39814 );
xor ( n39922 , n39921 , n39699 );
and ( n39923 , n39919 , n39922 );
and ( n39924 , n39915 , n39922 );
or ( n39925 , n39920 , n39923 , n39924 );
and ( n39926 , n39900 , n39925 );
xor ( n39927 , n39801 , n39818 );
xor ( n39928 , n39927 , n39821 );
and ( n39929 , n39925 , n39928 );
and ( n39930 , n39900 , n39928 );
or ( n39931 , n39926 , n39929 , n39930 );
xor ( n39932 , n39824 , n39828 );
xor ( n39933 , n39932 , n39831 );
and ( n39934 , n39931 , n39933 );
xor ( n39935 , n39868 , n39870 );
xor ( n39936 , n39935 , n39873 );
and ( n39937 , n39933 , n39936 );
and ( n39938 , n39931 , n39936 );
or ( n39939 , n39934 , n39937 , n39938 );
xor ( n39940 , n39876 , n39878 );
xor ( n39941 , n39940 , n39881 );
and ( n39942 , n39939 , n39941 );
xor ( n39943 , n39939 , n39941 );
xor ( n39944 , n39931 , n39933 );
xor ( n39945 , n39944 , n39936 );
xor ( n39946 , n39805 , n39809 );
and ( n39947 , n28810 , n28062 );
and ( n39948 , n28211 , n28060 );
nor ( n39949 , n39947 , n39948 );
xnor ( n39950 , n39949 , n27549 );
and ( n39951 , n29623 , n26990 );
not ( n39952 , n39951 );
and ( n39953 , n39952 , n26369 );
and ( n39954 , n39950 , n39953 );
and ( n39955 , n28211 , n28062 );
and ( n39956 , n27757 , n28060 );
nor ( n39957 , n39955 , n39956 );
xnor ( n39958 , n39957 , n27549 );
and ( n39959 , n39954 , n39958 );
and ( n39960 , n28700 , n27529 );
and ( n39961 , n28810 , n27527 );
nor ( n39962 , n39960 , n39961 );
xnor ( n39963 , n39962 , n27034 );
and ( n39964 , n39958 , n39963 );
and ( n39965 , n39954 , n39963 );
or ( n39966 , n39959 , n39964 , n39965 );
and ( n39967 , n39946 , n39966 );
and ( n39968 , n26851 , n29276 );
and ( n39969 , n26422 , n29274 );
nor ( n39970 , n39968 , n39969 );
xnor ( n39971 , n39970 , n28677 );
and ( n39972 , n39966 , n39971 );
and ( n39973 , n39946 , n39971 );
or ( n39974 , n39967 , n39972 , n39973 );
and ( n39975 , n27751 , n28628 );
and ( n39976 , n27352 , n28626 );
nor ( n39977 , n39975 , n39976 );
xnor ( n39978 , n39977 , n28096 );
and ( n39979 , n29318 , n26992 );
and ( n39980 , n29078 , n26990 );
nor ( n39981 , n39979 , n39980 );
xnor ( n39982 , n39981 , n26369 );
and ( n39983 , n39978 , n39982 );
and ( n39984 , n39982 , n39910 );
and ( n39985 , n39978 , n39910 );
or ( n39986 , n39983 , n39984 , n39985 );
and ( n39987 , n29623 , n26349 );
and ( n39988 , n29318 , n26347 );
nor ( n39989 , n39987 , n39988 );
xnor ( n39990 , n39989 , n25893 );
and ( n39991 , n39986 , n39990 );
xor ( n39992 , n39904 , n39908 );
xor ( n39993 , n39992 , n39912 );
and ( n39994 , n39990 , n39993 );
and ( n39995 , n39986 , n39993 );
or ( n39996 , n39991 , n39994 , n39995 );
and ( n39997 , n39974 , n39996 );
xor ( n39998 , n39890 , n39894 );
xor ( n39999 , n39998 , n39897 );
and ( n40000 , n39996 , n39999 );
and ( n40001 , n39974 , n39999 );
or ( n40002 , n39997 , n40000 , n40001 );
xor ( n40003 , n39858 , n39862 );
xor ( n40004 , n40003 , n39865 );
and ( n40005 , n40002 , n40004 );
xor ( n40006 , n39900 , n39925 );
xor ( n40007 , n40006 , n39928 );
and ( n40008 , n40004 , n40007 );
and ( n40009 , n40002 , n40007 );
or ( n40010 , n40005 , n40008 , n40009 );
and ( n40011 , n39945 , n40010 );
xor ( n40012 , n39945 , n40010 );
xor ( n40013 , n40002 , n40004 );
xor ( n40014 , n40013 , n40007 );
xor ( n40015 , n39950 , n39953 );
and ( n40016 , n27757 , n28628 );
and ( n40017 , n27751 , n28626 );
nor ( n40018 , n40016 , n40017 );
xnor ( n40019 , n40018 , n28096 );
and ( n40020 , n40015 , n40019 );
and ( n40021 , n29078 , n27529 );
and ( n40022 , n28700 , n27527 );
nor ( n40023 , n40021 , n40022 );
xnor ( n40024 , n40023 , n27034 );
and ( n40025 , n40019 , n40024 );
and ( n40026 , n40015 , n40024 );
or ( n40027 , n40020 , n40025 , n40026 );
and ( n40028 , n27135 , n29276 );
and ( n40029 , n26851 , n29274 );
nor ( n40030 , n40028 , n40029 );
xnor ( n40031 , n40030 , n28677 );
and ( n40032 , n40027 , n40031 );
xor ( n40033 , n39954 , n39958 );
xor ( n40034 , n40033 , n39963 );
and ( n40035 , n40031 , n40034 );
and ( n40036 , n40027 , n40034 );
or ( n40037 , n40032 , n40035 , n40036 );
and ( n40038 , n26319 , n29977 );
and ( n40039 , n25974 , n29974 );
nor ( n40040 , n40038 , n40039 );
xnor ( n40041 , n40040 , n28674 );
and ( n40042 , n40037 , n40041 );
xor ( n40043 , n39946 , n39966 );
xor ( n40044 , n40043 , n39971 );
and ( n40045 , n40041 , n40044 );
and ( n40046 , n40037 , n40044 );
or ( n40047 , n40042 , n40045 , n40046 );
xor ( n40048 , n39915 , n39919 );
xor ( n40049 , n40048 , n39922 );
and ( n40050 , n40047 , n40049 );
xor ( n40051 , n39974 , n39996 );
xor ( n40052 , n40051 , n39999 );
and ( n40053 , n40049 , n40052 );
and ( n40054 , n40047 , n40052 );
or ( n40055 , n40050 , n40053 , n40054 );
and ( n40056 , n40014 , n40055 );
xor ( n40057 , n40014 , n40055 );
xor ( n40058 , n40047 , n40049 );
xor ( n40059 , n40058 , n40052 );
and ( n40060 , n28211 , n28628 );
and ( n40061 , n27757 , n28626 );
nor ( n40062 , n40060 , n40061 );
xnor ( n40063 , n40062 , n28096 );
and ( n40064 , n28700 , n28062 );
and ( n40065 , n28810 , n28060 );
nor ( n40066 , n40064 , n40065 );
xnor ( n40067 , n40066 , n27549 );
and ( n40068 , n40063 , n40067 );
and ( n40069 , n40067 , n39951 );
and ( n40070 , n40063 , n39951 );
or ( n40071 , n40068 , n40069 , n40070 );
and ( n40072 , n27352 , n29276 );
and ( n40073 , n27135 , n29274 );
nor ( n40074 , n40072 , n40073 );
xnor ( n40075 , n40074 , n28677 );
and ( n40076 , n40071 , n40075 );
and ( n40077 , n29623 , n26992 );
and ( n40078 , n29318 , n26990 );
nor ( n40079 , n40077 , n40078 );
xnor ( n40080 , n40079 , n26369 );
and ( n40081 , n40075 , n40080 );
and ( n40082 , n40071 , n40080 );
or ( n40083 , n40076 , n40081 , n40082 );
and ( n40084 , n26422 , n29977 );
and ( n40085 , n26319 , n29974 );
nor ( n40086 , n40084 , n40085 );
xnor ( n40087 , n40086 , n28674 );
and ( n40088 , n40083 , n40087 );
xor ( n40089 , n39978 , n39982 );
xor ( n40090 , n40089 , n39910 );
and ( n40091 , n40087 , n40090 );
and ( n40092 , n40083 , n40090 );
or ( n40093 , n40088 , n40091 , n40092 );
xor ( n40094 , n39986 , n39990 );
xor ( n40095 , n40094 , n39993 );
and ( n40096 , n40093 , n40095 );
xor ( n40097 , n40037 , n40041 );
xor ( n40098 , n40097 , n40044 );
and ( n40099 , n40095 , n40098 );
and ( n40100 , n40093 , n40098 );
or ( n40101 , n40096 , n40099 , n40100 );
and ( n40102 , n40059 , n40101 );
xor ( n40103 , n40059 , n40101 );
and ( n40104 , n28810 , n28628 );
and ( n40105 , n28211 , n28626 );
nor ( n40106 , n40104 , n40105 );
xnor ( n40107 , n40106 , n28096 );
and ( n40108 , n29078 , n28062 );
and ( n40109 , n28700 , n28060 );
nor ( n40110 , n40108 , n40109 );
xnor ( n40111 , n40110 , n27549 );
and ( n40112 , n40107 , n40111 );
and ( n40113 , n27751 , n29276 );
and ( n40114 , n27352 , n29274 );
nor ( n40115 , n40113 , n40114 );
xnor ( n40116 , n40115 , n28677 );
and ( n40117 , n40112 , n40116 );
and ( n40118 , n29318 , n27529 );
and ( n40119 , n29078 , n27527 );
nor ( n40120 , n40118 , n40119 );
xnor ( n40121 , n40120 , n27034 );
and ( n40122 , n40116 , n40121 );
and ( n40123 , n40112 , n40121 );
or ( n40124 , n40117 , n40122 , n40123 );
and ( n40125 , n26851 , n29977 );
and ( n40126 , n26422 , n29974 );
nor ( n40127 , n40125 , n40126 );
xnor ( n40128 , n40127 , n28674 );
and ( n40129 , n40124 , n40128 );
xor ( n40130 , n40015 , n40019 );
xor ( n40131 , n40130 , n40024 );
and ( n40132 , n40128 , n40131 );
and ( n40133 , n40124 , n40131 );
or ( n40134 , n40129 , n40132 , n40133 );
xor ( n40135 , n40027 , n40031 );
xor ( n40136 , n40135 , n40034 );
and ( n40137 , n40134 , n40136 );
xor ( n40138 , n40083 , n40087 );
xor ( n40139 , n40138 , n40090 );
and ( n40140 , n40136 , n40139 );
and ( n40141 , n40134 , n40139 );
or ( n40142 , n40137 , n40140 , n40141 );
xor ( n40143 , n40093 , n40095 );
xor ( n40144 , n40143 , n40098 );
and ( n40145 , n40142 , n40144 );
xor ( n40146 , n40142 , n40144 );
xor ( n40147 , n40134 , n40136 );
xor ( n40148 , n40147 , n40139 );
xor ( n40149 , n40107 , n40111 );
and ( n40150 , n28700 , n28628 );
and ( n40151 , n28810 , n28626 );
nor ( n40152 , n40150 , n40151 );
xnor ( n40153 , n40152 , n28096 );
and ( n40154 , n29318 , n28062 );
and ( n40155 , n29078 , n28060 );
nor ( n40156 , n40154 , n40155 );
xnor ( n40157 , n40156 , n27549 );
and ( n40158 , n40153 , n40157 );
and ( n40159 , n29623 , n27527 );
and ( n40160 , n40157 , n40159 );
and ( n40161 , n40153 , n40159 );
or ( n40162 , n40158 , n40160 , n40161 );
and ( n40163 , n40149 , n40162 );
not ( n40164 , n40159 );
and ( n40165 , n40164 , n27034 );
and ( n40166 , n40162 , n40165 );
and ( n40167 , n40149 , n40165 );
or ( n40168 , n40163 , n40166 , n40167 );
and ( n40169 , n27135 , n29977 );
and ( n40170 , n26851 , n29974 );
nor ( n40171 , n40169 , n40170 );
xnor ( n40172 , n40171 , n28674 );
and ( n40173 , n40168 , n40172 );
xor ( n40174 , n40063 , n40067 );
xor ( n40175 , n40174 , n39951 );
and ( n40176 , n40172 , n40175 );
and ( n40177 , n40168 , n40175 );
or ( n40178 , n40173 , n40176 , n40177 );
xor ( n40179 , n40071 , n40075 );
xor ( n40180 , n40179 , n40080 );
and ( n40181 , n40178 , n40180 );
xor ( n40182 , n40124 , n40128 );
xor ( n40183 , n40182 , n40131 );
and ( n40184 , n40180 , n40183 );
and ( n40185 , n40178 , n40183 );
or ( n40186 , n40181 , n40184 , n40185 );
and ( n40187 , n40148 , n40186 );
xor ( n40188 , n40148 , n40186 );
xor ( n40189 , n40178 , n40180 );
xor ( n40190 , n40189 , n40183 );
and ( n40191 , n27757 , n29276 );
and ( n40192 , n27751 , n29274 );
nor ( n40193 , n40191 , n40192 );
xnor ( n40194 , n40193 , n28677 );
and ( n40195 , n29623 , n27529 );
and ( n40196 , n29318 , n27527 );
nor ( n40197 , n40195 , n40196 );
xnor ( n40198 , n40197 , n27034 );
and ( n40199 , n40194 , n40198 );
xor ( n40200 , n40149 , n40162 );
xor ( n40201 , n40200 , n40165 );
and ( n40202 , n40198 , n40201 );
and ( n40203 , n40194 , n40201 );
or ( n40204 , n40199 , n40202 , n40203 );
xor ( n40205 , n40112 , n40116 );
xor ( n40206 , n40205 , n40121 );
and ( n40207 , n40204 , n40206 );
xor ( n40208 , n40168 , n40172 );
xor ( n40209 , n40208 , n40175 );
and ( n40210 , n40206 , n40209 );
and ( n40211 , n40204 , n40209 );
or ( n40212 , n40207 , n40210 , n40211 );
and ( n40213 , n40190 , n40212 );
xor ( n40214 , n40190 , n40212 );
xor ( n40215 , n40204 , n40206 );
xor ( n40216 , n40215 , n40209 );
and ( n40217 , n29078 , n28628 );
and ( n40218 , n28700 , n28626 );
nor ( n40219 , n40217 , n40218 );
xnor ( n40220 , n40219 , n28096 );
and ( n40221 , n29623 , n28060 );
not ( n40222 , n40221 );
and ( n40223 , n40222 , n27549 );
and ( n40224 , n40220 , n40223 );
xor ( n40225 , n40220 , n40223 );
and ( n40226 , n28810 , n29276 );
and ( n40227 , n28211 , n29274 );
nor ( n40228 , n40226 , n40227 );
xnor ( n40229 , n40228 , n28677 );
and ( n40230 , n40225 , n40229 );
and ( n40231 , n29623 , n28062 );
and ( n40232 , n29318 , n28060 );
nor ( n40233 , n40231 , n40232 );
xnor ( n40234 , n40233 , n27549 );
and ( n40235 , n40229 , n40234 );
and ( n40236 , n40225 , n40234 );
or ( n40237 , n40230 , n40235 , n40236 );
and ( n40238 , n40224 , n40237 );
and ( n40239 , n28211 , n29276 );
and ( n40240 , n27757 , n29274 );
nor ( n40241 , n40239 , n40240 );
xnor ( n40242 , n40241 , n28677 );
and ( n40243 , n40237 , n40242 );
and ( n40244 , n40224 , n40242 );
or ( n40245 , n40238 , n40243 , n40244 );
and ( n40246 , n27352 , n29977 );
and ( n40247 , n27135 , n29974 );
nor ( n40248 , n40246 , n40247 );
xnor ( n40249 , n40248 , n28674 );
and ( n40250 , n40245 , n40249 );
xor ( n40251 , n40194 , n40198 );
xor ( n40252 , n40251 , n40201 );
and ( n40253 , n40249 , n40252 );
and ( n40254 , n40245 , n40252 );
or ( n40255 , n40250 , n40253 , n40254 );
and ( n40256 , n40216 , n40255 );
xor ( n40257 , n40216 , n40255 );
xor ( n40258 , n40245 , n40249 );
xor ( n40259 , n40258 , n40252 );
and ( n40260 , n27751 , n29977 );
and ( n40261 , n27352 , n29974 );
nor ( n40262 , n40260 , n40261 );
xnor ( n40263 , n40262 , n28674 );
xor ( n40264 , n40153 , n40157 );
xor ( n40265 , n40264 , n40159 );
and ( n40266 , n40263 , n40265 );
xor ( n40267 , n40224 , n40237 );
xor ( n40268 , n40267 , n40242 );
and ( n40269 , n40265 , n40268 );
and ( n40270 , n40263 , n40268 );
or ( n40271 , n40266 , n40269 , n40270 );
and ( n40272 , n40259 , n40271 );
xor ( n40273 , n40259 , n40271 );
and ( n40274 , n28700 , n29276 );
and ( n40275 , n28810 , n29274 );
nor ( n40276 , n40274 , n40275 );
xnor ( n40277 , n40276 , n28677 );
and ( n40278 , n29318 , n28628 );
and ( n40279 , n29078 , n28626 );
nor ( n40280 , n40278 , n40279 );
xnor ( n40281 , n40280 , n28096 );
and ( n40282 , n40277 , n40281 );
and ( n40283 , n40281 , n40221 );
and ( n40284 , n40277 , n40221 );
or ( n40285 , n40282 , n40283 , n40284 );
and ( n40286 , n27757 , n29977 );
and ( n40287 , n27751 , n29974 );
nor ( n40288 , n40286 , n40287 );
xnor ( n40289 , n40288 , n28674 );
and ( n40290 , n40285 , n40289 );
xor ( n40291 , n40225 , n40229 );
xor ( n40292 , n40291 , n40234 );
and ( n40293 , n40289 , n40292 );
and ( n40294 , n40285 , n40292 );
or ( n40295 , n40290 , n40293 , n40294 );
xor ( n40296 , n40263 , n40265 );
xor ( n40297 , n40296 , n40268 );
and ( n40298 , n40295 , n40297 );
xor ( n40299 , n40295 , n40297 );
and ( n40300 , n29078 , n29276 );
and ( n40301 , n28700 , n29274 );
nor ( n40302 , n40300 , n40301 );
xnor ( n40303 , n40302 , n28677 );
and ( n40304 , n29623 , n28626 );
not ( n40305 , n40304 );
and ( n40306 , n40305 , n28096 );
and ( n40307 , n40303 , n40306 );
and ( n40308 , n28211 , n29977 );
and ( n40309 , n27757 , n29974 );
nor ( n40310 , n40308 , n40309 );
xnor ( n40311 , n40310 , n28674 );
and ( n40312 , n40307 , n40311 );
xor ( n40313 , n40277 , n40281 );
xor ( n40314 , n40313 , n40221 );
and ( n40315 , n40311 , n40314 );
and ( n40316 , n40307 , n40314 );
or ( n40317 , n40312 , n40315 , n40316 );
xor ( n40318 , n40285 , n40289 );
xor ( n40319 , n40318 , n40292 );
and ( n40320 , n40317 , n40319 );
xor ( n40321 , n40317 , n40319 );
xor ( n40322 , n40307 , n40311 );
xor ( n40323 , n40322 , n40314 );
xor ( n40324 , n40303 , n40306 );
and ( n40325 , n28810 , n29977 );
and ( n40326 , n28211 , n29974 );
nor ( n40327 , n40325 , n40326 );
xnor ( n40328 , n40327 , n28674 );
and ( n40329 , n40324 , n40328 );
and ( n40330 , n29623 , n28628 );
and ( n40331 , n29318 , n28626 );
nor ( n40332 , n40330 , n40331 );
xnor ( n40333 , n40332 , n28096 );
and ( n40334 , n40328 , n40333 );
and ( n40335 , n40324 , n40333 );
or ( n40336 , n40329 , n40334 , n40335 );
and ( n40337 , n40323 , n40336 );
xor ( n40338 , n40323 , n40336 );
xor ( n40339 , n40324 , n40328 );
xor ( n40340 , n40339 , n40333 );
and ( n40341 , n29623 , n29274 );
not ( n40342 , n40341 );
and ( n40343 , n40342 , n28677 );
and ( n40344 , n29623 , n29276 );
and ( n40345 , n29318 , n29274 );
nor ( n40346 , n40344 , n40345 );
xnor ( n40347 , n40346 , n28677 );
and ( n40348 , n40343 , n40347 );
and ( n40349 , n29318 , n29276 );
and ( n40350 , n29078 , n29274 );
nor ( n40351 , n40349 , n40350 );
xnor ( n40352 , n40351 , n28677 );
and ( n40353 , n40348 , n40352 );
and ( n40354 , n40352 , n40304 );
and ( n40355 , n40348 , n40304 );
or ( n40356 , n40353 , n40354 , n40355 );
and ( n40357 , n40340 , n40356 );
xor ( n40358 , n40340 , n40356 );
and ( n40359 , n28700 , n29977 );
and ( n40360 , n28810 , n29974 );
nor ( n40361 , n40359 , n40360 );
xnor ( n40362 , n40361 , n28674 );
xor ( n40363 , n40348 , n40352 );
xor ( n40364 , n40363 , n40304 );
and ( n40365 , n40362 , n40364 );
xor ( n40366 , n40362 , n40364 );
and ( n40367 , n29078 , n29977 );
and ( n40368 , n28700 , n29974 );
nor ( n40369 , n40367 , n40368 );
xnor ( n40370 , n40369 , n28674 );
xor ( n40371 , n40343 , n40347 );
and ( n40372 , n40370 , n40371 );
xor ( n40373 , n40370 , n40371 );
and ( n40374 , n29318 , n29977 );
and ( n40375 , n29078 , n29974 );
nor ( n40376 , n40374 , n40375 );
xnor ( n40377 , n40376 , n28674 );
and ( n40378 , n40377 , n40341 );
xor ( n40379 , n40377 , n40341 );
and ( n40380 , n29623 , n29977 );
and ( n40381 , n29318 , n29974 );
nor ( n40382 , n40380 , n40381 );
xnor ( n40383 , n40382 , n28674 );
and ( n40384 , n29623 , n29974 );
not ( n40385 , n40384 );
and ( n40386 , n40385 , n28674 );
and ( n40387 , n40383 , n40386 );
and ( n40388 , n40379 , n40387 );
or ( n40389 , n40378 , n40388 );
and ( n40390 , n40373 , n40389 );
or ( n40391 , n40372 , n40390 );
and ( n40392 , n40366 , n40391 );
or ( n40393 , n40365 , n40392 );
and ( n40394 , n40358 , n40393 );
or ( n40395 , n40357 , n40394 );
and ( n40396 , n40338 , n40395 );
or ( n40397 , n40337 , n40396 );
and ( n40398 , n40321 , n40397 );
or ( n40399 , n40320 , n40398 );
and ( n40400 , n40299 , n40399 );
or ( n40401 , n40298 , n40400 );
and ( n40402 , n40273 , n40401 );
or ( n40403 , n40272 , n40402 );
and ( n40404 , n40257 , n40403 );
or ( n40405 , n40256 , n40404 );
and ( n40406 , n40214 , n40405 );
or ( n40407 , n40213 , n40406 );
and ( n40408 , n40188 , n40407 );
or ( n40409 , n40187 , n40408 );
and ( n40410 , n40146 , n40409 );
or ( n40411 , n40145 , n40410 );
and ( n40412 , n40103 , n40411 );
or ( n40413 , n40102 , n40412 );
and ( n40414 , n40057 , n40413 );
or ( n40415 , n40056 , n40414 );
and ( n40416 , n40012 , n40415 );
or ( n40417 , n40011 , n40416 );
and ( n40418 , n39943 , n40417 );
or ( n40419 , n39942 , n40418 );
and ( n40420 , n39886 , n40419 );
or ( n40421 , n39885 , n40420 );
and ( n40422 , n39852 , n40421 );
or ( n40423 , n39851 , n40422 );
and ( n40424 , n39783 , n40423 );
or ( n40425 , n39782 , n40424 );
and ( n40426 , n39682 , n40425 );
or ( n40427 , n39681 , n40426 );
and ( n40428 , n39626 , n40427 );
or ( n40429 , n39625 , n40428 );
and ( n40430 , n39538 , n40429 );
or ( n40431 , n39537 , n40430 );
and ( n40432 , n39471 , n40431 );
or ( n40433 , n39470 , n40432 );
and ( n40434 , n39353 , n40433 );
or ( n40435 , n39352 , n40434 );
and ( n40436 , n39266 , n40435 );
or ( n40437 , n39265 , n40436 );
and ( n40438 , n39144 , n40437 );
or ( n40439 , n39143 , n40438 );
and ( n40440 , n39047 , n40439 );
or ( n40441 , n39046 , n40440 );
and ( n40442 , n38951 , n40441 );
or ( n40443 , n38950 , n40442 );
and ( n40444 , n38861 , n40443 );
or ( n40445 , n38860 , n40444 );
and ( n40446 , n38706 , n40445 );
or ( n40447 , n38705 , n40446 );
and ( n40448 , n38583 , n40447 );
or ( n40449 , n38582 , n40448 );
and ( n40450 , n38420 , n40449 );
or ( n40451 , n38419 , n40450 );
and ( n40452 , n38398 , n40451 );
or ( n40453 , n38397 , n40452 );
and ( n40454 , n38226 , n40453 );
or ( n40455 , n38225 , n40454 );
and ( n40456 , n38070 , n40455 );
or ( n40457 , n38069 , n40456 );
and ( n40458 , n37954 , n40457 );
or ( n40459 , n37953 , n40458 );
and ( n40460 , n37829 , n40459 );
or ( n40461 , n37828 , n40460 );
and ( n40462 , n37707 , n40461 );
or ( n40463 , n37706 , n40462 );
and ( n40464 , n37554 , n40463 );
or ( n40465 , n37553 , n40464 );
and ( n40466 , n37338 , n40465 );
or ( n40467 , n37337 , n40466 );
and ( n40468 , n37122 , n40467 );
or ( n40469 , n37121 , n40468 );
and ( n40470 , n37023 , n40469 );
or ( n40471 , n37022 , n40470 );
and ( n40472 , n36766 , n40471 );
or ( n40473 , n36765 , n40472 );
and ( n40474 , n36708 , n40473 );
or ( n40475 , n36707 , n40474 );
and ( n40476 , n36503 , n40475 );
or ( n40477 , n36502 , n40476 );
and ( n40478 , n36231 , n40477 );
or ( n40479 , n36230 , n40478 );
and ( n40480 , n36052 , n40479 );
or ( n40481 , n36051 , n40480 );
and ( n40482 , n35897 , n40481 );
or ( n40483 , n35896 , n40482 );
and ( n40484 , n35647 , n40483 );
or ( n40485 , n35646 , n40484 );
and ( n40486 , n35531 , n40485 );
or ( n40487 , n35530 , n40486 );
and ( n40488 , n35176 , n40487 );
or ( n40489 , n35175 , n40488 );
and ( n40490 , n35011 , n40489 );
or ( n40491 , n35010 , n40490 );
and ( n40492 , n34743 , n40491 );
or ( n40493 , n34742 , n40492 );
and ( n40494 , n34663 , n40493 );
or ( n40495 , n34662 , n40494 );
and ( n40496 , n34264 , n40495 );
or ( n40497 , n34263 , n40496 );
and ( n40498 , n34038 , n40497 );
or ( n40499 , n34037 , n40498 );
and ( n40500 , n33794 , n40499 );
or ( n40501 , n33793 , n40500 );
and ( n40502 , n33549 , n40501 );
or ( n40503 , n33548 , n40502 );
and ( n40504 , n33411 , n40503 );
or ( n40505 , n33410 , n40504 );
and ( n40506 , n33104 , n40505 );
or ( n40507 , n33103 , n40506 );
and ( n40508 , n32965 , n40507 );
or ( n40509 , n32964 , n40508 );
and ( n40510 , n32514 , n40509 );
or ( n40511 , n32513 , n40510 );
and ( n40512 , n32264 , n40511 );
or ( n40513 , n32263 , n40512 );
and ( n40514 , n32004 , n40513 );
or ( n40515 , n32003 , n40514 );
and ( n40516 , n31724 , n40515 );
or ( n40517 , n31723 , n40516 );
and ( n40518 , n31367 , n40517 );
or ( n40519 , n31366 , n40518 );
and ( n40520 , n31142 , n40519 );
or ( n40521 , n31141 , n40520 );
and ( n40522 , n30775 , n40521 );
or ( n40523 , n30774 , n40522 );
and ( n40524 , n30525 , n40523 );
or ( n40525 , n30524 , n40524 );
and ( n40526 , n30188 , n40525 );
or ( n40527 , n30187 , n40526 );
and ( n40528 , n29815 , n40527 );
or ( n40529 , n29814 , n40528 );
and ( n40530 , n29545 , n40529 );
or ( n40531 , n29544 , n40530 );
and ( n40532 , n29229 , n40531 );
or ( n40533 , n29228 , n40532 );
and ( n40534 , n28955 , n40533 );
or ( n40535 , n28954 , n40534 );
and ( n40536 , n28590 , n40535 );
or ( n40537 , n28589 , n40536 );
and ( n40538 , n28301 , n40537 );
or ( n40539 , n28300 , n40538 );
and ( n40540 , n27977 , n40539 );
or ( n40541 , n27976 , n40540 );
and ( n40542 , n27684 , n40541 );
or ( n40543 , n27683 , n40542 );
and ( n40544 , n27410 , n40543 );
or ( n40545 , n27409 , n40544 );
and ( n40546 , n27123 , n40545 );
or ( n40547 , n27122 , n40546 );
and ( n40548 , n26839 , n40547 );
or ( n40549 , n26838 , n40548 );
and ( n40550 , n26572 , n40549 );
or ( n40551 , n26571 , n40550 );
and ( n40552 , n26216 , n40551 );
or ( n40553 , n26215 , n40552 );
and ( n40554 , n25962 , n40553 );
or ( n40555 , n25961 , n40554 );
and ( n40556 , n25737 , n40555 );
or ( n40557 , n25736 , n40556 );
and ( n40558 , n25444 , n40557 );
or ( n40559 , n25443 , n40558 );
and ( n40560 , n25222 , n40559 );
or ( n40561 , n25221 , n40560 );
and ( n40562 , n25009 , n40561 );
or ( n40563 , n25008 , n40562 );
and ( n40564 , n24749 , n40563 );
or ( n40565 , n24748 , n40564 );
and ( n40566 , n24354 , n40565 );
or ( n40567 , n24353 , n40566 );
and ( n40568 , n24217 , n40567 );
or ( n40569 , n24216 , n40568 );
and ( n40570 , n24033 , n40569 );
or ( n40571 , n24032 , n40570 );
and ( n40572 , n23783 , n40571 );
or ( n40573 , n23782 , n40572 );
and ( n40574 , n23543 , n40573 );
or ( n40575 , n23542 , n40574 );
and ( n40576 , n23337 , n40575 );
or ( n40577 , n23336 , n40576 );
and ( n40578 , n23091 , n40577 );
or ( n40579 , n23090 , n40578 );
and ( n40580 , n22795 , n40579 );
or ( n40581 , n22794 , n40580 );
and ( n40582 , n22676 , n40581 );
or ( n40583 , n22675 , n40582 );
and ( n40584 , n22533 , n40583 );
or ( n40585 , n22532 , n40584 );
and ( n40586 , n22341 , n40585 );
or ( n40587 , n22340 , n40586 );
and ( n40588 , n22042 , n40587 );
or ( n40589 , n22041 , n40588 );
and ( n40590 , n22012 , n40589 );
or ( n40591 , n22011 , n40590 );
and ( n40592 , n21836 , n40591 );
or ( n40593 , n21835 , n40592 );
and ( n40594 , n21682 , n40593 );
or ( n40595 , n21681 , n40594 );
and ( n40596 , n21423 , n40595 );
or ( n40597 , n21422 , n40596 );
and ( n40598 , n21274 , n40597 );
or ( n40599 , n21273 , n40598 );
and ( n40600 , n21132 , n40599 );
or ( n40601 , n21131 , n40600 );
and ( n40602 , n21060 , n40601 );
or ( n40603 , n21059 , n40602 );
and ( n40604 , n20916 , n40603 );
or ( n40605 , n20915 , n40604 );
and ( n40606 , n20773 , n40605 );
or ( n40607 , n20772 , n40606 );
and ( n40608 , n20654 , n40607 );
or ( n40609 , n20653 , n40608 );
and ( n40610 , n20535 , n40609 );
or ( n40611 , n20534 , n40610 );
and ( n40612 , n20423 , n40611 );
or ( n40613 , n20422 , n40612 );
and ( n40614 , n20256 , n40613 );
or ( n40615 , n20255 , n40614 );
and ( n40616 , n20168 , n40615 );
or ( n40617 , n20167 , n40616 );
and ( n40618 , n20110 , n40617 );
or ( n40619 , n20109 , n40618 );
and ( n40620 , n19990 , n40619 );
or ( n40621 , n19989 , n40620 );
and ( n40622 , n19934 , n40621 );
or ( n40623 , n19933 , n40622 );
and ( n40624 , n19851 , n40623 );
or ( n40625 , n19850 , n40624 );
and ( n40626 , n19743 , n40625 );
or ( n40627 , n19742 , n40626 );
and ( n40628 , n19684 , n40627 );
or ( n40629 , n19683 , n40628 );
and ( n40630 , n19625 , n40629 );
or ( n40631 , n19624 , n40630 );
and ( n40632 , n19575 , n40631 );
or ( n40633 , n19574 , n40632 );
and ( n40634 , n19538 , n40633 );
or ( n40635 , n19537 , n40634 );
and ( n40636 , n19482 , n40635 );
or ( n40637 , n19481 , n40636 );
xor ( n40638 , n19453 , n40637 );
buf ( n40639 , n40638 );
xor ( n40640 , n19482 , n40635 );
buf ( n40641 , n40640 );
xor ( n40642 , n19538 , n40633 );
buf ( n40643 , n40642 );
xor ( n40644 , n19575 , n40631 );
buf ( n40645 , n40644 );
xor ( n40646 , n19625 , n40629 );
buf ( n40647 , n40646 );
xor ( n40648 , n19684 , n40627 );
buf ( n40649 , n40648 );
xor ( n40650 , n19743 , n40625 );
buf ( n40651 , n40650 );
xor ( n40652 , n19851 , n40623 );
buf ( n40653 , n40652 );
xor ( n40654 , n19934 , n40621 );
buf ( n40655 , n40654 );
xor ( n40656 , n19990 , n40619 );
buf ( n40657 , n40656 );
xor ( n40658 , n20110 , n40617 );
buf ( n40659 , n40658 );
xor ( n40660 , n20168 , n40615 );
buf ( n40661 , n40660 );
xor ( n40662 , n20256 , n40613 );
buf ( n40663 , n40662 );
xor ( n40664 , n20423 , n40611 );
buf ( n40665 , n40664 );
xor ( n40666 , n20535 , n40609 );
buf ( n40667 , n40666 );
xor ( n40668 , n20654 , n40607 );
buf ( n40669 , n40668 );
xor ( n40670 , n20773 , n40605 );
buf ( n40671 , n40670 );
xor ( n40672 , n20916 , n40603 );
buf ( n40673 , n40672 );
xor ( n40674 , n21060 , n40601 );
buf ( n40675 , n40674 );
xor ( n40676 , n21132 , n40599 );
buf ( n40677 , n40676 );
xor ( n40678 , n21274 , n40597 );
buf ( n40679 , n40678 );
xor ( n40680 , n21423 , n40595 );
buf ( n40681 , n40680 );
xor ( n40682 , n21682 , n40593 );
buf ( n40683 , n40682 );
xor ( n40684 , n21836 , n40591 );
buf ( n40685 , n40684 );
xor ( n40686 , n22012 , n40589 );
buf ( n40687 , n40686 );
xor ( n40688 , n22042 , n40587 );
buf ( n40689 , n40688 );
xor ( n40690 , n22341 , n40585 );
buf ( n40691 , n40690 );
xor ( n40692 , n22533 , n40583 );
buf ( n40693 , n40692 );
xor ( n40694 , n22676 , n40581 );
buf ( n40695 , n40694 );
xor ( n40696 , n22795 , n40579 );
buf ( n40697 , n40696 );
xor ( n40698 , n23091 , n40577 );
buf ( n40699 , n40698 );
xor ( n40700 , n23337 , n40575 );
buf ( n40701 , n40700 );
xor ( n40702 , n23543 , n40573 );
buf ( n40703 , n40702 );
xor ( n40704 , n23783 , n40571 );
buf ( n40705 , n40704 );
xor ( n40706 , n24033 , n40569 );
buf ( n40707 , n40706 );
xor ( n40708 , n24217 , n40567 );
buf ( n40709 , n40708 );
xor ( n40710 , n24354 , n40565 );
buf ( n40711 , n40710 );
xor ( n40712 , n24749 , n40563 );
buf ( n40713 , n40712 );
xor ( n40714 , n25009 , n40561 );
buf ( n40715 , n40714 );
xor ( n40716 , n25222 , n40559 );
buf ( n40717 , n40716 );
xor ( n40718 , n25444 , n40557 );
buf ( n40719 , n40718 );
xor ( n40720 , n25737 , n40555 );
buf ( n40721 , n40720 );
xor ( n40722 , n25962 , n40553 );
buf ( n40723 , n40722 );
xor ( n40724 , n26216 , n40551 );
buf ( n40725 , n40724 );
xor ( n40726 , n26572 , n40549 );
buf ( n40727 , n40726 );
xor ( n40728 , n26839 , n40547 );
buf ( n40729 , n40728 );
xor ( n40730 , n27123 , n40545 );
buf ( n40731 , n40730 );
xor ( n40732 , n27410 , n40543 );
buf ( n40733 , n40732 );
xor ( n40734 , n27684 , n40541 );
buf ( n40735 , n40734 );
xor ( n40736 , n27977 , n40539 );
buf ( n40737 , n40736 );
xor ( n40738 , n28301 , n40537 );
buf ( n40739 , n40738 );
xor ( n40740 , n28590 , n40535 );
buf ( n40741 , n40740 );
xor ( n40742 , n28955 , n40533 );
buf ( n40743 , n40742 );
xor ( n40744 , n29229 , n40531 );
buf ( n40745 , n40744 );
xor ( n40746 , n29545 , n40529 );
buf ( n40747 , n40746 );
xor ( n40748 , n29815 , n40527 );
buf ( n40749 , n40748 );
xor ( n40750 , n30188 , n40525 );
buf ( n40751 , n40750 );
xor ( n40752 , n30525 , n40523 );
buf ( n40753 , n40752 );
xor ( n40754 , n30775 , n40521 );
buf ( n40755 , n40754 );
xor ( n40756 , n31142 , n40519 );
buf ( n40757 , n40756 );
xor ( n40758 , n31367 , n40517 );
buf ( n40759 , n40758 );
xor ( n40760 , n31724 , n40515 );
buf ( n40761 , n40760 );
xor ( n40762 , n32004 , n40513 );
buf ( n40763 , n40762 );
xor ( n40764 , n32264 , n40511 );
buf ( n40765 , n40764 );
xor ( n40766 , n32514 , n40509 );
buf ( n40767 , n40766 );
xor ( n40768 , n32965 , n40507 );
buf ( n40769 , n40768 );
xor ( n40770 , n33104 , n40505 );
buf ( n40771 , n40770 );
xor ( n40772 , n33411 , n40503 );
buf ( n40773 , n40772 );
xor ( n40774 , n33549 , n40501 );
buf ( n40775 , n40774 );
xor ( n40776 , n33794 , n40499 );
buf ( n40777 , n40776 );
xor ( n40778 , n34038 , n40497 );
buf ( n40779 , n40778 );
xor ( n40780 , n34264 , n40495 );
buf ( n40781 , n40780 );
xor ( n40782 , n34663 , n40493 );
buf ( n40783 , n40782 );
xor ( n40784 , n34743 , n40491 );
buf ( n40785 , n40784 );
xor ( n40786 , n35011 , n40489 );
buf ( n40787 , n40786 );
xor ( n40788 , n35176 , n40487 );
buf ( n40789 , n40788 );
xor ( n40790 , n35531 , n40485 );
buf ( n40791 , n40790 );
xor ( n40792 , n35647 , n40483 );
buf ( n40793 , n40792 );
xor ( n40794 , n35897 , n40481 );
buf ( n40795 , n40794 );
xor ( n40796 , n36052 , n40479 );
buf ( n40797 , n40796 );
xor ( n40798 , n36231 , n40477 );
buf ( n40799 , n40798 );
xor ( n40800 , n36503 , n40475 );
buf ( n40801 , n40800 );
xor ( n40802 , n36708 , n40473 );
buf ( n40803 , n40802 );
xor ( n40804 , n36766 , n40471 );
buf ( n40805 , n40804 );
xor ( n40806 , n37023 , n40469 );
buf ( n40807 , n40806 );
xor ( n40808 , n37122 , n40467 );
buf ( n40809 , n40808 );
xor ( n40810 , n37338 , n40465 );
buf ( n40811 , n40810 );
xor ( n40812 , n37554 , n40463 );
buf ( n40813 , n40812 );
xor ( n40814 , n37707 , n40461 );
buf ( n40815 , n40814 );
xor ( n40816 , n37829 , n40459 );
buf ( n40817 , n40816 );
xor ( n40818 , n37954 , n40457 );
buf ( n40819 , n40818 );
xor ( n40820 , n38070 , n40455 );
buf ( n40821 , n40820 );
xor ( n40822 , n38226 , n40453 );
buf ( n40823 , n40822 );
xor ( n40824 , n38398 , n40451 );
buf ( n40825 , n40824 );
xor ( n40826 , n38420 , n40449 );
buf ( n40827 , n40826 );
xor ( n40828 , n38583 , n40447 );
buf ( n40829 , n40828 );
xor ( n40830 , n38706 , n40445 );
buf ( n40831 , n40830 );
xor ( n40832 , n38861 , n40443 );
buf ( n40833 , n40832 );
xor ( n40834 , n38951 , n40441 );
buf ( n40835 , n40834 );
xor ( n40836 , n39047 , n40439 );
buf ( n40837 , n40836 );
xor ( n40838 , n39144 , n40437 );
buf ( n40839 , n40838 );
xor ( n40840 , n39266 , n40435 );
buf ( n40841 , n40840 );
xor ( n40842 , n39353 , n40433 );
buf ( n40843 , n40842 );
xor ( n40844 , n39471 , n40431 );
buf ( n40845 , n40844 );
xor ( n40846 , n39538 , n40429 );
buf ( n40847 , n40846 );
xor ( n40848 , n39626 , n40427 );
buf ( n40849 , n40848 );
xor ( n40850 , n39682 , n40425 );
buf ( n40851 , n40850 );
xor ( n40852 , n39783 , n40423 );
buf ( n40853 , n40852 );
xor ( n40854 , n39852 , n40421 );
buf ( n40855 , n40854 );
xor ( n40856 , n39886 , n40419 );
buf ( n40857 , n40856 );
xor ( n40858 , n39943 , n40417 );
buf ( n40859 , n40858 );
xor ( n40860 , n40012 , n40415 );
buf ( n40861 , n40860 );
xor ( n40862 , n40057 , n40413 );
buf ( n40863 , n40862 );
xor ( n40864 , n40103 , n40411 );
buf ( n40865 , n40864 );
xor ( n40866 , n40146 , n40409 );
buf ( n40867 , n40866 );
xor ( n40868 , n40188 , n40407 );
buf ( n40869 , n40868 );
xor ( n40870 , n40214 , n40405 );
buf ( n40871 , n40870 );
xor ( n40872 , n40257 , n40403 );
buf ( n40873 , n40872 );
xor ( n40874 , n40273 , n40401 );
buf ( n40875 , n40874 );
xor ( n40876 , n40299 , n40399 );
buf ( n40877 , n40876 );
xor ( n40878 , n40321 , n40397 );
buf ( n40879 , n40878 );
xor ( n40880 , n40338 , n40395 );
buf ( n40881 , n40880 );
xor ( n40882 , n40358 , n40393 );
buf ( n40883 , n40882 );
xor ( n40884 , n40366 , n40391 );
buf ( n40885 , n40884 );
xor ( n40886 , n40373 , n40389 );
buf ( n40887 , n40886 );
xor ( n40888 , n40379 , n40387 );
buf ( n40889 , n40888 );
xor ( n40890 , n40383 , n40386 );
buf ( n40891 , n40890 );
buf ( n40892 , n40384 );
buf ( n40893 , n40892 );
buf ( n40894 , n19282 );
buf ( n40895 , n19240 );
buf ( n40896 , n19186 );
buf ( n40897 , n19124 );
buf ( n40898 , n19050 );
buf ( n40899 , n18968 );
buf ( n40900 , n18874 );
buf ( n40901 , n18772 );
buf ( n40902 , n18658 );
buf ( n40903 , n18536 );
buf ( n40904 , n18402 );
buf ( n40905 , n18260 );
buf ( n40906 , n18106 );
buf ( n40907 , n17944 );
buf ( n40908 , n17770 );
buf ( n40909 , n17588 );
buf ( n40910 , n17394 );
buf ( n40911 , n17192 );
buf ( n40912 , n16978 );
buf ( n40913 , n16756 );
buf ( n40914 , n16522 );
buf ( n40915 , n16280 );
buf ( n40916 , n16026 );
buf ( n40917 , n15764 );
buf ( n40918 , n15490 );
buf ( n40919 , n15208 );
buf ( n40920 , n14914 );
buf ( n40921 , n14612 );
buf ( n40922 , n14298 );
buf ( n40923 , n13976 );
buf ( n40924 , n13646 );
buf ( n40925 , n13324 );
buf ( n40926 , n12996 );
buf ( n40927 , n12642 );
buf ( n40928 , n12316 );
buf ( n40929 , n11982 );
buf ( n40930 , n11676 );
buf ( n40931 , n11362 );
buf ( n40932 , n11076 );
buf ( n40933 , n10782 );
buf ( n40934 , n10516 );
buf ( n40935 , n10242 );
buf ( n40936 , n9996 );
buf ( n40937 , n9742 );
buf ( n40938 , n9516 );
buf ( n40939 , n9282 );
buf ( n40940 , n9076 );
buf ( n40941 , n8862 );
buf ( n40942 , n8676 );
buf ( n40943 , n8482 );
buf ( n40944 , n8316 );
buf ( n40945 , n8142 );
buf ( n40946 , n7996 );
buf ( n40947 , n7842 );
buf ( n40948 , n7716 );
buf ( n40949 , n7582 );
buf ( n40950 , n7476 );
buf ( n40951 , n7362 );
buf ( n40952 , n7276 );
buf ( n40953 , n6804 );
buf ( n40954 , n6806 );
buf ( n40955 , n6808 );
buf ( n40956 , n6810 );
buf ( n40957 , n6812 );
buf ( n40958 , n6814 );
buf ( n40959 , n6816 );
buf ( n40960 , n6818 );
buf ( n40961 , n6820 );
buf ( n40962 , n6822 );
buf ( n40963 , n6824 );
buf ( n40964 , n6826 );
buf ( n40965 , n6828 );
buf ( n40966 , n6830 );
buf ( n40967 , n6832 );
buf ( n40968 , n6834 );
buf ( n40969 , n6836 );
buf ( n40970 , n6838 );
buf ( n40971 , n6840 );
buf ( n40972 , n6842 );
buf ( n40973 , n6844 );
buf ( n40974 , n6846 );
buf ( n40975 , n6848 );
buf ( n40976 , n6850 );
buf ( n40977 , n6852 );
buf ( n40978 , n6854 );
buf ( n40979 , n6856 );
buf ( n40980 , n6858 );
buf ( n40981 , n6860 );
buf ( n40982 , n6862 );
buf ( n40983 , n6864 );
buf ( n40984 , n6866 );
buf ( n40985 , n6868 );
buf ( n40986 , n6870 );
buf ( n40987 , n6872 );
buf ( n40988 , n6874 );
buf ( n40989 , n6876 );
buf ( n40990 , n6878 );
buf ( n40991 , n6880 );
buf ( n40992 , n6882 );
buf ( n40993 , n6884 );
buf ( n40994 , n6886 );
buf ( n40995 , n6888 );
buf ( n40996 , n6890 );
buf ( n40997 , n6892 );
buf ( n40998 , n6894 );
buf ( n40999 , n6896 );
buf ( n41000 , n6898 );
buf ( n41001 , n6900 );
buf ( n41002 , n6902 );
buf ( n41003 , n6904 );
buf ( n41004 , n6906 );
buf ( n41005 , n6908 );
buf ( n41006 , n6910 );
buf ( n41007 , n6912 );
buf ( n41008 , n6914 );
buf ( n41009 , n6916 );
buf ( n41010 , n6918 );
buf ( n41011 , n6920 );
buf ( n41012 , n6922 );
buf ( n41013 , n6924 );
buf ( n41014 , n6926 );
buf ( n41015 , n6928 );
buf ( n41016 , n6930 );
and ( n41017 , n40894 , n40958 );
and ( n41018 , n40895 , n40959 );
and ( n41019 , n40896 , n40960 );
and ( n41020 , n40897 , n40961 );
and ( n41021 , n40898 , n40962 );
and ( n41022 , n40899 , n40963 );
and ( n41023 , n40900 , n40964 );
and ( n41024 , n40901 , n40965 );
and ( n41025 , n40902 , n40966 );
and ( n41026 , n40903 , n40967 );
and ( n41027 , n40904 , n40968 );
and ( n41028 , n40905 , n40969 );
and ( n41029 , n40906 , n40970 );
and ( n41030 , n40907 , n40971 );
and ( n41031 , n40908 , n40972 );
and ( n41032 , n40909 , n40973 );
and ( n41033 , n40910 , n40974 );
and ( n41034 , n40911 , n40975 );
and ( n41035 , n40912 , n40976 );
and ( n41036 , n40913 , n40977 );
and ( n41037 , n40914 , n40978 );
and ( n41038 , n40915 , n40979 );
and ( n41039 , n40916 , n40980 );
and ( n41040 , n40917 , n40981 );
and ( n41041 , n40918 , n40982 );
and ( n41042 , n40919 , n40983 );
and ( n41043 , n40920 , n40984 );
and ( n41044 , n40921 , n40985 );
and ( n41045 , n40922 , n40986 );
and ( n41046 , n40923 , n40987 );
and ( n41047 , n40924 , n40988 );
and ( n41048 , n40925 , n40989 );
and ( n41049 , n40926 , n40990 );
and ( n41050 , n40927 , n40991 );
and ( n41051 , n40928 , n40992 );
and ( n41052 , n40929 , n40993 );
and ( n41053 , n40930 , n40994 );
and ( n41054 , n40931 , n40995 );
and ( n41055 , n40932 , n40996 );
and ( n41056 , n40933 , n40997 );
and ( n41057 , n40934 , n40998 );
and ( n41058 , n40935 , n40999 );
and ( n41059 , n40936 , n41000 );
and ( n41060 , n40937 , n41001 );
and ( n41061 , n40938 , n41002 );
and ( n41062 , n40939 , n41003 );
and ( n41063 , n40940 , n41004 );
and ( n41064 , n40941 , n41005 );
and ( n41065 , n40942 , n41006 );
and ( n41066 , n40943 , n41007 );
and ( n41067 , n40944 , n41008 );
and ( n41068 , n40945 , n41009 );
and ( n41069 , n40946 , n41010 );
and ( n41070 , n40947 , n41011 );
and ( n41071 , n40948 , n41012 );
and ( n41072 , n40949 , n41013 );
and ( n41073 , n40950 , n41014 );
and ( n41074 , n40951 , n41015 );
and ( n41075 , n40952 , n41016 );
and ( n41076 , n41015 , n41075 );
and ( n41077 , n40951 , n41075 );
or ( n41078 , n41074 , n41076 , n41077 );
and ( n41079 , n41014 , n41078 );
and ( n41080 , n40950 , n41078 );
or ( n41081 , n41073 , n41079 , n41080 );
and ( n41082 , n41013 , n41081 );
and ( n41083 , n40949 , n41081 );
or ( n41084 , n41072 , n41082 , n41083 );
and ( n41085 , n41012 , n41084 );
and ( n41086 , n40948 , n41084 );
or ( n41087 , n41071 , n41085 , n41086 );
and ( n41088 , n41011 , n41087 );
and ( n41089 , n40947 , n41087 );
or ( n41090 , n41070 , n41088 , n41089 );
and ( n41091 , n41010 , n41090 );
and ( n41092 , n40946 , n41090 );
or ( n41093 , n41069 , n41091 , n41092 );
and ( n41094 , n41009 , n41093 );
and ( n41095 , n40945 , n41093 );
or ( n41096 , n41068 , n41094 , n41095 );
and ( n41097 , n41008 , n41096 );
and ( n41098 , n40944 , n41096 );
or ( n41099 , n41067 , n41097 , n41098 );
and ( n41100 , n41007 , n41099 );
and ( n41101 , n40943 , n41099 );
or ( n41102 , n41066 , n41100 , n41101 );
and ( n41103 , n41006 , n41102 );
and ( n41104 , n40942 , n41102 );
or ( n41105 , n41065 , n41103 , n41104 );
and ( n41106 , n41005 , n41105 );
and ( n41107 , n40941 , n41105 );
or ( n41108 , n41064 , n41106 , n41107 );
and ( n41109 , n41004 , n41108 );
and ( n41110 , n40940 , n41108 );
or ( n41111 , n41063 , n41109 , n41110 );
and ( n41112 , n41003 , n41111 );
and ( n41113 , n40939 , n41111 );
or ( n41114 , n41062 , n41112 , n41113 );
and ( n41115 , n41002 , n41114 );
and ( n41116 , n40938 , n41114 );
or ( n41117 , n41061 , n41115 , n41116 );
and ( n41118 , n41001 , n41117 );
and ( n41119 , n40937 , n41117 );
or ( n41120 , n41060 , n41118 , n41119 );
and ( n41121 , n41000 , n41120 );
and ( n41122 , n40936 , n41120 );
or ( n41123 , n41059 , n41121 , n41122 );
and ( n41124 , n40999 , n41123 );
and ( n41125 , n40935 , n41123 );
or ( n41126 , n41058 , n41124 , n41125 );
and ( n41127 , n40998 , n41126 );
and ( n41128 , n40934 , n41126 );
or ( n41129 , n41057 , n41127 , n41128 );
and ( n41130 , n40997 , n41129 );
and ( n41131 , n40933 , n41129 );
or ( n41132 , n41056 , n41130 , n41131 );
and ( n41133 , n40996 , n41132 );
and ( n41134 , n40932 , n41132 );
or ( n41135 , n41055 , n41133 , n41134 );
and ( n41136 , n40995 , n41135 );
and ( n41137 , n40931 , n41135 );
or ( n41138 , n41054 , n41136 , n41137 );
and ( n41139 , n40994 , n41138 );
and ( n41140 , n40930 , n41138 );
or ( n41141 , n41053 , n41139 , n41140 );
and ( n41142 , n40993 , n41141 );
and ( n41143 , n40929 , n41141 );
or ( n41144 , n41052 , n41142 , n41143 );
and ( n41145 , n40992 , n41144 );
and ( n41146 , n40928 , n41144 );
or ( n41147 , n41051 , n41145 , n41146 );
and ( n41148 , n40991 , n41147 );
and ( n41149 , n40927 , n41147 );
or ( n41150 , n41050 , n41148 , n41149 );
and ( n41151 , n40990 , n41150 );
and ( n41152 , n40926 , n41150 );
or ( n41153 , n41049 , n41151 , n41152 );
and ( n41154 , n40989 , n41153 );
and ( n41155 , n40925 , n41153 );
or ( n41156 , n41048 , n41154 , n41155 );
and ( n41157 , n40988 , n41156 );
and ( n41158 , n40924 , n41156 );
or ( n41159 , n41047 , n41157 , n41158 );
and ( n41160 , n40987 , n41159 );
and ( n41161 , n40923 , n41159 );
or ( n41162 , n41046 , n41160 , n41161 );
and ( n41163 , n40986 , n41162 );
and ( n41164 , n40922 , n41162 );
or ( n41165 , n41045 , n41163 , n41164 );
and ( n41166 , n40985 , n41165 );
and ( n41167 , n40921 , n41165 );
or ( n41168 , n41044 , n41166 , n41167 );
and ( n41169 , n40984 , n41168 );
and ( n41170 , n40920 , n41168 );
or ( n41171 , n41043 , n41169 , n41170 );
and ( n41172 , n40983 , n41171 );
and ( n41173 , n40919 , n41171 );
or ( n41174 , n41042 , n41172 , n41173 );
and ( n41175 , n40982 , n41174 );
and ( n41176 , n40918 , n41174 );
or ( n41177 , n41041 , n41175 , n41176 );
and ( n41178 , n40981 , n41177 );
and ( n41179 , n40917 , n41177 );
or ( n41180 , n41040 , n41178 , n41179 );
and ( n41181 , n40980 , n41180 );
and ( n41182 , n40916 , n41180 );
or ( n41183 , n41039 , n41181 , n41182 );
and ( n41184 , n40979 , n41183 );
and ( n41185 , n40915 , n41183 );
or ( n41186 , n41038 , n41184 , n41185 );
and ( n41187 , n40978 , n41186 );
and ( n41188 , n40914 , n41186 );
or ( n41189 , n41037 , n41187 , n41188 );
and ( n41190 , n40977 , n41189 );
and ( n41191 , n40913 , n41189 );
or ( n41192 , n41036 , n41190 , n41191 );
and ( n41193 , n40976 , n41192 );
and ( n41194 , n40912 , n41192 );
or ( n41195 , n41035 , n41193 , n41194 );
and ( n41196 , n40975 , n41195 );
and ( n41197 , n40911 , n41195 );
or ( n41198 , n41034 , n41196 , n41197 );
and ( n41199 , n40974 , n41198 );
and ( n41200 , n40910 , n41198 );
or ( n41201 , n41033 , n41199 , n41200 );
and ( n41202 , n40973 , n41201 );
and ( n41203 , n40909 , n41201 );
or ( n41204 , n41032 , n41202 , n41203 );
and ( n41205 , n40972 , n41204 );
and ( n41206 , n40908 , n41204 );
or ( n41207 , n41031 , n41205 , n41206 );
and ( n41208 , n40971 , n41207 );
and ( n41209 , n40907 , n41207 );
or ( n41210 , n41030 , n41208 , n41209 );
and ( n41211 , n40970 , n41210 );
and ( n41212 , n40906 , n41210 );
or ( n41213 , n41029 , n41211 , n41212 );
and ( n41214 , n40969 , n41213 );
and ( n41215 , n40905 , n41213 );
or ( n41216 , n41028 , n41214 , n41215 );
and ( n41217 , n40968 , n41216 );
and ( n41218 , n40904 , n41216 );
or ( n41219 , n41027 , n41217 , n41218 );
and ( n41220 , n40967 , n41219 );
and ( n41221 , n40903 , n41219 );
or ( n41222 , n41026 , n41220 , n41221 );
and ( n41223 , n40966 , n41222 );
and ( n41224 , n40902 , n41222 );
or ( n41225 , n41025 , n41223 , n41224 );
and ( n41226 , n40965 , n41225 );
and ( n41227 , n40901 , n41225 );
or ( n41228 , n41024 , n41226 , n41227 );
and ( n41229 , n40964 , n41228 );
and ( n41230 , n40900 , n41228 );
or ( n41231 , n41023 , n41229 , n41230 );
and ( n41232 , n40963 , n41231 );
and ( n41233 , n40899 , n41231 );
or ( n41234 , n41022 , n41232 , n41233 );
and ( n41235 , n40962 , n41234 );
and ( n41236 , n40898 , n41234 );
or ( n41237 , n41021 , n41235 , n41236 );
and ( n41238 , n40961 , n41237 );
and ( n41239 , n40897 , n41237 );
or ( n41240 , n41020 , n41238 , n41239 );
and ( n41241 , n40960 , n41240 );
and ( n41242 , n40896 , n41240 );
or ( n41243 , n41019 , n41241 , n41242 );
and ( n41244 , n40959 , n41243 );
and ( n41245 , n40895 , n41243 );
or ( n41246 , n41018 , n41244 , n41245 );
and ( n41247 , n40958 , n41246 );
and ( n41248 , n40894 , n41246 );
or ( n41249 , n41017 , n41247 , n41248 );
and ( n41250 , n40957 , n41249 );
and ( n41251 , n40956 , n41250 );
and ( n41252 , n40955 , n41251 );
and ( n41253 , n40954 , n41252 );
xor ( n41254 , n40953 , n41253 );
buf ( n41255 , n41254 );
xor ( n41256 , n40954 , n41252 );
buf ( n41257 , n41256 );
xor ( n41258 , n40955 , n41251 );
buf ( n41259 , n41258 );
xor ( n41260 , n40956 , n41250 );
buf ( n41261 , n41260 );
xor ( n41262 , n40957 , n41249 );
buf ( n41263 , n41262 );
xor ( n41264 , n40894 , n40958 );
xor ( n41265 , n41264 , n41246 );
buf ( n41266 , n41265 );
xor ( n41267 , n40895 , n40959 );
xor ( n41268 , n41267 , n41243 );
buf ( n41269 , n41268 );
xor ( n41270 , n40896 , n40960 );
xor ( n41271 , n41270 , n41240 );
buf ( n41272 , n41271 );
xor ( n41273 , n40897 , n40961 );
xor ( n41274 , n41273 , n41237 );
buf ( n41275 , n41274 );
xor ( n41276 , n40898 , n40962 );
xor ( n41277 , n41276 , n41234 );
buf ( n41278 , n41277 );
xor ( n41279 , n40899 , n40963 );
xor ( n41280 , n41279 , n41231 );
buf ( n41281 , n41280 );
xor ( n41282 , n40900 , n40964 );
xor ( n41283 , n41282 , n41228 );
buf ( n41284 , n41283 );
xor ( n41285 , n40901 , n40965 );
xor ( n41286 , n41285 , n41225 );
buf ( n41287 , n41286 );
xor ( n41288 , n40902 , n40966 );
xor ( n41289 , n41288 , n41222 );
buf ( n41290 , n41289 );
xor ( n41291 , n40903 , n40967 );
xor ( n41292 , n41291 , n41219 );
buf ( n41293 , n41292 );
xor ( n41294 , n40904 , n40968 );
xor ( n41295 , n41294 , n41216 );
buf ( n41296 , n41295 );
xor ( n41297 , n40905 , n40969 );
xor ( n41298 , n41297 , n41213 );
buf ( n41299 , n41298 );
xor ( n41300 , n40906 , n40970 );
xor ( n41301 , n41300 , n41210 );
buf ( n41302 , n41301 );
xor ( n41303 , n40907 , n40971 );
xor ( n41304 , n41303 , n41207 );
buf ( n41305 , n41304 );
xor ( n41306 , n40908 , n40972 );
xor ( n41307 , n41306 , n41204 );
buf ( n41308 , n41307 );
xor ( n41309 , n40909 , n40973 );
xor ( n41310 , n41309 , n41201 );
buf ( n41311 , n41310 );
xor ( n41312 , n40910 , n40974 );
xor ( n41313 , n41312 , n41198 );
buf ( n41314 , n41313 );
xor ( n41315 , n40911 , n40975 );
xor ( n41316 , n41315 , n41195 );
buf ( n41317 , n41316 );
xor ( n41318 , n40912 , n40976 );
xor ( n41319 , n41318 , n41192 );
buf ( n41320 , n41319 );
xor ( n41321 , n40913 , n40977 );
xor ( n41322 , n41321 , n41189 );
buf ( n41323 , n41322 );
xor ( n41324 , n40914 , n40978 );
xor ( n41325 , n41324 , n41186 );
buf ( n41326 , n41325 );
xor ( n41327 , n40915 , n40979 );
xor ( n41328 , n41327 , n41183 );
buf ( n41329 , n41328 );
xor ( n41330 , n40916 , n40980 );
xor ( n41331 , n41330 , n41180 );
buf ( n41332 , n41331 );
xor ( n41333 , n40917 , n40981 );
xor ( n41334 , n41333 , n41177 );
buf ( n41335 , n41334 );
xor ( n41336 , n40918 , n40982 );
xor ( n41337 , n41336 , n41174 );
buf ( n41338 , n41337 );
xor ( n41339 , n40919 , n40983 );
xor ( n41340 , n41339 , n41171 );
buf ( n41341 , n41340 );
xor ( n41342 , n40920 , n40984 );
xor ( n41343 , n41342 , n41168 );
buf ( n41344 , n41343 );
xor ( n41345 , n40921 , n40985 );
xor ( n41346 , n41345 , n41165 );
buf ( n41347 , n41346 );
xor ( n41348 , n40922 , n40986 );
xor ( n41349 , n41348 , n41162 );
buf ( n41350 , n41349 );
xor ( n41351 , n40923 , n40987 );
xor ( n41352 , n41351 , n41159 );
buf ( n41353 , n41352 );
xor ( n41354 , n40924 , n40988 );
xor ( n41355 , n41354 , n41156 );
buf ( n41356 , n41355 );
xor ( n41357 , n40925 , n40989 );
xor ( n41358 , n41357 , n41153 );
buf ( n41359 , n41358 );
xor ( n41360 , n40926 , n40990 );
xor ( n41361 , n41360 , n41150 );
buf ( n41362 , n41361 );
xor ( n41363 , n40927 , n40991 );
xor ( n41364 , n41363 , n41147 );
buf ( n41365 , n41364 );
xor ( n41366 , n40928 , n40992 );
xor ( n41367 , n41366 , n41144 );
buf ( n41368 , n41367 );
xor ( n41369 , n40929 , n40993 );
xor ( n41370 , n41369 , n41141 );
buf ( n41371 , n41370 );
xor ( n41372 , n40930 , n40994 );
xor ( n41373 , n41372 , n41138 );
buf ( n41374 , n41373 );
xor ( n41375 , n40931 , n40995 );
xor ( n41376 , n41375 , n41135 );
buf ( n41377 , n41376 );
xor ( n41378 , n40932 , n40996 );
xor ( n41379 , n41378 , n41132 );
buf ( n41380 , n41379 );
xor ( n41381 , n40933 , n40997 );
xor ( n41382 , n41381 , n41129 );
buf ( n41383 , n41382 );
xor ( n41384 , n40934 , n40998 );
xor ( n41385 , n41384 , n41126 );
buf ( n41386 , n41385 );
xor ( n41387 , n40935 , n40999 );
xor ( n41388 , n41387 , n41123 );
buf ( n41389 , n41388 );
xor ( n41390 , n40936 , n41000 );
xor ( n41391 , n41390 , n41120 );
buf ( n41392 , n41391 );
xor ( n41393 , n40937 , n41001 );
xor ( n41394 , n41393 , n41117 );
buf ( n41395 , n41394 );
xor ( n41396 , n40938 , n41002 );
xor ( n41397 , n41396 , n41114 );
buf ( n41398 , n41397 );
xor ( n41399 , n40939 , n41003 );
xor ( n41400 , n41399 , n41111 );
buf ( n41401 , n41400 );
xor ( n41402 , n40940 , n41004 );
xor ( n41403 , n41402 , n41108 );
buf ( n41404 , n41403 );
xor ( n41405 , n40941 , n41005 );
xor ( n41406 , n41405 , n41105 );
buf ( n41407 , n41406 );
xor ( n41408 , n40942 , n41006 );
xor ( n41409 , n41408 , n41102 );
buf ( n41410 , n41409 );
xor ( n41411 , n40943 , n41007 );
xor ( n41412 , n41411 , n41099 );
buf ( n41413 , n41412 );
xor ( n41414 , n40944 , n41008 );
xor ( n41415 , n41414 , n41096 );
buf ( n41416 , n41415 );
xor ( n41417 , n40945 , n41009 );
xor ( n41418 , n41417 , n41093 );
buf ( n41419 , n41418 );
xor ( n41420 , n40946 , n41010 );
xor ( n41421 , n41420 , n41090 );
buf ( n41422 , n41421 );
xor ( n41423 , n40947 , n41011 );
xor ( n41424 , n41423 , n41087 );
buf ( n41425 , n41424 );
xor ( n41426 , n40948 , n41012 );
xor ( n41427 , n41426 , n41084 );
buf ( n41428 , n41427 );
xor ( n41429 , n40949 , n41013 );
xor ( n41430 , n41429 , n41081 );
buf ( n41431 , n41430 );
xor ( n41432 , n40950 , n41014 );
xor ( n41433 , n41432 , n41078 );
buf ( n41434 , n41433 );
xor ( n41435 , n40951 , n41015 );
xor ( n41436 , n41435 , n41075 );
buf ( n41437 , n41436 );
xor ( n41438 , n40952 , n41016 );
buf ( n41439 , n41438 );
buf ( n41440 , n19278 );
buf ( n41441 , n19236 );
buf ( n41442 , n19182 );
buf ( n41443 , n19120 );
buf ( n41444 , n19046 );
buf ( n41445 , n18964 );
buf ( n41446 , n18870 );
buf ( n41447 , n18768 );
buf ( n41448 , n18654 );
buf ( n41449 , n18532 );
buf ( n41450 , n18398 );
buf ( n41451 , n18256 );
buf ( n41452 , n18102 );
buf ( n41453 , n17940 );
buf ( n41454 , n17766 );
buf ( n41455 , n17584 );
buf ( n41456 , n17390 );
buf ( n41457 , n17188 );
buf ( n41458 , n16974 );
buf ( n41459 , n16752 );
buf ( n41460 , n16518 );
buf ( n41461 , n16276 );
buf ( n41462 , n16022 );
buf ( n41463 , n15760 );
buf ( n41464 , n15486 );
buf ( n41465 , n15204 );
buf ( n41466 , n14910 );
buf ( n41467 , n14608 );
buf ( n41468 , n14294 );
buf ( n41469 , n13972 );
buf ( n41470 , n13642 );
buf ( n41471 , n13320 );
buf ( n41472 , n12992 );
buf ( n41473 , n12638 );
buf ( n41474 , n12312 );
buf ( n41475 , n11978 );
buf ( n41476 , n11672 );
buf ( n41477 , n11358 );
buf ( n41478 , n11072 );
buf ( n41479 , n10778 );
buf ( n41480 , n10512 );
buf ( n41481 , n10238 );
buf ( n41482 , n9992 );
buf ( n41483 , n9738 );
buf ( n41484 , n9512 );
buf ( n41485 , n9278 );
buf ( n41486 , n9072 );
buf ( n41487 , n8858 );
buf ( n41488 , n8672 );
buf ( n41489 , n8478 );
buf ( n41490 , n8312 );
buf ( n41491 , n8138 );
buf ( n41492 , n7992 );
buf ( n41493 , n7838 );
buf ( n41494 , n7712 );
buf ( n41495 , n7578 );
buf ( n41496 , n7472 );
buf ( n41497 , n7358 );
buf ( n41498 , n7272 );
buf ( n41499 , n19282 );
buf ( n41500 , n19240 );
buf ( n41501 , n19186 );
buf ( n41502 , n19124 );
buf ( n41503 , n19050 );
buf ( n41504 , n18968 );
buf ( n41505 , n18874 );
buf ( n41506 , n18772 );
buf ( n41507 , n18658 );
buf ( n41508 , n18536 );
buf ( n41509 , n18402 );
buf ( n41510 , n18260 );
buf ( n41511 , n18106 );
buf ( n41512 , n17944 );
buf ( n41513 , n17770 );
buf ( n41514 , n17588 );
buf ( n41515 , n17394 );
buf ( n41516 , n17192 );
buf ( n41517 , n16978 );
buf ( n41518 , n16756 );
buf ( n41519 , n16522 );
buf ( n41520 , n16280 );
buf ( n41521 , n16026 );
buf ( n41522 , n15764 );
buf ( n41523 , n15490 );
buf ( n41524 , n15208 );
buf ( n41525 , n14914 );
buf ( n41526 , n14612 );
buf ( n41527 , n14298 );
buf ( n41528 , n13976 );
buf ( n41529 , n13646 );
buf ( n41530 , n13324 );
buf ( n41531 , n12996 );
buf ( n41532 , n12642 );
buf ( n41533 , n12316 );
buf ( n41534 , n11982 );
buf ( n41535 , n11676 );
buf ( n41536 , n11362 );
buf ( n41537 , n11076 );
buf ( n41538 , n10782 );
buf ( n41539 , n10516 );
buf ( n41540 , n10242 );
buf ( n41541 , n9996 );
buf ( n41542 , n9742 );
buf ( n41543 , n9516 );
buf ( n41544 , n9282 );
buf ( n41545 , n9076 );
buf ( n41546 , n8862 );
buf ( n41547 , n8676 );
buf ( n41548 , n8482 );
buf ( n41549 , n8316 );
buf ( n41550 , n8142 );
buf ( n41551 , n7996 );
buf ( n41552 , n7842 );
buf ( n41553 , n7716 );
buf ( n41554 , n7582 );
buf ( n41555 , n7476 );
buf ( n41556 , n7362 );
buf ( n41557 , n7276 );
buf ( n41558 , n7182 );
buf ( n41559 , n7116 );
buf ( n41560 , n7042 );
buf ( n41561 , n6996 );
buf ( n41562 , n6952 );
and ( n41563 , n41440 , n41504 );
and ( n41564 , n41441 , n41505 );
and ( n41565 , n41442 , n41506 );
and ( n41566 , n41443 , n41507 );
and ( n41567 , n41444 , n41508 );
and ( n41568 , n41445 , n41509 );
and ( n41569 , n41446 , n41510 );
and ( n41570 , n41447 , n41511 );
and ( n41571 , n41448 , n41512 );
and ( n41572 , n41449 , n41513 );
and ( n41573 , n41450 , n41514 );
and ( n41574 , n41451 , n41515 );
and ( n41575 , n41452 , n41516 );
and ( n41576 , n41453 , n41517 );
and ( n41577 , n41454 , n41518 );
and ( n41578 , n41455 , n41519 );
and ( n41579 , n41456 , n41520 );
and ( n41580 , n41457 , n41521 );
and ( n41581 , n41458 , n41522 );
and ( n41582 , n41459 , n41523 );
and ( n41583 , n41460 , n41524 );
and ( n41584 , n41461 , n41525 );
and ( n41585 , n41462 , n41526 );
and ( n41586 , n41463 , n41527 );
and ( n41587 , n41464 , n41528 );
and ( n41588 , n41465 , n41529 );
and ( n41589 , n41466 , n41530 );
and ( n41590 , n41467 , n41531 );
and ( n41591 , n41468 , n41532 );
and ( n41592 , n41469 , n41533 );
and ( n41593 , n41470 , n41534 );
and ( n41594 , n41471 , n41535 );
and ( n41595 , n41472 , n41536 );
and ( n41596 , n41473 , n41537 );
and ( n41597 , n41474 , n41538 );
and ( n41598 , n41475 , n41539 );
and ( n41599 , n41476 , n41540 );
and ( n41600 , n41477 , n41541 );
and ( n41601 , n41478 , n41542 );
and ( n41602 , n41479 , n41543 );
and ( n41603 , n41480 , n41544 );
and ( n41604 , n41481 , n41545 );
and ( n41605 , n41482 , n41546 );
and ( n41606 , n41483 , n41547 );
and ( n41607 , n41484 , n41548 );
and ( n41608 , n41485 , n41549 );
and ( n41609 , n41486 , n41550 );
and ( n41610 , n41487 , n41551 );
and ( n41611 , n41488 , n41552 );
and ( n41612 , n41489 , n41553 );
and ( n41613 , n41490 , n41554 );
and ( n41614 , n41491 , n41555 );
and ( n41615 , n41492 , n41556 );
and ( n41616 , n41493 , n41557 );
and ( n41617 , n41494 , n41558 );
and ( n41618 , n41495 , n41559 );
and ( n41619 , n41496 , n41560 );
and ( n41620 , n41497 , n41561 );
and ( n41621 , n41498 , n41562 );
and ( n41622 , n41561 , n41621 );
and ( n41623 , n41497 , n41621 );
or ( n41624 , n41620 , n41622 , n41623 );
and ( n41625 , n41560 , n41624 );
and ( n41626 , n41496 , n41624 );
or ( n41627 , n41619 , n41625 , n41626 );
and ( n41628 , n41559 , n41627 );
and ( n41629 , n41495 , n41627 );
or ( n41630 , n41618 , n41628 , n41629 );
and ( n41631 , n41558 , n41630 );
and ( n41632 , n41494 , n41630 );
or ( n41633 , n41617 , n41631 , n41632 );
and ( n41634 , n41557 , n41633 );
and ( n41635 , n41493 , n41633 );
or ( n41636 , n41616 , n41634 , n41635 );
and ( n41637 , n41556 , n41636 );
and ( n41638 , n41492 , n41636 );
or ( n41639 , n41615 , n41637 , n41638 );
and ( n41640 , n41555 , n41639 );
and ( n41641 , n41491 , n41639 );
or ( n41642 , n41614 , n41640 , n41641 );
and ( n41643 , n41554 , n41642 );
and ( n41644 , n41490 , n41642 );
or ( n41645 , n41613 , n41643 , n41644 );
and ( n41646 , n41553 , n41645 );
and ( n41647 , n41489 , n41645 );
or ( n41648 , n41612 , n41646 , n41647 );
and ( n41649 , n41552 , n41648 );
and ( n41650 , n41488 , n41648 );
or ( n41651 , n41611 , n41649 , n41650 );
and ( n41652 , n41551 , n41651 );
and ( n41653 , n41487 , n41651 );
or ( n41654 , n41610 , n41652 , n41653 );
and ( n41655 , n41550 , n41654 );
and ( n41656 , n41486 , n41654 );
or ( n41657 , n41609 , n41655 , n41656 );
and ( n41658 , n41549 , n41657 );
and ( n41659 , n41485 , n41657 );
or ( n41660 , n41608 , n41658 , n41659 );
and ( n41661 , n41548 , n41660 );
and ( n41662 , n41484 , n41660 );
or ( n41663 , n41607 , n41661 , n41662 );
and ( n41664 , n41547 , n41663 );
and ( n41665 , n41483 , n41663 );
or ( n41666 , n41606 , n41664 , n41665 );
and ( n41667 , n41546 , n41666 );
and ( n41668 , n41482 , n41666 );
or ( n41669 , n41605 , n41667 , n41668 );
and ( n41670 , n41545 , n41669 );
and ( n41671 , n41481 , n41669 );
or ( n41672 , n41604 , n41670 , n41671 );
and ( n41673 , n41544 , n41672 );
and ( n41674 , n41480 , n41672 );
or ( n41675 , n41603 , n41673 , n41674 );
and ( n41676 , n41543 , n41675 );
and ( n41677 , n41479 , n41675 );
or ( n41678 , n41602 , n41676 , n41677 );
and ( n41679 , n41542 , n41678 );
and ( n41680 , n41478 , n41678 );
or ( n41681 , n41601 , n41679 , n41680 );
and ( n41682 , n41541 , n41681 );
and ( n41683 , n41477 , n41681 );
or ( n41684 , n41600 , n41682 , n41683 );
and ( n41685 , n41540 , n41684 );
and ( n41686 , n41476 , n41684 );
or ( n41687 , n41599 , n41685 , n41686 );
and ( n41688 , n41539 , n41687 );
and ( n41689 , n41475 , n41687 );
or ( n41690 , n41598 , n41688 , n41689 );
and ( n41691 , n41538 , n41690 );
and ( n41692 , n41474 , n41690 );
or ( n41693 , n41597 , n41691 , n41692 );
and ( n41694 , n41537 , n41693 );
and ( n41695 , n41473 , n41693 );
or ( n41696 , n41596 , n41694 , n41695 );
and ( n41697 , n41536 , n41696 );
and ( n41698 , n41472 , n41696 );
or ( n41699 , n41595 , n41697 , n41698 );
and ( n41700 , n41535 , n41699 );
and ( n41701 , n41471 , n41699 );
or ( n41702 , n41594 , n41700 , n41701 );
and ( n41703 , n41534 , n41702 );
and ( n41704 , n41470 , n41702 );
or ( n41705 , n41593 , n41703 , n41704 );
and ( n41706 , n41533 , n41705 );
and ( n41707 , n41469 , n41705 );
or ( n41708 , n41592 , n41706 , n41707 );
and ( n41709 , n41532 , n41708 );
and ( n41710 , n41468 , n41708 );
or ( n41711 , n41591 , n41709 , n41710 );
and ( n41712 , n41531 , n41711 );
and ( n41713 , n41467 , n41711 );
or ( n41714 , n41590 , n41712 , n41713 );
and ( n41715 , n41530 , n41714 );
and ( n41716 , n41466 , n41714 );
or ( n41717 , n41589 , n41715 , n41716 );
and ( n41718 , n41529 , n41717 );
and ( n41719 , n41465 , n41717 );
or ( n41720 , n41588 , n41718 , n41719 );
and ( n41721 , n41528 , n41720 );
and ( n41722 , n41464 , n41720 );
or ( n41723 , n41587 , n41721 , n41722 );
and ( n41724 , n41527 , n41723 );
and ( n41725 , n41463 , n41723 );
or ( n41726 , n41586 , n41724 , n41725 );
and ( n41727 , n41526 , n41726 );
and ( n41728 , n41462 , n41726 );
or ( n41729 , n41585 , n41727 , n41728 );
and ( n41730 , n41525 , n41729 );
and ( n41731 , n41461 , n41729 );
or ( n41732 , n41584 , n41730 , n41731 );
and ( n41733 , n41524 , n41732 );
and ( n41734 , n41460 , n41732 );
or ( n41735 , n41583 , n41733 , n41734 );
and ( n41736 , n41523 , n41735 );
and ( n41737 , n41459 , n41735 );
or ( n41738 , n41582 , n41736 , n41737 );
and ( n41739 , n41522 , n41738 );
and ( n41740 , n41458 , n41738 );
or ( n41741 , n41581 , n41739 , n41740 );
and ( n41742 , n41521 , n41741 );
and ( n41743 , n41457 , n41741 );
or ( n41744 , n41580 , n41742 , n41743 );
and ( n41745 , n41520 , n41744 );
and ( n41746 , n41456 , n41744 );
or ( n41747 , n41579 , n41745 , n41746 );
and ( n41748 , n41519 , n41747 );
and ( n41749 , n41455 , n41747 );
or ( n41750 , n41578 , n41748 , n41749 );
and ( n41751 , n41518 , n41750 );
and ( n41752 , n41454 , n41750 );
or ( n41753 , n41577 , n41751 , n41752 );
and ( n41754 , n41517 , n41753 );
and ( n41755 , n41453 , n41753 );
or ( n41756 , n41576 , n41754 , n41755 );
and ( n41757 , n41516 , n41756 );
and ( n41758 , n41452 , n41756 );
or ( n41759 , n41575 , n41757 , n41758 );
and ( n41760 , n41515 , n41759 );
and ( n41761 , n41451 , n41759 );
or ( n41762 , n41574 , n41760 , n41761 );
and ( n41763 , n41514 , n41762 );
and ( n41764 , n41450 , n41762 );
or ( n41765 , n41573 , n41763 , n41764 );
and ( n41766 , n41513 , n41765 );
and ( n41767 , n41449 , n41765 );
or ( n41768 , n41572 , n41766 , n41767 );
and ( n41769 , n41512 , n41768 );
and ( n41770 , n41448 , n41768 );
or ( n41771 , n41571 , n41769 , n41770 );
and ( n41772 , n41511 , n41771 );
and ( n41773 , n41447 , n41771 );
or ( n41774 , n41570 , n41772 , n41773 );
and ( n41775 , n41510 , n41774 );
and ( n41776 , n41446 , n41774 );
or ( n41777 , n41569 , n41775 , n41776 );
and ( n41778 , n41509 , n41777 );
and ( n41779 , n41445 , n41777 );
or ( n41780 , n41568 , n41778 , n41779 );
and ( n41781 , n41508 , n41780 );
and ( n41782 , n41444 , n41780 );
or ( n41783 , n41567 , n41781 , n41782 );
and ( n41784 , n41507 , n41783 );
and ( n41785 , n41443 , n41783 );
or ( n41786 , n41566 , n41784 , n41785 );
and ( n41787 , n41506 , n41786 );
and ( n41788 , n41442 , n41786 );
or ( n41789 , n41565 , n41787 , n41788 );
and ( n41790 , n41505 , n41789 );
and ( n41791 , n41441 , n41789 );
or ( n41792 , n41564 , n41790 , n41791 );
and ( n41793 , n41504 , n41792 );
and ( n41794 , n41440 , n41792 );
or ( n41795 , n41563 , n41793 , n41794 );
and ( n41796 , n41503 , n41795 );
and ( n41797 , n41502 , n41796 );
and ( n41798 , n41501 , n41797 );
and ( n41799 , n41500 , n41798 );
xor ( n41800 , n41499 , n41799 );
buf ( n41801 , n41800 );
xor ( n41802 , n41500 , n41798 );
buf ( n41803 , n41802 );
xor ( n41804 , n41501 , n41797 );
buf ( n41805 , n41804 );
xor ( n41806 , n41502 , n41796 );
buf ( n41807 , n41806 );
xor ( n41808 , n41503 , n41795 );
buf ( n41809 , n41808 );
xor ( n41810 , n41440 , n41504 );
xor ( n41811 , n41810 , n41792 );
buf ( n41812 , n41811 );
xor ( n41813 , n41441 , n41505 );
xor ( n41814 , n41813 , n41789 );
buf ( n41815 , n41814 );
xor ( n41816 , n41442 , n41506 );
xor ( n41817 , n41816 , n41786 );
buf ( n41818 , n41817 );
xor ( n41819 , n41443 , n41507 );
xor ( n41820 , n41819 , n41783 );
buf ( n41821 , n41820 );
xor ( n41822 , n41444 , n41508 );
xor ( n41823 , n41822 , n41780 );
buf ( n41824 , n41823 );
xor ( n41825 , n41445 , n41509 );
xor ( n41826 , n41825 , n41777 );
buf ( n41827 , n41826 );
xor ( n41828 , n41446 , n41510 );
xor ( n41829 , n41828 , n41774 );
buf ( n41830 , n41829 );
xor ( n41831 , n41447 , n41511 );
xor ( n41832 , n41831 , n41771 );
buf ( n41833 , n41832 );
xor ( n41834 , n41448 , n41512 );
xor ( n41835 , n41834 , n41768 );
buf ( n41836 , n41835 );
xor ( n41837 , n41449 , n41513 );
xor ( n41838 , n41837 , n41765 );
buf ( n41839 , n41838 );
xor ( n41840 , n41450 , n41514 );
xor ( n41841 , n41840 , n41762 );
buf ( n41842 , n41841 );
xor ( n41843 , n41451 , n41515 );
xor ( n41844 , n41843 , n41759 );
buf ( n41845 , n41844 );
xor ( n41846 , n41452 , n41516 );
xor ( n41847 , n41846 , n41756 );
buf ( n41848 , n41847 );
xor ( n41849 , n41453 , n41517 );
xor ( n41850 , n41849 , n41753 );
buf ( n41851 , n41850 );
xor ( n41852 , n41454 , n41518 );
xor ( n41853 , n41852 , n41750 );
buf ( n41854 , n41853 );
xor ( n41855 , n41455 , n41519 );
xor ( n41856 , n41855 , n41747 );
buf ( n41857 , n41856 );
xor ( n41858 , n41456 , n41520 );
xor ( n41859 , n41858 , n41744 );
buf ( n41860 , n41859 );
xor ( n41861 , n41457 , n41521 );
xor ( n41862 , n41861 , n41741 );
buf ( n41863 , n41862 );
xor ( n41864 , n41458 , n41522 );
xor ( n41865 , n41864 , n41738 );
buf ( n41866 , n41865 );
xor ( n41867 , n41459 , n41523 );
xor ( n41868 , n41867 , n41735 );
buf ( n41869 , n41868 );
xor ( n41870 , n41460 , n41524 );
xor ( n41871 , n41870 , n41732 );
buf ( n41872 , n41871 );
xor ( n41873 , n41461 , n41525 );
xor ( n41874 , n41873 , n41729 );
buf ( n41875 , n41874 );
xor ( n41876 , n41462 , n41526 );
xor ( n41877 , n41876 , n41726 );
buf ( n41878 , n41877 );
xor ( n41879 , n41463 , n41527 );
xor ( n41880 , n41879 , n41723 );
buf ( n41881 , n41880 );
xor ( n41882 , n41464 , n41528 );
xor ( n41883 , n41882 , n41720 );
buf ( n41884 , n41883 );
xor ( n41885 , n41465 , n41529 );
xor ( n41886 , n41885 , n41717 );
buf ( n41887 , n41886 );
xor ( n41888 , n41466 , n41530 );
xor ( n41889 , n41888 , n41714 );
buf ( n41890 , n41889 );
xor ( n41891 , n41467 , n41531 );
xor ( n41892 , n41891 , n41711 );
buf ( n41893 , n41892 );
xor ( n41894 , n41468 , n41532 );
xor ( n41895 , n41894 , n41708 );
buf ( n41896 , n41895 );
xor ( n41897 , n41469 , n41533 );
xor ( n41898 , n41897 , n41705 );
buf ( n41899 , n41898 );
xor ( n41900 , n41470 , n41534 );
xor ( n41901 , n41900 , n41702 );
buf ( n41902 , n41901 );
xor ( n41903 , n41471 , n41535 );
xor ( n41904 , n41903 , n41699 );
buf ( n41905 , n41904 );
xor ( n41906 , n41472 , n41536 );
xor ( n41907 , n41906 , n41696 );
buf ( n41908 , n41907 );
xor ( n41909 , n41473 , n41537 );
xor ( n41910 , n41909 , n41693 );
buf ( n41911 , n41910 );
xor ( n41912 , n41474 , n41538 );
xor ( n41913 , n41912 , n41690 );
buf ( n41914 , n41913 );
xor ( n41915 , n41475 , n41539 );
xor ( n41916 , n41915 , n41687 );
buf ( n41917 , n41916 );
xor ( n41918 , n41476 , n41540 );
xor ( n41919 , n41918 , n41684 );
buf ( n41920 , n41919 );
xor ( n41921 , n41477 , n41541 );
xor ( n41922 , n41921 , n41681 );
buf ( n41923 , n41922 );
xor ( n41924 , n41478 , n41542 );
xor ( n41925 , n41924 , n41678 );
buf ( n41926 , n41925 );
xor ( n41927 , n41479 , n41543 );
xor ( n41928 , n41927 , n41675 );
buf ( n41929 , n41928 );
xor ( n41930 , n41480 , n41544 );
xor ( n41931 , n41930 , n41672 );
buf ( n41932 , n41931 );
xor ( n41933 , n41481 , n41545 );
xor ( n41934 , n41933 , n41669 );
buf ( n41935 , n41934 );
xor ( n41936 , n41482 , n41546 );
xor ( n41937 , n41936 , n41666 );
buf ( n41938 , n41937 );
xor ( n41939 , n41483 , n41547 );
xor ( n41940 , n41939 , n41663 );
buf ( n41941 , n41940 );
xor ( n41942 , n41484 , n41548 );
xor ( n41943 , n41942 , n41660 );
buf ( n41944 , n41943 );
xor ( n41945 , n41485 , n41549 );
xor ( n41946 , n41945 , n41657 );
buf ( n41947 , n41946 );
xor ( n41948 , n41486 , n41550 );
xor ( n41949 , n41948 , n41654 );
buf ( n41950 , n41949 );
xor ( n41951 , n41487 , n41551 );
xor ( n41952 , n41951 , n41651 );
buf ( n41953 , n41952 );
xor ( n41954 , n41488 , n41552 );
xor ( n41955 , n41954 , n41648 );
buf ( n41956 , n41955 );
xor ( n41957 , n41489 , n41553 );
xor ( n41958 , n41957 , n41645 );
buf ( n41959 , n41958 );
xor ( n41960 , n41490 , n41554 );
xor ( n41961 , n41960 , n41642 );
buf ( n41962 , n41961 );
xor ( n41963 , n41491 , n41555 );
xor ( n41964 , n41963 , n41639 );
buf ( n41965 , n41964 );
xor ( n41966 , n41492 , n41556 );
xor ( n41967 , n41966 , n41636 );
buf ( n41968 , n41967 );
xor ( n41969 , n41493 , n41557 );
xor ( n41970 , n41969 , n41633 );
buf ( n41971 , n41970 );
xor ( n41972 , n41494 , n41558 );
xor ( n41973 , n41972 , n41630 );
buf ( n41974 , n41973 );
xor ( n41975 , n41495 , n41559 );
xor ( n41976 , n41975 , n41627 );
buf ( n41977 , n41976 );
xor ( n41978 , n41496 , n41560 );
xor ( n41979 , n41978 , n41624 );
buf ( n41980 , n41979 );
xor ( n41981 , n41497 , n41561 );
xor ( n41982 , n41981 , n41621 );
buf ( n41983 , n41982 );
xor ( n41984 , n41498 , n41562 );
buf ( n41985 , n41984 );
endmodule
