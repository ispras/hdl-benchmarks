module mul_11_11_1(a, b, c);
  input [10:0] a;
  input [10:0] b;
  output c;
  assign c = a * b;
endmodule
