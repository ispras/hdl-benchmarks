//NOTE: no-implementation module stub

module GTECH_NOT (
    output Z,
    input A
);

endmodule
