//NOTE: no-implementation module stub

module Delaya (
    input wire DSack,
    output reg delDSack
);

endmodule
