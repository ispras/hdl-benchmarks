// IWLS benchmark module "i10" printed on Wed May 29 16:34:21 2002
module i10(\V32(0) , \V32(1) , \V32(2) , \V32(3) , \V56(0) , \V289(0) , \V10(0) , \V13(0) , \V35(0) , \V203(0) , \V288(6) , \V288(7) , \V248(0) , \V249(0) , \V62(0) , \V59(0) , \V174(0) , \V215(0) , \V66(0) , \V70(0) , \V43(0) , \V214(0) , \V37(0) , \V271(0) , \V40(0) , \V45(0) , \V149(7) , \V149(6) , \V149(5) , \V149(4) , \V1(0) , \V7(0) , \V34(0) , \V243(0) , \V244(0) , \V245(0) , \V246(0) , \V247(0) , \V293(0) , \V302(0) , \V270(0) , \V269(0) , \V274(0) , \V202(0) , \V275(0) , \V257(7) , \V257(5) , \V257(3) , \V257(1) , \V257(2) , \V257(4) , \V257(6) , \V9(0) , \V149(0) , \V149(1) , \V149(2) , \V149(3) , \V169(1) , \V165(0) , \V165(2) , \V165(4) , \V165(5) , \V165(6) , \V165(7) , \V165(1) , \V88(2) , \V88(3) , \V55(0) , \V169(0) , \V52(0) , \V5(0) , \V6(0) , \V12(0) , \V11(0) , \V4(0) , \V165(3) , \V51(0) , \V65(0) , \V290(0) , \V279(0) , \V280(0) , \V288(4) , \V288(2) , \V288(0) , \V258(0) , \V229(5) , \V229(4) , \V229(3) , \V229(2) , \V229(1) , \V229(0) , \V223(5) , \V223(4) , \V223(3) , \V223(2) , \V223(1) , \V223(0) , \V189(5) , \V189(4) , \V189(3) , \V189(2) , \V189(1) , \V189(0) , \V183(5) , \V183(4) , \V183(3) , \V183(2) , \V183(1) , \V183(0) , \V239(4) , \V239(3) , \V239(2) , \V239(1) , \V239(0) , \V234(4) , \V234(3) , \V234(2) , \V234(1) , \V234(0) , \V199(4) , \V199(3) , \V199(2) , \V199(1) , \V199(0) , \V194(4) , \V194(3) , \V194(2) , \V194(1) , \V194(0) , \V257(0) , \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(11) , \V32(10) , \V32(9) , \V88(1) , \V88(0) , \V84(5) , \V84(4) , \V84(3) , \V84(2) , \V84(1) , \V84(0) , \V78(5) , \V78(4) , \V2(0) , \V3(0) , \V14(0) , \V213(0) , \V213(5) , \V213(4) , \V213(3) , \V213(2) , \V213(1) , \V268(5) , \V268(3) , \V268(1) , \V268(2) , \V268(4) , \V8(0) , \V60(0) , \V53(0) , \V57(0) , \V109(0) , \V277(0) , \V278(0) , \V259(0) , \V260(0) , \V67(0) , \V68(0) , \V69(0) , \V216(0) , \V175(0) , \V177(0) , \V172(0) , \V171(0) , \V50(0) , \V63(0) , \V71(0) , \V292(0) , \V291(0) , \V91(0) , \V91(1) , \V294(0) , \V207(0) , \V295(0) , \V204(0) , \V205(0) , \V261(0) , \V262(0) , \V100(0) , \V100(5) , \V100(4) , \V100(3) , \V100(2) , \V100(1) , \V240(0) , \V242(0) , \V241(0) , \V33(0) , \V16(0) , \V15(0) , \V101(0) , \V268(0) , \V288(1) , \V288(3) , \V288(5) , \V301(0) , \V108(0) , \V108(1) , \V108(2) , \V108(3) , \V108(4) , \V108(5) , \V124(5) , \V124(4) , \V124(3) , \V124(2) , \V124(1) , \V124(0) , \V132(7) , \V132(6) , \V132(5) , \V132(4) , \V132(3) , \V132(2) , \V132(1) , \V132(0) , \V118(5) , \V118(4) , \V118(3) , \V118(2) , \V118(1) , \V118(0) , \V118(7) , \V118(6) , \V46(0) , \V48(0) , \V102(0) , \V110(0) , \V134(1) , \V134(0) , \V272(0) , \V78(2) , \V78(3) , \V39(0) , \V38(0) , \V42(0) , \V44(0) , \V41(0) , \V78(1) , \V78(0) , \V94(0) , \V94(1) , \V321(2) , V356, V357, V373, \V375(0) , V377, \V393(0) , \V398(0) , \V410(0) , \V423(0) , V432, \V435(0) , \V500(0) , \V508(0) , \V511(0) , V512, V527, V537, V538, V539, V540, V541, V542, V543, V544, V545, V546, V547, V548, \V572(9) , \V572(8) , \V572(7) , \V572(6) , \V572(5) , \V572(4) , \V572(3) , \V572(2) , \V572(1) , \V572(0) , \V585(0) , V587, \V591(0) , \V597(0) , \V603(0) , \V609(0) , V620, V621, V630, \V634(0) , \V640(0) , V657, V707, V763, V775, V778, V779, V780, V781, V782, V783, V784, V787, V789, \V798(0) , V801, \V802(0) , \V821(0) , \V826(0) , V966, V986, \V1213(11) , \V1213(10) , \V1213(9) , \V1213(8) , \V1213(7) , \V1213(6) , \V1213(5) , \V1213(4) , \V1213(3) , \V1213(2) , \V1213(1) , \V1213(0) , \V1243(9) , \V1243(8) , \V1243(7) , \V1243(6) , \V1243(5) , \V1243(4) , \V1243(3) , \V1243(2) , \V1243(1) , \V1243(0) , V1256, V1257, V1258, V1259, V1260, V1261, V1262, V1263, V1264, V1265, V1266, V1267, \V1274(0) , \V1281(0) , \V1297(4) , \V1297(3) , \V1297(2) , \V1297(1) , \V1297(0) , V1365, V1375, V1378, V1380, V1382, V1384, V1386, V1387, \V1392(0) , V1423, V1426, V1428, V1429, V1431, V1432, \V1439(0) , \V1440(0) , \V1451(0) , \V1459(0) , \V1467(0) , V1470, \V1480(0) , \V1481(0) , \V1492(0) , \V1495(0) , \V1512(3) , \V1512(2) , \V1512(1) , \V1536(0) , V1537, V1539, \V1552(1) , \V1552(0) , \V1613(0) , \V1613(1) , \V1620(0) , \V1629(0) , \V1645(0) , \V1652(0) , V1669, \V1671(0) , \V1679(0) , \V1693(0) , \V1709(4) , \V1709(3) , \V1709(2) , \V1709(1) , \V1709(0) , \V1717(0) , V1719, \V1726(0) , V1736, \V1741(0) , \V1745(0) , \V1757(0) , \V1758(0) , \V1759(0) , \V1760(0) , \V1771(1) , \V1771(0) , \V1781(1) , \V1781(0) , \V1829(9) , \V1829(8) , \V1829(7) , \V1829(6) , \V1829(5) , \V1829(4) , \V1829(3) , \V1829(2) , \V1829(1) , \V1829(0) , V1832, \V1833(0) , \V1863(0) , \V1864(0) , \V1896(0) , \V1897(0) , \V1898(0) , \V1899(0) , \V1900(0) , \V1901(0) , \V1921(5) , \V1921(4) , \V1921(3) , \V1921(2) , \V1921(1) , \V1921(0) , \V1953(1) , \V1953(7) , \V1953(6) , \V1953(5) , \V1953(4) , \V1953(3) , \V1953(2) , \V1953(0) , \V1960(1) , \V1960(0) , \V1968(0) , \V1992(1) , \V1992(0) , V650, V651, V652, V653, V654, V655, V656, V1370, V1371, V1372, V1373, V1374);
input
  \V223(1) ,
  \V223(0) ,
  \V100(3) ,
  \V100(2) ,
  \V100(5) ,
  \V100(4) ,
  \V100(1) ,
  \V100(0) ,
  \V60(0) ,
  \V247(0) ,
  \V7(0) ,
  \V124(3) ,
  \V124(2) ,
  \V124(5) ,
  \V124(4) ,
  \V11(0) ,
  \V124(1) ,
  \V124(0) ,
  \V259(0) ,
  \V84(0) ,
  \V84(1) ,
  \V84(2) ,
  \V84(3) ,
  \V84(4) ,
  \V84(5) ,
  \V35(0) ,
  \V302(0) ,
  \V59(0) ,
  \V240(0) ,
  \V203(0) ,
  \V288(3) ,
  \V215(0) ,
  \V288(2) ,
  \V288(5) ,
  \V288(4) ,
  \V40(0) ,
  \V288(1) ,
  \V288(0) ,
  \V165(3) ,
  \V165(2) ,
  \V165(5) ,
  \V165(4) ,
  \V239(3) ,
  \V288(7) ,
  \V239(2) ,
  \V288(6) ,
  \V52(0) ,
  \V165(1) ,
  \V239(4) ,
  \V165(0) ,
  \V239(1) ,
  \V239(0) ,
  \V165(7) ,
  \V165(6) ,
  \V177(0) ,
  \V189(3) ,
  \V189(2) ,
  \V189(5) ,
  \V189(4) ,
  \V189(1) ,
  \V189(0) ,
  \V15(0) ,
  \V88(0) ,
  \V88(1) ,
  \V88(2) ,
  \V88(3) ,
  \V39(0) ,
  \V293(0) ,
  \V244(0) ,
  \V4(0) ,
  \V194(3) ,
  \V194(2) ,
  \V194(4) ,
  \V268(3) ,
  \V268(2) ,
  \V268(5) ,
  \V194(1) ,
  \V268(4) ,
  \V194(0) ,
  \V268(1) ,
  \V268(0) ,
  \V207(0) ,
  \V32(0) ,
  \V32(1) ,
  \V32(2) ,
  \V32(3) ,
  \V32(4) ,
  \V32(5) ,
  \V32(6) ,
  \V32(7) ,
  \V32(8) ,
  \V44(0) ,
  \V32(9) ,
  \V108(3) ,
  \V108(2) ,
  \V56(0) ,
  \V108(5) ,
  \V108(4) ,
  \V169(1) ,
  \V169(0) ,
  \V108(1) ,
  \V108(0) ,
  \V68(0) ,
  \V261(0) ,
  \V101(0) ,
  \V174(0) ,
  \V248(0) ,
  \V8(0) ,
  \V12(0) ,
  \V149(3) ,
  \V149(2) ,
  \V149(5) ,
  \V149(4) ,
  \V149(1) ,
  \V149(0) ,
  \V149(7) ,
  \V149(6) ,
  \V48(0) ,
  \V290(0) ,
  \V32(11) ,
  \V32(10) ,
  \V241(0) ,
  \V1(0) ,
  \V204(0) ,
  \V277(0) ,
  \V216(0) ,
  \V41(0) ,
  \V289(0) ,
  \V53(0) ,
  \V65(0) ,
  \V16(0) ,
  \V270(0) ,
  \V294(0) ,
  \V171(0) ,
  \V183(3) ,
  \V110(0) ,
  \V183(2) ,
  \V245(0) ,
  \V183(5) ,
  \V5(0) ,
  \V183(4) ,
  \V257(3) ,
  \V257(2) ,
  \V70(0) ,
  \V257(5) ,
  \V183(1) ,
  \V257(4) ,
  \V183(0) ,
  \V257(1) ,
  \V257(0) ,
  \V257(7) ,
  \V257(6) ,
  \V134(1) ,
  \V134(0) ,
  \V269(0) ,
  \V94(0) ,
  \V94(1) ,
  \V33(0) ,
  \V45(0) ,
  \V57(0) ,
  \V109(0) ,
  \V69(0) ,
  \V262(0) ,
  \V213(3) ,
  \V213(2) ,
  \V213(5) ,
  \V213(4) ,
  \V274(0) ,
  \V213(1) ,
  \V213(0) ,
  \V50(0) ,
  \V102(0) ,
  \V62(0) ,
  \V175(0) ,
  \V249(0) ,
  \V9(0) ,
  \V13(0) ,
  \V199(3) ,
  \V199(2) ,
  \V199(4) ,
  \V199(1) ,
  \V199(0) ,
  \V37(0) ,
  \V291(0) ,
  \V242(0) ,
  \V2(0) ,
  \V205(0) ,
  \V91(0) ,
  \V91(1) ,
  \V278(0) ,
  \V229(3) ,
  \V229(2) ,
  \V42(0) ,
  \V229(5) ,
  \V229(4) ,
  \V229(1) ,
  \V229(0) ,
  \V118(3) ,
  \V118(2) ,
  \V66(0) ,
  \V118(5) ,
  \V118(4) ,
  \V118(1) ,
  \V118(0) ,
  \V78(0) ,
  \V78(1) ,
  \V118(7) ,
  \V78(2) ,
  \V118(6) ,
  \V78(3) ,
  \V78(4) ,
  \V78(5) ,
  \V271(0) ,
  \V234(3) ,
  \V234(2) ,
  \V234(4) ,
  \V295(0) ,
  \V234(1) ,
  \V234(0) ,
  \V172(0) ,
  \V246(0) ,
  \V6(0) ,
  \V71(0) ,
  \V10(0) ,
  \V258(0) ,
  \V34(0) ,
  \V46(0) ,
  \V301(0) ,
  \V202(0) ,
  \V275(0) ,
  \V214(0) ,
  \V51(0) ,
  \V63(0) ,
  \V14(0) ,
  \V38(0) ,
  \V280(0) ,
  \V292(0) ,
  \V243(0) ,
  \V3(0) ,
  \V132(3) ,
  \V132(2) ,
  \V132(5) ,
  \V132(4) ,
  \V132(1) ,
  \V132(0) ,
  \V132(7) ,
  \V132(6) ,
  \V279(0) ,
  \V43(0) ,
  \V55(0) ,
  \V67(0) ,
  \V260(0) ,
  \V272(0) ,
  \V223(3) ,
  \V223(2) ,
  \V223(5) ,
  \V223(4) ;
output
  \V1243(7) ,
  \V500(0) ,
  \V1243(6) ,
  \V1243(9) ,
  \V1243(8) ,
  \V1243(1) ,
  \V1243(0) ,
  \V1717(0) ,
  \V1243(3) ,
  \V1243(2) ,
  \V1243(5) ,
  \V1243(4) ,
  \V585(0) ,
  \V597(0) ,
  \V1679(0) ,
  \V1833(0) ,
  \V1968(0) ,
  \V1771(1) ,
  \V1771(0) ,
  \V640(0) ,
  \V375(0) ,
  \V603(0) ,
  \V1758(0) ,
  \V1900(0) ,
  \V1709(1) ,
  \V1709(0) ,
  \V1709(3) ,
  \V1709(2) ,
  \V1709(4) ,
  \V1512(1) ,
  \V1512(3) ,
  \V1512(2) ,
  \V1536(0) ,
  \V1898(0) ,
  \V1652(0) ,
  \V1726(0) ,
  \V1953(7) ,
  \V1953(6) ,
  \V410(0) ,
  \V1953(1) ,
  \V1953(0) ,
  \V1953(3) ,
  \V1953(2) ,
  \V1953(5) ,
  \V1953(4) ,
  \V508(0) ,
  \V1392(0) ,
  \V1829(7) ,
  \V1829(6) ,
  \V1829(9) ,
  \V1829(8) ,
  \V1281(0) ,
  \V1620(0) ,
  \V1829(1) ,
  \V1829(0) ,
  \V1829(3) ,
  \V1829(2) ,
  \V1693(0) ,
  \V1829(5) ,
  \V1829(4) ,
  \V1921(1) ,
  \V1921(0) ,
  \V1921(3) ,
  \V1921(2) ,
  \V1921(5) ,
  \V1921(4) ,
  \V802(0) ,
  \V826(0) ,
  \V1213(10) ,
  \V1213(11) ,
  \V1760(0) ,
  \V1495(0) ,
  \V591(0) ,
  \V1759(0) ,
  \V1901(0) ,
  \V1297(1) ,
  \V1297(0) ,
  \V1297(3) ,
  \V1297(2) ,
  \V1297(4) ,
  \V1451(0) ,
  \V1863(0) ,
  \V393(0) ,
  \V1899(0) ,
  \V1480(0) ,
  \V423(0) ,
  \V1492(0) ,
  \V435(0) ,
  \V1781(1) ,
  \V1781(0) ,
  V1256,
  V1257,
  V1258,
  V1259,
  V1260,
  V1261,
  V1262,
  V1263,
  V1264,
  V1265,
  V1266,
  V1267,
  \V1467(0) ,
  V1365,
  V1370,
  V1371,
  V1372,
  V1373,
  V1374,
  V1375,
  V1378,
  V1380,
  V1382,
  V1384,
  V1386,
  V1387,
  V1423,
  V1426,
  V1428,
  V1429,
  V1431,
  V1432,
  V1470,
  \V1645(0) ,
  V1537,
  V1539,
  V1669,
  V1719,
  \V1896(0) ,
  V1736,
  V1832,
  \V1459(0) ,
  \V1213(7) ,
  \V1213(6) ,
  \V1213(9) ,
  \V1213(8) ,
  \V1613(1) ,
  \V1274(0) ,
  \V1613(0) ,
  \V1213(1) ,
  \V1213(0) ,
  \V1213(3) ,
  \V1213(2) ,
  \V1213(5) ,
  \V1213(4) ,
  \V1440(0) ,
  \V321(2) ,
  \V1864(0) ,
  \V1741(0) ,
  \V572(3) ,
  \V572(2) ,
  \V634(0) ,
  \V572(5) ,
  \V572(4) ,
  \V1439(0) ,
  \V572(1) ,
  \V572(0) ,
  \V511(0) ,
  \V572(7) ,
  \V572(6) ,
  \V572(9) ,
  \V572(8) ,
  \V1992(1) ,
  \V1992(0) ,
  \V609(0) ,
  \V1481(0) ,
  \V1629(0) ,
  \V798(0) ,
  \V398(0) ,
  \V1671(0) ,
  \V1745(0) ,
  \V1757(0) ,
  \V1960(1) ,
  \V1960(0) ,
  V356,
  V357,
  V373,
  V377,
  \V1897(0) ,
  V432,
  V512,
  V527,
  V537,
  V538,
  V539,
  V540,
  V541,
  V542,
  V543,
  V544,
  V545,
  V546,
  V547,
  V548,
  V587,
  V620,
  V621,
  V630,
  V650,
  V651,
  V652,
  V653,
  V654,
  V655,
  V656,
  V657,
  \V821(0) ,
  \V1552(1) ,
  \V1552(0) ,
  V707,
  V763,
  V775,
  V778,
  V779,
  V780,
  V781,
  V782,
  V783,
  V784,
  V787,
  V789,
  V801,
  V966,
  V986;
wire
  \V758(0) ,
  \V1354(0) ,
  \V1631(0) ,
  \V709(1) ,
  \V709(0) ,
  \V912(0) ,
  \V985(0) ,
  \V450(0) ,
  \V924(0) ,
  \V659(0) ,
  \V1255(1) ,
  \V1255(0) ,
  \V1255(3) ,
  \V862(0) ,
  \V1255(2) ,
  \V536(0) ,
  \[200] ,
  \[201] ,
  \[202] ,
  \V874(0) ,
  \[203] ,
  \V1124(12) ,
  \[204] ,
  \V1124(13) ,
  \[205] ,
  \V813(0) ,
  \[206] ,
  \[207] ,
  \V413(0) ,
  \[208] ,
  \[209] ,
  \V1124(10) ,
  \V1124(11) ,
  \V1421(0) ,
  \[210] ,
  \[211] ,
  \V2033(0) ,
  \[212] ,
  \[213] ,
  \[214] ,
  \[215] ,
  \[216] ,
  \V363(0) ,
  \[217] ,
  \V837(0) ,
  \[218] ,
  \[219] ,
  \[220] ,
  \[221] ,
  \[222] ,
  \[223] ,
  \V1857(0) ,
  \V1069(7) ,
  \V1069(6) ,
  \V1069(9) ,
  \V1069(8) ,
  \V2008(0) ,
  \V1395(0) ,
  \V399(0) ,
  \V676(5) ,
  \V1334(0) ,
  \V676(4) ,
  \V1408(0) ,
  \V1069(5) ,
  \V1746(0) ,
  \V1069(4) ,
  \V676(7) ,
  \V676(6) ,
  \V1684(0) ,
  \V1623(0) ,
  \V965(0) ,
  \V904(0) ,
  \V504(0) ,
  \V639(0) ,
  \V842(0) ,
  \V1647(0) ,
  \V1124(7) ,
  \V1124(6) ,
  \V1124(9) ,
  \V1124(8) ,
  \V380(0) ,
  \V854(0) ,
  \V528(0) ,
  \V1124(1) ,
  \V1862(0) ,
  \V1124(3) ,
  \V731(0) ,
  \V1124(2) ,
  \V1124(5) ,
  \V1597(0) ,
  \V1124(4) ,
  \V405(0) ,
  \V681(3) ,
  \V681(5) ,
  \V681(4) ,
  \V817(0) ,
  \V1351(0) ,
  \V681(7) ,
  \V681(6) ,
  \V1086(1) ,
  \V1086(0) ,
  \V1086(3) ,
  \V1086(2) ,
  \V1763(1) ,
  \V1763(0) ,
  \V1498(0) ,
  \V1837(0) ,
  \V367(0) ,
  \V1437(0) ,
  \V982(0) ,
  \V933(0) ,
  \V533(0) ,
  \V1399(0) ,
  \V945(0) ,
  \V883(0) ,
  \V822(0) ,
  \V957(0) ,
  \V1553(0) ,
  \V895(0) ,
  \V1965(0) ,
  \V834(0) ,
  \V1565(0) ,
  \V1177(7) ,
  \V434(0) ,
  \V1177(6) ,
  \V1177(9) ,
  \V1177(8) ,
  \[10] ,
  \[11] ,
  \V1977(0) ,
  \[12] ,
  \[13] ,
  \V1442(0) ,
  \[14] ,
  \[15] ,
  \V1177(1) ,
  \[16] ,
  \V1177(0) ,
  \[17] ,
  \V1177(3) ,
  \[18] ,
  \V1177(2) ,
  \[19] ,
  \V1177(5) ,
  \V1854(0) ,
  \V1177(4) ,
  \V384(0) ,
  \[20] ,
  \[21] ,
  \[22] ,
  \V1866(0) ,
  \[23] ,
  \V396(0) ,
  \[24] ,
  \[25] ,
  \V1331(0) ,
  \[26] ,
  \V2078(0) ,
  \[27] ,
  \[28] ,
  \[29] ,
  \V612(0) ,
  \[30] ,
  \[31] ,
  \V1417(0) ,
  \V1681(0) ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \V759(0) ,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  \V1767(1) ,
  \V1632(0) ,
  \V1767(0) ,
  \[40] ,
  \[41] ,
  \[42] ,
  \V1306(0) ,
  \[43] ,
  \[44] ,
  \V913(0) ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \V1718(0) ,
  \V925(0) ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \V863(0) ,
  \[54] ,
  \[55] ,
  \[56] ,
  \V598(0) ,
  \V937(0) ,
  \[57] ,
  \[58] ,
  \[59] ,
  \V2010(0) ,
  \V1268(0) ,
  \V875(0) ,
  \V1471(0) ,
  \V1069(10) ,
  \[60] ,
  \V1069(11) ,
  \V1410(0) ,
  \[61] ,
  \V414(0) ,
  \[62] ,
  \V2022(0) ,
  \[63] ,
  \[64] ,
  \[65] ,
  \V887(0) ,
  \[66] ,
  \[67] ,
  \V487(0) ,
  \[68] ,
  \[69] ,
  \V1422(0) ,
  \V764(0) ,
  \V1360(0) ,
  \[70] ,
  \V364(0) ,
  \[71] ,
  \[72] ,
  \[73] ,
  \[74] ,
  \[75] ,
  \[76] ,
  \V641(0) ,
  \[77] ,
  \[78] ,
  \V1711(0) ,
  \[79] ,
  \V376(0) ,
  \V1311(0) ,
  \V1446(0) ,
  \V2058(0) ,
  \V788(0) ,
  \[80] ,
  \[81] ,
  \[82] ,
  \V1858(0) ,
  \V1809(7) ,
  \[83] ,
  \V1809(6) ,
  \[84] ,
  \[85] ,
  \[86] ,
  \[87] ,
  \[88] ,
  \[89] ,
  \V1396(0) ,
  \V604(0) ,
  \V1809(1) ,
  \V1809(0) ,
  \V1809(3) ,
  \V942(0) ,
  \V1809(2) ,
  \[90] ,
  \V1409(0) ,
  \V1809(5) ,
  \[91] ,
  \V1809(4) ,
  \[92] ,
  \[93] ,
  \V1747(0) ,
  \[94] ,
  \[95] ,
  \[96] ,
  \[97] ,
  \[98] ,
  \[99] ,
  \V1685(0) ,
  \V892(0) ,
  \V905(0) ,
  \V843(0) ,
  \V917(0) ,
  \V381(0) ,
  \V855(0) ,
  \V2002(0) ,
  \V1998(0) ,
  \V867(0) ,
  \V1463(0) ,
  \V467(0) ,
  \V1340(0) ,
  \V1475(0) ,
  \V2087(0) ,
  \V694(2) ,
  \V694(5) ,
  \V694(4) ,
  \V1690(1) ,
  \V694(0) ,
  \V2038(0) ,
  \V633(0) ,
  \V694(7) ,
  \V368(0) ,
  \V694(6) ,
  \V1641(0) ,
  \V510(0) ,
  \V583(0) ,
  \V922(0) ,
  \V1653(0) ,
  \V1388(0) ,
  \V1727(0) ,
  \V934(0) ,
  \V872(0) ,
  V1000,
  V1002,
  V1004,
  V1006,
  V1008,
  \V1277(0) ,
  V1010,
  V1012,
  V1014,
  V1016,
  V1018,
  V1020,
  V1022,
  V1024,
  \V884(0) ,
  V1025,
  V1026,
  V1027,
  V1028,
  V1029,
  V1030,
  V1031,
  V1032,
  V1033,
  V1034,
  V1036,
  V1038,
  V1040,
  V1042,
  V1044,
  V1046,
  V1048,
  V1050,
  V1052,
  V1054,
  V1055,
  \V958(0) ,
  V1056,
  V1057,
  V1058,
  V1059,
  V1060,
  V1061,
  \V1554(0) ,
  V1070,
  V1071,
  \V1689(0) ,
  V1072,
  V1073,
  V1074,
  V1075,
  V1076,
  V1077,
  V1078,
  V1079,
  V1081,
  V1083,
  V1085,
  V1087,
  V1088,
  V1089,
  V1090,
  V1092,
  V1093,
  V1094,
  V1095,
  V1096,
  V1097,
  V1098,
  V1099,
  \V1831(0) ,
  \V361(0) ,
  \V496(0) ,
  \V835(0) ,
  V1100,
  V1101,
  V1103,
  V1105,
  V1107,
  V1109,
  V1111,
  V1113,
  V1115,
  V1117,
  V1119,
  V1121,
  V1123,
  V1125,
  V1127,
  V1128,
  V1129,
  V1130,
  V1131,
  V1132,
  V1133,
  V1134,
  V1136,
  V1138,
  V1140,
  V1142,
  V1144,
  V1146,
  V1148,
  V1149,
  V1150,
  V1151,
  V1152,
  V1153,
  V1154,
  V1155,
  V1156,
  V1157,
  V1158,
  V1160,
  V1162,
  V1164,
  V1166,
  V1168,
  V1170,
  \V847(0) ,
  V1172,
  V1174,
  V1176,
  V1178,
  V1179,
  V1180,
  V1181,
  V1182,
  V1183,
  V1184,
  V1185,
  V1186,
  V1187,
  V1188,
  V1189,
  V1190,
  V1192,
  V1194,
  V1196,
  V1198,
  \V1720(0) ,
  \V1855(0) ,
  \V385(0) ,
  V1200,
  V1202,
  V1204,
  V1206,
  V1208,
  V1210,
  V1212,
  V1214,
  V1215,
  V1216,
  V1217,
  V1218,
  V1219,
  \V1455(0) ,
  V1220,
  V1221,
  V1222,
  V1223,
  V1224,
  V1226,
  V1228,
  \V2067(0) ,
  V1230,
  V1232,
  V1234,
  V1236,
  V1238,
  V1240,
  V1242,
  V1244,
  V1245,
  V1246,
  V1247,
  V1248,
  V1250,
  V1252,
  V1254,
  V1269,
  V1270,
  V1271,
  V1272,
  V1273,
  V1276,
  V1279,
  V1280,
  V1283,
  V1284,
  V1285,
  V1286,
  V1287,
  V1288,
  V1290,
  V1292,
  V1294,
  V1296,
  V1298,
  V1299,
  \V336(0) ,
  \V1670(0) ,
  \V2018(0) ,
  V1300,
  V1301,
  V1302,
  V1303,
  V1304,
  V1305,
  V1307,
  V1308,
  V1309,
  \V686(3) ,
  V1310,
  V1312,
  V1313,
  V1314,
  V1315,
  V1316,
  V1317,
  V1318,
  V1319,
  V1320,
  V1321,
  V1322,
  V1323,
  V1324,
  V1325,
  V1326,
  V1327,
  V1328,
  V1329,
  \V686(5) ,
  V1330,
  V1332,
  V1333,
  V1335,
  V1336,
  V1338,
  V1339,
  \V686(4) ,
  V1341,
  V1342,
  V1343,
  V1344,
  V1345,
  V1346,
  V1347,
  V1348,
  V1349,
  V1350,
  V1352,
  V1353,
  V1355,
  V1356,
  V1358,
  V1359,
  V1361,
  V1362,
  V1363,
  V1364,
  V1366,
  V1367,
  V1368,
  V1369,
  V1376,
  V1377,
  V1379,
  V1381,
  V1383,
  \V1282(1) ,
  V1385,
  V1390,
  V1391,
  V1393,
  \V686(7) ,
  \V686(6) ,
  \V1694(1) ,
  V1400,
  V1401,
  V1402,
  V1403,
  V1404,
  V1405,
  V1406,
  V1407,
  \V902(0) ,
  V1411,
  V1412,
  V1413,
  V1414,
  V1416,
  V1418,
  V1419,
  V1420,
  V1424,
  V1425,
  V1427,
  V1430,
  V1433,
  V1434,
  V1435,
  V1436,
  V1438,
  V1443,
  V1445,
  V1448,
  V1449,
  V1450,
  V1453,
  V1454,
  V1456,
  V1457,
  V1458,
  V1461,
  V1462,
  V1464,
  V1465,
  V1466,
  V1469,
  V1473,
  V1474,
  V1476,
  V1477,
  V1478,
  V1479,
  V1482,
  V1483,
  V1484,
  V1485,
  V1486,
  V1487,
  V1488,
  V1489,
  V1490,
  V1491,
  V1494,
  V1497,
  V1499,
  \V914(0) ,
  \V1983(0) ,
  \V852(0) ,
  \V987(0) ,
  V1500,
  V1501,
  V1503,
  V1504,
  V1505,
  V1506,
  V1507,
  V1509,
  V1511,
  V1513,
  V1515,
  V1516,
  V1517,
  V1518,
  V1519,
  V1520,
  V1521,
  V1522,
  V1523,
  V1524,
  V1525,
  V1526,
  V1527,
  V1528,
  V1529,
  V1530,
  V1531,
  V1532,
  V1533,
  V1534,
  V1535,
  V1540,
  V1541,
  V1542,
  V1543,
  V1544,
  V1545,
  V1547,
  V1548,
  V1549,
  V1551,
  V1555,
  V1556,
  V1557,
  V1558,
  V1559,
  V1560,
  V1561,
  V1562,
  V1563,
  V1564,
  V1566,
  V1567,
  V1568,
  V1569,
  V1570,
  V1571,
  V1572,
  V1573,
  V1574,
  V1575,
  V1576,
  V1577,
  V1578,
  V1579,
  \V1860(0) ,
  V1580,
  V1581,
  V1582,
  V1583,
  V1584,
  V1585,
  V1586,
  V1587,
  V1588,
  V1589,
  \V864(0) ,
  V1590,
  V1591,
  V1592,
  V1593,
  V1594,
  V1598,
  V1599,
  \V1460(0) ,
  \V803(0) ,
  \V2011(0) ,
  V1600,
  V1601,
  V1602,
  V1603,
  V1604,
  V1605,
  V1606,
  V1607,
  V1608,
  V1609,
  V1610,
  V1611,
  V1614,
  V1615,
  V1616,
  V1617,
  V1618,
  V1619,
  V1621,
  V1622,
  V1624,
  V1625,
  V1626,
  V1627,
  V1628,
  \V1472(0) ,
  V1633,
  V1634,
  V1635,
  V1636,
  V1637,
  V1638,
  V1639,
  V1640,
  \V476(0) ,
  V1643,
  V1644,
  V1646,
  \V2084(0) ,
  V1648,
  V1650,
  V1651,
  V1654,
  V1655,
  V1656,
  V1657,
  V1658,
  V1659,
  V1660,
  V1661,
  V1662,
  V1663,
  \V1546(0) ,
  V1664,
  V1665,
  V1666,
  V1667,
  V1668,
  \V1023(7) ,
  V1672,
  V1673,
  V1675,
  V1676,
  V1677,
  V1678,
  \V1023(6) ,
  V1682,
  V1683,
  V1686,
  V1688,
  \V1023(9) ,
  V1691,
  V1692,
  V1695,
  V1696,
  V1697,
  V1698,
  V1699,
  \V1023(8) ,
  \V1023(10) ,
  \V1023(11) ,
  \V827(0) ,
  V1700,
  V1702,
  V1704,
  V1706,
  V1708,
  \V1023(1) ,
  V1710,
  V1712,
  V1713,
  V1714,
  V1715,
  V1716,
  \V1023(0) ,
  V1721,
  V1722,
  V1723,
  V1724,
  V1725,
  \V1761(0) ,
  V1729,
  \V1023(3) ,
  V1730,
  V1731,
  V1732,
  V1733,
  V1734,
  \V765(0) ,
  V1735,
  V1737,
  V1738,
  V1739,
  \V1023(2) ,
  V1740,
  V1742,
  V1743,
  V1744,
  V1748,
  V1749,
  \V1023(5) ,
  V1750,
  \V1496(0) ,
  V1751,
  V1752,
  V1754,
  V1755,
  V1756,
  \V1835(0) ,
  \V1023(4) ,
  \V365(0) ,
  V1764,
  V1765,
  V1768,
  V1770,
  V1774,
  V1775,
  V1778,
  V1780,
  V1782,
  V1792,
  V1793,
  V1794,
  V1795,
  V1796,
  V1797,
  V1798,
  V1799,
  \V1773(1) ,
  \V1773(0) ,
  \V642(0) ,
  \V777(0) ,
  V1800,
  V1801,
  \V1447(0) ,
  V1810,
  V1812,
  V1814,
  V1816,
  V1818,
  V1820,
  V1822,
  V1824,
  V1826,
  V1828,
  V1830,
  V1834,
  V1836,
  V1838,
  V1839,
  V1840,
  V1841,
  V1842,
  V1843,
  V1844,
  V1845,
  V1846,
  V1847,
  V1848,
  V1849,
  V1850,
  V1851,
  V1852,
  V1867,
  V1868,
  V1869,
  V1870,
  V1871,
  V1872,
  V1873,
  V1874,
  \V1859(0) ,
  V1875,
  V1876,
  V1877,
  V1878,
  V1879,
  V1880,
  V1881,
  V1882,
  V1883,
  V1884,
  V1885,
  V1886,
  V1887,
  V1888,
  \[0] ,
  V1889,
  V1890,
  V1891,
  V1892,
  V1893,
  V1894,
  V1895,
  \[1] ,
  \[2] ,
  \V592(0) ,
  \[3] ,
  \[4] ,
  \[5] ,
  \[6] ,
  \[7] ,
  \V1397(0) ,
  V1902,
  V1904,
  V1905,
  V1906,
  V1907,
  V1908,
  \[8] ,
  V1909,
  V1910,
  V1912,
  V1914,
  V1916,
  V1918,
  \[9] ,
  V1920,
  V1922,
  V1923,
  V1924,
  V1925,
  V1926,
  V1927,
  V1928,
  V1929,
  V1930,
  V1931,
  V1932,
  V1933,
  V1934,
  V1935,
  V1936,
  V1937,
  V1938,
  V1940,
  V1941,
  V1943,
  \V943(0) ,
  V1945,
  V1947,
  V1949,
  V1951,
  V1954,
  V1955,
  V1956,
  V1957,
  V1959,
  \V1674(0) ,
  V1961,
  V1962,
  V1966,
  V1967,
  V1969,
  V1970,
  V1971,
  V1972,
  V1973,
  V1974,
  V1978,
  V1979,
  V1980,
  V1981,
  V1982,
  V1985,
  V1986,
  V1987,
  V1988,
  V1989,
  V1991,
  V1993,
  V1994,
  V1995,
  V1996,
  V1997,
  \V629(0) ,
  \V893(0) ,
  \V1963(0) ,
  \V493(0) ,
  \V832(0) ,
  \V967(0) ,
  \V1502(0) ,
  \V1975(0) ,
  \V370(0) ,
  \V844(0) ,
  \V1514(0) ,
  \V1649(0) ,
  \V382(0) ,
  \V1452(0) ,
  \V2064(0) ,
  \V1126(1) ,
  \V1999(0) ,
  \V394(0) ,
  \V733(0) ,
  \V807(0) ,
  \V1538(0) ,
  \V610(0) ,
  \V1415(0) ,
  \V1753(0) ,
  \V622(0) ,
  \V1630(0) ,
  \V369(0) ,
  \V1777(1) ,
  \V1642(0) ,
  \V1777(0) ,
  \V584(0) ,
  \V923(0) ,
  \V658(0) ,
  \V1389(0) ,
  \V1728(0) ,
  \V800(0) ,
  \V935(0) ,
  \[100] ,
  \[101] ,
  \[102] ,
  \V873(0) ,
  \[103] ,
  \[104] ,
  \V473(0) ,
  \[105] ,
  \V2081(0) ,
  \V812(0) ,
  \V947(0) ,
  \[106] ,
  \[107] ,
  \V412(0) ,
  \[108] ,
  \V2020(0) ,
  \V1278(1) ,
  \[109] ,
  V2000,
  V2001,
  V2003,
  V2005,
  V2006,
  V2009,
  V2012,
  V2013,
  V2014,
  V2015,
  V2016,
  V2017,
  V2021,
  V2023,
  \V885(0) ,
  V2025,
  V2026,
  V2027,
  V2028,
  V2029,
  V2030,
  V2031,
  V2032,
  V2034,
  V2035,
  V2036,
  V2037,
  V2039,
  V2040,
  V2041,
  V2042,
  V2043,
  V2044,
  V2045,
  V2046,
  V2047,
  V2048,
  V2049,
  V2050,
  V2051,
  V2052,
  V2053,
  V2054,
  V2055,
  \V959(0) ,
  V2056,
  V2057,
  V2059,
  V2060,
  V2062,
  V2063,
  V2065,
  V2066,
  V2068,
  V2069,
  \[110] ,
  V2070,
  V2071,
  V2072,
  V2073,
  V2074,
  V2075,
  V2076,
  V2077,
  V2079,
  \V424(0) ,
  \[111] ,
  V2080,
  V2082,
  V2083,
  V2085,
  V2086,
  V2088,
  V2089,
  \[112] ,
  V2090,
  V2091,
  V2092,
  V2093,
  V2094,
  V2095,
  V2096,
  V2097,
  V2098,
  V2099,
  \[113] ,
  \[114] ,
  \V762(0) ,
  \V897(0) ,
  \[115] ,
  \V1493(0) ,
  \[116] ,
  \V362(0) ,
  \[117] ,
  \[118] ,
  \[119] ,
  V2100,
  V2101,
  V2102,
  V2103,
  V2104,
  V2105,
  V2106,
  V2107,
  V2108,
  V2109,
  \V436(0) ,
  V2110,
  V2111,
  V2112,
  V2113,
  V2114,
  V2115,
  V2116,
  V2117,
  V2118,
  V2119,
  V2120,
  V2121,
  V2122,
  V2123,
  V2124,
  V2125,
  V2126,
  V2127,
  V2128,
  V2129,
  V2130,
  V2131,
  V2132,
  V2133,
  V2134,
  V2135,
  V2136,
  V2137,
  V2138,
  V2139,
  V2140,
  V2141,
  V2142,
  V2143,
  V2144,
  V2145,
  V2146,
  V2147,
  V2148,
  V2149,
  V2150,
  V2151,
  V2152,
  V2153,
  V2154,
  V2155,
  V2156,
  V2157,
  V2158,
  V2159,
  V2160,
  V2161,
  V2162,
  V2163,
  V2164,
  V2165,
  V2166,
  V2167,
  V2168,
  V2169,
  \V374(0) ,
  \[120] ,
  V2170,
  V2171,
  V2172,
  V2173,
  V2174,
  V2175,
  V2176,
  V2177,
  V2178,
  V2179,
  \[121] ,
  V2180,
  V2181,
  V2182,
  V2183,
  V2184,
  V2185,
  V2186,
  V2187,
  V2188,
  V2189,
  \V1444(0) ,
  \[122] ,
  V2190,
  V2191,
  V2192,
  V2193,
  V2194,
  V2195,
  V2196,
  V2197,
  V2198,
  V2199,
  \[123] ,
  \[124] ,
  \[125] ,
  \[126] ,
  \[127] ,
  \[128] ,
  \V1856(0) ,
  \V386(0) ,
  \[129] ,
  V2200,
  V2201,
  V2202,
  V2203,
  V2204,
  V2205,
  V2206,
  V2207,
  V2208,
  V2209,
  V2210,
  V2211,
  V2212,
  V2213,
  V2214,
  V2215,
  V2216,
  V2217,
  V2218,
  V2219,
  V2220,
  V2221,
  V2222,
  V2223,
  V2224,
  V2225,
  V2226,
  V2227,
  V2228,
  V2229,
  V2230,
  V2231,
  V2232,
  V2233,
  V2234,
  V2235,
  V2236,
  V2237,
  V2238,
  V2239,
  V2240,
  V2241,
  V2242,
  V2243,
  V2244,
  V2245,
  V2246,
  V2247,
  V2248,
  V2249,
  V2250,
  V2251,
  V2252,
  V2253,
  V2254,
  V2255,
  V2256,
  V2257,
  V2258,
  V2259,
  \V2007(0) ,
  V2260,
  V2261,
  V2262,
  V2263,
  V2264,
  V2265,
  V2266,
  V2267,
  V2268,
  V2269,
  \[130] ,
  V2270,
  V2271,
  V2272,
  V2273,
  V2274,
  V2275,
  V2276,
  V2277,
  V2278,
  \V1394(0) ,
  V2279,
  \[131] ,
  V2280,
  V2281,
  V2282,
  V2283,
  V2284,
  V2285,
  V2286,
  V2287,
  V2288,
  V2289,
  \[132] ,
  V2290,
  V2291,
  V2292,
  V2293,
  V2294,
  V2295,
  V2296,
  V2297,
  V2298,
  V2299,
  \[133] ,
  \V1468(0) ,
  \[134] ,
  \[135] ,
  \[136] ,
  \[137] ,
  \V2019(0) ,
  \[138] ,
  \[139] ,
  V2300,
  V2301,
  V2302,
  V2303,
  V2304,
  V2305,
  V2306,
  V2307,
  V2308,
  V2309,
  V2310,
  V2311,
  V2312,
  V2313,
  V2314,
  V2315,
  V2316,
  V2317,
  V2318,
  V2319,
  V2320,
  V2321,
  V2322,
  V2323,
  V2324,
  V2325,
  V2326,
  V2327,
  V2328,
  V2329,
  V2330,
  V2331,
  V2332,
  V2333,
  V2334,
  V2335,
  V2336,
  V2337,
  V2338,
  V2339,
  V2340,
  V2341,
  V2342,
  V2343,
  V2344,
  V2345,
  V2346,
  V2347,
  V2348,
  V2349,
  V2350,
  V2351,
  V2352,
  V2353,
  V2354,
  V2355,
  V2356,
  V2357,
  V2358,
  V2359,
  V2360,
  V2361,
  V2362,
  V2363,
  V2364,
  V2365,
  V2366,
  V2367,
  V2368,
  V2369,
  \[140] ,
  V2370,
  V2371,
  V2372,
  V2373,
  V2374,
  V2375,
  V2376,
  V2377,
  V2378,
  V2379,
  \[141] ,
  V2380,
  V2381,
  V2382,
  V2383,
  V2384,
  V2385,
  V2386,
  V2387,
  V2388,
  V2389,
  \[142] ,
  V2390,
  V2391,
  V2392,
  V2393,
  V2394,
  V2395,
  V2396,
  V2397,
  V2398,
  V2399,
  \[143] ,
  \[144] ,
  \[145] ,
  \V1357(0) ,
  \[146] ,
  \V490(0) ,
  \[147] ,
  \[148] ,
  \[149] ,
  V2400,
  V2401,
  V2402,
  V2403,
  V2404,
  V2405,
  V2406,
  V2407,
  V2408,
  V2409,
  \V699(0) ,
  \V903(0) ,
  V2410,
  V2411,
  V2412,
  V2413,
  V2414,
  V2415,
  V2416,
  V2417,
  V2418,
  V2419,
  V2420,
  V2421,
  V2422,
  V2423,
  V2424,
  V2425,
  V2426,
  V2427,
  V2428,
  V2429,
  V2430,
  V2431,
  V2432,
  V2433,
  V2434,
  V2435,
  V2436,
  \V503(0) ,
  V2437,
  V2438,
  V2439,
  V2440,
  V2441,
  V2442,
  V2443,
  V2444,
  V2445,
  V2446,
  V2447,
  V2448,
  V2449,
  V2450,
  V2451,
  V2452,
  V2453,
  V2454,
  V2455,
  V2456,
  V2457,
  V2458,
  V2459,
  V2460,
  V2461,
  V2462,
  V2463,
  V2464,
  V2465,
  V2466,
  V2467,
  V2468,
  V2469,
  \[150] ,
  V2470,
  V2471,
  V2472,
  V2473,
  V2474,
  V2475,
  V2476,
  V2477,
  V2478,
  V2479,
  \[151] ,
  V2480,
  V2481,
  V2482,
  V2483,
  V2484,
  V2485,
  V2486,
  V2487,
  V2488,
  V2489,
  \[152] ,
  V2490,
  V2491,
  V2492,
  V2493,
  V2494,
  V2495,
  V2496,
  V2497,
  V2498,
  V2499,
  \V915(0) ,
  \[153] ,
  \[154] ,
  \[155] ,
  \[156] ,
  \[157] ,
  \V1984(0) ,
  \[158] ,
  \V853(0) ,
  \[159] ,
  V2500,
  V2501,
  V2502,
  V2503,
  V2504,
  V2505,
  V2506,
  V2507,
  V2508,
  V2509,
  V2510,
  V2511,
  V2512,
  V2513,
  V2514,
  V2515,
  V2516,
  V2517,
  V2518,
  V2519,
  V2520,
  V2521,
  V2522,
  V2523,
  V2524,
  V2525,
  \V588(0) ,
  V2526,
  V2527,
  V2528,
  \V2061(0) ,
  V2529,
  \V927(0) ,
  V2530,
  V2531,
  V2532,
  V2533,
  V2534,
  V2535,
  V2536,
  V2537,
  V2538,
  V2539,
  V2540,
  V2541,
  V2542,
  V2543,
  V2544,
  V2545,
  V2546,
  V2547,
  V2548,
  V2549,
  V2550,
  V2551,
  V2552,
  V2553,
  V2554,
  V2555,
  V2556,
  V2557,
  V2558,
  V2559,
  V2560,
  V2561,
  V2562,
  V2563,
  V2564,
  V2565,
  V2566,
  V2567,
  V2568,
  V2569,
  \[160] ,
  V2570,
  V2571,
  V2572,
  V2573,
  V2574,
  V2575,
  V2576,
  V2577,
  V2578,
  V2579,
  \V1861(0) ,
  \[161] ,
  V2580,
  V2581,
  \V391(0) ,
  V2582,
  V2583,
  V2584,
  V2585,
  V2586,
  V2587,
  \V730(0) ,
  V2588,
  V2589,
  \V865(0) ,
  \[162] ,
  V2590,
  V2591,
  V2592,
  V2593,
  V2594,
  V2595,
  \V1596(1) ,
  V2596,
  V2597,
  V2598,
  V2599,
  \[163] ,
  \V1596(0) ,
  \[164] ,
  \[165] ,
  \[166] ,
  \V1147(7) ,
  \[167] ,
  \V404(0) ,
  \V1147(6) ,
  \[168] ,
  \V1147(9) ,
  \[169] ,
  V2600,
  V2601,
  V2602,
  V2603,
  V2604,
  V2605,
  V2606,
  V2607,
  V2608,
  V2609,
  \V1147(8) ,
  V2610,
  V2611,
  V2612,
  V2613,
  V2614,
  V2615,
  V2616,
  V2617,
  V2618,
  \V877(0) ,
  V2619,
  V2620,
  V2621,
  V2622,
  V2623,
  V2624,
  V2625,
  V2626,
  V2627,
  V2628,
  V2629,
  V2630,
  V2631,
  V2632,
  V2633,
  V2634,
  V2635,
  V2636,
  V2637,
  V2638,
  V2639,
  \V342(0) ,
  V2640,
  V2641,
  V2642,
  V322,
  V2643,
  V323,
  V2644,
  V324,
  V2645,
  V325,
  V2646,
  V326,
  V2647,
  V327,
  V2648,
  V328,
  V2649,
  V329,
  V2650,
  V330,
  V2651,
  V331,
  V2652,
  V332,
  V2653,
  V333,
  V2654,
  V334,
  V2655,
  V335,
  V2656,
  V2657,
  V337,
  V2658,
  V338,
  V2659,
  V339,
  V2660,
  V340,
  V2661,
  V341,
  V2662,
  V2663,
  V343,
  V2664,
  V344,
  V2665,
  V345,
  V2666,
  V2667,
  V347,
  V2668,
  V348,
  V2669,
  V349,
  \[170] ,
  V2670,
  V350,
  V2671,
  V351,
  V2672,
  V352,
  V2673,
  V353,
  V2674,
  V354,
  V2675,
  \V2024(0) ,
  V355,
  V2676,
  V2677,
  V2678,
  V358,
  V2679,
  V359,
  \[171] ,
  V2680,
  V360,
  V2681,
  V2682,
  V2683,
  V2684,
  V2685,
  V2686,
  V2687,
  V2688,
  V2689,
  \[172] ,
  V2690,
  V2691,
  V2692,
  V372,
  V2693,
  V2694,
  V2695,
  V2696,
  V2697,
  V2698,
  V2699,
  V379,
  \[173] ,
  V387,
  V388,
  V389,
  \[174] ,
  V390,
  V392,
  V395,
  V397,
  \V1147(5) ,
  \[175] ,
  \[176] ,
  \[177] ,
  \[178] ,
  \[179] ,
  V2700,
  V2701,
  V2702,
  V2703,
  V2704,
  V2705,
  V2706,
  V2707,
  V2708,
  V2709,
  V2710,
  V2711,
  V2712,
  V2713,
  V2714,
  V2715,
  V2716,
  V2717,
  V2718,
  V2719,
  V2720,
  V400,
  V2721,
  V401,
  V2722,
  V402,
  V2723,
  V403,
  V2724,
  V2725,
  V2726,
  V406,
  V2727,
  V407,
  V2728,
  V2729,
  V409,
  V2730,
  V2731,
  V411,
  V2732,
  V2733,
  V2734,
  V2735,
  V415,
  V2736,
  V416,
  V2737,
  V417,
  V2738,
  V418,
  V2739,
  V419,
  V2740,
  V420,
  V2741,
  V421,
  V2742,
  V422,
  V2743,
  V2744,
  V2745,
  V425,
  V2746,
  V426,
  V2747,
  V427,
  V2748,
  V428,
  V2749,
  V429,
  V2750,
  V430,
  V2751,
  V431,
  V2752,
  V2753,
  V433,
  V2754,
  V2755,
  V2756,
  V2757,
  V437,
  V2758,
  V438,
  V2759,
  V439,
  \V366(0) ,
  V2760,
  V440,
  V2761,
  V441,
  V2762,
  V442,
  V2763,
  V443,
  V2764,
  V444,
  V2765,
  V2766,
  V446,
  V2767,
  V447,
  V2768,
  V448,
  V2769,
  V449,
  \[180] ,
  V2770,
  V2771,
  V451,
  V2772,
  V452,
  V2773,
  V453,
  V2774,
  V454,
  V2775,
  V455,
  V2776,
  V456,
  V2777,
  V457,
  V2778,
  V458,
  V2779,
  V459,
  \[181] ,
  V2780,
  V460,
  V2781,
  V461,
  V2782,
  V462,
  V2783,
  V463,
  V2784,
  V464,
  V2785,
  V465,
  V2786,
  V466,
  V2787,
  V2788,
  V468,
  V2789,
  V469,
  \[182] ,
  V2790,
  V2791,
  V471,
  V2792,
  V472,
  V2793,
  V2794,
  V474,
  V2795,
  V475,
  V2796,
  V2797,
  V477,
  V2798,
  V478,
  V2799,
  V479,
  \[183] ,
  V480,
  V481,
  V482,
  V483,
  V484,
  V485,
  V486,
  V488,
  V489,
  \[184] ,
  V491,
  V492,
  V494,
  V495,
  V497,
  V498,
  V499,
  \[185] ,
  \[186] ,
  \V1147(10) ,
  \[187] ,
  \V1147(11) ,
  \V378(0) ,
  \[188] ,
  \[189] ,
  V2800,
  V2801,
  V2802,
  V2803,
  V2804,
  V2805,
  V2806,
  V2807,
  V2808,
  V2809,
  V2810,
  V2811,
  V2812,
  V2813,
  V2814,
  V2815,
  V2816,
  V2817,
  V501,
  V502,
  V505,
  V506,
  V507,
  V509,
  V513,
  V514,
  V515,
  V516,
  V517,
  V518,
  V519,
  V520,
  V521,
  V522,
  V523,
  V524,
  V525,
  V526,
  V529,
  V530,
  V531,
  V534,
  V535,
  V549,
  \[190] ,
  \V667(3) ,
  V550,
  V551,
  V552,
  V553,
  V555,
  V557,
  V559,
  \[191] ,
  \V667(2) ,
  \V729(0) ,
  V561,
  V563,
  V565,
  V567,
  V569,
  \[192] ,
  \V667(5) ,
  V571,
  V573,
  V574,
  V575,
  V576,
  V577,
  V578,
  V579,
  \[193] ,
  \V667(4) ,
  V580,
  V581,
  V582,
  V586,
  V589,
  \[194] ,
  V590,
  V593,
  \V932(0) ,
  V594,
  V595,
  V596,
  V599,
  \[195] ,
  \[196] ,
  \V667(1) ,
  \V532(0) ,
  \[197] ,
  \V667(0) ,
  \[198] ,
  \V1398(0) ,
  \[199] ,
  V600,
  V601,
  V602,
  V605,
  V606,
  V607,
  V608,
  \V1337(0) ,
  \V667(7) ,
  V611,
  V613,
  V614,
  V615,
  V616,
  V617,
  V618,
  V619,
  \V470(0) ,
  \V667(6) ,
  \V944(0) ,
  V623,
  V624,
  V625,
  V626,
  V627,
  V628,
  V631,
  V632,
  V635,
  V636,
  V637,
  V638,
  V643,
  V644,
  V645,
  V646,
  V647,
  V648,
  V649,
  \V1275(0) ,
  \V882(0) ,
  V687,
  V688,
  V695,
  V696,
  V697,
  V698,
  \V956(0) ,
  \V1687(0) ,
  V700,
  V701,
  V702,
  V703,
  V704,
  V705,
  V706,
  \V894(0) ,
  V710,
  V711,
  V712,
  V713,
  V714,
  V715,
  V716,
  V717,
  V718,
  V719,
  V720,
  V721,
  V722,
  V723,
  V724,
  V725,
  V726,
  V727,
  V728,
  \V1964(0) ,
  V732,
  V734,
  V735,
  V736,
  V737,
  V738,
  V739,
  \V833(0) ,
  V740,
  V741,
  V742,
  V743,
  V744,
  V745,
  V746,
  V747,
  V748,
  V749,
  V750,
  V751,
  V752,
  V753,
  V754,
  V755,
  V756,
  V757,
  V760,
  V761,
  V766,
  V767,
  V768,
  V769,
  \V907(0) ,
  V770,
  V771,
  V772,
  V773,
  V774,
  V776,
  V785,
  V786,
  V790,
  V791,
  V792,
  V793,
  V794,
  V795,
  V796,
  V797,
  V799,
  \V1903(4) ,
  \V1976(0) ,
  \V371(0) ,
  \V845(0) ,
  \V1441(0) ,
  \V1053(7) ,
  \V445(0) ,
  \V1791(7) ,
  \V1053(6) ,
  V804,
  V805,
  V806,
  V808,
  V809,
  \V1791(6) ,
  \V1053(9) ,
  V810,
  V811,
  V814,
  V815,
  V816,
  V818,
  V819,
  \V1053(8) ,
  V820,
  V823,
  V824,
  V825,
  V828,
  V829,
  \V1791(8) ,
  V830,
  V831,
  V836,
  V838,
  V839,
  V840,
  V841,
  V846,
  V848,
  V849,
  \V1853(0) ,
  V850,
  V851,
  \V383(0) ,
  V856,
  V858,
  V859,
  \V857(0) ,
  V860,
  V861,
  V866,
  V868,
  V869,
  V870,
  V871,
  V876,
  V878,
  V879,
  V880,
  V881,
  V886,
  V888,
  V889,
  \V1053(1) ,
  V890,
  V891,
  V896,
  V898,
  V899,
  \V1791(1) ,
  \V1053(0) ,
  \V1791(0) ,
  \V1053(3) ,
  \V2004(0) ,
  \V1791(3) ,
  \V1053(2) ,
  \V1791(2) ,
  \V1053(5) ,
  \V672(3) ,
  \V1791(5) ,
  \V1865(0) ,
  \V1053(4) ,
  \V1791(4) ,
  \V672(5) ,
  V900,
  V901,
  V906,
  \V672(4) ,
  V908,
  V909,
  V910,
  V911,
  V916,
  V918,
  V919,
  V920,
  V921,
  V926,
  V928,
  V929,
  V930,
  V931,
  V936,
  V938,
  V939,
  V940,
  V941,
  \V408(0) ,
  V946,
  V948,
  V949,
  V950,
  V951,
  V952,
  V953,
  V954,
  V955,
  V960,
  V961,
  V962,
  V963,
  V964,
  V968,
  V969,
  V970,
  V971,
  V972,
  V973,
  V974,
  V975,
  V976,
  V977,
  V978,
  V979,
  V980,
  V981,
  V983,
  V984,
  V988,
  V989,
  V990,
  V991,
  V992,
  V993,
  V994,
  V995,
  V996,
  V997,
  \V672(7) ,
  V998,
  V999,
  \V346(0) ,
  \V672(6) ,
  \V1680(0) ;
assign
  \V758(0)  = V756 | (V755 | V757),
  \V1354(0)  = V1353 | V1352,
  \V1631(0)  = V766 | V769,
  \V1243(7)  = \[84] ,
  \V500(0)  = \[12] ,
  \V1243(6)  = \[85] ,
  \V1243(9)  = \[82] ,
  \V709(1)  = ~\V88(3) ,
  \V1243(8)  = \[83] ,
  \V709(0)  = ~\V88(2) ,
  \V912(0)  = ~V908,
  \V1243(1)  = \[90] ,
  \V1243(0)  = \[91] ,
  \V1717(0)  = \[159] ,
  \V1243(3)  = \[88] ,
  \V985(0)  = V983 | (V978 | V984),
  \V1243(2)  = \[89] ,
  \V1243(5)  = \[86] ,
  \V1243(4)  = \[87] ,
  \V450(0)  = V448 | (V447 | V449),
  \V585(0)  = \[39] ,
  \V924(0)  = ~V920,
  \V659(0)  = ~\V9(0) ,
  \V1255(1)  = V1252 | V1246,
  \V1255(0)  = V1254 | V1247,
  \V1255(3)  = V1248 | V1244,
  \V862(0)  = ~V858,
  \V1255(2)  = V1250 | V1245,
  \V597(0)  = \[42] ,
  \V536(0)  = V534 | V535,
  \[200]  = V1941 | V1933,
  \[201]  = V1943 | V1934,
  \[202]  = V1945 | V1935,
  \V874(0)  = ~V870,
  \[203]  = V1947 | V1936,
  \V1124(12)  = V1103 | V1093,
  \[204]  = V1949 | V1937,
  \V1124(13)  = V1101 | V1092,
  \[205]  = V1951 | V1938,
  \V813(0)  = \V807(0)  | V697,
  \[206]  = V1954 | V1940,
  \[207]  = V1957 | V1955,
  \V1679(0)  = \[152] ,
  \V413(0)  = \V174(0)  | (V502 | (V411 | \V404(0) )),
  \[208]  = V1959 | V1956,
  \[209]  = V1966 | V1967,
  \V1124(10)  = V1107 | V1095,
  \V1124(11)  = V1105 | V1094,
  \V1421(0)  = V1404 | (V1403 | V1418),
  \[210]  = V1989 | V1987,
  \[211]  = V1991 | V1988,
  \V2033(0)  = V2031 | (V2030 | V2032),
  \[212]  = V2293 | V2292,
  \[213]  = V2297 | V2296,
  \[214]  = V2301 | V2300,
  \[215]  = V2305 | V2304,
  \[216]  = V2309 | V2308,
  \V1833(0)  = \[184] ,
  \V1968(0)  = \[209] ,
  \V363(0)  = ~V350,
  \[217]  = V2313 | V2312,
  \V837(0)  = ~V836,
  \[218]  = V2317 | V2316,
  \[219]  = V2573 | V2572,
  \V1771(1)  = \[169] ,
  \V1771(0)  = \[170] ,
  \V640(0)  = \[49] ,
  \V375(0)  = \[4] ,
  \[220]  = V2577 | V2576,
  \[221]  = V2581 | V2580,
  \[222]  = V2585 | V2584,
  \[223]  = V2589 | V2588,
  \V1857(0)  = ~V1842,
  \V1069(7)  = V1074 | V1058,
  \V1069(6)  = V1075 | V1059,
  \V1069(9)  = V1072 | V1056,
  \V1069(8)  = V1073 | V1057,
  \V2008(0)  = ~V2005,
  \V1395(0)  = V700 | V701,
  \V399(0)  = ~\V249(0) ,
  \V603(0)  = \[43] ,
  \V676(5)  = ~\V667(5) ,
  \V1334(0)  = V1333 | V1332,
  \V676(4)  = ~\V667(4) ,
  \V1408(0)  = ~V1402,
  \V1069(5)  = V1076 | V1060,
  \V1746(0)  = ~\[163] ,
  \V1069(4)  = V1077 | V1061,
  \V676(7)  = ~\V667(7) ,
  \V676(6)  = ~\V667(6) ,
  \V1684(0)  = ~V1683,
  \V1623(0)  = V1621 | V1622,
  \V1758(0)  = \[166] ,
  \V965(0)  = V962 | (V960 | (V961 | V963)),
  \V1900(0)  = \[191] ,
  \V904(0)  = ~V900,
  \V504(0)  = V740 | V741,
  \V639(0)  = ~V637,
  \V1709(1)  = \[157] ,
  \V1709(0)  = \[158] ,
  \V1709(3)  = \[155] ,
  \V842(0)  = ~V838,
  \V1709(2)  = \[156] ,
  \V1709(4)  = \[154] ,
  \V1512(1)  = \[138] ,
  \V1647(0)  = V727 | (V769 | V726),
  \V1124(7)  = V1113 | V1098,
  \V1512(3)  = \[136] ,
  \V1124(6)  = V1115 | V1099,
  \V1512(2)  = \[137] ,
  \V1124(9)  = V1109 | V1096,
  \V1124(8)  = V1111 | V1097,
  \V380(0)  = V379 | V721,
  \V854(0)  = ~V850,
  \V528(0)  = ~\V43(0) ,
  \V1124(1)  = V1402 & V2124,
  \V1862(0)  = ~V1852,
  \V1124(3)  = V1121 | \V1124(1) ,
  \V731(0)  = V723 | (V722 | V724),
  \V1124(2)  = V1123 | \V1124(1) ,
  \V1124(5)  = V1117 | V1100,
  \V1597(0)  = \V1596(0)  | \V1596(1) ,
  \V1124(4)  = V1119 | \V1124(1) ,
  \V1536(0)  = \[139] ,
  \V405(0)  = V734 | (V515 | \V731(0) ),
  \V681(3)  = ~\V149(3) ,
  \V681(5)  = ~\V149(5) ,
  \V681(4)  = ~\V149(4) ,
  \V817(0)  = V696 | (\V214(0)  | (V815 | (V814 | (\V289(0)  | (\V302(0)  | V816))))),
  \V1351(0)  = V1350 | V1349,
  \V681(7)  = ~\V149(7) ,
  \V681(6)  = ~\V149(6) ,
  \V1086(1)  = V1083 | V1089,
  \V1086(0)  = V1090 | (V1085 | V1078),
  \V1086(3)  = V1079 | V1087,
  \V1086(2)  = V1081 | V1088,
  \V1763(1)  = ~\V88(3) ,
  \V1763(0)  = ~\V88(2) ,
  \V1898(0)  = \[189] ,
  \V1498(0)  = ~V1497,
  \V1837(0)  = ~V1836,
  \V367(0)  = ~V354,
  \V1437(0)  = V1436 | \V1442(0) ,
  \V982(0)  = V501 | (\V2011(0)  | V721),
  \V1652(0)  = \[149] ,
  \V1726(0)  = \[161] ,
  \V933(0)  = ~V929,
  \V533(0)  = ~V531,
  \V1399(0)  = V721 | V769,
  \V1953(7)  = \[200] ,
  \V1953(6)  = \[201] ,
  \V945(0)  = ~V941,
  \V410(0)  = \[8] ,
  \V883(0)  = ~V879,
  \V1953(1)  = \[199] ,
  \V1953(0)  = \[206] ,
  \V822(0)  = ~\V279(0) ,
  \V957(0)  = ~V953,
  \V1953(3)  = \[204] ,
  \V1953(2)  = \[205] ,
  \V1553(0)  = \V60(0)  | \V63(0) ,
  \V1953(5)  = \[202] ,
  \V1953(4)  = \[203] ,
  \V895(0)  = ~V891,
  \V1965(0)  = ~V1962,
  \V834(0)  = ~V830,
  \V1565(0)  = ~V1564,
  \V1177(7)  = V1162 | V1150,
  \V434(0)  = ~V433,
  \V1177(6)  = V1164 | V1151,
  \V1177(9)  = V1158 | V1148,
  \V1177(8)  = V1160 | V1149,
  \V508(0)  = \[13] ,
  \[10]  = V1578 & (V1576 & (V1574 & (V1573 & (V1575 & (V1577 & (\[9]  & (V428 & (V337 & (V426 & (V403 & (V427 & (V429 & (\V1685(0)  & (V430 & V431)))))))))))))),
  \[11]  = \[10]  | \[47] ,
  \V1977(0)  = V700 | V702,
  \[12]  = ~V499,
  \[13]  = V506 | (V613 | (V505 | V507)),
  \V1442(0)  = ~\V278(0) ,
  \[14]  = \V40(0)  | V529,
  \[15]  = \V510(0)  & \V532(0) ,
  \V1177(1)  = V1174 | V1156,
  \[16]  = V430 & (V338 & (V526 & (V431 & V428))),
  \V1177(0)  = V1176 | V1157,
  \[17]  = V769 & \[81] ,
  \V1177(3)  = V1170 | V1154,
  \[18]  = V769 & \[80] ,
  \V1177(2)  = V1172 | V1155,
  \[19]  = V769 & \[79] ,
  \V1177(5)  = V1166 | V1152,
  \V1854(0)  = \V288(2)  | \V288(3) ,
  \V1177(4)  = V1168 | V1153,
  \V384(0)  = \V363(0)  | \V364(0) ,
  \[20]  = V769 & \[78] ,
  \[21]  = V769 & \[77] ,
  \[22]  = V769 & \[76] ,
  \V1392(0)  = \[119] ,
  \V1866(0)  = ~\V16(0) ,
  \[23]  = V769 & \[75] ,
  \V396(0)  = V395 | \[9] ,
  \[24]  = V769 & \[74] ,
  \[25]  = V769 & \[73] ,
  \V1331(0)  = V1330 | V1329,
  \[26]  = V769 & \[72] ,
  \V2078(0)  = V2077 | V2076,
  \[27]  = V769 & \[71] ,
  \[28]  = V769 & \[70] ,
  \[29]  = V553 | V573,
  \V612(0)  = V611 | V502,
  \V1829(7)  = \[175] ,
  \V1829(6)  = \[176] ,
  \V1829(9)  = \[173] ,
  \V1829(8)  = \[174] ,
  \[30]  = V555 | V574,
  \[31]  = V557 | V575,
  \V1417(0)  = V1416 | (V1406 | V745),
  \V1681(0)  = \V262(0)  | \V1674(0) ,
  \[32]  = V559 | V576,
  \[33]  = V561 | V577,
  \[34]  = V563 | V578,
  \V1281(0)  = \[105] ,
  \V1620(0)  = \[146] ,
  \[35]  = V579 | (V565 | V549),
  \V759(0)  = V747 | V748,
  \[36]  = V580 | (V567 | V550),
  \V1829(1)  = \[181] ,
  \[37]  = V581 | (V569 | V551),
  \V1829(0)  = \[182] ,
  \[38]  = V582 | (V571 | V552),
  \V1829(3)  = \[179] ,
  \[39]  = ~\V34(0) ,
  \V1829(2)  = \[180] ,
  \V1693(0)  = \[153] ,
  \V1829(5)  = \[177] ,
  \V1829(4)  = \[178] ,
  \V1767(1)  = ~\V134(1) ,
  \V1632(0)  = V739 | (V741 | (V740 | V768)),
  \V1767(0)  = ~\V134(0) ,
  \[40]  = V586 & \V588(0) ,
  \[41]  = V589 | V590,
  \[42]  = V594 | V596,
  \V1306(0)  = V1304 | (V1303 | V1305),
  \[43]  = V600 | V602,
  \[44]  = V606 | V608,
  \V913(0)  = ~V909,
  \[45]  = V618 & (V617 & V619),
  \[46]  = \V293(0)  & \V533(0) ,
  \[47]  = V625 & (V624 & \V629(0) ),
  \[48]  = ~\V633(0) ,
  \[49]  = ~V638,
  \V1718(0)  = ~\V240(0) ,
  \V1921(1)  = \[197] ,
  \V1921(0)  = \[198] ,
  \V925(0)  = ~V921,
  \V1921(3)  = \[195] ,
  \V1921(2)  = \[196] ,
  \V1921(5)  = \[193] ,
  \[50]  = ~\V257(7) ,
  \V1921(4)  = \[194] ,
  \[51]  = V766 & \V667(3) ,
  \[52]  = V1619 & (V1617 & (V1618 & (\V762(0)  & \V169(0) ))),
  \[53]  = V498 & (V964 & (\[52]  & (\V1674(0)  & \V70(0) ))),
  \V863(0)  = ~V859,
  \[54]  = \V9(0)  & \V5(0) ,
  \[55]  = \V6(0)  & V372,
  \[56]  = \V6(0)  & \V9(0) ,
  \V598(0)  = ~\V245(0) ,
  \V802(0)  = \[65] ,
  \V937(0)  = ~V936,
  \[57]  = \V6(0)  & (\V12(0)  & \V777(0) ),
  \[58]  = \V7(0)  & V372,
  \[59]  = \V11(0)  & \V5(0) ,
  \V2010(0)  = ~V2009,
  \V1268(0)  = V721 | (V726 | (V400 | (V501 | (V769 | (V727 | V728))))),
  \V875(0)  = ~V871,
  \V1471(0)  = V769 | (V766 | V701),
  \V1069(10)  = V1071 | V1055,
  \[60]  = \V11(0)  & \V7(0) ,
  \V1069(11)  = V1070 | V1054,
  \V1410(0)  = ~V1407,
  \[61]  = V785 & V786,
  \V414(0)  = \V1681(0)  | \V405(0) ,
  \[62]  = \V4(0)  & (\V788(0)  & \V9(0) ),
  \V2022(0)  = ~V2021,
  \[63]  = ~V797,
  \[64]  = V799 & \V800(0) ,
  \[65]  = \V51(0)  | \V52(0) ,
  \V887(0)  = ~V886,
  \[66]  = V818 | V820,
  \[67]  = V824 | (V823 | V825),
  \V487(0)  = V486 | V485,
  \[68]  = V498 & (V964 & \V965(0) ),
  \V826(0)  = \[67] ,
  \[69]  = V498 & (V964 & \V985(0) ),
  \V1422(0)  = V1419 | V1420,
  \V1213(10)  = \[71] ,
  \V1213(11)  = \[70] ,
  \V1760(0)  = \[168] ,
  \V764(0)  = ~\[52] ,
  \V1360(0)  = V1359 | V1358,
  \V1495(0)  = \[135] ,
  \[70]  = V1190 | V1178,
  \V364(0)  = ~V351,
  \[71]  = V1192 | V1179,
  \[72]  = V1194 | V1180,
  \[73]  = V1196 | V1181,
  \[74]  = V1198 | V1182,
  \[75]  = V1200 | V1183,
  \[76]  = V1202 | V1184,
  \V641(0)  = ~\V271(0) ,
  \[77]  = V1204 | V1185,
  \[78]  = V1206 | V1186,
  \V1711(0)  = V421 | V721,
  \[79]  = V1208 | V1187,
  \V376(0)  = V697 | \V35(0) ,
  \V1311(0)  = V1309 | (V1308 | V1310),
  \V1446(0)  = ~V1445,
  \V2058(0)  = V2057 | V2056,
  \V788(0)  = \V1565(0)  | \V13(0) ,
  \[80]  = V1210 | V1188,
  \[81]  = V1212 | V1189,
  \[82]  = V1224 | V1214,
  \V1858(0)  = ~V1844,
  \V1809(7)  = ~\[70] ,
  \[83]  = V1226 | V1215,
  \V1809(6)  = ~\[71] ,
  \[84]  = V1228 | V1216,
  \[85]  = V1230 | V1217,
  \V591(0)  = \[41] ,
  \[86]  = V1232 | V1218,
  \[87]  = V1234 | V1219,
  \[88]  = V1236 | V1220,
  \[89]  = V1238 | V1221,
  \V1396(0)  = \V60(0)  | \V59(0) ,
  \V604(0)  = ~\V246(0) ,
  \V1809(1)  = ~\[76] ,
  \V1809(0)  = ~\[77] ,
  \V1809(3)  = ~\[74] ,
  \V942(0)  = ~V938,
  \V1809(2)  = ~\[75] ,
  \[90]  = V1240 | V1222,
  \V1409(0)  = V726 | (\V1395(0)  | V769),
  \V1809(5)  = ~\[72] ,
  \[91]  = V1242 | V1223,
  \V1809(4)  = ~\[73] ,
  \[92]  = V372 & \V2(0) ,
  \[93]  = V1563 & (V1561 & (V1559 & (V1560 & (V1562 & (\V12(0)  & \V2(0) ))))),
  \V1747(0)  = ~\V290(0) ,
  \[94]  = \V9(0)  & \V2(0) ,
  \[95]  = \V9(0)  & \V3(0) ,
  \[96]  = \V11(0)  & \V3(0) ,
  \[97]  = \[96]  & \V1275(0) ,
  \[98]  = V372 & \V4(0) ,
  \[99]  = \V9(0)  & \V4(0) ,
  \V1685(0)  = ~\V1681(0) ,
  \V1759(0)  = \[167] ,
  \V892(0)  = ~V888,
  \V1901(0)  = \[192] ,
  \V905(0)  = ~V901,
  \V1297(1)  = \[109] ,
  \V1297(0)  = \[110] ,
  \V1297(3)  = \[107] ,
  \V1297(2)  = \[108] ,
  \V1297(4)  = \[106] ,
  \V843(0)  = ~V839,
  \V917(0)  = ~V916,
  \V381(0)  = ~\V380(0) ,
  \V855(0)  = ~V851,
  \V1451(0)  = \[128] ,
  \V2002(0)  = V2001 | (V1996 | (V2000 | (\V1999(0)  | V1997))),
  \V1863(0)  = \[185] ,
  \V1998(0)  = ~V1996,
  \V393(0)  = \[6] ,
  \V867(0)  = ~V866,
  \V1463(0)  = V1461 | V1462,
  \V467(0)  = V466 | V465,
  \V1340(0)  = V1339 | V1338,
  \V1475(0)  = V1473 | V1474,
  \V2087(0)  = V2086 | V2085,
  \V694(2)  = ~\V165(2) ,
  \V694(5)  = ~\V165(5) ,
  \V694(4)  = ~\V165(4) ,
  \V1690(1)  = ~\V1983(0) ,
  \V694(0)  = ~\V165(0) ,
  \V2038(0)  = V2036 | (V2035 | V2037),
  \V1899(0)  = \[190] ,
  \V633(0)  = V631 | V632,
  \V694(7)  = ~\V165(7) ,
  \V368(0)  = ~V355,
  \V694(6)  = ~\V165(6) ,
  \V1641(0)  = V1636 | (V1634 | (V1633 | (V1635 | V1637))),
  \V510(0)  = ~V509,
  \V583(0)  = ~\V1(0) ,
  \V922(0)  = ~V918,
  \V1653(0)  = V746 | (V743 | (V736 | (V735 | (V742 | (V744 | \V1687(0) ))))),
  \V1388(0)  = ~V401,
  \V1727(0)  = ~V1721,
  \V934(0)  = ~V930,
  \V872(0)  = ~V868,
  V1000 = \V2011(0)  & (V2111 & \V189(5) ),
  V1002 = \V2011(0)  & (V2111 & \V189(4) ),
  V1004 = \V2011(0)  & (V2111 & \V189(3) ),
  V1006 = \V2011(0)  & (V2111 & \V189(2) ),
  V1008 = \V2011(0)  & (V2111 & \V189(1) ),
  \V1277(0)  = ~V1276,
  V1010 = \V2011(0)  & (V2111 & \V189(0) ),
  V1012 = \V2011(0)  & (V2111 & \V183(5) ),
  V1014 = \V2011(0)  & (V2111 & \V183(4) ),
  V1016 = \V2011(0)  & (V2111 & \V183(3) ),
  V1018 = \V2011(0)  & (V2111 & \V183(2) ),
  V1020 = \V2011(0)  & (V2111 & \V183(1) ),
  V1022 = \V2011(0)  & (V2111 & \V183(0) ),
  V1024 = V2112 & (\V1395(0)  & \V239(4) ),
  \V884(0)  = ~V880,
  V1025 = V2112 & (\V1395(0)  & \V239(3) ),
  V1026 = V2112 & (\V1395(0)  & \V239(2) ),
  V1027 = V2112 & (\V1395(0)  & \V239(1) ),
  V1028 = V2112 & (\V1395(0)  & \V239(0) ),
  V1029 = V2112 & (\V1395(0)  & \V234(4) ),
  V1030 = V2112 & (\V1395(0)  & \V234(3) ),
  V1031 = V2112 & (\V1395(0)  & \V234(2) ),
  V1032 = V2112 & (\V1395(0)  & \V234(1) ),
  V1033 = V2112 & (\V1395(0)  & \V234(0) ),
  V1034 = \V2011(0)  & (V2113 & \V199(4) ),
  V1036 = \V2011(0)  & (V2113 & \V199(3) ),
  V1038 = \V2011(0)  & (V2113 & \V199(2) ),
  \V1480(0)  = \[132] ,
  V1040 = \V2011(0)  & (V2113 & \V199(1) ),
  V1042 = \V2011(0)  & (V2113 & \V199(0) ),
  V1044 = \V2011(0)  & (V2113 & \V194(4) ),
  V1046 = \V2011(0)  & (V2113 & \V194(3) ),
  V1048 = \V2011(0)  & (V2113 & \V194(2) ),
  V1050 = \V2011(0)  & (V2113 & \V194(1) ),
  V1052 = \V2011(0)  & (V2113 & \V194(0) ),
  V1054 = V2114 & (V2115 & (\V1681(0)  & \V257(6) )),
  V1055 = V2114 & (V2115 & (\V1681(0)  & \V257(5) )),
  \V958(0)  = ~V954,
  V1056 = V2114 & (V2115 & (\V1681(0)  & \V257(4) )),
  V1057 = V2114 & (V2115 & (\V1681(0)  & \V257(3) )),
  V1058 = V2114 & (V2115 & (\V1681(0)  & \V257(2) )),
  V1059 = V2114 & (V2115 & (\V1681(0)  & \V257(1) )),
  V1060 = V2114 & (V2115 & (\V1681(0)  & \V257(0) )),
  V1061 = V2114 & (V2115 & (\V1681(0)  & \V257(6) )),
  \V1554(0)  = V769 | (\V731(0)  | (V710 | (\V729(0)  | (V721 | \V730(0) )))),
  V1070 = \V1421(0)  & (V2116 & (V2117 & \V1023(11) )),
  V1071 = \V1421(0)  & (V2116 & (V2117 & \V1023(10) )),
  \V1689(0)  = ~V1688,
  V1072 = \V1421(0)  & (V2116 & (V2117 & \V1023(9) )),
  V1073 = \V1421(0)  & (V2116 & (V2117 & \V1023(8) )),
  V1074 = \V1421(0)  & (V2116 & (V2117 & \V1023(7) )),
  V1075 = \V1421(0)  & (V2116 & (V2117 & \V1023(6) )),
  V1076 = \V1421(0)  & (V2116 & (V2117 & \V1023(5) )),
  V1077 = \V1421(0)  & (V2116 & (V2117 & \V1023(4) )),
  V1078 = V2118 & (V2119 & (\V1681(0)  & \V257(7) )),
  V1079 = V2120 & (V2121 & (V727 & (\V1446(0)  & (\V987(0)  & \V149(7) )))),
  \V423(0)  = \[9] ,
  V1081 = V2120 & (V2121 & (V727 & (\V1446(0)  & (\V987(0)  & \V149(6) )))),
  V1083 = V2120 & (V2121 & (V727 & (\V1446(0)  & (\V987(0)  & \V149(5) )))),
  V1085 = V2120 & (V2121 & (V727 & (\V1446(0)  & (\V987(0)  & \V149(4) )))),
  V1087 = \V1421(0)  & (V2122 & (V2123 & \V1053(3) )),
  V1088 = \V1421(0)  & (V2122 & (V2123 & \V1053(2) )),
  V1089 = \V1421(0)  & (V2122 & (V2123 & \V1053(1) )),
  V1090 = \V1421(0)  & (V2122 & (V2123 & \V1053(0) )),
  V1092 = \V32(8)  & \V1124(1) ,
  V1093 = \V32(7)  & \V1124(1) ,
  V1094 = \V32(6)  & \V1124(1) ,
  V1095 = \V32(5)  & \V1124(1) ,
  V1096 = \V32(4)  & \V1124(1) ,
  V1097 = \V32(3)  & \V1124(1) ,
  V1098 = \V32(2)  & \V1124(1) ,
  V1099 = \V32(1)  & \V1124(1) ,
  \V1492(0)  = \[134] ,
  \V1831(0)  = V1830 | V1834,
  \V361(0)  = ~V348,
  \V496(0)  = V495 | V494,
  \V835(0)  = ~V831,
  V1100 = \V32(0)  & \V1124(1) ,
  V1101 = \V1408(0)  & (V2125 & \V32(11) ),
  V1103 = \V1408(0)  & (V2125 & \V32(10) ),
  V1105 = \V1408(0)  & (V2125 & \V32(9) ),
  V1107 = \V1408(0)  & (V2125 & \V32(8) ),
  V1109 = \V1408(0)  & (V2125 & \V32(7) ),
  \V435(0)  = \[11] ,
  V1111 = \V1408(0)  & (V2125 & \V32(6) ),
  V1113 = \V1408(0)  & (V2125 & \V32(5) ),
  V1115 = \V1408(0)  & (V2125 & \V32(4) ),
  V1117 = \V1408(0)  & (V2125 & \V32(3) ),
  V1119 = \V1408(0)  & (V2125 & \V32(2) ),
  V1121 = \V1408(0)  & (V2125 & \V32(1) ),
  V1123 = \V1408(0)  & (V2125 & \V32(0) ),
  V1125 = \[52]  & \V1685(0) ,
  V1127 = V2126 & (\V1126(1)  & \V1069(11) ),
  V1128 = V2126 & (\V1126(1)  & \V1069(10) ),
  V1129 = V2126 & (\V1126(1)  & \V1069(9) ),
  V1130 = V2126 & (\V1126(1)  & \V1069(8) ),
  V1131 = V2126 & (\V1126(1)  & \V1069(7) ),
  V1132 = V2126 & (\V1126(1)  & \V1069(6) ),
  V1133 = V2126 & (\V1126(1)  & \V1069(5) ),
  V1134 = V1125 & (V2127 & \V1124(6) ),
  V1136 = V1125 & (V2127 & \V1124(5) ),
  V1138 = V1125 & (V2127 & \V1124(4) ),
  V1140 = V1125 & (V2127 & \V1124(3) ),
  V1142 = V1125 & (V2127 & \V1124(2) ),
  V1144 = V1125 & (V2127 & \V1124(1) ),
  V1146 = V1125 & (V2127 & (V2125 & \V1408(0) )),
  V1148 = V2128 & (\V1126(1)  & (V2122 & (V2123 & (\V1053(9)  & \V1421(0) )))),
  V1149 = V2128 & (\V1126(1)  & (V2122 & (V2123 & (\V1053(8)  & \V1421(0) )))),
  V1150 = V2128 & (\V1126(1)  & (V2122 & (V2123 & (\V1053(7)  & \V1421(0) )))),
  V1151 = V2128 & (\V1126(1)  & (V2122 & (V2123 & (\V1053(6)  & \V1421(0) )))),
  V1152 = V2128 & (\V1126(1)  & (V2122 & (V2123 & (\V1053(5)  & \V1421(0) )))),
  V1153 = V2128 & (\V1126(1)  & (V2122 & (V2123 & (\V1053(4)  & \V1421(0) )))),
  V1154 = V2128 & (\V1126(1)  & \V1086(3) ),
  V1155 = V2128 & (\V1126(1)  & \V1086(2) ),
  V1156 = V2128 & (\V1126(1)  & \V1086(1) ),
  V1157 = V2128 & (\V1126(1)  & \V1086(0) ),
  V1158 = V1125 & (V2129 & (\V32(11)  & \V1124(1) )),
  V1160 = V1125 & (V2129 & (\V32(10)  & \V1124(1) )),
  V1162 = V1125 & (V2129 & (\V32(9)  & \V1124(1) )),
  V1164 = V1125 & (V2129 & \V1124(13) ),
  V1166 = V1125 & (V2129 & \V1124(12) ),
  V1168 = V1125 & (V2129 & \V1124(11) ),
  V1170 = V1125 & (V2129 & \V1124(10) ),
  \V847(0)  = ~V846,
  V1172 = V1125 & (V2129 & \V1124(9) ),
  V1174 = V1125 & (V2129 & \V1124(8) ),
  V1176 = V1125 & (V2129 & \V1124(7) ),
  V1178 = V2130 & (\V1422(0)  & \V1147(11) ),
  V1179 = V2130 & (\V1422(0)  & \V1147(10) ),
  V1180 = V2130 & (\V1422(0)  & \V1147(9) ),
  V1181 = V2130 & (\V1422(0)  & \V1147(8) ),
  V1182 = V2130 & (\V1422(0)  & \V1147(7) ),
  V1183 = V2130 & (\V1422(0)  & \V1147(6) ),
  V1184 = V2130 & (\V1422(0)  & \V1147(5) ),
  V1185 = V2130 & (\V1422(0)  & (\V1126(1)  & (\V1069(4)  & V2126))),
  V1186 = V2130 & (\V1422(0)  & (\V1126(1)  & (V2116 & (V2117 & (\V1023(3)  & (\V1421(0)  & V2126)))))),
  V1187 = V2130 & (\V1422(0)  & (\V1126(1)  & (V2116 & (V2117 & (\V1023(2)  & (\V1421(0)  & V2126)))))),
  V1188 = V2130 & (\V1422(0)  & (\V1126(1)  & (V2116 & (V2117 & (\V1023(1)  & (\V1421(0)  & V2126)))))),
  V1189 = V2130 & (\V1422(0)  & (\V1126(1)  & (V2116 & (V2117 & (\V1023(0)  & (\V1421(0)  & V2126)))))),
  V1190 = \V1417(0)  & (V2131 & \V32(11) ),
  V1192 = \V1417(0)  & (V2131 & \V32(10) ),
  V1194 = \V1417(0)  & (V2131 & \V32(9) ),
  V1196 = \V1417(0)  & (V2131 & \V32(8) ),
  V1198 = \V1417(0)  & (V2131 & \V32(7) ),
  \V1781(1)  = \[171] ,
  \V1781(0)  = \[172] ,
  \V1720(0)  = ~\[160] ,
  \V1855(0)  = \V288(4)  | \V288(5) ,
  \V385(0)  = \V365(0)  | \V366(0) ,
  V1200 = \V1417(0)  & (V2131 & \V32(6) ),
  V1202 = \V1417(0)  & (V2131 & \V32(5) ),
  V1204 = \V1417(0)  & (V2131 & \V32(4) ),
  V1206 = \V1417(0)  & (V2131 & \V32(3) ),
  V1208 = \V1417(0)  & (V2131 & \V32(2) ),
  V1210 = \V1417(0)  & (V2131 & \V32(1) ),
  V1212 = \V1417(0)  & (V2131 & \V32(0) ),
  V1214 = V2132 & (\V1422(0)  & \V1177(9) ),
  V1215 = V2132 & (\V1422(0)  & \V1177(8) ),
  V1216 = V2132 & (\V1422(0)  & \V1177(7) ),
  V1217 = V2132 & (\V1422(0)  & \V1177(6) ),
  V1218 = V2132 & (\V1422(0)  & \V1177(5) ),
  V1219 = V2132 & (\V1422(0)  & \V1177(4) ),
  \V1455(0)  = V1453 | V1454,
  V1220 = V2132 & (\V1422(0)  & \V1177(3) ),
  V1221 = V2132 & (\V1422(0)  & \V1177(2) ),
  V1222 = V2132 & (\V1422(0)  & \V1177(1) ),
  V1223 = V2132 & (\V1422(0)  & \V1177(0) ),
  V1224 = \V1417(0)  & (V2133 & \V88(1) ),
  V1226 = \V1417(0)  & (V2133 & \V88(0) ),
  V1228 = \V1417(0)  & (V2133 & \V84(5) ),
  \V2067(0)  = V2066 | V2065,
  V1230 = \V1417(0)  & (V2133 & \V84(4) ),
  V1232 = \V1417(0)  & (V2133 & \V84(3) ),
  V1234 = \V1417(0)  & (V2133 & \V84(2) ),
  V1236 = \V1417(0)  & (V2133 & \V84(1) ),
  V1238 = \V1417(0)  & (V2133 & \V84(0) ),
  V1240 = \V1417(0)  & (V2133 & \V78(5) ),
  V1242 = \V1417(0)  & (V2133 & \V78(4) ),
  V1244 = V2134 & (\V1422(0)  & (\V1126(1)  & (V2116 & (V2117 & (\V1023(3)  & (\V1421(0)  & V2126)))))),
  V1245 = V2134 & (\V1422(0)  & (\V1126(1)  & (V2116 & (V2117 & (\V1023(2)  & (\V1421(0)  & V2126)))))),
  V1246 = V2134 & (\V1422(0)  & (\V1126(1)  & (V2116 & (V2117 & (\V1023(1)  & (\V1421(0)  & V2126)))))),
  V1247 = V2134 & (\V1422(0)  & (\V1126(1)  & (V2116 & (V2117 & (\V1023(0)  & (\V1421(0)  & V2126)))))),
  V1248 = \V1417(0)  & (V2135 & \V32(3) ),
  V1250 = \V1417(0)  & (V2135 & \V32(2) ),
  V1252 = \V1417(0)  & (V2135 & \V32(1) ),
  V1254 = \V1417(0)  & (V2135 & \V32(0) ),
  V1256 = \[92] ,
  V1257 = \[93] ,
  V1258 = \[94] ,
  V1259 = \[95] ,
  V1260 = \[96] ,
  V1261 = \[97] ,
  V1262 = \[98] ,
  V1263 = \[99] ,
  V1264 = \[100] ,
  V1265 = \[101] ,
  V1266 = \[102] ,
  V1267 = \[103] ,
  V1269 = ~\V1268(0) ,
  V1270 = ~V767,
  V1271 = ~V768,
  V1272 = \V62(0)  & (V502 & (V964 & V498)),
  V1273 = V498 & (V964 & (V754 & (V1270 & (V1269 & (V1271 & (\V59(0)  & \V1720(0) )))))),
  V1276 = \V56(0)  & V735,
  V1279 = V2136 & (\V1278(1)  & (\V213(0)  & (\V14(0)  & \V1277(0) ))),
  V1280 = \V1984(0)  & (V2137 & \V1546(0) ),
  V1283 = V2138 & (\V1282(1)  & (\V213(5)  & (\V14(0)  & \V1277(0) ))),
  V1284 = V2138 & (\V1282(1)  & (\V213(4)  & (\V14(0)  & \V1277(0) ))),
  V1285 = V2138 & (\V1282(1)  & (\V213(3)  & (\V14(0)  & \V1277(0) ))),
  V1286 = V2138 & (\V1282(1)  & (\V213(2)  & (\V14(0)  & \V1277(0) ))),
  V1287 = V2138 & (\V1282(1)  & (\V213(1)  & (\V14(0)  & \V1277(0) ))),
  V1288 = V1979 & (V2139 & \V165(7) ),
  V1290 = V1979 & (V2139 & \V165(6) ),
  V1292 = V1979 & (V2139 & \V165(5) ),
  V1294 = V1979 & (V2139 & \V165(4) ),
  V1296 = V1979 & (V2139 & \V165(3) ),
  V1298 = V2513 | V2512,
  V1299 = V2025 & V1846,
  \V1467(0)  = \[130] ,
  \V336(0)  = V332 | (V323 | (V329 | V335)),
  \V1670(0)  = ~\V204(0) ,
  \V2018(0)  = V2013 | (V2012 | V2014),
  V1300 = V2517 | V2516,
  V1301 = V2521 | V2520,
  V1302 = V2525 | V2524,
  V1303 = V1299 & V1848,
  V1304 = V1299 & V2029,
  V1305 = V1848 & V2029,
  V1307 = V2529 | V2528,
  V1308 = \V1306(0)  & V1839,
  V1309 = \V1306(0)  & V2034,
  \V686(3)  = ~\V667(3) ,
  V1310 = V1839 & V2034,
  V1312 = V2533 | V2532,
  V1313 = ~V1298,
  V1314 = ~V1302,
  V1315 = ~V1307,
  V1316 = V2537 | V2536,
  V1317 = V1313 & V1314,
  V1318 = V2541 | V2540,
  V1319 = V1317 & V1315,
  V1320 = V2545 | V2544,
  V1321 = ~V1313,
  V1322 = ~V1316,
  V1323 = ~V1318,
  V1324 = V2549 | V2548,
  V1325 = V1321 & V1322,
  V1326 = V2553 | V2552,
  V1327 = V1325 & V1323,
  V1328 = V2557 | V2556,
  V1329 = V2140 & (V1848 & V1312),
  \V686(5)  = ~\V667(5) ,
  V1330 = \V1860(0)  & (V2141 & V1328),
  V1332 = V2142 & (V1848 & V1307),
  V1333 = \V1860(0)  & (V2143 & V1326),
  V1335 = V2144 & (V1848 & V1302),
  V1336 = \V1860(0)  & (V2145 & V1324),
  V1338 = V2146 & (V1848 & V1298),
  V1339 = \V1860(0)  & (V2147 & V1321),
  \V686(4)  = ~\V667(4) ,
  V1341 = ~\V1340(0) ,
  V1342 = ~\V1337(0) ,
  V1343 = ~\V1334(0) ,
  V1344 = V2561 | V2560,
  V1345 = V1341 & V1342,
  V1346 = V2565 | V2564,
  V1347 = V1345 & V1343,
  V1348 = V2569 | V2568,
  V1349 = V2148 & (V1846 & V1312),
  V1350 = \V1859(0)  & (V2149 & V1348),
  V1352 = V2150 & (V1846 & V1307),
  V1353 = \V1859(0)  & (V2151 & V1346),
  V1355 = V2152 & (V1846 & V1302),
  V1356 = \V1859(0)  & (V2153 & V1344),
  V1358 = V2154 & (V1846 & V1298),
  V1359 = \V1859(0)  & (V2155 & V1341),
  V1361 = ~V734,
  V1362 = ~V515,
  V1363 = ~\V731(0) ,
  V1364 = ~V738,
  V1365 = \[111] ,
  V1366 = \V268(4)  & (\V268(2)  & (\V268(1)  & (\V268(3)  & \V268(5) ))),
  V1367 = \V268(4)  & (\V268(2)  & (\V268(3)  & \V268(5) )),
  V1368 = \V268(4)  & (\V268(3)  & \V268(5) ),
  V1369 = \V268(4)  & \V268(5) ,
  V1370 = \[219] ,
  V1371 = \[220] ,
  V1372 = \[221] ,
  V1373 = \[222] ,
  V1374 = \[223] ,
  V1375 = \[112] ,
  V1376 = ~\V2010(0) ,
  V1377 = ~\V374(0) ,
  V1378 = \[113] ,
  V1379 = ~\V2020(0) ,
  V1380 = \[114] ,
  V1381 = ~\V381(0) ,
  V1382 = \[115] ,
  V1383 = ~\V342(0) ,
  V1384 = \[116] ,
  \V1282(1)  = ~V1979,
  V1385 = ~\V1837(0) ,
  V1386 = \[117] ,
  V1387 = \[118] ,
  V1390 = \V1388(0)  & (\V65(0)  & (\V1389(0)  & (V964 & V498))),
  V1391 = \V70(0)  & (\V165(6)  & (\V694(4)  & (\V165(3)  & (\V694(5)  & (\[52]  & (V964 & V498)))))),
  V1393 = \V1446(0)  & V769,
  \V686(7)  = ~\V667(7) ,
  \V686(6)  = ~\V667(6) ,
  \V1694(1)  = ~V1978,
  V1400 = ~V727,
  V1401 = ~V726,
  V1402 = \V1394(0)  & \[52] ,
  V1403 = V1445 & V727,
  V1404 = \V1396(0)  & (\V1446(0)  & V727),
  V1405 = ~\V1415(0) ,
  V1406 = \V1398(0)  & (\V1397(0)  & V1405),
  V1407 = \V1399(0)  & \V60(0) ,
  \V902(0)  = ~V898,
  V1411 = V502 & \V56(0) ,
  V1412 = V502 & \V60(0) ,
  V1413 = V411 & \V56(0) ,
  V1414 = V411 & \V60(0) ,
  V1416 = \V967(0)  & (\V53(0)  & (V1400 & (V1401 & V793))),
  V1418 = \V1409(0)  & \V765(0) ,
  V1419 = ~\V1417(0) ,
  V1420 = ~\V1410(0) ,
  V1423 = \[120] ,
  V1424 = ~\V583(0) ,
  V1425 = V1424 & V786,
  V1426 = \[121] ,
  V1427 = \V109(0)  & \V658(0) ,
  V1428 = \[122] ,
  V1429 = \[123] ,
  V1430 = ~V1427,
  V1431 = \[124] ,
  V1432 = \[125] ,
  V1433 = ~V769,
  V1434 = ~\V1441(0) ,
  V1435 = V498 & (V1433 & V1434),
  V1436 = V769 & \V277(0) ,
  V1438 = \V1437(0)  & \V14(0) ,
  V1443 = \V277(0)  & V769,
  V1445 = \V1444(0)  & \V278(0) ,
  V1448 = \V1452(0)  & (\V14(0)  & \V1447(0) ),
  V1449 = ~\V1447(0) ,
  V1450 = \V258(0)  & (\V14(0)  & V1449),
  V1453 = \V258(0)  & V1830,
  V1454 = \V1452(0)  & V1836,
  V1456 = \V14(0)  & (\V1455(0)  & \V1460(0) ),
  V1457 = ~\V1455(0) ,
  V1458 = \V14(0)  & (V1457 & \V259(0) ),
  V1461 = \V259(0)  & V1453,
  V1462 = \V1460(0)  & V1454,
  V1464 = \V14(0)  & (\V1463(0)  & \V1468(0) ),
  V1465 = ~\V1463(0) ,
  V1466 = \V14(0)  & (V1465 & \V260(0) ),
  V1469 = ~V737,
  V1470 = \[131] ,
  V1473 = \V1471(0)  & \[65] ,
  V1474 = \V1472(0)  & \V56(0) ,
  V1476 = \V1475(0)  & \V1597(0) ,
  V1477 = ~V701,
  V1478 = \[165]  & V1477,
  V1479 = V701 & (\[165]  & \[65] ),
  V1482 = ~\V66(0) ,
  V1483 = ~\V68(0) ,
  V1484 = ~\V69(0) ,
  V1485 = ~\V70(0) ,
  V1486 = V1484 & (V1482 & (V1483 & V1485)),
  V1487 = ~V1486,
  V1488 = ~\V1999(0) ,
  V1489 = ~\V1493(0) ,
  V1490 = V1488 & (V1487 & (V498 & V1489)),
  V1491 = \V66(0)  & \V215(0) ,
  V1494 = \V216(0)  & \[133] ,
  V1497 = \V536(0)  & (\V1496(0)  & \V346(0) ),
  V1499 = ~\V2002(0) ,
  \V914(0)  = ~V910,
  \V1645(0)  = \[148] ,
  \V1983(0)  = V1981 | V1978,
  \V852(0)  = ~V848,
  \V987(0)  = ~\V59(0) ,
  V1500 = ~\V346(0) ,
  V1501 = V1499 & V1500,
  V1503 = \V1496(0)  & \[139] ,
  V1504 = \V1498(0)  & \[139] ,
  V1505 = \V1502(0)  & \[139] ,
  V1506 = ~\[139] ,
  V1507 = \V371(0)  & V1506,
  V1509 = \V370(0)  & V1506,
  V1511 = \V369(0)  & V1506,
  V1513 = \V278(0)  & \V2011(0) ,
  V1515 = ~\V274(0) ,
  V1516 = V497 & V1515,
  V1517 = \V172(0)  & \V56(0) ,
  V1518 = \V171(0)  & (\V1395(0)  & \V56(0) ),
  V1519 = ~\V1514(0) ,
  V1520 = ~\V248(0) ,
  V1521 = ~V1513,
  V1522 = ~V1517,
  V1523 = ~V1518,
  V1524 = V1522 & (V1520 & (V1519 & (V1521 & V1523))),
  V1525 = ~\V172(0) ,
  V1526 = V406 & V1525,
  V1527 = V515 & \V59(0) ,
  V1528 = ~V1516,
  V1529 = ~V1524,
  V1530 = ~V1526,
  V1531 = ~V1527,
  V1532 = V1530 & (V1528 & (V1529 & V1531)),
  V1533 = ~V1532,
  V1534 = ~\V536(0) ,
  V1535 = V1534 & (V1533 & V1499),
  V1537 = \[140] ,
  V1539 = \[141] ,
  V1540 = ~\V165(3) ,
  V1541 = ~\V165(4) ,
  V1542 = ~\V165(5) ,
  V1543 = ~\V165(6) ,
  V1544 = ~\V165(7) ,
  V1545 = V1543 & (V1541 & (V1540 & (V1542 & V1544))),
  V1547 = V2156 & (V721 & (\V803(0)  & V1985)),
  V1548 = V2156 & (V721 & (\V803(0)  & V1986)),
  V1549 = V379 & (V2157 & \[82] ),
  V1551 = V379 & (V2157 & \[83] ),
  V1555 = \V1554(0)  & \V57(0) ,
  V1556 = ~\V57(0) ,
  V1557 = V739 & V1556,
  V1558 = V745 & \V1553(0) ,
  V1559 = ~V1555,
  V1560 = ~V1557,
  V1561 = ~V1558,
  V1562 = ~\V174(0) ,
  V1563 = ~\V35(0) ,
  V1564 = \V71(0)  & \V202(0) ,
  V1566 = ~\[186] ,
  V1567 = ~\V1720(0) ,
  V1568 = V1566 & V1567,
  V1569 = V697 & \[160] ,
  V1570 = \[160]  & V698,
  V1571 = \[160]  & (V1867 & \V394(0) ),
  V1572 = \V247(0)  & (\[160]  & (V605 & \V394(0) )),
  V1573 = ~V1571,
  V1574 = ~V392,
  V1575 = ~V1568,
  V1576 = ~V1569,
  V1577 = ~V1570,
  V1578 = ~V1572,
  V1579 = V2593 | V2592,
  \V1860(0)  = ~V1848,
  V1580 = V2597 | V2596,
  V1581 = V2601 | V2600,
  V1582 = V2605 | V2604,
  V1583 = V2609 | V2608,
  V1584 = V2613 | V2612,
  V1585 = V2617 | V2616,
  V1586 = V2621 | V2620,
  V1587 = V2625 | V2624,
  V1588 = V2629 | V2628,
  V1589 = V2633 | V2632,
  \V864(0)  = ~V860,
  V1590 = V2637 | V2636,
  V1591 = V2641 | V2640,
  V1592 = V2645 | V2644,
  V1593 = V2649 | V2648,
  V1594 = V2653 | V2652,
  V1598 = V2657 | V2656,
  V1599 = V2661 | V2660,
  \V1460(0)  = ~\V259(0) ,
  \V803(0)  = ~\[65] ,
  \V2011(0)  = \V2007(0)  | V726,
  V1600 = V2665 | V2664,
  V1601 = V2669 | V2668,
  V1602 = V2673 | V2672,
  V1603 = V2677 | V2676,
  V1604 = V2681 | V2680,
  V1605 = V2685 | V2684,
  V1606 = V2689 | V2688,
  V1607 = V2693 | V2692,
  V1608 = V2697 | V2696,
  V1609 = V2701 | V2700,
  V1610 = V2705 | V2704,
  V1611 = V2709 | V2708,
  V1614 = \[186]  & \V292(0) ,
  V1615 = \V174(0)  & V695,
  V1616 = \V174(0)  & \V2002(0) ,
  V1617 = ~V799,
  V1618 = ~\V291(0) ,
  V1619 = ~\V292(0) ,
  V1621 = \V91(0)  & \V59(0) ,
  V1622 = \V91(1)  & \V62(0) ,
  V1624 = \V1623(0)  & V739,
  V1625 = ~\V294(0) ,
  V1626 = ~V611,
  V1627 = ~V741,
  V1628 = V1626 & (V1625 & V1627),
  \V1472(0)  = V744 | (V745 | V739),
  V1633 = \V764(0)  & (\V1631(0)  & \[65] ),
  V1634 = \[65]  & V701,
  V1635 = V737 & \V66(0) ,
  V1636 = \V1632(0)  & \V56(0) ,
  V1637 = \V66(0)  & \[52] ,
  V1638 = \V149(7)  & (V701 & \[65] ),
  V1639 = V766 & V687,
  V1640 = V701 & \[186] ,
  \V476(0)  = V475 | V474,
  V1643 = \V1641(0)  & \V336(0) ,
  V1644 = V338 & (V1646 & (\V1642(0)  & (V344 & \V14(0) ))),
  V1646 = V1522 & \V207(0) ,
  \V2084(0)  = V2083 | V2082,
  V1648 = \V1647(0)  & V1445,
  V1650 = ~\V290(0) ,
  V1651 = V1650 & (\V295(0)  & (\V1649(0)  & (\V399(0)  & (\V1685(0)  & V344)))),
  V1654 = ~\V1653(0) ,
  V1655 = ~\V1687(0) ,
  V1656 = V1627 & (V1655 & (V1654 & (V804 & V805))),
  V1657 = ~V1656,
  V1658 = ~\V812(0) ,
  V1659 = ~V696,
  V1660 = V1659 & (V1657 & (V1499 & (V1658 & V344))),
  V1661 = ~\V1746(0) ,
  V1662 = V1661 & (V1654 & V344),
  V1663 = \V803(0)  & (V698 & V344),
  \V1546(0)  = V1545 | V1646,
  V1664 = \V66(0)  & V737,
  V1665 = ~V1660,
  V1666 = ~V1662,
  V1667 = ~V1663,
  V1668 = ~V1664,
  V1669 = \[150] ,
  \V1023(7)  = V1008 | V992,
  V1672 = \V165(2)  & (\V165(1)  & (\V165(0)  & (\V1670(0)  & (\V261(0)  & (\V165(4)  & (\V165(3)  & (\V165(5)  & (\V165(6)  & \V165(7) )))))))),
  V1673 = \[52]  & (\V165(2)  & (\V165(1)  & (\V165(0)  & (\V165(6)  & (\V165(4)  & (\V165(3)  & (\V165(5)  & (\V261(0)  & (\V165(7)  & \V70(0) ))))))))),
  V1675 = \V258(0)  & (\V1468(0)  & (\V1460(0)  & \V987(0) )),
  V1676 = ~\V1680(0) ,
  V1677 = ~V1675,
  V1678 = V1677 & (V1676 & V498),
  \V1023(6)  = V1010 | V993,
  V1682 = ~V1678,
  V1683 = \V1835(0)  & (V1682 & V1676),
  V1686 = \V262(0)  & V1678,
  V1688 = \V56(0)  & V736,
  \V1023(9)  = V1004 | V990,
  V1691 = V2158 & (\V1690(1)  & (\V100(0)  & (\V14(0)  & \V1689(0) ))),
  V1692 = \V1983(0)  & (V2159 & \V1546(0) ),
  V1695 = V2160 & (\V1694(1)  & (\V100(5)  & (\V14(0)  & \V1689(0) ))),
  V1696 = V2160 & (\V1694(1)  & (\V100(4)  & (\V14(0)  & \V1689(0) ))),
  V1697 = V2160 & (\V1694(1)  & (\V100(3)  & (\V14(0)  & \V1689(0) ))),
  V1698 = V2160 & (\V1694(1)  & (\V100(2)  & (\V14(0)  & \V1689(0) ))),
  V1699 = V2160 & (\V1694(1)  & (\V100(1)  & (\V14(0)  & \V1689(0) ))),
  \V1023(8)  = V1006 | V991,
  \V1023(10)  = V1002 | V989,
  \V1023(11)  = V1000 | V988,
  \V827(0)  = ~\V280(0) ,
  V1700 = V1978 & (V2161 & \V165(7) ),
  V1702 = V1978 & (V2161 & \V165(6) ),
  V1704 = V1978 & (V2161 & \V165(5) ),
  V1706 = V1978 & (V2161 & \V165(4) ),
  V1708 = V1978 & (V2161 & \V165(3) ),
  \V1023(1)  = V1020 | V998,
  V1710 = V721 & \V827(0) ,
  V1712 = \V1711(0)  & \[65] ,
  V1713 = ~V1710,
  V1714 = ~\V1718(0) ,
  V1715 = ~V697,
  V1716 = V1525 & (V1714 & (V1713 & (V964 & (V1715 & V338)))),
  V1719 = \[160] ,
  \V1023(0)  = V1022 | V999,
  V1721 = V1867 & \V194(0) ,
  V1722 = ~\[139] ,
  V1723 = V1722 & (V1721 & \V2011(0) ),
  V1724 = ~\V2007(0) ,
  V1725 = V1724 & (\V242(0)  & V498),
  \V1761(0)  = ~V745,
  \V1896(0)  = \[187] ,
  V1729 = \V1728(0)  & \V241(0) ,
  \V1023(3)  = V1016 | V996,
  V1730 = \V733(0)  & (V1364 & (V1271 & (V1646 & V1477))),
  V1731 = \V59(0)  & (V1646 & (V687 & V1477)),
  V1732 = V768 & (V1646 & (\V59(0)  & V1477)),
  V1733 = \V62(0)  & (V1646 & (V738 & V1477)),
  V1734 = ~V1729,
  \V765(0)  = ~\V174(0) ,
  V1735 = V1734 & V1401,
  V1736 = \[162] ,
  V1737 = ~V1735,
  V1738 = V1730 & V338,
  V1739 = V1731 & V338,
  \V1023(2)  = V1018 | V997,
  V1740 = V338 & V1732,
  V1742 = ~V725,
  V1743 = ~V747,
  V1744 = V1742 & (\V289(0)  & (\V33(0)  & V1743)),
  V1748 = \V290(0)  & V695,
  V1749 = V751 & \V56(0) ,
  \V1023(5)  = V1012 | V994,
  V1750 = \V15(0)  & \V16(0) ,
  \V1496(0)  = ~\V2002(0) ,
  V1751 = \V15(0)  & \V1866(0) ,
  V1752 = \V1865(0)  & \V16(0) ,
  V1754 = V1752 & V700,
  V1755 = \V14(0)  & (\V1753(0)  & \V101(0) ),
  V1756 = V1752 & V725,
  \V1835(0)  = \V62(0)  | (\V56(0)  | \V50(0) ),
  \V1023(4)  = V1014 | V995,
  \V365(0)  = ~V352,
  V1764 = V2162 & (V745 & \V1763(1) ),
  V1765 = V2162 & (V745 & \V1763(0) ),
  V1768 = \V1761(0)  & (V2163 & \V1767(1) ),
  V1770 = \V1761(0)  & (V2163 & \V1767(0) ),
  V1774 = V2164 & (\V1761(0)  & \V1773(1) ),
  V1775 = V2164 & (\V1761(0)  & \V1773(0) ),
  V1778 = V745 & (V2165 & \V1777(1) ),
  V1780 = V745 & (V2165 & \V1777(0) ),
  V1782 = ~\[79] ,
  V1792 = V2166 & (\V37(0)  & \V1791(8) ),
  V1793 = V2166 & (\V37(0)  & \V1791(7) ),
  V1794 = V2166 & (\V37(0)  & \V1791(6) ),
  V1795 = V2166 & (\V37(0)  & \V1791(5) ),
  V1796 = V2166 & (\V37(0)  & \V1791(4) ),
  V1797 = V2166 & (\V37(0)  & \V1791(3) ),
  V1798 = V2166 & (\V37(0)  & \V1791(2) ),
  V1799 = V2166 & (\V37(0)  & \V1791(1) ),
  \V1773(1)  = ~\[70] ,
  \V1773(0)  = ~\[71] ,
  \V642(0)  = ~\V274(0) ,
  \V777(0)  = \V52(0)  | V776,
  V1800 = V2166 & (\V37(0)  & \V1791(0) ),
  V1801 = V2166 & (\V37(0)  & V1782),
  \V1447(0)  = V1830 | V1836,
  V1810 = \V436(0)  & (V2167 & \[0] ),
  V1812 = \V436(0)  & (V2167 & \V1809(7) ),
  V1814 = \V436(0)  & (V2167 & \V1809(6) ),
  V1816 = \V436(0)  & (V2167 & \V1809(5) ),
  V1818 = \V436(0)  & (V2167 & \V1809(4) ),
  V1820 = \V436(0)  & (V2167 & \V1809(3) ),
  V1822 = \V436(0)  & (V2167 & \V1809(2) ),
  V1824 = \V436(0)  & (V2167 & \V1809(1) ),
  V1826 = \V436(0)  & (V2167 & \V1809(0) ),
  V1828 = \V436(0)  & (V2167 & \[0] ),
  V1830 = V1366 & \V268(0) ,
  V1832 = \[183] ,
  V1834 = \V261(0)  & \V1684(0) ,
  V1836 = \V1835(0)  & \V1681(0) ,
  V1838 = \V288(0)  & \V288(1) ,
  V1839 = \V288(2)  & \V288(3) ,
  V1840 = \V288(4)  & \V288(5) ,
  V1841 = ~\V288(4) ,
  V1842 = V1841 & \V288(5) ,
  V1843 = ~\V288(5) ,
  V1844 = \V288(4)  & V1843,
  V1845 = ~\V288(2) ,
  V1846 = V1845 & \V288(3) ,
  V1847 = ~\V288(3) ,
  V1848 = \V288(2)  & V1847,
  V1849 = ~\V288(0) ,
  V1850 = V1849 & \V288(1) ,
  V1851 = ~\V288(1) ,
  V1852 = \V288(0)  & V1851,
  V1867 = \V199(3)  & (\V199(1)  & (\V194(4)  & (\V194(2)  & (\V194(1)  & (\V194(3)  & (\V199(0)  & (\V199(2)  & \V199(4) ))))))),
  V1868 = \V199(3)  & (\V199(1)  & (\V194(4)  & (\V194(2)  & (\V194(3)  & (\V199(0)  & (\V199(2)  & \V199(4) )))))),
  V1869 = \V199(3)  & (\V199(1)  & (\V194(4)  & (\V194(3)  & (\V199(0)  & (\V199(2)  & \V199(4) ))))),
  V1870 = \V199(3)  & (\V199(1)  & (\V194(4)  & (\V199(0)  & (\V199(2)  & \V199(4) )))),
  V1871 = \V199(3)  & (\V199(1)  & (\V199(0)  & (\V199(2)  & \V199(4) ))),
  V1872 = \V199(3)  & (\V199(1)  & (\V199(2)  & \V199(4) )),
  V1873 = \V199(3)  & (\V199(2)  & \V199(4) ),
  V1874 = \V199(3)  & \V199(4) ,
  \V1859(0)  = ~V1846,
  V1875 = V2713 | V2712,
  V1876 = V2717 | V2716,
  V1877 = V2721 | V2720,
  V1878 = V2725 | V2724,
  V1879 = V2729 | V2728,
  V1880 = V2733 | V2732,
  V1881 = V2737 | V2736,
  V1882 = V2741 | V2740,
  V1883 = V2745 | V2744,
  V1884 = ~\V199(4) ,
  V1885 = V1476 & V769,
  V1886 = V1995 & V725,
  V1887 = V1995 & V700,
  V1888 = ~V1902,
  \[0]  = ~\[91] ,
  V1889 = V1888 & \V108(0) ,
  V1890 = V1888 & \V108(1) ,
  V1891 = V1888 & \V108(2) ,
  V1892 = V1888 & \V108(3) ,
  V1893 = V1888 & \V108(4) ,
  V1894 = ~V1749,
  V1895 = V1894 & \V108(5) ,
  \[1]  = \V937(0)  & (\V897(0)  & (\V857(0)  & (\V958(0)  & (\V956(0)  & (\V837(0)  & (\V877(0)  & (\V917(0)  & V347))))))),
  \V1459(0)  = \[129] ,
  \[2]  = \V947(0)  & (\V907(0)  & (\V867(0)  & (\V959(0)  & (\V957(0)  & (\V847(0)  & (\V887(0)  & (\V927(0)  & \V1685(0) ))))))),
  \V592(0)  = ~\V244(0) ,
  \[3]  = \V10(0)  & \V13(0) ,
  \[4]  = \[120]  | (V1425 | (\[94]  | (\[124]  | (\[61]  | (\[54]  | (\[56]  | (\[118]  | (\[95]  | (\[99]  | \[62] ))))))))),
  \[5]  = \V376(0)  & \V203(0) ,
  \[6]  = V1571 | (V392 | V1572),
  \[7]  = ~V397,
  \V1397(0)  = V721 | (\V729(0)  | (V710 | (\V731(0)  | V1393))),
  V1902 = V750 & \V56(0) ,
  V1904 = V2168 & (V2169 & (V2170 & (V736 & \V100(5) ))),
  V1905 = V2168 & (V2169 & (V2170 & (V736 & \V100(4) ))),
  V1906 = V2168 & (V2169 & (V2170 & (V736 & \V100(3) ))),
  V1907 = V2168 & (V2169 & (V2170 & (V736 & \V100(2) ))),
  \V1213(7)  = \[74] ,
  V1908 = V2168 & (V2169 & (V2170 & (V736 & \V100(1) ))),
  \[8]  = ~V409,
  V1909 = V2168 & (V2169 & (V2170 & (V736 & \V100(0) ))),
  V1910 = V2171 & (V2172 & (V735 & (V2173 & \V213(5) ))),
  V1912 = V2171 & (V2172 & (V735 & (V2173 & \V213(4) ))),
  V1914 = V2171 & (V2172 & (V735 & (V2173 & \V213(3) ))),
  V1916 = V2171 & (V2172 & (V735 & (V2173 & \V213(2) ))),
  \V1213(6)  = \[75] ,
  V1918 = V2171 & (V2172 & (V735 & (V2173 & \V213(1) ))),
  \[9]  = V420 | (V402 | (V417 | (V415 | (V416 | (V419 | (\[160]  | V422)))))),
  V1920 = V2171 & (V2172 & (V735 & (V2173 & \V213(0) ))),
  V1922 = V2174 & (V742 & (V2175 & (V2176 & \V124(5) ))),
  V1923 = V2174 & (V742 & (V2175 & (V2176 & \V124(4) ))),
  V1924 = V2174 & (V742 & (V2175 & (V2176 & \V124(3) ))),
  V1925 = V2174 & (V742 & (V2175 & (V2176 & \V124(2) ))),
  V1926 = V2174 & (V742 & (V2175 & (V2176 & \V124(1) ))),
  V1927 = V2174 & (V742 & (V2175 & (V2176 & \V124(0) ))),
  \V1213(9)  = \[72] ,
  V1928 = V750 & (V2177 & (V2178 & (V2179 & \V108(4) ))),
  V1929 = V750 & (V2177 & (V2178 & (V2179 & \V108(3) ))),
  V1930 = V750 & (V2177 & (V2178 & (V2179 & \V108(2) ))),
  V1931 = V750 & (V2177 & (V2178 & (V2179 & \V108(1) ))),
  V1932 = V750 & (V2177 & (V2178 & (V2179 & \V108(0) ))),
  V1933 = V2180 & (V2181 & (V742 & \V132(7) )),
  V1934 = V2180 & (V2181 & (V742 & \V132(6) )),
  V1935 = V2180 & (V2181 & (V742 & \V132(5) )),
  V1936 = V2180 & (V2181 & (V742 & \V132(4) )),
  V1937 = V2180 & (V2181 & (V742 & \V132(3) )),
  \V1213(8)  = \[73] ,
  V1938 = V2180 & (V2181 & (V742 & \V132(2) )),
  V1940 = V2180 & (V2181 & (V742 & \V132(0) )),
  V1941 = V2182 & (V743 & (V2183 & \V118(5) )),
  V1943 = V2182 & (V743 & (V2183 & \V118(4) )),
  \V943(0)  = ~V939,
  V1945 = V2182 & (V743 & (V2183 & \V118(3) )),
  V1947 = V2182 & (V743 & (V2183 & \V118(2) )),
  V1949 = V2182 & (V743 & (V2183 & \V118(1) )),
  V1951 = V2182 & (V743 & (V2183 & \V118(0) )),
  V1954 = V751 & (V2184 & (V2185 & \V108(5) )),
  V1955 = V2186 & (V743 & \V118(7) ),
  V1956 = V2186 & (V743 & \V118(6) ),
  V1957 = \V382(0)  & (V2187 & \V46(0) ),
  V1959 = \V382(0)  & (V2187 & \V48(0) ),
  \V1674(0)  = V1672 | V1673,
  V1961 = V743 & \V56(0) ,
  V1962 = \V101(0)  & (V1751 & \V1903(4) ),
  V1966 = V700 & (\V1963(0)  & V1969),
  V1967 = \V14(0)  & (\V1964(0)  & (\V1965(0)  & \V110(0) )),
  V1969 = ~\V110(0) ,
  V1970 = ~\V288(6) ,
  V1971 = ~\V288(7) ,
  V1972 = V1970 & V1971,
  V1973 = V2749 | V2748,
  V1974 = V1970 & \V288(7) ,
  V1978 = \V290(0)  & (\V1977(0)  & V695),
  V1979 = V725 & (\V290(0)  & V695),
  \V1613(1)  = \[145] ,
  V1980 = ~V1644,
  V1981 = V1743 & (V1980 & (V1646 & (V338 & \V1977(0) ))),
  V1982 = V1743 & (V1980 & (V1646 & (V338 & V725))),
  V1985 = ~\V239(4) ,
  V1986 = V2753 | V2752,
  V1987 = V2188 & (V2006 & (\V2010(0)  & V1993)),
  V1988 = V2188 & (V2006 & (\V2010(0)  & V1994)),
  \V1274(0)  = \[104] ,
  V1989 = V2189 & (V2016 & (V2017 & \V134(1) )),
  \V1613(0)  = \[144] ,
  V1991 = V2189 & (V2016 & (V2017 & \V134(0) )),
  V1993 = ~\V134(1) ,
  V1994 = V2757 | V2756,
  V1995 = \V215(0)  & (\V172(0)  & \V67(0) ),
  V1996 = \V803(0)  & (V1737 & (\V261(0)  & \V1446(0) )),
  V1997 = V1445 & (V643 & (\V272(0)  & (\V803(0)  & (V1737 & \V261(0) )))),
  \V1213(1)  = \[80] ,
  \V1213(0)  = \[81] ,
  \V1213(3)  = \[78] ,
  \V1213(2)  = \[79] ,
  \V1213(5)  = \[76] ,
  \V1213(4)  = \[77] ,
  \V629(0)  = \V270(0)  | (V626 | (V627 | V628)),
  \V893(0)  = ~V889,
  \V1963(0)  = \[166]  | \V102(0) ,
  \V493(0)  = V492 | V491,
  \V832(0)  = ~V828,
  \V967(0)  = ~\V56(0) ,
  \V1502(0)  = ~V1501,
  \V1975(0)  = ~V1973,
  \V370(0)  = ~V359,
  \V844(0)  = ~V840,
  \V1440(0)  = \[127] ,
  \V1514(0)  = ~\V177(0) ,
  \V1649(0)  = ~V1648,
  \V321(2)  = \[0] ,
  \V382(0)  = V740 | V741,
  \V1452(0)  = ~\V258(0) ,
  \V2064(0)  = V2063 | V2062,
  \V1126(1)  = ~V1125,
  \V1864(0)  = \[186] ,
  \V1999(0)  = V1732 | (V1730 | (V1995 | (\V214(0)  | (V1731 | V1733)))),
  \V394(0)  = ~\V248(0) ,
  \V733(0)  = V732 | V688,
  \V807(0)  = \V2002(0)  | (V698 | (\V302(0)  | V696)),
  \V1538(0)  = \V69(0)  | \V50(0) ,
  \V1741(0)  = \[163] ,
  \V610(0)  = ~\V247(0) ,
  \V1415(0)  = V1413 | (V1411 | (V1412 | V1414)),
  \V1753(0)  = ~V1749,
  \V622(0)  = ~\V533(0) ,
  \V572(3)  = \[35] ,
  \V1630(0)  = ~\V14(0) ,
  \V572(2)  = \[36] ,
  \V634(0)  = \[48] ,
  \V572(5)  = \[33] ,
  \V572(4)  = \[34] ,
  \V369(0)  = ~V358,
  \V1439(0)  = \[126] ,
  \V572(1)  = \[37] ,
  \V572(0)  = \[38] ,
  \V1777(1)  = ~\V78(3) ,
  \V1642(0)  = V738 | (V1639 | (V768 | V1640)),
  \V1777(0)  = ~\V78(2) ,
  \V511(0)  = \[14] ,
  \V572(7)  = \[31] ,
  \V572(6)  = \[32] ,
  \V572(9)  = \[29] ,
  \V572(8)  = \[30] ,
  \V584(0)  = ~\V7(0) ,
  \V923(0)  = ~V919,
  \V658(0)  = ~\V13(0) ,
  \V1992(1)  = \[210] ,
  \V1389(0)  = ~V741,
  \V1728(0)  = V769 | V727,
  \V1992(0)  = \[211] ,
  \V800(0)  = ~\V759(0) ,
  \V935(0)  = ~V931,
  \[100]  = \V12(0)  & \V4(0) ,
  \[101]  = \[100]  & \V52(0) ,
  \[102]  = \V11(0)  & \V4(0) ,
  \V609(0)  = \[44] ,
  \V873(0)  = ~V869,
  \[103]  = \V11(0)  & \V2(0) ,
  \[104]  = V1273 | V1272,
  \V473(0)  = V472 | V471,
  \[105]  = V1280 | V1279,
  \V2081(0)  = V2080 | V2079,
  \V812(0)  = V811 | (V808 | V981),
  \V947(0)  = ~V946,
  \[106]  = V1288 | V1283,
  \[107]  = V1290 | V1284,
  \V412(0)  = V721 | (\V729(0)  | (V710 | (\V1681(0)  | \V731(0) ))),
  \[108]  = V1292 | V1285,
  \V2020(0)  = ~\V2018(0) ,
  \V1278(1)  = ~\V1984(0) ,
  \[109]  = V1294 | V1286,
  V2000 = \V2011(0)  & (\V803(0)  & (\V242(0)  & (\V1446(0)  & \V2004(0) ))),
  V2001 = V1445 & (V643 & (\V272(0)  & (\V803(0)  & (\V242(0)  & (\V134(0)  & \V134(1) ))))),
  V2003 = \V56(0)  & \V2007(0) ,
  V2005 = V1445 & \V803(0) ,
  V2006 = \V642(0)  & (\V271(0)  & \V1761(0) ),
  V2009 = \V2007(0)  & \[65] ,
  V2012 = \V2024(0)  & (\V2008(0)  & (\V2007(0)  & (\V2022(0)  & \V1998(0) ))),
  V2013 = \V1727(0)  & (V726 & (\V803(0)  & (\V1446(0)  & (\V2024(0)  & \V1998(0) )))),
  V2014 = \V134(1)  & (\V134(0)  & (V1445 & (V2006 & \V1727(0) ))),
  V2015 = \V2011(0)  & (\V1446(0)  & \V803(0) ),
  V2016 = ~V2009,
  V2017 = ~V2006,
  V2021 = V1721 & \V803(0) ,
  V2023 = \V248(0)  & \V803(0) ,
  \V885(0)  = ~V881,
  V2025 = V2761 | V2760,
  V2026 = \V1976(0)  & V1842,
  V2027 = V2765 | V2764,
  V2028 = V2769 | V2768,
  V2029 = V2773 | V2772,
  V2030 = V2026 & V1844,
  V2031 = V2026 & \V1975(0) ,
  V2032 = V1844 & \V1975(0) ,
  V2034 = V2777 | V2776,
  V2035 = \V2033(0)  & V1840,
  V2036 = \V2033(0)  & V1972,
  V2037 = V1840 & V1972,
  V2039 = V2781 | V2780,
  \V1481(0)  = \[133] ,
  V2040 = ~V2025,
  V2041 = ~V2029,
  V2042 = ~V2034,
  V2043 = V2785 | V2784,
  V2044 = V2040 & V2041,
  V2045 = V2789 | V2788,
  V2046 = V2044 & V2042,
  V2047 = V2793 | V2792,
  V2048 = ~V2040,
  V2049 = ~V2043,
  V2050 = ~V2045,
  V2051 = V2797 | V2796,
  V2052 = V2048 & V2049,
  V2053 = V2801 | V2800,
  V2054 = V2052 & V2050,
  V2055 = V2805 | V2804,
  \V959(0)  = ~V955,
  V2056 = V2190 & (V1844 & V2039),
  V2057 = \V1858(0)  & (V2191 & V2055),
  V2059 = V2192 & (V1844 & V2034),
  V2060 = \V1858(0)  & (V2193 & V2053),
  V2062 = V2194 & (V1844 & V2029),
  V2063 = \V1858(0)  & (V2195 & V2051),
  V2065 = V2196 & (V1844 & V2025),
  V2066 = \V1858(0)  & (V2197 & V2048),
  V2068 = ~\V2067(0) ,
  V2069 = ~\V2064(0) ,
  \[110]  = V1296 | V1287,
  V2070 = ~\V2061(0) ,
  V2071 = V2809 | V2808,
  V2072 = V2068 & V2069,
  V2073 = V2813 | V2812,
  V2074 = V2072 & V2070,
  V2075 = V2817 | V2816,
  V2076 = V2198 & (V1842 & V2039),
  V2077 = \V1857(0)  & (V2199 & V2075),
  V2079 = V2200 & (V1842 & V2034),
  \V424(0)  = \[52]  | V687,
  \[111]  = \V62(0)  & (V804 & (V1363 & (V1361 & (V793 & (V1362 & (V1364 & (V805 & (V964 & V498)))))))),
  V2080 = \V1857(0)  & (V2201 & V2073),
  V2082 = V2202 & (V1842 & V2029),
  V2083 = \V1857(0)  & (V2203 & V2071),
  V2085 = V2204 & (V1842 & V2025),
  V2086 = \V1857(0)  & (V2205 & V2068),
  V2088 = ~\V1862(0) ,
  V2089 = ~V1852,
  \[112]  = ~\V268(5) ,
  V2090 = ~\V1862(0) ,
  V2091 = ~V1852,
  V2092 = ~\V1862(0) ,
  V2093 = ~V1852,
  V2094 = ~\V1862(0) ,
  V2095 = ~V1852,
  V2096 = ~\V1861(0) ,
  V2097 = ~V1850,
  V2098 = ~\V1861(0) ,
  V2099 = ~V1850,
  \[113]  = V1376 & (V785 & V1377),
  \V1629(0)  = \[147] ,
  \[114]  = V1379 & (V785 & V1377),
  \V762(0)  = V761 | (V700 | V725),
  \V897(0)  = ~V896,
  \[115]  = V1377 & (V785 & V1381),
  \V1493(0)  = ~\V215(0) ,
  \[116]  = V1377 & (V785 & V1383),
  \V362(0)  = ~V349,
  \[117]  = V1377 & (V785 & V1385),
  \[118]  = \V8(0)  & \V9(0) ,
  \[119]  = V1390 | V1391,
  V2100 = ~\V1861(0) ,
  V2101 = ~V1850,
  V2102 = ~\V1861(0) ,
  V2103 = ~V1850,
  V2104 = ~\[65]  | ~V769,
  V2105 = ~\V2019(0) ,
  V2106 = ~\[65]  | ~V769,
  V2107 = ~\[65]  | ~V727,
  V2108 = ~\V2019(0) ,
  V2109 = ~\[65]  | ~V727,
  \V436(0)  = ~\V37(0) ,
  V2110 = ~\V2011(0) ,
  V2111 = ~\V1395(0) ,
  V2112 = ~\V2011(0) ,
  V2113 = ~\V1395(0) ,
  V2114 = ~\V1421(0) ,
  V2115 = ~\V987(0)  | (~\V1446(0)  | ~V727),
  V2116 = ~\V987(0)  | (~\V1446(0)  | ~V727),
  V2117 = ~\V1681(0) ,
  V2118 = ~\V1421(0) ,
  V2119 = ~\V987(0)  | (~\V1446(0)  | ~V727),
  V2120 = ~\V1421(0) ,
  V2121 = ~\V1681(0) ,
  V2122 = ~\V987(0)  | (~\V1446(0)  | ~V727),
  V2123 = ~\V1681(0) ,
  V2124 = ~\V1408(0) ,
  V2125 = ~V1402,
  V2126 = ~V1125,
  V2127 = ~\V1126(1) ,
  V2128 = ~V1125,
  V2129 = ~\V1126(1) ,
  V2130 = ~\V1417(0) ,
  V2131 = ~\V1422(0) ,
  V2132 = ~\V1417(0) ,
  V2133 = ~\V1422(0) ,
  V2134 = ~\V1417(0) ,
  V2135 = ~\V1422(0) ,
  V2136 = ~\V1984(0) ,
  V2137 = ~\V1278(1) ,
  V2138 = ~V1979,
  V2139 = ~\V1282(1) ,
  V2140 = ~\V1860(0) ,
  V2141 = ~V1848,
  V2142 = ~\V1860(0) ,
  V2143 = ~V1848,
  V2144 = ~\V1860(0) ,
  V2145 = ~V1848,
  V2146 = ~\V1860(0) ,
  V2147 = ~V1848,
  V2148 = ~\V1859(0) ,
  V2149 = ~V1846,
  V2150 = ~\V1859(0) ,
  V2151 = ~V1846,
  V2152 = ~\V1859(0) ,
  V2153 = ~V1846,
  V2154 = ~\V1859(0) ,
  V2155 = ~V1846,
  V2156 = ~V379,
  V2157 = ~\V803(0)  | ~V721,
  V2158 = ~\V1983(0) ,
  V2159 = ~\V1690(1) ,
  V2160 = ~V1978,
  V2161 = ~\V1694(1) ,
  V2162 = ~\V1761(0) ,
  V2163 = ~V745,
  V2164 = ~V745,
  V2165 = ~\V1761(0) ,
  V2166 = ~\V436(0) ,
  V2167 = ~\V37(0) ,
  V2168 = ~V750,
  V2169 = ~V742,
  \V374(0)  = ~V372,
  \[120]  = \V9(0)  & \V1(0) ,
  V2170 = ~V735,
  V2171 = ~V750,
  V2172 = ~V742,
  V2173 = ~V736,
  V2174 = ~V750,
  V2175 = ~V735,
  V2176 = ~V736,
  V2177 = ~V742,
  V2178 = ~V735,
  V2179 = ~V736,
  \[121]  = V1377 & V1424,
  V2180 = ~V751,
  V2181 = ~V743,
  V2182 = ~V751,
  V2183 = ~V742,
  V2184 = ~V743,
  V2185 = ~V742,
  V2186 = ~\V382(0) ,
  V2187 = ~V743,
  V2188 = ~V2017 | ~V2016,
  V2189 = ~\V2010(0)  | ~V2006,
  \V1444(0)  = ~V1443,
  \[122]  = \V1(0)  & \V11(0) ,
  V2190 = ~\V1858(0) ,
  V2191 = ~V1844,
  V2192 = ~\V1858(0) ,
  V2193 = ~V1844,
  V2194 = ~\V1858(0) ,
  V2195 = ~V1844,
  V2196 = ~\V1858(0) ,
  V2197 = ~V1844,
  V2198 = ~\V1857(0) ,
  V2199 = ~V1842,
  \[123]  = \V1(0)  & \V12(0) ,
  \[124]  = V1430 & (V1424 & V786),
  \[125]  = V498 & (V964 & \V66(0) ),
  \[126]  = V1435 | V746,
  \[127]  = ~V1438,
  \[128]  = V1448 | V1450,
  \V1856(0)  = \V288(6)  | \V288(7) ,
  \V386(0)  = \V367(0)  | \V368(0) ,
  \[129]  = V1456 | V1458,
  V2200 = ~\V1857(0) ,
  V2201 = ~V1842,
  V2202 = ~\V1857(0) ,
  V2203 = ~V1842,
  V2204 = ~\V1857(0) ,
  V2205 = ~V1842,
  V2206 = ~V451,
  V2207 = ~\V32(0) ,
  V2208 = V2207 & V451,
  V2209 = \V32(0)  & V2206,
  V2210 = ~V446,
  V2211 = ~\V32(1) ,
  V2212 = V2211 & V446,
  V2213 = \V32(1)  & V2210,
  V2214 = ~V441,
  V2215 = ~\V32(2) ,
  V2216 = V2215 & V441,
  V2217 = \V32(2)  & V2214,
  V2218 = ~V1850,
  V2219 = ~V1298,
  V2220 = V2219 & V1850,
  V2221 = V1298 & V2218,
  V2222 = ~V1852,
  V2223 = ~V1302,
  V2224 = V2223 & V1852,
  V2225 = V1302 & V2222,
  V2226 = ~V1838,
  V2227 = ~V1307,
  V2228 = V2227 & V1838,
  V2229 = V1307 & V2226,
  V2230 = ~V439,
  V2231 = ~V438,
  V2232 = V2231 & V439,
  V2233 = V438 & V2230,
  V2234 = ~\V445(0) ,
  V2235 = ~V440,
  V2236 = V2235 & \V445(0) ,
  V2237 = V440 & V2234,
  V2238 = ~V1312,
  V2239 = ~\V450(0) ,
  V2240 = V2239 & V1312,
  V2241 = \V450(0)  & V2238,
  V2242 = ~V441,
  V2243 = ~V333,
  V2244 = V2243 & V441,
  V2245 = V333 & V2242,
  V2246 = ~V446,
  V2247 = ~V453,
  V2248 = V2247 & V446,
  V2249 = V453 & V2246,
  V2250 = ~V451,
  V2251 = ~V455,
  V2252 = V2251 & V451,
  V2253 = V455 & V2250,
  V2254 = ~V452,
  V2255 = ~V457,
  V2256 = V2255 & V452,
  V2257 = V457 & V2254,
  V2258 = ~V454,
  V2259 = ~V461,
  \V2007(0)  = V769 | V727,
  \V798(0)  = \[63] ,
  V2260 = V2259 & V454,
  V2261 = V461 & V2258,
  V2262 = ~V456,
  V2263 = ~V463,
  V2264 = V2263 & V456,
  V2265 = V463 & V2262,
  V2266 = ~\V473(0) ,
  V2267 = ~V477,
  V2268 = V2267 & \V473(0) ,
  V2269 = V477 & V2266,
  \[130]  = V1464 | V1466,
  V2270 = ~\V470(0) ,
  V2271 = ~V481,
  V2272 = V2271 & \V470(0) ,
  V2273 = V481 & V2270,
  V2274 = ~\V467(0) ,
  V2275 = ~V483,
  V2276 = V2275 & \V467(0) ,
  V2277 = V483 & V2274,
  V2278 = ~\V39(0) ,
  \V1394(0)  = \V60(0)  | (\V56(0)  | \V59(0) ),
  V2279 = ~\V38(0) ,
  \[131]  = \V67(0)  & (V964 & (V498 & V1469)),
  V2280 = V2279 & \V39(0) ,
  V2281 = \V38(0)  & V2278,
  V2282 = ~\V42(0) ,
  V2283 = ~\V44(0) ,
  V2284 = V2283 & \V42(0) ,
  V2285 = \V44(0)  & V2282,
  V2286 = ~\V41(0) ,
  V2287 = ~\V45(0) ,
  \V398(0)  = \[7] ,
  V2288 = V2287 & \V41(0) ,
  V2289 = \V45(0)  & V2286,
  \[132]  = V1478 | (V1476 | V1479),
  V2290 = ~\V257(0) ,
  V2291 = ~V644,
  V2292 = V2291 & \V257(0) ,
  V2293 = V644 & V2290,
  V2294 = ~\V257(1) ,
  V2295 = ~V645,
  V2296 = V2295 & \V257(1) ,
  V2297 = V645 & V2294,
  V2298 = ~\V257(2) ,
  V2299 = ~V646,
  \[133]  = ~\V214(0) ,
  \V1468(0)  = ~\V260(0) ,
  \[134]  = V1490 | V1494,
  \[135]  = ~\V175(0) ,
  \[136]  = V1507 | V1503,
  \V1671(0)  = \[151] ,
  \[137]  = V1509 | V1504,
  \V2019(0)  = V2014 | V2015,
  \[138]  = V1511 | V1505,
  \[139]  = ~V1535,
  V2300 = V2299 & \V257(2) ,
  V2301 = V646 & V2298,
  V2302 = ~\V257(3) ,
  V2303 = ~V647,
  V2304 = V2303 & \V257(3) ,
  V2305 = V647 & V2302,
  V2306 = ~\V257(4) ,
  V2307 = ~V648,
  V2308 = V2307 & \V257(4) ,
  V2309 = V648 & V2306,
  \V1745(0)  = \[164] ,
  V2310 = ~\V257(5) ,
  V2311 = ~V649,
  V2312 = V2311 & \V257(5) ,
  V2313 = V649 & V2310,
  V2314 = ~\V257(6) ,
  V2315 = ~\V257(7) ,
  V2316 = V2315 & \V257(6) ,
  V2317 = \V257(7)  & V2314,
  V2318 = ~\V2078(0) ,
  V2319 = ~\V1255(0) ,
  V2320 = V2319 & \V2078(0) ,
  V2321 = \V1255(0)  & V2318,
  V2322 = ~\V2081(0) ,
  V2323 = ~\V1255(1) ,
  V2324 = V2323 & \V2081(0) ,
  V2325 = \V1255(1)  & V2322,
  V2326 = ~\V2084(0) ,
  V2327 = ~\V1255(2) ,
  V2328 = V2327 & \V2084(0) ,
  V2329 = \V1255(2)  & V2326,
  V2330 = ~\V2087(0) ,
  V2331 = ~\V1255(3) ,
  V2332 = V2331 & \V2087(0) ,
  V2333 = \V1255(3)  & V2330,
  V2334 = ~\V2058(0) ,
  V2335 = ~\V1255(0) ,
  V2336 = V2335 & \V2058(0) ,
  V2337 = \V1255(0)  & V2334,
  V2338 = ~\V2061(0) ,
  V2339 = ~\V1255(1) ,
  V2340 = V2339 & \V2061(0) ,
  V2341 = \V1255(1)  & V2338,
  V2342 = ~\V2064(0) ,
  V2343 = ~\V1255(2) ,
  V2344 = V2343 & \V2064(0) ,
  V2345 = \V1255(2)  & V2342,
  V2346 = ~\V2067(0) ,
  V2347 = ~\V1255(3) ,
  V2348 = V2347 & \V2067(0) ,
  V2349 = \V1255(3)  & V2346,
  V2350 = ~V2047,
  V2351 = ~\V1255(0) ,
  V2352 = V2351 & V2047,
  V2353 = \V1255(0)  & V2350,
  V2354 = ~V2045,
  V2355 = ~\V1255(1) ,
  V2356 = V2355 & V2045,
  V2357 = \V1255(1)  & V2354,
  V2358 = ~V2043,
  V2359 = ~\V1255(2) ,
  V2360 = V2359 & V2043,
  V2361 = \V1255(2)  & V2358,
  V2362 = ~V2040,
  V2363 = ~\V1255(3) ,
  V2364 = V2363 & V2040,
  V2365 = \V1255(3)  & V2362,
  V2366 = ~V2039,
  V2367 = ~\V1255(0) ,
  V2368 = V2367 & V2039,
  V2369 = \V1255(0)  & V2366,
  \[140]  = V498 & (V964 & \V68(0) ),
  V2370 = ~V2034,
  V2371 = ~\V1255(1) ,
  V2372 = V2371 & V2034,
  V2373 = \V1255(1)  & V2370,
  V2374 = ~V2029,
  V2375 = ~\V1255(2) ,
  V2376 = V2375 & V2029,
  V2377 = \V1255(2)  & V2374,
  V2378 = ~V2025,
  V2379 = ~\V1255(3) ,
  \[141]  = V498 & (V964 & \V1538(0) ),
  V2380 = V2379 & V2025,
  V2381 = \V1255(3)  & V2378,
  V2382 = ~\V1351(0) ,
  V2383 = ~\V1255(0) ,
  V2384 = V2383 & \V1351(0) ,
  V2385 = \V1255(0)  & V2382,
  V2386 = ~\V1354(0) ,
  V2387 = ~\V1255(1) ,
  V2388 = V2387 & \V1354(0) ,
  V2389 = \V1255(1)  & V2386,
  \[142]  = V1549 | V1547,
  V2390 = ~\V1357(0) ,
  V2391 = ~\V1255(2) ,
  V2392 = V2391 & \V1357(0) ,
  V2393 = \V1255(2)  & V2390,
  V2394 = ~\V1360(0) ,
  V2395 = ~\V1255(3) ,
  V2396 = V2395 & \V1360(0) ,
  V2397 = \V1255(3)  & V2394,
  V2398 = ~\V1331(0) ,
  V2399 = ~\V1255(0) ,
  \V1757(0)  = \[165] ,
  \[143]  = V1551 | V1548,
  \[144]  = ~V1610,
  \[145]  = ~V1611,
  \V1960(1)  = \[207] ,
  \V1357(0)  = V1356 | V1355,
  \[146]  = V1616 | (V1614 | (V1615 | V799)),
  \V1960(0)  = \[208] ,
  \V490(0)  = V489 | V488,
  \[147]  = V1628 | (V1624 | \V622(0) ),
  \[148]  = V1643 | (V1644 | V1638),
  \[149]  = ~V1651,
  V2400 = V2399 & \V1331(0) ,
  V2401 = \V1255(0)  & V2398,
  V2402 = ~\V1334(0) ,
  V2403 = ~\V1255(1) ,
  V2404 = V2403 & \V1334(0) ,
  V2405 = \V1255(1)  & V2402,
  V2406 = ~\V1337(0) ,
  V2407 = ~\V1255(2) ,
  V2408 = V2407 & \V1337(0) ,
  V2409 = \V1255(2)  & V2406,
  \V699(0)  = ~V698,
  \V903(0)  = ~V899,
  V2410 = ~\V1340(0) ,
  V2411 = ~\V1255(3) ,
  V2412 = V2411 & \V1340(0) ,
  V2413 = \V1255(3)  & V2410,
  V2414 = ~V1320,
  V2415 = ~\V1255(0) ,
  V2416 = V2415 & V1320,
  V2417 = \V1255(0)  & V2414,
  V2418 = ~V1318,
  V2419 = ~\V1255(1) ,
  V2420 = V2419 & V1318,
  V2421 = \V1255(1)  & V2418,
  V2422 = ~V1316,
  V2423 = ~\V1255(2) ,
  V2424 = V2423 & V1316,
  V2425 = \V1255(2)  & V2422,
  V2426 = ~V1313,
  V2427 = ~\V1255(3) ,
  V2428 = V2427 & V1313,
  V2429 = \V1255(3)  & V2426,
  V2430 = ~V1312,
  V2431 = ~\V1255(0) ,
  V2432 = V2431 & V1312,
  V2433 = \V1255(0)  & V2430,
  V2434 = ~V1307,
  V2435 = ~\V1255(1) ,
  V2436 = V2435 & V1307,
  \V503(0)  = V727 | (V721 | (V501 | (V769 | V611))),
  V2437 = \V1255(1)  & V2434,
  V2438 = ~V1302,
  V2439 = ~\V1255(2) ,
  V2440 = V2439 & V1302,
  V2441 = \V1255(2)  & V2438,
  V2442 = ~V1298,
  V2443 = ~\V1255(3) ,
  V2444 = V2443 & V1298,
  V2445 = \V1255(3)  & V2442,
  V2446 = ~\V487(0) ,
  V2447 = ~\V1255(0) ,
  V2448 = V2447 & \V487(0) ,
  V2449 = \V1255(0)  & V2446,
  V2450 = ~\V490(0) ,
  V2451 = ~\V1255(1) ,
  V2452 = V2451 & \V490(0) ,
  V2453 = \V1255(1)  & V2450,
  V2454 = ~\V493(0) ,
  V2455 = ~\V1255(2) ,
  V2456 = V2455 & \V493(0) ,
  V2457 = \V1255(2)  & V2454,
  V2458 = ~\V496(0) ,
  V2459 = ~\V1255(3) ,
  V2460 = V2459 & \V496(0) ,
  V2461 = \V1255(3)  & V2458,
  V2462 = ~\V467(0) ,
  V2463 = ~\V1255(0) ,
  V2464 = V2463 & \V467(0) ,
  V2465 = \V1255(0)  & V2462,
  V2466 = ~\V470(0) ,
  V2467 = ~\V1255(1) ,
  V2468 = V2467 & \V470(0) ,
  V2469 = \V1255(1)  & V2466,
  \[150]  = V1667 & (V1665 & (V1666 & V1668)),
  V2470 = ~\V473(0) ,
  V2471 = ~\V1255(2) ,
  V2472 = V2471 & \V473(0) ,
  V2473 = \V1255(2)  & V2470,
  V2474 = ~\V476(0) ,
  V2475 = ~\V1255(3) ,
  V2476 = V2475 & \V476(0) ,
  V2477 = \V1255(3)  & V2474,
  V2478 = ~V456,
  V2479 = ~\V1255(0) ,
  \[151]  = ~\V205(0) ,
  V2480 = V2479 & V456,
  V2481 = \V1255(0)  & V2478,
  V2482 = ~V454,
  V2483 = ~\V1255(1) ,
  V2484 = V2483 & V454,
  V2485 = \V1255(1)  & V2482,
  V2486 = ~V452,
  V2487 = ~\V1255(2) ,
  V2488 = V2487 & V452,
  V2489 = \V1255(2)  & V2486,
  \[152]  = \V1674(0)  | V1678,
  V2490 = ~V333,
  V2491 = ~\V1255(3) ,
  V2492 = V2491 & V333,
  V2493 = \V1255(3)  & V2490,
  V2494 = ~V451,
  V2495 = ~\V1255(0) ,
  V2496 = V2495 & V451,
  V2497 = \V1255(0)  & V2494,
  V2498 = ~V446,
  V2499 = ~\V1255(1) ,
  \V915(0)  = ~V911,
  \[153]  = V1692 | V1691,
  \[154]  = V1700 | V1695,
  \[155]  = V1702 | V1696,
  \[156]  = V1704 | V1697,
  \[157]  = V1706 | V1698,
  \V1984(0)  = V1979 | V1982,
  \[158]  = V1708 | V1699,
  \V853(0)  = ~V849,
  \[159]  = V1712 | V1716,
  V2500 = V2499 & V446,
  V2501 = \V1255(1)  & V2498,
  V2502 = ~V441,
  V2503 = ~\V1255(2) ,
  V2504 = V2503 & V441,
  V2505 = \V1255(2)  & V2502,
  V2506 = ~V437,
  V2507 = ~\V1255(3) ,
  V2508 = V2507 & V437,
  V2509 = \V1255(3)  & V2506,
  V2510 = ~V1846,
  V2511 = ~V2025,
  V2512 = V2511 & V1846,
  V2513 = V2025 & V2510,
  V2514 = ~V1848,
  V2515 = ~V2029,
  V2516 = V2515 & V1848,
  V2517 = V2029 & V2514,
  V2518 = ~V1839,
  V2519 = ~V2034,
  V2520 = V2519 & V1839,
  V2521 = V2034 & V2518,
  V2522 = ~V1300,
  V2523 = ~V1299,
  V2524 = V2523 & V1300,
  V2525 = V1299 & V2522,
  \V588(0)  = ~\V243(0) ,
  V2526 = ~\V1306(0) ,
  V2527 = ~V1301,
  V2528 = V2527 & \V1306(0) ,
  \V2061(0)  = V2060 | V2059,
  V2529 = V1301 & V2526,
  \V927(0)  = ~V926,
  V2530 = ~V2039,
  V2531 = ~\V1311(0) ,
  V2532 = V2531 & V2039,
  V2533 = \V1311(0)  & V2530,
  V2534 = ~V1302,
  V2535 = ~V1313,
  V2536 = V2535 & V1302,
  V2537 = V1313 & V2534,
  V2538 = ~V1307,
  V2539 = ~V1317,
  V2540 = V2539 & V1307,
  V2541 = V1317 & V2538,
  V2542 = ~V1312,
  V2543 = ~V1319,
  V2544 = V2543 & V1312,
  V2545 = V1319 & V2542,
  V2546 = ~V1316,
  V2547 = ~V1321,
  V2548 = V2547 & V1316,
  V2549 = V1321 & V2546,
  V2550 = ~V1318,
  V2551 = ~V1325,
  V2552 = V2551 & V1318,
  V2553 = V1325 & V2550,
  V2554 = ~V1320,
  V2555 = ~V1327,
  V2556 = V2555 & V1320,
  V2557 = V1327 & V2554,
  V2558 = ~\V1337(0) ,
  V2559 = ~V1341,
  V2560 = V2559 & \V1337(0) ,
  V2561 = V1341 & V2558,
  V2562 = ~\V1334(0) ,
  V2563 = ~V1345,
  V2564 = V2563 & \V1334(0) ,
  V2565 = V1345 & V2562,
  V2566 = ~\V1331(0) ,
  V2567 = ~V1347,
  V2568 = V2567 & \V1331(0) ,
  V2569 = V1347 & V2566,
  \[160]  = V1525 & (\V240(0)  & V338),
  V2570 = ~\V268(0) ,
  V2571 = ~V1366,
  V2572 = V2571 & \V268(0) ,
  V2573 = V1366 & V2570,
  V2574 = ~\V268(1) ,
  V2575 = ~V1367,
  V2576 = V2575 & \V268(1) ,
  V2577 = V1367 & V2574,
  V2578 = ~\V268(2) ,
  V2579 = ~V1368,
  \V1861(0)  = ~V1850,
  \[161]  = V1723 | V1725,
  V2580 = V2579 & \V268(2) ,
  V2581 = V1368 & V2578,
  \V391(0)  = V389 | (V387 | (V388 | V390)),
  V2582 = ~\V268(3) ,
  V2583 = ~V1369,
  V2584 = V2583 & \V268(3) ,
  V2585 = V1369 & V2582,
  V2586 = ~\V268(4) ,
  V2587 = ~\V268(5) ,
  \V730(0)  = V719 | V720,
  V2588 = V2587 & \V268(4) ,
  V2589 = \V268(5)  & V2586,
  \V865(0)  = ~V861,
  \[162]  = \V1747(0)  & (\V803(0)  & (V1735 & (V698 & V344))),
  V2590 = ~\V78(1) ,
  V2591 = ~\V78(0) ,
  V2592 = V2591 & \V78(1) ,
  V2593 = \V78(0)  & V2590,
  V2594 = ~\V78(3) ,
  V2595 = ~\V78(2) ,
  \V1596(1)  = ~V1594,
  V2596 = V2595 & \V78(3) ,
  V2597 = \V78(2)  & V2594,
  V2598 = ~\V78(5) ,
  V2599 = ~\V78(4) ,
  \[163]  = V1740 | (V1738 | (V1748 | (V1739 | V1733))),
  \V1596(0)  = ~V1593,
  \[164]  = ~V1744,
  \[165]  = V1750 | V1751,
  \[166]  = V1751 | V1752,
  \V1147(7)  = V1142 | V1131,
  \[167]  = V1755 | (V1754 | V1756),
  \V404(0)  = V400 | V728,
  \V1147(6)  = V1144 | V1132,
  \[168]  = ~\V101(0) ,
  \V1147(9)  = V1138 | V1129,
  \[169]  = V1768 | V1764,
  V2600 = V2599 & \V78(5) ,
  V2601 = \V78(4)  & V2598,
  V2602 = ~\V84(1) ,
  V2603 = ~\V84(0) ,
  V2604 = V2603 & \V84(1) ,
  V2605 = \V84(0)  & V2602,
  V2606 = ~\V84(3) ,
  V2607 = ~\V84(2) ,
  V2608 = V2607 & \V84(3) ,
  V2609 = \V84(2)  & V2606,
  \V1147(8)  = V1140 | V1130,
  V2610 = ~\V84(5) ,
  V2611 = ~\V84(4) ,
  V2612 = V2611 & \V84(5) ,
  V2613 = \V84(4)  & V2610,
  V2614 = ~\V88(1) ,
  V2615 = ~\V88(0) ,
  V2616 = V2615 & \V88(1) ,
  V2617 = \V88(0)  & V2614,
  V2618 = ~\V88(3) ,
  \V877(0)  = ~V876,
  V2619 = ~\V88(2) ,
  V2620 = V2619 & \V88(3) ,
  V2621 = \V88(2)  & V2618,
  V2622 = ~V1580,
  V2623 = ~V1579,
  V2624 = V2623 & V1580,
  V2625 = V1579 & V2622,
  V2626 = ~V1582,
  V2627 = ~V1581,
  V2628 = V2627 & V1582,
  V2629 = V1581 & V2626,
  V2630 = ~V1584,
  V2631 = ~V1583,
  V2632 = V2631 & V1584,
  V2633 = V1583 & V2630,
  V2634 = ~V1586,
  V2635 = ~V1585,
  V2636 = V2635 & V1586,
  V2637 = V1585 & V2634,
  V2638 = ~V1588,
  V2639 = ~V1587,
  \V342(0)  = ~V339,
  V2640 = V2639 & V1588,
  V2641 = V1587 & V2638,
  V2642 = ~V1590,
  V322 = ~V451,
  V2643 = ~V1589,
  V323 = \V32(0)  & V322,
  V2644 = V2643 & V1590,
  V324 = V2209 | V2208,
  V2645 = V1589 & V2642,
  V325 = V2213 | V2212,
  V2646 = ~\V94(0) ,
  V326 = V2217 | V2216,
  V2647 = ~V1591,
  V327 = ~V446,
  V2648 = V2647 & \V94(0) ,
  V328 = ~V324,
  V2649 = V1591 & V2646,
  V329 = V327 & (\V32(1)  & V328),
  V2650 = ~\V94(1) ,
  V330 = ~V441,
  V2651 = ~V1592,
  V331 = ~V325,
  V2652 = V2651 & \V94(1) ,
  V332 = V328 & (\V32(2)  & (V330 & V331)),
  V2653 = V1592 & V2650,
  V333 = ~V437,
  V2654 = ~\[197] ,
  V334 = ~V326,
  V2655 = ~\[198] ,
  V335 = V331 & (V333 & (\V32(3)  & (V328 & V334))),
  V2656 = V2655 & \[197] ,
  V2657 = \[198]  & V2654,
  V337 = ~V1476,
  V2658 = ~\[195] ,
  V338 = ~V695,
  V2659 = ~\[196] ,
  V339 = V337 & (V744 & (\V56(0)  & V338)),
  V2660 = V2659 & \[195] ,
  V340 = V721 & \[65] ,
  V2661 = \[196]  & V2658,
  V341 = \[65]  & \V2011(0) ,
  V2662 = ~\[193] ,
  V2663 = ~\[194] ,
  V343 = ~\[65] ,
  V2664 = V2663 & \[193] ,
  V344 = ~\V289(0) ,
  V2665 = \[194]  & V2662,
  V345 = \V759(0)  & \V56(0) ,
  V2666 = ~\[199] ,
  V2667 = ~\[206] ,
  V347 = \V1685(0)  & \V434(0) ,
  V2668 = V2667 & \[199] ,
  V348 = \V947(0)  & (\V937(0)  & \V1685(0) ),
  V2669 = \[206]  & V2666,
  V349 = \V927(0)  & (\V917(0)  & \V1685(0) ),
  \[170]  = V1770 | V1765,
  V2670 = ~\[204] ,
  V350 = \V907(0)  & (\V897(0)  & \V1685(0) ),
  V2671 = ~\[205] ,
  V351 = \V887(0)  & (\V877(0)  & \V1685(0) ),
  V2672 = V2671 & \[204] ,
  V352 = \V867(0)  & (\V857(0)  & \V1685(0) ),
  V2673 = \[205]  & V2670,
  V353 = \V847(0)  & (\V837(0)  & \V1685(0) ),
  V2674 = ~\[202] ,
  V354 = \V959(0)  & (\V958(0)  & \V1685(0) ),
  V2675 = ~\[203] ,
  \V2024(0)  = ~V2023,
  V355 = \V957(0)  & (\V956(0)  & \V1685(0) ),
  V2676 = V2675 & \[202] ,
  V356 = \[1] ,
  V2677 = \[203]  & V2674,
  V357 = \[2] ,
  V2678 = ~\[200] ,
  V358 = \V937(0)  & (\V917(0)  & (\V897(0)  & (\V877(0)  & (\V887(0)  & (\V907(0)  & (\V927(0)  & \V947(0) )))))),
  V2679 = ~\[201] ,
  V359 = \V937(0)  & (\V917(0)  & (\V857(0)  & (\V837(0)  & (\V847(0)  & (\V867(0)  & (\V927(0)  & \V947(0) )))))),
  \[171]  = V1778 | V1774,
  V2680 = V2679 & \[200] ,
  V360 = \V937(0)  & (\V897(0)  & (\V857(0)  & (\V958(0)  & (\V959(0)  & (\V867(0)  & (\V907(0)  & \V947(0) )))))),
  V2681 = \[201]  & V2678,
  V2682 = ~\[207] ,
  V2683 = ~\[208] ,
  V2684 = V2683 & \[207] ,
  V2685 = \[208]  & V2682,
  V2686 = ~V1599,
  V2687 = ~V1598,
  V2688 = V2687 & V1599,
  V2689 = V1598 & V2686,
  \[172]  = V1780 | V1775,
  V2690 = ~V1601,
  V2691 = ~V1600,
  V2692 = V2691 & V1601,
  V372 = \V10(0)  & \V658(0) ,
  V2693 = V1600 & V2690,
  V373 = \[3] ,
  V2694 = ~V1603,
  V2695 = ~V1602,
  V2696 = V2695 & V1603,
  V2697 = V1602 & V2694,
  V377 = \[5] ,
  V2698 = ~V1605,
  V2699 = ~V1604,
  V379 = \V378(0)  & \[65] ,
  \[173]  = V1810 | V1792,
  V387 = V1838 & \V383(0) ,
  V388 = V1839 & \V384(0) ,
  V389 = V1840 & \V385(0) ,
  \[174]  = V1812 | V1793,
  V390 = \V288(7)  & (\V288(6)  & \V386(0) ),
  V392 = \[160]  & (\[82]  & (\[84]  & (\[83]  & (\V391(0)  & \V394(0) )))),
  V395 = \V248(0)  & \[160] ,
  V397 = V1578 & (V1576 & (V1574 & (V1573 & (V1575 & (V1577 & (V430 & (\V396(0)  & (V426 & V431)))))))),
  \V1147(5)  = V1146 | V1133,
  \[175]  = V1814 | V1794,
  \[176]  = V1816 | V1795,
  \[177]  = V1818 | V1796,
  \[178]  = V1820 | V1797,
  \[179]  = V1822 | V1798,
  V2700 = V2699 & V1605,
  V2701 = V1604 & V2698,
  V2702 = ~V1607,
  V2703 = ~V1606,
  V2704 = V2703 & V1607,
  V2705 = V1606 & V2702,
  V2706 = ~V1609,
  V2707 = ~V1608,
  V2708 = V2707 & V1609,
  V2709 = V1608 & V2706,
  V2710 = ~\V194(0) ,
  V2711 = ~V1867,
  V2712 = V2711 & \V194(0) ,
  V2713 = V1867 & V2710,
  V2714 = ~\V194(1) ,
  V2715 = ~V1868,
  V2716 = V2715 & \V194(1) ,
  V2717 = V1868 & V2714,
  V2718 = ~\V194(2) ,
  V2719 = ~V1869,
  V2720 = V2719 & \V194(2) ,
  V400 = \V730(0)  & \V733(0) ,
  V2721 = V1869 & V2718,
  V401 = \V729(0)  & V687,
  V2722 = ~\V194(3) ,
  V402 = V401 & \V62(0) ,
  V2723 = ~V1870,
  V403 = ~\[165] ,
  V2724 = V2723 & \V194(3) ,
  V2725 = V1870 & V2722,
  V2726 = ~\V194(4) ,
  V406 = \V404(0)  & \V56(0) ,
  V2727 = ~V1871,
  \V1897(0)  = \[188] ,
  V407 = \V405(0)  & \V59(0) ,
  V2728 = V2727 & \V194(4) ,
  V2729 = V1871 & V2726,
  V409 = V403 & (V338 & \V408(0) ),
  V2730 = ~\V199(0) ,
  V2731 = ~V1872,
  V411 = V687 & \V729(0) ,
  V2732 = V2731 & \V199(0) ,
  V2733 = V1872 & V2730,
  V2734 = ~\V199(1) ,
  V2735 = ~V1873,
  V415 = \V412(0)  & \[65] ,
  V2736 = V2735 & \V199(1) ,
  V416 = \V413(0)  & \V56(0) ,
  V2737 = V1873 & V2734,
  V417 = \V414(0)  & \V59(0) ,
  V2738 = ~\V199(2) ,
  V418 = ~\V215(0) ,
  V2739 = ~V1874,
  V419 = V418 & (\[52]  & (\V66(0)  & V338)),
  V2740 = V2739 & \V199(2) ,
  V420 = \V1681(0)  & \V70(0) ,
  V2741 = V1874 & V2738,
  V421 = \V2011(0)  & \V1446(0) ,
  V2742 = ~\V199(3) ,
  V422 = V421 & \[65] ,
  V2743 = ~\V199(4) ,
  V2744 = V2743 & \V199(3) ,
  V2745 = \V199(4)  & V2742,
  V425 = \V424(0)  & \[65] ,
  V2746 = ~\V288(7) ,
  V426 = ~V425,
  V2747 = ~\V288(6) ,
  V427 = ~V1643,
  V2748 = V2747 & \V288(7) ,
  V428 = ~V1646,
  V2749 = \V288(6)  & V2746,
  V429 = ~V1491,
  V2750 = ~\V239(4) ,
  V430 = ~\V43(0) ,
  V2751 = ~\V239(3) ,
  V431 = ~\V214(0) ,
  V2752 = V2751 & \V239(4) ,
  V432 = \[10] ,
  V2753 = \V239(3)  & V2750,
  V433 = V749 & \V803(0) ,
  V2754 = ~\V134(1) ,
  V2755 = ~\V134(0) ,
  V2756 = V2755 & \V134(1) ,
  V2757 = \V134(0)  & V2754,
  V437 = V2221 | V2220,
  V2758 = ~V1842,
  V438 = V1298 & V1850,
  V2759 = ~\V1976(0) ,
  V439 = V2225 | V2224,
  \V366(0)  = ~V353,
  V2760 = V2759 & V1842,
  V440 = V2229 | V2228,
  V2761 = \V1976(0)  & V2758,
  V441 = V2233 | V2232,
  V2762 = ~V1844,
  V442 = V438 & V1852,
  V2763 = ~\V1975(0) ,
  V443 = V438 & V1302,
  V2764 = V2763 & V1844,
  V444 = V1852 & V1302,
  V2765 = \V1975(0)  & V2762,
  V2766 = ~V1840,
  V446 = V2237 | V2236,
  V2767 = ~V1972,
  V447 = \V445(0)  & V1838,
  V2768 = V2767 & V1840,
  V448 = \V445(0)  & V1307,
  V2769 = V1972 & V2766,
  V449 = V1838 & V1307,
  \[180]  = V1824 | V1799,
  V2770 = ~V2027,
  V2771 = ~V2026,
  V451 = V2241 | V2240,
  V2772 = V2771 & V2027,
  V452 = V2245 | V2244,
  V2773 = V2026 & V2770,
  V453 = V333 & V330,
  V2774 = ~\V2033(0) ,
  V454 = V2249 | V2248,
  V2775 = ~V2028,
  V455 = V453 & V327,
  V2776 = V2775 & \V2033(0) ,
  V456 = V2253 | V2252,
  V2777 = V2028 & V2774,
  V457 = ~V333,
  V2778 = ~V1972,
  V458 = ~V452,
  V2779 = ~\V2038(0) ,
  V459 = ~V454,
  \[181]  = V1826 | V1800,
  V2780 = V2779 & V1972,
  V460 = V2257 | V2256,
  V2781 = \V2038(0)  & V2778,
  V461 = V457 & V458,
  V2782 = ~V2029,
  V462 = V2261 | V2260,
  V2783 = ~V2040,
  V463 = V461 & V459,
  V2784 = V2783 & V2029,
  V464 = V2265 | V2264,
  V2785 = V2040 & V2782,
  V465 = V2088 & (V1852 & V451),
  V2786 = ~V2034,
  V466 = \V1862(0)  & (V2089 & V464),
  V2787 = ~V2044,
  V2788 = V2787 & V2034,
  V468 = V2090 & (V1852 & V446),
  V2789 = V2044 & V2786,
  V469 = \V1862(0)  & (V2091 & V462),
  \[182]  = V1828 | V1801,
  V2790 = ~V2039,
  V2791 = ~V2046,
  V471 = V2092 & (V1852 & V441),
  V2792 = V2791 & V2039,
  V472 = \V1862(0)  & (V2093 & V460),
  V2793 = V2046 & V2790,
  V2794 = ~V2043,
  V474 = V2094 & (V1852 & V437),
  V2795 = ~V2048,
  V475 = \V1862(0)  & (V2095 & V457),
  V2796 = V2795 & V2043,
  V2797 = V2048 & V2794,
  V477 = ~\V476(0) ,
  V2798 = ~V2045,
  V478 = ~\V473(0) ,
  V2799 = ~V2052,
  V479 = ~\V470(0) ,
  \[183]  = \V1831(0)  & \V14(0) ,
  V480 = V2269 | V2268,
  V481 = V477 & V478,
  V482 = V2273 | V2272,
  V483 = V481 & V479,
  V484 = V2277 | V2276,
  V485 = V2096 & (V1850 & V451),
  V486 = \V1861(0)  & (V2097 & V484),
  V488 = V2098 & (V1850 & V446),
  V489 = \V1861(0)  & (V2099 & V482),
  \[184]  = ~\V261(0) ,
  V491 = V2100 & (V1850 & V441),
  V492 = \V1861(0)  & (V2101 & V480),
  V494 = V2102 & (V1850 & V437),
  V495 = \V1861(0)  & (V2103 & V477),
  V497 = ~\V271(0) ,
  V498 = ~\V1630(0) ,
  V499 = V497 & V498,
  \[185]  = ~\V301(0) ,
  \[186]  = ~\V302(0) ,
  \V1147(10)  = V1136 | V1128,
  \[187]  = V1750 | (V1476 | V1889),
  \V1147(11)  = V1134 | V1127,
  \V378(0)  = V766 | V701,
  \[188]  = V1890 | V1885,
  \[189]  = V1891 | V1886,
  V2800 = V2799 & V2045,
  V2801 = V2052 & V2798,
  V2802 = ~V2047,
  V2803 = ~V2054,
  V2804 = V2803 & V2047,
  V2805 = V2054 & V2802,
  V2806 = ~\V2064(0) ,
  V2807 = ~V2068,
  V2808 = V2807 & \V2064(0) ,
  V2809 = V2068 & V2806,
  V2810 = ~\V2061(0) ,
  V2811 = ~V2072,
  V2812 = V2811 & \V2061(0) ,
  V2813 = V2072 & V2810,
  V2814 = ~\V2058(0) ,
  V2815 = ~V2074,
  V2816 = V2815 & \V2058(0) ,
  V2817 = V2074 & V2814,
  V501 = V710 & \V733(0) ,
  V502 = V710 & V687,
  V505 = \V503(0)  & \V56(0) ,
  V506 = \V504(0)  & \V56(0) ,
  V507 = \V59(0)  & V502,
  V509 = V2281 | V2280,
  V512 = \[15] ,
  V513 = V400 & \V56(0) ,
  V514 = \V56(0)  & V728,
  V515 = \V730(0)  & V687,
  V516 = V515 & \V59(0) ,
  V517 = \V729(0)  & (\V59(0)  & \V733(0) ),
  V518 = \V59(0)  & \V731(0) ,
  V519 = ~V513,
  V520 = ~V514,
  V521 = ~V516,
  V522 = ~V517,
  V523 = ~V518,
  V524 = ~V402,
  V525 = V523 & (V521 & (V519 & (V520 & (V522 & V524)))),
  V526 = ~V525,
  V527 = \[16] ,
  V529 = \V528(0)  & \V45(0) ,
  V530 = V2285 | V2284,
  V531 = V2289 | V2288,
  V534 = \V149(7)  & (V701 & \V56(0) ),
  V535 = V701 & V1646,
  V537 = \[17] ,
  V538 = \[18] ,
  V539 = \[19] ,
  V540 = \[20] ,
  V541 = \[21] ,
  V542 = \[22] ,
  V543 = \[23] ,
  V544 = \[24] ,
  V545 = \[25] ,
  V546 = \[26] ,
  V547 = \[27] ,
  V548 = \[28] ,
  V549 = V2104 & (V2105 & (V727 & (\[65]  & \V149(7) ))),
  \[190]  = V1892 | V1887,
  \V667(3)  = ~\V149(3) ,
  V550 = V2104 & (V2105 & (V727 & (\[65]  & \V149(6) ))),
  V551 = V2104 & (V2105 & (V727 & (\[65]  & \V149(5) ))),
  V552 = V2104 & (V2105 & (V727 & (\[65]  & \V149(4) ))),
  V553 = V2106 & (\V2019(0)  & (V2107 & V1884)),
  V555 = V2106 & (\V2019(0)  & (V2107 & V1883)),
  V557 = V2106 & (\V2019(0)  & (V2107 & V1882)),
  V559 = V2106 & (\V2019(0)  & (V2107 & V1881)),
  \[191]  = V1893 | V1751,
  \V667(2)  = ~\V149(2) ,
  \V729(0)  = V717 | (V715 | (V713 | (V711 | (V712 | (V714 | (V716 | V718)))))),
  V561 = V2106 & (\V2019(0)  & (V2107 & V1880)),
  V563 = V2106 & (\V2019(0)  & (V2107 & V1879)),
  V565 = V2106 & (\V2019(0)  & (V2107 & V1878)),
  V567 = V2106 & (\V2019(0)  & (V2107 & V1877)),
  V569 = V2106 & (\V2019(0)  & (V2107 & V1876)),
  \[192]  = V1895 | V1752,
  \V667(5)  = ~\V149(5) ,
  V571 = V2106 & (\V2019(0)  & (V2107 & V1875)),
  V573 = V2109 & (V2108 & (V769 & (\[65]  & \[82] ))),
  V574 = V2109 & (V2108 & (V769 & (\[65]  & \[83] ))),
  V575 = V2109 & (V2108 & (V769 & (\[65]  & \[84] ))),
  V576 = V2109 & (V2108 & (V769 & (\[65]  & \[85] ))),
  V577 = V2109 & (V2108 & (V769 & (\[65]  & \[86] ))),
  V578 = V2109 & (V2108 & (V769 & (\[65]  & \[87] ))),
  V579 = V2109 & (V2108 & (V769 & (\[65]  & \[88] ))),
  \[193]  = V1922 | (V1910 | V1904),
  \V667(4)  = ~\V149(4) ,
  V580 = V2109 & (V2108 & (V769 & (\[65]  & \[89] ))),
  V581 = V2109 & (V2108 & (V769 & (\[65]  & \[90] ))),
  V582 = V2109 & (V2108 & (V769 & (\[65]  & \[91] ))),
  V586 = ~V341,
  V587 = \[40] ,
  V589 = V586 & (\V243(0)  & \V592(0) ),
  \[194]  = V1928 | (V1923 | (V1912 | V1905)),
  V590 = V586 & (\V588(0)  & \V244(0) ),
  V593 = \V244(0)  & \V243(0) ,
  \V932(0)  = ~V928,
  V594 = V586 & (V593 & \V598(0) ),
  V595 = ~V593,
  V596 = V586 & (V595 & \V245(0) ),
  V599 = \V245(0)  & V593,
  \[195]  = V1929 | (V1924 | (V1914 | V1906)),
  \[196]  = V1930 | (V1925 | (V1916 | V1907)),
  \V667(1)  = ~\V149(1) ,
  \V532(0)  = ~V530,
  \[197]  = V1931 | (V1926 | (V1918 | V1908)),
  \V667(0)  = ~\V149(0) ,
  \[198]  = V1932 | (V1927 | (V1920 | V1909)),
  \V1398(0)  = \V57(0)  | (\V53(0)  | \V56(0) ),
  \[199]  = V2180 & (V2181 & (V742 & \V132(1) )),
  V600 = V586 & (V599 & \V604(0) ),
  V601 = ~V599,
  V602 = V586 & (V601 & \V246(0) ),
  V605 = \V246(0)  & V599,
  V606 = V586 & (V605 & \V610(0) ),
  V607 = ~V605,
  V608 = V586 & (V607 & \V247(0) ),
  \V1337(0)  = V1336 | V1335,
  \V667(7)  = ~\V149(7) ,
  V611 = V739 & V337,
  V613 = \V62(0)  & V741,
  V614 = \[133]  & (V505 & (V338 & V428)),
  V615 = V338 & (\V612(0)  & (\V59(0)  & \[133] )),
  V616 = V338 & (V741 & (\V62(0)  & \[133] )),
  V617 = ~V614,
  V618 = ~V615,
  V619 = ~V616,
  \V470(0)  = V469 | V468,
  \V667(6)  = ~\V149(6) ,
  V620 = \[45] ,
  V621 = \[46] ,
  \V944(0)  = ~V940,
  V623 = \V62(0)  & V745,
  V624 = ~\V302(0) ,
  V625 = ~V623,
  V626 = \[65]  & (\V1647(0)  & V1445),
  V627 = V1737 & (V1445 & \V59(0) ),
  V628 = \V56(0)  & V745,
  V630 = \[47] ,
  V631 = \V269(0)  & (\V639(0)  & \V271(0) ),
  V632 = \V274(0)  & (\V639(0)  & \V641(0) ),
  V635 = ~\V202(0) ,
  V636 = ~\V642(0) ,
  V637 = V497 & (V635 & V636),
  V638 = \V641(0)  & \V639(0) ,
  V643 = ~\V275(0) ,
  V644 = \V257(6)  & (\V257(4)  & (\V257(2)  & (\V257(1)  & (\V257(3)  & (\V257(5)  & \V257(7) ))))),
  V645 = \V257(6)  & (\V257(4)  & (\V257(2)  & (\V257(3)  & (\V257(5)  & \V257(7) )))),
  V646 = \V257(6)  & (\V257(4)  & (\V257(3)  & (\V257(5)  & \V257(7) ))),
  V647 = \V257(6)  & (\V257(4)  & (\V257(5)  & \V257(7) )),
  V648 = \V257(6)  & (\V257(5)  & \V257(7) ),
  V649 = \V257(6)  & \V257(7) ,
  V650 = \[212] ,
  V651 = \[213] ,
  V652 = \[214] ,
  V653 = \[215] ,
  V654 = \[216] ,
  V655 = \[217] ,
  V656 = \[218] ,
  V657 = \[50] ,
  \V1275(0)  = ~\V62(0) ,
  \V882(0)  = ~V878,
  V687 = \V169(1)  & \V1395(0) ,
  V688 = ~V687,
  V695 = \V165(1)  & (\V165(0)  & \V694(2) ),
  V696 = \V165(7)  & (V695 & \V1747(0) ),
  V697 = \V165(2)  & (\V694(0)  & (\V165(1)  & \V203(0) )),
  V698 = V695 & \V694(7) ,
  \V821(0)  = \[66] ,
  \V956(0)  = ~V952,
  \V1552(1)  = \[142] ,
  \V1552(0)  = \[143] ,
  \V1687(0)  = V1686 | \V1674(0) ,
  V700 = \V667(1)  & (\V667(0)  & \V667(2) ),
  V701 = \V667(0)  & (\V149(2)  & \V667(1) ),
  V702 = \V667(0)  & (\V149(1)  & \V667(2) ),
  V703 = \V149(2)  & (\V149(0)  & \V667(1) ),
  V704 = \V149(1)  & (\V149(0)  & \V149(2) ),
  V705 = ~\V149(2) ,
  V706 = \V149(1)  & (\V149(0)  & V705),
  V707 = \[51] ,
  \V894(0)  = ~V890,
  V710 = V766 & \V149(3) ,
  V711 = \V149(4)  & (\[51]  & \V667(5) ),
  V712 = \V149(4)  & (\[51]  & \V149(5) ),
  V713 = \V88(3)  & (\V709(0)  & (\[51]  & (\V667(4)  & \V667(5) ))),
  V714 = \V709(1)  & (\V88(2)  & (\[51]  & (\V667(4)  & \V667(5) ))),
  V715 = \V88(3)  & (\V88(2)  & (\[51]  & (\V667(4)  & \V667(5) ))),
  V716 = \V709(1)  & (\V709(0)  & (\V149(5)  & (V766 & (\V667(3)  & \V667(4) )))),
  V717 = \V88(3)  & (\V709(0)  & (\V149(5)  & (V766 & (\V667(3)  & \V667(4) )))),
  V718 = \V709(1)  & (\V88(2)  & (\V149(5)  & (V766 & (\V667(3)  & \V667(4) )))),
  V719 = \V709(1)  & (\V709(0)  & (\[51]  & (\V667(4)  & \V667(5) ))),
  V720 = \V88(3)  & (\V88(2)  & (\V149(5)  & (V766 & (\V667(3)  & \V667(4) )))),
  V721 = V701 & \V149(3) ,
  V722 = \V667(4)  & (V701 & (\V667(3)  & \V667(5) )),
  V723 = \V667(4)  & (V701 & (\V667(3)  & \V149(5) )),
  V724 = \V149(4)  & (V701 & (\V667(3)  & \V667(5) )),
  V725 = \V667(3)  & (\V149(2)  & (\V149(1)  & (\V667(0)  & \V149(4) ))),
  V726 = \V667(3)  & (\V149(2)  & (\V149(1)  & (\V667(0)  & \V667(4) ))),
  V727 = \V667(0)  & (\V149(1)  & (\V149(2)  & \V149(3) )),
  V728 = \V149(4)  & (V701 & (\V667(3)  & \V149(5) )),
  \V1964(0)  = ~V1961,
  V732 = ~V687,
  V734 = \V733(0)  & \V729(0) ,
  V735 = \V672(6)  & (\V672(4)  & (V702 & (\V672(3)  & (\V672(5)  & \V676(7) )))),
  V736 = \V676(6)  & (\V672(4)  & (V702 & (\V672(3)  & (\V672(5)  & \V672(7) )))),
  V737 = \V676(6)  & (\V672(4)  & (V702 & (\V672(3)  & (\V672(5)  & \V676(7) )))),
  V738 = \V672(6)  & (\V672(4)  & (V702 & (\V672(3)  & (\V676(5)  & \V672(7) )))),
  V739 = \V672(6)  & (\V672(4)  & (V702 & (\V672(3)  & (\V676(5)  & \V676(7) )))),
  \V833(0)  = ~V829,
  V740 = \V676(6)  & (\V672(4)  & (V702 & (\V672(3)  & (\V676(5)  & \V672(7) )))),
  V741 = \V676(6)  & (\V672(4)  & (V702 & (\V672(3)  & (\V676(5)  & \V676(7) )))),
  V742 = \V672(6)  & (\V676(4)  & (V702 & (\V672(3)  & (\V672(5)  & \V672(7) )))),
  V743 = \V681(6)  & (\V686(4)  & (V702 & (\V681(3)  & (\V681(5)  & \V686(7) )))),
  V744 = \V686(6)  & (\V686(4)  & (V702 & (\V681(3)  & (\V681(5)  & \V681(7) )))),
  V745 = \V686(6)  & (\V686(4)  & (V702 & (\V681(3)  & (\V681(5)  & \V686(7) )))),
  V746 = \V681(6)  & (\V686(4)  & (V702 & (\V681(3)  & (\V686(5)  & \V686(7) )))),
  V747 = \V686(6)  & (\V686(4)  & (V702 & (\V681(3)  & (\V686(5)  & \V681(7) )))),
  V748 = \V686(6)  & (\V686(4)  & (V702 & (\V681(3)  & (\V686(5)  & \V686(7) )))),
  V749 = \V681(6)  & (\V681(4)  & (V702 & (\V686(3)  & (\V681(5)  & \V681(7) )))),
  V750 = \V681(6)  & (\V681(4)  & (V702 & (\V686(3)  & (\V681(5)  & \V686(7) )))),
  V751 = \V686(6)  & (\V681(4)  & (V702 & (\V686(3)  & (\V681(5)  & \V681(7) )))),
  V752 = ~V750,
  V753 = ~V751,
  V754 = ~V749,
  V755 = V753 & (\V686(3)  & (V702 & (V752 & V754))),
  V756 = \V681(6)  & (\V681(4)  & (V702 & (\V681(3)  & (\V681(5)  & \V681(7) )))),
  V757 = \V681(6)  & (\V686(5)  & (V702 & (\V686(4)  & (\V681(3)  & \V681(7) )))),
  V760 = ~\V55(0) ,
  V761 = V343 & (\V759(0)  & V760),
  V763 = \[52] ,
  V766 = \V765(0)  & V700,
  V767 = \V765(0)  & V747,
  V768 = \V765(0)  & V748,
  V769 = \V765(0)  & V725,
  \V907(0)  = ~V906,
  V770 = ~\V758(0) ,
  V771 = ~V703,
  V772 = ~V706,
  V773 = ~V704,
  V774 = V772 & (V770 & (V771 & V773)),
  V775 = \[53] ,
  V776 = V345 & \V765(0) ,
  V778 = \[54] ,
  V779 = \[55] ,
  V780 = \[56] ,
  V781 = \[57] ,
  V782 = \[58] ,
  V783 = \[59] ,
  V784 = \[60] ,
  V785 = ~\V584(0) ,
  V786 = ~\V659(0) ,
  V787 = \[61] ,
  V789 = \[62] ,
  V790 = \V758(0)  & \[186] ,
  V791 = ~V790,
  V792 = ~V774,
  V793 = ~\V1681(0) ,
  V794 = V792 & (V791 & V793),
  V795 = ~V794,
  V796 = ~\V817(0) ,
  V797 = V796 & (V795 & V498),
  V799 = \V694(6)  & (\V694(4)  & (\V165(3)  & (\V694(5)  & \V70(0) ))),
  \V1903(4)  = ~\V108(4) ,
  \V1976(0)  = ~V1974,
  \V371(0)  = ~V360,
  \V845(0)  = ~V841,
  \V1441(0)  = ~\V277(0) ,
  \V1053(7)  = V1038 | V1026,
  \V445(0)  = V443 | (V442 | V444),
  \V1791(7)  = ~\[83] ,
  \V1053(6)  = V1040 | V1027,
  V801 = \[64] ,
  V804 = ~V740,
  V805 = ~V739,
  V806 = V804 & V805,
  V808 = V741 & \V65(0) ,
  V809 = ~V806,
  \V1791(6)  = ~\[84] ,
  \V1053(9)  = V1034 | V1024,
  V810 = ~\V1275(0) ,
  V811 = V809 & V810,
  V814 = \V1746(0)  & (\V812(0)  & \V699(0) ),
  V815 = \V813(0)  & V1737,
  V816 = \V290(0)  & V338,
  V818 = V340 & \V149(5) ,
  V819 = ~V340,
  \V1053(8)  = V1036 | V1025,
  V820 = V819 & \V822(0) ,
  V823 = V340 & \V149(4) ,
  V824 = V820 & \V827(0) ,
  V825 = \V279(0)  & (V819 & \V280(0) ),
  V828 = V2321 | V2320,
  V829 = V2325 | V2324,
  \V1791(8)  = ~\[82] ,
  V830 = V2329 | V2328,
  V831 = V2333 | V2332,
  V836 = \V1855(0)  & (\V834(0)  & (\V832(0)  & (\V833(0)  & (\V835(0)  & \V434(0) )))),
  V838 = V2337 | V2336,
  V839 = V2341 | V2340,
  V840 = V2345 | V2344,
  V841 = V2349 | V2348,
  V846 = \V288(4)  & (\V844(0)  & (\V842(0)  & (\V843(0)  & (\V845(0)  & \V434(0) )))),
  V848 = V2353 | V2352,
  V849 = V2357 | V2356,
  \V1853(0)  = \V288(0)  | \V288(1) ,
  V850 = V2361 | V2360,
  V851 = V2365 | V2364,
  \V383(0)  = \V361(0)  | \V362(0) ,
  V856 = V1840 & (\V854(0)  & (\V852(0)  & (\V853(0)  & (\V855(0)  & \V434(0) )))),
  V858 = V2369 | V2368,
  V859 = V2373 | V2372,
  \V857(0)  = ~V856,
  V860 = V2377 | V2376,
  V861 = V2381 | V2380,
  V866 = V1840 & (\V864(0)  & (\V862(0)  & (\V863(0)  & (\V865(0)  & \V434(0) )))),
  V868 = V2385 | V2384,
  V869 = V2389 | V2388,
  V870 = V2393 | V2392,
  V871 = V2397 | V2396,
  V876 = \V1854(0)  & (\V874(0)  & (\V872(0)  & (\V873(0)  & (\V875(0)  & \V434(0) )))),
  V878 = V2401 | V2400,
  V879 = V2405 | V2404,
  V880 = V2409 | V2408,
  V881 = V2413 | V2412,
  V886 = \V288(2)  & (\V884(0)  & (\V882(0)  & (\V883(0)  & (\V885(0)  & \V434(0) )))),
  V888 = V2417 | V2416,
  V889 = V2421 | V2420,
  \V1053(1)  = V1050 | V1032,
  V890 = V2425 | V2424,
  V891 = V2429 | V2428,
  V896 = V1839 & (\V894(0)  & (\V892(0)  & (\V893(0)  & (\V895(0)  & \V434(0) )))),
  V898 = V2433 | V2432,
  V899 = V2437 | V2436,
  \V1791(1)  = ~\[89] ,
  \V1053(0)  = V1052 | V1033,
  \V1791(0)  = ~\[90] ,
  \V1053(3)  = V1046 | V1030,
  \V2004(0)  = ~V2003,
  \V1791(3)  = ~\[87] ,
  \V1053(2)  = V1048 | V1031,
  \V1791(2)  = ~\[88] ,
  \V1053(5)  = V1042 | V1028,
  \V672(3)  = ~\V149(3) ,
  \V1791(5)  = ~\[85] ,
  \V1865(0)  = ~\V15(0) ,
  \V1053(4)  = V1044 | V1029,
  \V1791(4)  = ~\[86] ,
  \V672(5)  = ~\V149(5) ,
  V900 = V2441 | V2440,
  V901 = V2445 | V2444,
  V906 = V1839 & (\V904(0)  & (\V902(0)  & (\V903(0)  & (\V905(0)  & \V434(0) )))),
  \V672(4)  = ~\V149(4) ,
  V908 = V2449 | V2448,
  V909 = V2453 | V2452,
  V910 = V2457 | V2456,
  V911 = V2461 | V2460,
  V916 = \V1853(0)  & (\V914(0)  & (\V912(0)  & (\V913(0)  & (\V915(0)  & \V434(0) )))),
  V918 = V2465 | V2464,
  V919 = V2469 | V2468,
  V920 = V2473 | V2472,
  V921 = V2477 | V2476,
  V926 = \V288(0)  & (\V924(0)  & (\V922(0)  & (\V923(0)  & (\V925(0)  & \V434(0) )))),
  V928 = V2481 | V2480,
  V929 = V2485 | V2484,
  V930 = V2489 | V2488,
  V931 = V2493 | V2492,
  V936 = V1838 & (\V934(0)  & (\V932(0)  & (\V933(0)  & (\V935(0)  & \V434(0) )))),
  V938 = V2497 | V2496,
  V939 = V2501 | V2500,
  V940 = V2505 | V2504,
  V941 = V2509 | V2508,
  \V408(0)  = V407 | (V406 | V402),
  V946 = V1838 & (\V944(0)  & (\V942(0)  & (\V943(0)  & (\V945(0)  & \V434(0) )))),
  V948 = ~\V1255(0) ,
  V949 = ~\V1255(1) ,
  V950 = ~\V1255(2) ,
  V951 = ~\V1255(3) ,
  V952 = \V1856(0)  & (V950 & (V948 & (V949 & (V951 & \V434(0) )))),
  V953 = \V288(6)  & (V950 & (V948 & (V949 & (\V1255(3)  & \V434(0) )))),
  V954 = \V288(7)  & (\V288(6)  & (V951 & (V948 & (V949 & (\V1255(2)  & \V434(0) ))))),
  V955 = \V288(7)  & (\V288(6)  & (\V1255(3)  & (\V1255(2)  & (V948 & (V949 & \V434(0) ))))),
  V960 = V795 & \[65] ,
  V961 = \V777(0)  & (\V759(0)  & (\[52]  & \V56(0) )),
  V962 = \V758(0)  & \V56(0) ,
  V963 = \V759(0)  & V799,
  V964 = ~\V807(0) ,
  V966 = \[68] ,
  V968 = \V258(0)  & (\V1468(0)  & (\V1460(0)  & (\V1681(0)  & \V987(0) ))),
  V969 = ~V968,
  V970 = ~V736,
  V971 = ~V742,
  V972 = ~V743,
  V973 = ~V744,
  V974 = ~V735,
  V975 = ~V746,
  V976 = V974 & (V972 & (V970 & (V969 & (V971 & (V973 & V975))))),
  V977 = ~V961,
  V978 = V977 & (V976 & (V770 & \V56(0) )),
  V979 = ~V976,
  V980 = ~\V967(0) ,
  V981 = V979 & V980,
  V983 = \V982(0)  & \V59(0) ,
  V984 = \V1681(0)  & \V62(0) ,
  V986 = \[69] ,
  V988 = V2110 & (\V1395(0)  & \V229(5) ),
  V989 = V2110 & (\V1395(0)  & \V229(4) ),
  V990 = V2110 & (\V1395(0)  & \V229(3) ),
  V991 = V2110 & (\V1395(0)  & \V229(2) ),
  V992 = V2110 & (\V1395(0)  & \V229(1) ),
  V993 = V2110 & (\V1395(0)  & \V229(0) ),
  V994 = V2110 & (\V1395(0)  & \V223(5) ),
  V995 = V2110 & (\V1395(0)  & \V223(4) ),
  V996 = V2110 & (\V1395(0)  & \V223(3) ),
  V997 = V2110 & (\V1395(0)  & \V223(2) ),
  \V672(7)  = ~\V149(7) ,
  V998 = V2110 & (\V1395(0)  & \V223(1) ),
  V999 = V2110 & (\V1395(0)  & \V223(0) ),
  \V346(0)  = ~V345,
  \V672(6)  = ~\V149(6) ,
  \V1680(0)  = ~\V262(0) ;
endmodule

