// IWLS benchmark module "i6" printed on Wed May 29 17:26:47 2002
module i6(\V138(0) , \V138(2) , \V32(27) , \V32(26) , \V32(25) , \V32(24) , \V32(23) , \V32(22) , \V32(21) , \V32(20) , \V32(19) , \V32(18) , \V32(17) , \V32(16) , \V32(15) , \V32(14) , \V32(13) , \V32(12) , \V32(11) , \V32(10) , \V32(9) , \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(3) , \V32(2) , \V32(1) , \V32(0) , \V64(27) , \V64(26) , \V64(25) , \V64(24) , \V64(23) , \V64(22) , \V64(21) , \V64(20) , \V64(19) , \V64(18) , \V64(17) , \V64(16) , \V64(15) , \V64(14) , \V64(13) , \V64(12) , \V64(11) , \V64(10) , \V64(9) , \V64(8) , \V64(7) , \V64(6) , \V64(5) , \V64(4) , \V64(3) , \V64(2) , \V64(1) , \V64(0) , \V96(27) , \V138(4) , \V96(26) , \V96(25) , \V96(24) , \V96(23) , \V96(22) , \V96(21) , \V96(20) , \V96(19) , \V96(18) , \V96(17) , \V96(16) , \V96(15) , \V96(14) , \V96(13) , \V96(12) , \V96(11) , \V96(10) , \V96(9) , \V96(8) , \V96(7) , \V96(6) , \V96(5) , \V96(4) , \V96(3) , \V96(2) , \V96(1) , \V96(0) , \V32(31) , \V32(30) , \V32(29) , \V32(28) , \V131(27) , \V131(26) , \V131(25) , \V131(24) , \V131(23) , \V131(22) , \V131(21) , \V131(20) , \V131(19) , \V131(18) , \V131(17) , \V131(16) , \V131(15) , \V131(14) , \V131(13) , \V131(12) , \V131(11) , \V131(10) , \V131(9) , \V131(8) , \V131(7) , \V131(6) , \V131(5) , \V131(4) , \V131(3) , \V131(2) , \V131(1) , \V131(0) , \V64(31) , \V64(30) , \V64(29) , \V64(28) , \V99(0) , \V138(3) , \V98(0) , \V97(0) , \V96(31) , \V96(30) , \V96(29) , \V96(28) , \V134(0) , \V133(1) , \V133(0) , \V131(31) , \V131(30) , \V131(29) , \V131(28) , \V166(27) , \V166(26) , \V166(25) , \V166(24) , \V166(23) , \V166(22) , \V166(21) , \V166(20) , \V166(19) , \V166(18) , \V166(17) , \V166(16) , \V166(15) , \V166(14) , \V166(13) , \V166(12) , \V166(11) , \V166(10) , \V166(9) , \V166(8) , \V166(7) , \V166(6) , \V166(5) , \V166(4) , \V166(3) , \V166(2) , \V166(1) , \V166(0) , \V198(31) , \V198(30) , \V198(29) , \V198(28) , \V198(27) , \V198(26) , \V198(25) , \V198(24) , \V198(23) , \V198(22) , \V198(21) , \V198(20) , \V198(19) , \V198(18) , \V198(17) , \V198(16) , \V198(15) , \V198(14) , \V198(13) , \V198(12) , \V198(11) , \V198(10) , \V198(9) , \V198(8) , \V198(7) , \V198(6) , \V198(5) , \V198(4) , \V198(3) , \V198(2) , \V198(1) , \V198(0) , \V205(6) , \V205(5) , \V205(4) , \V205(3) , \V205(2) , \V205(1) , \V205(0) );
input
  \V32(30) ,
  \V138(3) ,
  \V138(2) ,
  \V138(4) ,
  \V138(0) ,
  \V32(0) ,
  \V32(1) ,
  \V32(2) ,
  \V32(3) ,
  \V32(4) ,
  \V32(5) ,
  \V131(27) ,
  \V32(6) ,
  \V131(26) ,
  \V32(7) ,
  \V131(29) ,
  \V32(8) ,
  \V131(28) ,
  \V32(9) ,
  \V96(0) ,
  \V96(1) ,
  \V131(21) ,
  \V96(2) ,
  \V131(20) ,
  \V96(3) ,
  \V131(23) ,
  \V96(4) ,
  \V96(13) ,
  \V131(22) ,
  \V96(5) ,
  \V96(12) ,
  \V131(25) ,
  \V96(6) ,
  \V97(0) ,
  \V96(15) ,
  \V131(24) ,
  \V96(7) ,
  \V96(14) ,
  \V131(17) ,
  \V96(8) ,
  \V131(16) ,
  \V96(9) ,
  \V131(19) ,
  \V96(11) ,
  \V131(18) ,
  \V96(10) ,
  \V98(0) ,
  \V96(17) ,
  \V96(16) ,
  \V131(11) ,
  \V96(19) ,
  \V131(10) ,
  \V99(0) ,
  \V96(18) ,
  \V131(13) ,
  \V96(23) ,
  \V131(12) ,
  \V96(22) ,
  \V131(15) ,
  \V64(13) ,
  \V96(25) ,
  \V131(14) ,
  \V64(12) ,
  \V96(24) ,
  \V64(15) ,
  \V64(14) ,
  \V96(21) ,
  \V96(20) ,
  \V64(11) ,
  \V64(10) ,
  \V96(27) ,
  \V96(26) ,
  \V64(17) ,
  \V96(29) ,
  \V64(16) ,
  \V96(28) ,
  \V131(3) ,
  \V64(19) ,
  \V131(2) ,
  \V64(18) ,
  \V131(5) ,
  \V64(23) ,
  \V131(4) ,
  \V64(22) ,
  \V32(13) ,
  \V64(25) ,
  \V32(12) ,
  \V64(24) ,
  \V32(15) ,
  \V131(1) ,
  \V32(14) ,
  \V96(31) ,
  \V131(0) ,
  \V96(30) ,
  \V64(21) ,
  \V64(20) ,
  \V32(11) ,
  \V32(10) ,
  \V131(7) ,
  \V131(6) ,
  \V131(9) ,
  \V131(31) ,
  \V64(27) ,
  \V131(8) ,
  \V131(30) ,
  \V64(26) ,
  \V32(17) ,
  \V64(29) ,
  \V32(16) ,
  \V64(28) ,
  \V32(19) ,
  \V32(18) ,
  \V133(1) ,
  \V32(23) ,
  \V133(0) ,
  \V64(0) ,
  \V32(22) ,
  \V64(1) ,
  \V32(25) ,
  \V64(2) ,
  \V32(24) ,
  \V64(3) ,
  \V64(4) ,
  \V64(31) ,
  \V64(5) ,
  \V64(30) ,
  \V32(21) ,
  \V64(6) ,
  \V134(0) ,
  \V32(20) ,
  \V64(7) ,
  \V64(8) ,
  \V64(9) ,
  \V32(27) ,
  \V32(26) ,
  \V32(29) ,
  \V32(28) ,
  \V32(31) ;
output
  \V198(7) ,
  \V198(6) ,
  \V198(9) ,
  \V198(8) ,
  \V166(3) ,
  \V166(2) ,
  \V166(5) ,
  \V166(4) ,
  \V166(1) ,
  \V166(0) ,
  \V166(7) ,
  \V166(6) ,
  \V166(9) ,
  \V198(27) ,
  \V166(8) ,
  \V205(3) ,
  \V198(26) ,
  \V205(2) ,
  \V198(29) ,
  \V205(5) ,
  \V198(28) ,
  \V205(4) ,
  \V205(1) ,
  \V205(0) ,
  \V198(21) ,
  \V198(20) ,
  \V198(23) ,
  \V198(22) ,
  \V205(6) ,
  \V198(25) ,
  \V198(24) ,
  \V198(17) ,
  \V198(16) ,
  \V166(27) ,
  \V198(19) ,
  \V166(26) ,
  \V198(18) ,
  \V198(11) ,
  \V198(10) ,
  \V166(21) ,
  \V198(13) ,
  \V166(20) ,
  \V198(12) ,
  \V166(23) ,
  \V198(15) ,
  \V166(22) ,
  \V198(14) ,
  \V166(25) ,
  \V166(24) ,
  \V166(17) ,
  \V166(16) ,
  \V166(19) ,
  \V166(18) ,
  \V166(11) ,
  \V166(10) ,
  \V166(13) ,
  \V166(12) ,
  \V166(15) ,
  \V166(14) ,
  \V198(3) ,
  \V198(2) ,
  \V198(5) ,
  \V198(4) ,
  \V198(31) ,
  \V198(30) ,
  \V198(1) ,
  \V198(0) ;
wire
  \[60] ,
  \[61] ,
  \[62] ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[66] ,
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[5] ,
  \[6] ,
  \[7] ,
  \[8] ,
  \[9] ,
  V208,
  V209,
  V210,
  V211,
  V212,
  V213,
  V214,
  V215,
  V216,
  V217,
  V218,
  V219,
  V220,
  V221,
  V222,
  V223,
  V224,
  V225,
  V226,
  V227,
  V228,
  V229,
  V230,
  V231,
  V232,
  V233,
  V234,
  V235,
  V236,
  V237,
  V238,
  V239,
  V240,
  V241,
  V242,
  V243,
  V244,
  V245,
  V246,
  V247,
  V248,
  V249,
  V250,
  V251,
  V252,
  V253,
  V254,
  V255,
  V256,
  V257,
  V258,
  V259,
  V260,
  V261,
  V262,
  V263,
  V292,
  V293,
  V294,
  V295,
  V296,
  V297,
  V298,
  V299,
  V300,
  V301,
  V302,
  V303,
  V304,
  V305,
  V306,
  V307,
  V308,
  V309,
  V310,
  V311,
  V312,
  V313,
  V314,
  V315,
  V316,
  V317,
  V318,
  V319,
  V322,
  V323,
  V324,
  V325,
  V326,
  V327,
  V328,
  V329,
  \[10] ,
  V330,
  V331,
  V332,
  V333,
  V334,
  V335,
  V336,
  V337,
  V338,
  V339,
  \[11] ,
  V340,
  V341,
  V342,
  V343,
  V344,
  V345,
  V346,
  V347,
  V348,
  V349,
  \[12] ,
  V350,
  V351,
  V352,
  V353,
  V354,
  V355,
  V356,
  V357,
  V358,
  V359,
  \[13] ,
  V360,
  V361,
  V362,
  V363,
  V364,
  V365,
  V366,
  V367,
  V368,
  V369,
  \[14] ,
  V370,
  V371,
  V372,
  V373,
  V374,
  V375,
  V376,
  V377,
  V378,
  V379,
  \[15] ,
  V380,
  V381,
  V382,
  V383,
  V384,
  V385,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  V418,
  V419,
  V420,
  V421,
  V422,
  V423,
  V424,
  V425,
  V426,
  V427,
  V428,
  V429,
  \[20] ,
  V430,
  V431,
  V432,
  V433,
  V434,
  V435,
  V436,
  V437,
  V438,
  V439,
  \[21] ,
  V440,
  V441,
  V442,
  V443,
  V444,
  V445,
  V446,
  V447,
  V448,
  V449,
  \[22] ,
  V451,
  V454,
  V455,
  V456,
  V457,
  V458,
  V459,
  \[23] ,
  V460,
  V461,
  V462,
  V463,
  V464,
  V465,
  V466,
  V467,
  \[24] ,
  V474,
  V475,
  V476,
  V477,
  V478,
  V479,
  \[25] ,
  V480,
  V482,
  \[26] ,
  \[27] ,
  \[28] ,
  \[29] ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ;
assign
  \[60]  = V474 | (V461 | V454),
  \[61]  = V482 | (V475 | (V462 | V455)),
  \[62]  = V482 | (V476 | (V463 | V456)),
  \V198(7)  = \[52] ,
  \[63]  = V482 | (V477 | (V464 | V457)),
  \V198(6)  = \[53] ,
  \[64]  = V482 | (V478 | (V465 | V458)),
  \V198(9)  = \[50] ,
  \[65]  = V482 | (V479 | (V466 | V459)),
  \V198(8)  = \[51] ,
  \[66]  = V482 | (V480 | (V467 | V460)),
  \[0]  = V292 | (V236 | V208),
  \[1]  = V293 | (V237 | V209),
  \[2]  = V294 | (V238 | V210),
  \[3]  = V295 | (V239 | V211),
  \[4]  = V296 | (V240 | V212),
  \[5]  = V297 | (V241 | V213),
  \[6]  = V298 | (V242 | V214),
  \[7]  = V299 | (V243 | V215),
  \[8]  = V300 | (V244 | V216),
  \[9]  = V301 | (V245 | V217),
  V208 = \V32(27)  & (~\V138(2)  & ~\V138(0) ),
  V209 = \V32(26)  & (~\V138(2)  & ~\V138(0) ),
  V210 = \V32(25)  & (~\V138(2)  & ~\V138(0) ),
  V211 = \V32(24)  & (~\V138(2)  & ~\V138(0) ),
  V212 = \V32(23)  & (~\V138(2)  & ~\V138(0) ),
  V213 = \V32(22)  & (~\V138(2)  & ~\V138(0) ),
  V214 = \V32(21)  & (~\V138(2)  & ~\V138(0) ),
  V215 = \V32(20)  & (~\V138(2)  & ~\V138(0) ),
  V216 = \V32(19)  & (~\V138(2)  & ~\V138(0) ),
  V217 = \V32(18)  & (~\V138(2)  & ~\V138(0) ),
  V218 = \V32(17)  & (~\V138(2)  & ~\V138(0) ),
  V219 = \V32(16)  & (~\V138(2)  & ~\V138(0) ),
  V220 = \V32(15)  & (~\V138(2)  & ~\V138(0) ),
  V221 = \V32(14)  & (~\V138(2)  & ~\V138(0) ),
  V222 = \V32(13)  & (~\V138(2)  & ~\V138(0) ),
  V223 = \V32(12)  & (~\V138(2)  & ~\V138(0) ),
  V224 = \V32(11)  & (~\V138(2)  & ~\V138(0) ),
  V225 = \V32(10)  & (~\V138(2)  & ~\V138(0) ),
  V226 = \V32(9)  & (~\V138(2)  & ~\V138(0) ),
  V227 = \V32(8)  & (~\V138(2)  & ~\V138(0) ),
  V228 = \V32(7)  & (~\V138(2)  & ~\V138(0) ),
  V229 = \V32(6)  & (~\V138(2)  & ~\V138(0) ),
  V230 = \V32(5)  & (~\V138(2)  & ~\V138(0) ),
  V231 = \V32(4)  & (~\V138(2)  & ~\V138(0) ),
  V232 = \V32(3)  & (~\V138(2)  & ~\V138(0) ),
  V233 = \V32(2)  & (~\V138(2)  & ~\V138(0) ),
  V234 = \V32(1)  & (~\V138(2)  & ~\V138(0) ),
  V235 = \V32(0)  & (~\V138(2)  & ~\V138(0) ),
  V236 = \V64(27)  & (~\V138(2)  & \V138(0) ),
  V237 = \V64(26)  & (~\V138(2)  & \V138(0) ),
  V238 = \V64(25)  & (~\V138(2)  & \V138(0) ),
  V239 = \V64(24)  & (~\V138(2)  & \V138(0) ),
  V240 = \V64(23)  & (~\V138(2)  & \V138(0) ),
  V241 = \V64(22)  & (~\V138(2)  & \V138(0) ),
  V242 = \V64(21)  & (~\V138(2)  & \V138(0) ),
  V243 = \V64(20)  & (~\V138(2)  & \V138(0) ),
  V244 = \V64(19)  & (~\V138(2)  & \V138(0) ),
  V245 = \V64(18)  & (~\V138(2)  & \V138(0) ),
  V246 = \V64(17)  & (~\V138(2)  & \V138(0) ),
  V247 = \V64(16)  & (~\V138(2)  & \V138(0) ),
  V248 = \V64(15)  & (~\V138(2)  & \V138(0) ),
  V249 = \V64(14)  & (~\V138(2)  & \V138(0) ),
  V250 = \V64(13)  & (~\V138(2)  & \V138(0) ),
  V251 = \V64(12)  & (~\V138(2)  & \V138(0) ),
  V252 = \V64(11)  & (~\V138(2)  & \V138(0) ),
  V253 = \V64(10)  & (~\V138(2)  & \V138(0) ),
  V254 = \V64(9)  & (~\V138(2)  & \V138(0) ),
  V255 = \V64(8)  & (~\V138(2)  & \V138(0) ),
  V256 = \V64(7)  & (~\V138(2)  & \V138(0) ),
  V257 = \V64(6)  & (~\V138(2)  & \V138(0) ),
  V258 = \V64(5)  & (~\V138(2)  & \V138(0) ),
  V259 = \V64(4)  & (~\V138(2)  & \V138(0) ),
  V260 = \V64(3)  & (~\V138(2)  & \V138(0) ),
  V261 = \V64(2)  & (~\V138(2)  & \V138(0) ),
  V262 = \V64(1)  & (~\V138(2)  & \V138(0) ),
  V263 = \V64(0)  & (~\V138(2)  & \V138(0) ),
  V292 = ~\V64(27)  & (\V138(2)  & \V138(0) ),
  V293 = ~\V64(26)  & (\V138(2)  & \V138(0) ),
  V294 = ~\V64(25)  & (\V138(2)  & \V138(0) ),
  V295 = ~\V64(24)  & (\V138(2)  & \V138(0) ),
  V296 = ~\V64(23)  & (\V138(2)  & \V138(0) ),
  V297 = ~\V64(22)  & (\V138(2)  & \V138(0) ),
  V298 = ~\V64(21)  & (\V138(2)  & \V138(0) ),
  V299 = ~\V64(20)  & (\V138(2)  & \V138(0) ),
  V300 = ~\V64(19)  & (\V138(2)  & \V138(0) ),
  V301 = ~\V64(18)  & (\V138(2)  & \V138(0) ),
  V302 = ~\V64(17)  & (\V138(2)  & \V138(0) ),
  V303 = ~\V64(16)  & (\V138(2)  & \V138(0) ),
  V304 = ~\V64(15)  & (\V138(2)  & \V138(0) ),
  V305 = ~\V64(14)  & (\V138(2)  & \V138(0) ),
  V306 = ~\V64(13)  & (\V138(2)  & \V138(0) ),
  V307 = ~\V64(12)  & (\V138(2)  & \V138(0) ),
  V308 = ~\V64(11)  & (\V138(2)  & \V138(0) ),
  V309 = ~\V64(10)  & (\V138(2)  & \V138(0) ),
  V310 = ~\V64(9)  & (\V138(2)  & \V138(0) ),
  V311 = ~\V64(8)  & (\V138(2)  & \V138(0) ),
  V312 = ~\V64(7)  & (\V138(2)  & \V138(0) ),
  V313 = ~\V64(6)  & (\V138(2)  & \V138(0) ),
  V314 = ~\V64(5)  & (\V138(2)  & \V138(0) ),
  V315 = ~\V64(4)  & (\V138(2)  & \V138(0) ),
  V316 = ~\V64(3)  & (\V138(2)  & \V138(0) ),
  V317 = ~\V64(2)  & (\V138(2)  & \V138(0) ),
  V318 = ~\V64(1)  & (\V138(2)  & \V138(0) ),
  V319 = ~\V64(0)  & (\V138(2)  & \V138(0) ),
  V322 = \V138(4)  & (\V96(27)  & (~\V138(2)  & ~\V138(0) )),
  V323 = \V96(26)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V324 = \V96(25)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V325 = \V96(24)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V326 = \V96(23)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V327 = \V96(22)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V328 = \V96(21)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V329 = \V96(20)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  \[10]  = V302 | (V246 | V218),
  V330 = \V96(19)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V331 = \V96(18)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V332 = \V96(17)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V333 = \V96(16)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V334 = \V96(15)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V335 = \V96(14)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V336 = \V96(13)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V337 = \V96(12)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V338 = \V96(11)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V339 = \V96(10)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  \[11]  = V303 | (V247 | V219),
  \V166(3)  = \[24] ,
  V340 = \V96(9)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V341 = \V96(8)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V342 = \V96(7)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V343 = \V96(6)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V344 = \V96(5)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V345 = \V96(4)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V346 = \V96(3)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V347 = \V96(2)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V348 = \V96(1)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V349 = \V96(0)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  \[12]  = V304 | (V248 | V220),
  \V166(2)  = \[25] ,
  V350 = \V32(31)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V351 = \V32(30)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V352 = \V32(29)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V353 = \V32(28)  & (\V138(4)  & (~\V138(2)  & ~\V138(0) )),
  V354 = \V131(27)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V355 = \V131(26)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V356 = \V131(25)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V357 = \V131(24)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V358 = \V131(23)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V359 = \V131(22)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  \[13]  = V305 | (V249 | V221),
  \V166(5)  = \[22] ,
  V360 = \V131(21)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V361 = \V131(20)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V362 = \V131(19)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V363 = \V131(18)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V364 = \V131(17)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V365 = \V131(16)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V366 = \V131(15)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V367 = \V131(14)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V368 = \V131(13)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V369 = \V131(12)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  \[14]  = V306 | (V250 | V222),
  \V166(4)  = \[23] ,
  V370 = \V131(11)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V371 = \V131(10)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V372 = \V131(9)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V373 = \V131(8)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V374 = \V131(7)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V375 = \V131(6)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V376 = \V131(5)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V377 = \V131(4)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V378 = \V131(3)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V379 = \V131(2)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  \[15]  = V307 | (V251 | V223),
  V380 = \V131(1)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V381 = \V131(0)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V382 = \V64(31)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V383 = \V64(30)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V384 = \V64(29)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  V385 = \V64(28)  & (\V138(4)  & (~\V138(2)  & \V138(0) )),
  \[16]  = V308 | (V252 | V224),
  \[17]  = V309 | (V253 | V225),
  \V166(1)  = \[26] ,
  \[18]  = V310 | (V254 | V226),
  \V166(0)  = \[27] ,
  \[19]  = V311 | (V255 | V227),
  \V166(7)  = \[20] ,
  \V166(6)  = \[21] ,
  V418 = ~\V131(27)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V419 = ~\V131(26)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  \V166(9)  = \[18] ,
  V420 = ~\V131(25)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V421 = ~\V131(24)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V422 = ~\V131(23)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V423 = ~\V131(22)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V424 = ~\V131(21)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  \V198(27)  = \[32] ,
  V425 = ~\V131(20)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V426 = ~\V131(19)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V427 = ~\V131(18)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V428 = ~\V131(17)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V429 = ~\V131(16)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  \[20]  = V312 | (V256 | V228),
  \V166(8)  = \[19] ,
  \V205(3)  = \[63] ,
  V430 = ~\V131(15)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V431 = ~\V131(14)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V432 = ~\V131(13)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V433 = ~\V131(12)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V434 = ~\V131(11)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  \V198(26)  = \[33] ,
  V435 = ~\V131(10)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V436 = ~\V131(9)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V437 = ~\V131(8)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V438 = ~\V131(7)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V439 = ~\V131(6)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  \[21]  = V313 | (V257 | V229),
  \V205(2)  = \[64] ,
  V440 = ~\V131(5)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V441 = ~\V131(4)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V442 = ~\V131(3)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V443 = ~\V131(2)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V444 = ~\V131(1)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  \V198(29)  = \[30] ,
  V445 = ~\V131(0)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V446 = ~\V64(31)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V447 = ~\V64(30)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V448 = ~\V64(29)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  V449 = ~\V64(28)  & (\V138(4)  & (\V138(2)  & \V138(0) )),
  \[22]  = V314 | (V258 | V230),
  \V205(5)  = \[61] ,
  V451 = ~\V138(4)  & \V138(2) ,
  V454 = \V138(3)  & (\V99(0)  & (~\V138(2)  & ~\V138(0) )),
  \V198(28)  = \[31] ,
  V455 = \V98(0)  & (\V138(3)  & (~\V138(2)  & ~\V138(0) )),
  V456 = \V97(0)  & (\V138(3)  & (~\V138(2)  & ~\V138(0) )),
  V457 = \V96(31)  & (\V138(3)  & (~\V138(2)  & ~\V138(0) )),
  V458 = \V96(30)  & (\V138(3)  & (~\V138(2)  & ~\V138(0) )),
  V459 = \V96(29)  & (\V138(3)  & (~\V138(2)  & ~\V138(0) )),
  \[23]  = V315 | (V259 | V231),
  \V205(4)  = \[62] ,
  V460 = \V96(28)  & (\V138(3)  & (~\V138(2)  & ~\V138(0) )),
  V461 = \V134(0)  & (\V138(3)  & (~\V138(2)  & \V138(0) )),
  V462 = \V133(1)  & (\V138(3)  & (~\V138(2)  & \V138(0) )),
  V463 = \V133(0)  & (\V138(3)  & (~\V138(2)  & \V138(0) )),
  V464 = \V131(31)  & (\V138(3)  & (~\V138(2)  & \V138(0) )),
  V465 = \V131(30)  & (\V138(3)  & (~\V138(2)  & \V138(0) )),
  V466 = \V131(29)  & (\V138(3)  & (~\V138(2)  & \V138(0) )),
  V467 = \V131(28)  & (\V138(3)  & (~\V138(2)  & \V138(0) )),
  \[24]  = V316 | (V260 | V232),
  V474 = \V138(3)  & (\V138(2)  & (\V138(0)  & \V134(0) )),
  V475 = ~\V133(1)  & (\V138(3)  & (\V138(2)  & \V138(0) )),
  V476 = ~\V133(0)  & (\V138(3)  & (\V138(2)  & \V138(0) )),
  V477 = ~\V131(31)  & (\V138(3)  & (\V138(2)  & \V138(0) )),
  V478 = ~\V131(30)  & (\V138(3)  & (\V138(2)  & \V138(0) )),
  V479 = ~\V131(29)  & (\V138(3)  & (\V138(2)  & \V138(0) )),
  \[25]  = V317 | (V261 | V233),
  V480 = ~\V131(28)  & (\V138(3)  & (\V138(2)  & \V138(0) )),
  V482 = ~\V138(3)  & \V138(2) ,
  \[26]  = V318 | (V262 | V234),
  \V205(1)  = \[65] ,
  \[27]  = V319 | (V263 | V235),
  \V205(0)  = \[66] ,
  \[28]  = V451 | (V418 | (V354 | V322)),
  \[29]  = V451 | (V419 | (V355 | V323)),
  \V198(21)  = \[38] ,
  \V198(20)  = \[39] ,
  \V198(23)  = \[36] ,
  \V198(22)  = \[37] ,
  \V205(6)  = \[60] ,
  \V198(25)  = \[34] ,
  \V198(24)  = \[35] ,
  \V198(17)  = \[42] ,
  \[30]  = V451 | (V420 | (V356 | V324)),
  \V198(16)  = \[43] ,
  \V166(27)  = \[0] ,
  \[31]  = V451 | (V421 | (V357 | V325)),
  \V198(19)  = \[40] ,
  \V166(26)  = \[1] ,
  \[32]  = V451 | (V422 | (V358 | V326)),
  \V198(18)  = \[41] ,
  \[33]  = V451 | (V423 | (V359 | V327)),
  \[34]  = V451 | (V424 | (V360 | V328)),
  \[35]  = V451 | (V425 | (V361 | V329)),
  \[36]  = V451 | (V426 | (V362 | V330)),
  \[37]  = V451 | (V427 | (V363 | V331)),
  \[38]  = V451 | (V428 | (V364 | V332)),
  \[39]  = V451 | (V429 | (V365 | V333)),
  \V198(11)  = \[48] ,
  \V198(10)  = \[49] ,
  \V166(21)  = \[6] ,
  \V198(13)  = \[46] ,
  \V166(20)  = \[7] ,
  \V198(12)  = \[47] ,
  \V166(23)  = \[4] ,
  \V198(15)  = \[44] ,
  \V166(22)  = \[5] ,
  \V198(14)  = \[45] ,
  \V166(25)  = \[2] ,
  \V166(24)  = \[3] ,
  \[40]  = V451 | (V430 | (V366 | V334)),
  \V166(17)  = \[10] ,
  \[41]  = V451 | (V431 | (V367 | V335)),
  \V166(16)  = \[11] ,
  \[42]  = V451 | (V432 | (V368 | V336)),
  \V166(19)  = \[8] ,
  \[43]  = V451 | (V433 | (V369 | V337)),
  \V166(18)  = \[9] ,
  \[44]  = V451 | (V434 | (V370 | V338)),
  \[45]  = V451 | (V435 | (V371 | V339)),
  \[46]  = V451 | (V436 | (V372 | V340)),
  \[47]  = V451 | (V437 | (V373 | V341)),
  \[48]  = V451 | (V438 | (V374 | V342)),
  \[49]  = V451 | (V439 | (V375 | V343)),
  \V166(11)  = \[16] ,
  \V166(10)  = \[17] ,
  \V166(13)  = \[14] ,
  \V166(12)  = \[15] ,
  \V166(15)  = \[12] ,
  \V166(14)  = \[13] ,
  \[50]  = V451 | (V440 | (V376 | V344)),
  \[51]  = V451 | (V441 | (V377 | V345)),
  \[52]  = V451 | (V442 | (V378 | V346)),
  \[53]  = V451 | (V443 | (V379 | V347)),
  \[54]  = V451 | (V444 | (V380 | V348)),
  \[55]  = V451 | (V445 | (V381 | V349)),
  \[56]  = V451 | (V446 | (V382 | V350)),
  \V198(3)  = \[56] ,
  \[57]  = V451 | (V447 | (V383 | V351)),
  \V198(2)  = \[57] ,
  \[58]  = V451 | (V448 | (V384 | V352)),
  \V198(5)  = \[54] ,
  \[59]  = V451 | (V449 | (V385 | V353)),
  \V198(4)  = \[55] ,
  \V198(31)  = \[28] ,
  \V198(30)  = \[29] ,
  \V198(1)  = \[58] ,
  \V198(0)  = \[59] ;
endmodule

