// IWLS benchmark module "i5" printed on Wed May 29 17:26:47 2002
module i5(\V4(0) , \V2(1) , \V4(1) , \V2(0) , \V28(1) , \V16(2) , \V28(2) , \V16(3) , \V28(3) , \V28(5) , \V16(6) , \V28(6) , \V16(7) , \V28(7) , \V28(9) , \V16(10) , \V28(10) , \V16(11) , \V28(11) , \V28(13) , \V16(14) , \V28(14) , \V16(15) , \V28(15) , \V16(1) , \V16(5) , \V16(9) , \V16(13) , \V52(1) , \V40(2) , \V52(2) , \V40(3) , \V52(3) , \V52(5) , \V40(6) , \V52(6) , \V40(7) , \V52(7) , \V52(9) , \V40(10) , \V52(10) , \V40(11) , \V52(11) , \V52(13) , \V40(14) , \V52(14) , \V40(15) , \V52(15) , \V40(1) , \V40(5) , \V40(9) , \V40(13) , \V76(1) , \V64(2) , \V76(2) , \V64(3) , \V76(3) , \V76(5) , \V64(6) , \V76(6) , \V64(7) , \V76(7) , \V76(9) , \V64(10) , \V76(10) , \V64(11) , \V76(11) , \V76(13) , \V64(14) , \V76(14) , \V64(15) , \V76(15) , \V64(1) , \V64(5) , \V64(9) , \V64(13) , \V100(1) , \V88(2) , \V100(2) , \V88(3) , \V100(3) , \V100(5) , \V88(6) , \V100(6) , \V88(7) , \V100(7) , \V100(9) , \V88(10) , \V100(10) , \V88(11) , \V100(11) , \V100(13) , \V88(14) , \V100(14) , \V88(15) , \V133(0) , \V100(15) , \V88(1) , \V88(5) , \V88(9) , \V88(13) , \V106(1) , \V103(2) , \V106(2) , \V103(3) , \V106(3) , \V112(1) , \V109(2) , \V112(2) , \V109(3) , \V112(3) , \V118(1) , \V115(2) , \V118(2) , \V115(3) , \V118(3) , \V124(1) , \V121(2) , \V124(2) , \V121(3) , \V124(3) , \V103(1) , \V109(1) , \V115(1) , \V121(1) , \V132(0) , \V128(1) , \V132(1) , \V128(2) , \V132(2) , \V128(3) , \V132(3) , \V128(0) , \V135(0) , \V135(1) , \V151(1) , \V151(2) , \V151(3) , \V151(5) , \V151(6) , \V151(7) , \V151(9) , \V151(10) , \V151(11) , \V151(13) , \V151(14) , \V151(15) , \V167(1) , \V167(2) , \V167(3) , \V167(5) , \V167(6) , \V167(7) , \V167(9) , \V167(10) , \V167(11) , \V167(13) , \V167(14) , \V167(15) , \V183(1) , \V183(2) , \V183(3) , \V183(5) , \V183(6) , \V183(7) , \V183(9) , \V183(10) , \V183(11) , \V183(13) , \V183(14) , \V183(15) , \V199(1) , \V199(2) , \V199(3) , \V199(5) , \V199(6) , \V199(7) , \V199(9) , \V199(10) , \V199(11) , \V199(13) , \V199(14) , \V199(15) , \V151(4) , \V151(8) , \V151(12) , \V167(4) , \V167(8) , \V167(12) , \V183(4) , \V183(8) , \V183(12) , \V199(4) , \V199(8) , \V199(12) , \V151(0) , \V167(0) , \V183(0) , \V199(0) );
input
  \V64(3) ,
  \V28(13) ,
  \V52(11) ,
  \V52(10) ,
  \V64(5) ,
  \V28(15) ,
  \V109(3) ,
  \V64(6) ,
  \V28(14) ,
  \V109(2) ,
  \V132(1) ,
  \V64(7) ,
  \V132(0) ,
  \V64(9) ,
  \V28(11) ,
  \V115(3) ,
  \V28(10) ,
  \V115(2) ,
  \V88(1) ,
  \V109(1) ,
  \V16(1) ,
  \V88(2) ,
  \V121(3) ,
  \V16(2) ,
  \V88(3) ,
  \V121(2) ,
  \V16(3) ,
  \V64(13) ,
  \V115(1) ,
  \V88(5) ,
  \V16(5) ,
  \V88(6) ,
  \V16(6) ,
  \V64(15) ,
  \V88(7) ,
  \V16(7) ,
  \V64(14) ,
  \V121(1) ,
  \V88(9) ,
  \V16(9) ,
  \V100(3) ,
  \V100(2) ,
  \V64(11) ,
  \V100(5) ,
  \V64(10) ,
  \V4(0) ,
  \V100(1) ,
  \V4(1) ,
  \V118(3) ,
  \V118(2) ,
  \V52(1) ,
  \V52(2) ,
  \V124(3) ,
  \V52(3) ,
  \V124(2) ,
  \V128(3) ,
  \V100(7) ,
  \V76(13) ,
  \V128(2) ,
  \V100(6) ,
  \V118(1) ,
  \V52(5) ,
  \V100(9) ,
  \V76(15) ,
  \V52(6) ,
  \V76(14) ,
  \V52(7) ,
  \V100(11) ,
  \V124(1) ,
  \V100(10) ,
  \V52(9) ,
  \V128(1) ,
  \V103(3) ,
  \V100(13) ,
  \V76(11) ,
  \V128(0) ,
  \V103(2) ,
  \V76(10) ,
  \V100(15) ,
  \V76(1) ,
  \V100(14) ,
  \V76(2) ,
  \V76(3) ,
  \V103(1) ,
  \V76(5) ,
  \V76(6) ,
  \V76(7) ,
  \V76(9) ,
  \V40(13) ,
  \V88(13) ,
  \V40(15) ,
  \V28(1) ,
  \V40(14) ,
  \V88(15) ,
  \V28(2) ,
  \V88(14) ,
  \V28(3) ,
  \V16(13) ,
  \V40(11) ,
  \V28(5) ,
  \V40(10) ,
  \V16(15) ,
  \V88(11) ,
  \V106(3) ,
  \V28(6) ,
  \V16(14) ,
  \V88(10) ,
  \V106(2) ,
  \V28(7) ,
  \V40(1) ,
  \V2(0) ,
  \V133(0) ,
  \V28(9) ,
  \V40(2) ,
  \V112(3) ,
  \V16(11) ,
  \V2(1) ,
  \V40(3) ,
  \V112(2) ,
  \V16(10) ,
  \V106(1) ,
  \V40(5) ,
  \V40(6) ,
  \V40(7) ,
  \V112(1) ,
  \V52(13) ,
  \V40(9) ,
  \V52(15) ,
  \V132(3) ,
  \V52(14) ,
  \V64(1) ,
  \V132(2) ,
  \V64(2) ;
output
  \V167(4) ,
  \V167(1) ,
  \V167(0) ,
  \V183(3) ,
  \V183(2) ,
  \V183(5) ,
  \V183(4) ,
  \V167(7) ,
  \V151(11) ,
  \V167(6) ,
  \V151(10) ,
  \V199(11) ,
  \V167(9) ,
  \V183(1) ,
  \V151(13) ,
  \V199(10) ,
  \V167(8) ,
  \V183(0) ,
  \V151(12) ,
  \V199(13) ,
  \V151(15) ,
  \V199(12) ,
  \V151(14) ,
  \V199(15) ,
  \V199(14) ,
  \V183(7) ,
  \V183(6) ,
  \V183(9) ,
  \V183(8) ,
  \V135(1) ,
  \V135(0) ,
  \V151(3) ,
  \V151(2) ,
  \V151(5) ,
  \V151(4) ,
  \V151(1) ,
  \V151(0) ,
  \V151(7) ,
  \V151(6) ,
  \V151(9) ,
  \V151(8) ,
  \V183(11) ,
  \V183(10) ,
  \V183(13) ,
  \V183(12) ,
  \V167(11) ,
  \V199(3) ,
  \V183(15) ,
  \V167(10) ,
  \V199(2) ,
  \V183(14) ,
  \V167(13) ,
  \V199(5) ,
  \V167(12) ,
  \V199(4) ,
  \V167(15) ,
  \V167(14) ,
  \V199(1) ,
  \V199(0) ,
  \V199(7) ,
  \V199(6) ,
  \V199(9) ,
  \V199(8) ,
  \V167(3) ,
  \V167(2) ,
  \V167(5) ;
wire
  \[59] ,
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  \[60] ,
  \[61] ,
  \[62] ,
  \[0] ,
  \[63] ,
  \[1] ,
  \[64] ,
  \[20] ,
  \[2] ,
  \[65] ,
  \[21] ,
  \[3] ,
  \[22] ,
  \[4] ,
  \[23] ,
  \[5] ,
  \[24] ,
  \[6] ,
  \[25] ,
  \[7] ,
  \[26] ,
  \[8] ,
  \[27] ,
  \[9] ,
  \[28] ,
  \[29] ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[10] ,
  \[55] ,
  \[11] ,
  \[56] ,
  \[12] ,
  \[57] ,
  \[13] ,
  \[58] ,
  \[14] ;
assign
  \[59]  = (\[60]  & \V124(1) ) | \V121(1) ,
  \[15]  = (\[16]  & \V52(2) ) | \V40(2) ,
  \V167(4)  = \[53] ,
  \[16]  = (\[53]  & \V52(3) ) | \V40(3) ,
  \[17]  = (\[18]  & \V52(5) ) | \V40(5) ,
  \[18]  = (\[19]  & \V52(6) ) | \V40(6) ,
  \V167(1)  = \[14] ,
  \[19]  = (\[54]  & \V52(7) ) | \V40(7) ,
  \V167(0)  = \[63] ,
  \V183(3)  = \[28] ,
  \V183(2)  = \[27] ,
  \[60]  = (\[61]  & \V124(2) ) | \V121(2) ,
  \V183(5)  = \[29] ,
  \[61]  = (\V124(3)  & \V133(0) ) | \V121(3) ,
  \V183(4)  = \[56] ,
  \[62]  = (\[63]  & \V132(0) ) | \V128(0) ,
  \V167(7)  = \[19] ,
  \[0]  = (\[1]  & \V4(0) ) | \V2(0) ,
  \V151(11)  = \[10] ,
  \[63]  = (\[64]  & \V132(1) ) | \V128(1) ,
  \V167(6)  = \[18] ,
  \[1]  = (\[62]  & \V4(1) ) | \V2(1) ,
  \V151(10)  = \[9] ,
  \V199(11)  = \[46] ,
  \[64]  = (\[65]  & \V132(2) ) | \V128(2) ,
  \[20]  = (\[21]  & \V52(9) ) | \V40(9) ,
  \V167(9)  = \[20] ,
  \[2]  = (\[3]  & \V28(1) ) | \V16(1) ,
  \V183(1)  = \[26] ,
  \V151(13)  = \[11] ,
  \V199(10)  = \[45] ,
  \[65]  = (\V132(3)  & \V133(0) ) | \V128(3) ,
  \[21]  = (\[22]  & \V52(10) ) | \V40(10) ,
  \V167(8)  = \[54] ,
  \[3]  = (\[4]  & \V28(2) ) | \V16(2) ,
  \V183(0)  = \[64] ,
  \V151(12)  = \[52] ,
  \V199(13)  = \[47] ,
  \[22]  = (\[55]  & \V52(11) ) | \V40(11) ,
  \[4]  = (\[50]  & \V28(3) ) | \V16(3) ,
  \V151(15)  = \[13] ,
  \V199(12)  = \[61] ,
  \[23]  = (\[24]  & \V52(13) ) | \V40(13) ,
  \[5]  = (\[6]  & \V28(5) ) | \V16(5) ,
  \V151(14)  = \[12] ,
  \V199(15)  = \[49] ,
  \[24]  = (\[25]  & \V52(14) ) | \V40(14) ,
  \[6]  = (\[7]  & \V28(6) ) | \V16(6) ,
  \V199(14)  = \[48] ,
  \[25]  = (\[64]  & \V52(15) ) | \V40(15) ,
  \[7]  = (\[51]  & \V28(7) ) | \V16(7) ,
  \[26]  = (\[27]  & \V76(1) ) | \V64(1) ,
  \[8]  = (\[9]  & \V28(9) ) | \V16(9) ,
  \V183(7)  = \[31] ,
  \[27]  = (\[28]  & \V76(2) ) | \V64(2) ,
  \[9]  = (\[10]  & \V28(10) ) | \V16(10) ,
  \V183(6)  = \[30] ,
  \[28]  = (\[56]  & \V76(3) ) | \V64(3) ,
  \V183(9)  = \[32] ,
  \[29]  = (\[30]  & \V76(5) ) | \V64(5) ,
  \V183(8)  = \[57] ,
  \V135(1)  = \[1] ,
  \V135(0)  = \[0] ,
  \V151(3)  = \[4] ,
  \V151(2)  = \[3] ,
  \V151(5)  = \[5] ,
  \[30]  = (\[31]  & \V76(6) ) | \V64(6) ,
  \V151(4)  = \[50] ,
  \[31]  = (\[57]  & \V76(7) ) | \V64(7) ,
  \[32]  = (\[33]  & \V76(9) ) | \V64(9) ,
  \[33]  = (\[34]  & \V76(10) ) | \V64(10) ,
  \V151(1)  = \[2] ,
  \[34]  = (\[58]  & \V76(11) ) | \V64(11) ,
  \V151(0)  = \[62] ,
  \[35]  = (\[36]  & \V76(13) ) | \V64(13) ,
  \[36]  = (\[37]  & \V76(14) ) | \V64(14) ,
  \[37]  = (\[65]  & \V76(15) ) | \V64(15) ,
  \[38]  = (\[39]  & \V100(1) ) | \V88(1) ,
  \[39]  = (\[40]  & \V100(2) ) | \V88(2) ,
  \V151(7)  = \[7] ,
  \V151(6)  = \[6] ,
  \V151(9)  = \[8] ,
  \V151(8)  = \[51] ,
  \V183(11)  = \[34] ,
  \[40]  = (\[59]  & \V100(3) ) | \V88(3) ,
  \V183(10)  = \[33] ,
  \[41]  = (\[42]  & \V100(5) ) | \V88(5) ,
  \V183(13)  = \[35] ,
  \[42]  = (\[43]  & \V100(6) ) | \V88(6) ,
  \V183(12)  = \[58] ,
  \V167(11)  = \[22] ,
  \V199(3)  = \[40] ,
  \[43]  = (\[60]  & \V100(7) ) | \V88(7) ,
  \V183(15)  = \[37] ,
  \V167(10)  = \[21] ,
  \V199(2)  = \[39] ,
  \[44]  = (\[45]  & \V100(9) ) | \V88(9) ,
  \V183(14)  = \[36] ,
  \V167(13)  = \[23] ,
  \V199(5)  = \[41] ,
  \[45]  = (\[46]  & \V100(10) ) | \V88(10) ,
  \V167(12)  = \[55] ,
  \V199(4)  = \[59] ,
  \[46]  = (\[61]  & \V100(11) ) | \V88(11) ,
  \V167(15)  = \[25] ,
  \[47]  = (\[48]  & \V100(13) ) | \V88(13) ,
  \V167(14)  = \[24] ,
  \[48]  = (\[49]  & \V100(14) ) | \V88(14) ,
  \V199(1)  = \[38] ,
  \[49]  = (\V100(15)  & \V133(0) ) | \V88(15) ,
  \V199(0)  = \[65] ,
  \V199(7)  = \[43] ,
  \V199(6)  = \[42] ,
  \[50]  = (\[51]  & \V106(1) ) | \V103(1) ,
  \V199(9)  = \[44] ,
  \[51]  = (\[52]  & \V106(2) ) | \V103(2) ,
  \V199(8)  = \[60] ,
  \[52]  = (\[63]  & \V106(3) ) | \V103(3) ,
  \[53]  = (\[54]  & \V112(1) ) | \V109(1) ,
  \[54]  = (\[55]  & \V112(2) ) | \V109(2) ,
  \[10]  = (\[52]  & \V28(11) ) | \V16(11) ,
  \[55]  = (\[64]  & \V112(3) ) | \V109(3) ,
  \[11]  = (\[12]  & \V28(13) ) | \V16(13) ,
  \[56]  = (\[57]  & \V118(1) ) | \V115(1) ,
  \[12]  = (\[13]  & \V28(14) ) | \V16(14) ,
  \V167(3)  = \[16] ,
  \[57]  = (\[58]  & \V118(2) ) | \V115(2) ,
  \[13]  = (\[63]  & \V28(15) ) | \V16(15) ,
  \V167(2)  = \[15] ,
  \[58]  = (\[65]  & \V118(3) ) | \V115(3) ,
  \[14]  = (\[15]  & \V52(1) ) | \V40(1) ,
  \V167(5)  = \[17] ;
endmodule

