// IWLS benchmark module "t481" printed on Wed May 29 17:28:13 2002
module t481(v0, v1, v2, v3, v4, v5, v6, v7, v8, v9, v10, v11, v12, v13, v14, v15, \v16.0 );
input
  v10,
  v11,
  v12,
  v13,
  v14,
  v15,
  v0,
  v1,
  v2,
  v3,
  v4,
  v5,
  v6,
  v7,
  v8,
  v9;
output
  \v16.0 ;
wire
  \[8612] ,
  \[12396] ,
  \[11535] ,
  \[10348] ,
  \[14053] ,
  \[4566] ,
  \[14056] ,
  \[6956] ,
  \[13200] ,
  \[4900] ,
  \[12737] ,
  \[13597] ,
  \[10344] ,
  \[9477] ,
  \[3375] ,
  \[8281] ,
  \[4905] ,
  \[5765] ,
  \[12005] ,
  \[1322] ,
  \[5037] ,
  \[12740] ,
  \[10352] ,
  \[12012] ,
  \[7427] ,
  \[13937] ,
  \[7090] ,
  \[6231] ,
  \[8620] ,
  \[8289] ,
  \[3715] ,
  \[584] ,
  \[4575] ,
  \[11545] ,
  \[6964] ,
  \[13206] ,
  \[1329] ,
  \[14065] ,
  \[9484] ,
  \[4910] ,
  \[11552] ,
  \[7098] ,
  \[6239] ,
  \[12749] ,
  \[14072] ,
  \[14071] ,
  \[5773] ,
  \[3385] ,
  \[2526] ,
  \[8629] ,
  \[21807] ,
  \[12745] ,
  \[21471] ,
  \[926] ,
  \[21809] ,
  \[12020] ,
  \[13948] ,
  \[2193] ,
  \[21803] ,
  \[12752] ,
  \[13219] ,
  \[21805] ,
  \[8299] ,
  \[3725] ,
  \[21477] ,
  \[4585] ,
  \[13216] ,
  \[21479] ,
  \[21811] ,
  \[12028] ,
  \[2531] ,
  \[597] ,
  \[10702] ,
  \[14075] ,
  \[21473] ,
  \[11561] ,
  \[4922] ,
  \[6249] ,
  \[14082] ,
  \[21475] ,
  \[3394] ,
  \[14081] ,
  \[5783] ,
  \[933] ,
  \[8639] ,
  \[204] ,
  \[21817] ,
  \[5055] ,
  \[205] ,
  \[11568] ,
  \[206] ,
  \[3000] ,
  \[21481] ,
  \[21819] ,
  \[4927] ,
  \[12760] ,
  \[207] ,
  \[13958] ,
  \[13227] ,
  \[21813] ,
  \[1344] ,
  \[3733] ,
  \[9107] ,
  \[4593] ,
  \[21815] ,
  \[6982] ,
  \[21487] ,
  \[10378] ,
  \[3008] ,
  \[21489] ,
  \[21821] ,
  \[14085] ,
  \[12037] ,
  \[6257] ,
  \[10711] ,
  \[21483] ,
  \[940] ,
  \[4931] ,
  \[2543] ,
  \[11571] ,
  \[211] ,
  \[5791] ,
  \[8647] ,
  \[12769] ,
  \[212] ,
  \[11904] ,
  \[21485] ,
  \[213] ,
  \[10376] ,
  \[214] ,
  \[21827] ,
  \[9841] ,
  \[215] ,
  \[216] ,
  \[21491] ,
  \[21829] ,
  \[7455] ,
  \[217] ,
  \[9844] ,
  \[13968] ,
  \[218] ,
  \[4209] ,
  \[21823] ,
  \[11579] ,
  \[12041] ,
  \[3743] ,
  \[21825] ,
  \[13969] ,
  \[11576] ,
  \[21497] ,
  \[13963] ,
  \[5405] ,
  \[14093] ,
  \[10387] ,
  \[3018] ,
  \[6995] ,
  \[14096] ,
  \[21499] ,
  \[13235] ,
  \[21831] ,
  \[2551] ,
  \[6267] ,
  \[21493] ,
  \[11581] ,
  \[8657] ,
  \[13972] ,
  \[12779] ,
  \[10383] ,
  \[11914] ,
  \[21495] ,
  \[223] ,
  \[4944] ,
  \[224] ,
  \[954] ,
  \[12776] ,
  \[225] ,
  \[10728] ,
  \[1361] ,
  \[4217] ,
  \[12050] ,
  \[11587] ,
  \[13248] ,
  \[3751] ,
  \[13978] ,
  \[6607] ,
  \[4949] ,
  \[11921] ,
  \[10724] ,
  \[6272] ,
  \[13979] ,
  \[13244] ,
  \[3026] ,
  \[7803] ,
  \[22307] ,
  \[13245] ,
  \[2561] ,
  \[6276] ,
  \[22309] ,
  \[11591] ,
  \[13982] ,
  \[12789] ,
  \[11924] ,
  \[12784] ,
  \[9130] ,
  \[4954] ,
  \[12056] ,
  \[9861] ,
  \[10738] ,
  \[7474] ,
  \[10007] ,
  \[6615] ,
  \[11930] ,
  \[21849] ,
  \[2569] ,
  \[22311] ,
  \[3761] ,
  \[11202] ,
  \[2902] ,
  \[13988] ,
  \[1374] ,
  \[12792] ,
  \[10733] ,
  \[13989] ,
  \[11593] ,
  \[13254] ,
  \[3036] ,
  \[10735] ,
  \[9869] ,
  \[1710] ,
  \[22317] ,
  \[13256] ,
  \[11208] ,
  \[11938] ,
  \[21851] ,
  \[12068] ,
  \[8674] ,
  \[12400] ,
  \[22319] ,
  \[5427] ,
  \[10741] ,
  \[22313] ,
  \[971] ,
  \[13262] ,
  \[6289] ,
  \[13992] ,
  \[22315] ,
  \[5094] ,
  \[7483] ,
  \[12796] ,
  \[12065] ,
  \[1381] ,
  \[11210] ,
  \[6625] ,
  \[4237] ,
  \[10747] ,
  \[9143] ,
  \[3770] ,
  \[2579] ,
  \[12408] ,
  \[22321] ,
  \[11212] ,
  \[13998] ,
  \[10749] ,
  \[21853] ,
  \[12071] ,
  \[12409] ,
  \[3044] ,
  \[21855] ,
  \[13264] ,
  \[1388] ,
  \[6294] ,
  \[7823] ,
  \[22327] ,
  \[11218] ,
  \[2918] ,
  \[1721] ,
  \[11948] ,
  \[3778] ,
  \[22329] ,
  \[10752] ,
  \[13270] ,
  \[12077] ,
  \[8685] ,
  \[10021] ,
  \[4971] ,
  \[12412] ,
  \[6298] ,
  \[22323] ,
  \[12079] ,
  \[22325] ,
  \[6633] ,
  \[21867] ,
  \[2587] ,
  \[7493] ,
  \[10028] ,
  \[10758] ,
  \[985] ,
  \[256] ,
  \[21869] ,
  \[13605] ,
  \[12418] ,
  \[257] ,
  \[22331] ,
  \[13610] ,
  \[258] ,
  \[21863] ,
  \[259] ,
  \[12419] ,
  \[3054] ,
  \[21865] ,
  \[7833] ,
  \[22337] ,
  \[3787] ,
  \[11958] ,
  \[21871] ,
  \[12088] ,
  \[1732] ,
  \[22339] ,
  \[10762] ,
  \[260] ,
  \[12422] ,
  \[261] ,
  \[22333] ,
  \[5449] ,
  \[7108] ,
  \[11224] ,
  \[262] ,
  \[992] ,
  \[263] ,
  \[22335] ,
  \[1737] ,
  \[9161] ,
  \[21877] ,
  \[2597] ,
  \[12085] ,
  \[2931] ,
  \[22341] ,
  \[268] ,
  \[4259] ,
  \[3062] ,
  \[21873] ,
  \[269] ,
  \[10764] ,
  \[999] ,
  \[13622] ,
  \[12429] ,
  \[21875] ,
  \[7841] ,
  \[604] ,
  \[13283] ,
  \[12098] ,
  \[12430] ,
  \[1742] ,
  \[11967] ,
  \[7116] ,
  \[270] ,
  \[3402] ,
  \[13627] ,
  \[13291] ,
  \[4993] ,
  \[8310] ,
  \[12094] ,
  \[11233] ,
  \[6653] ,
  \[11966] ,
  \[21887] ,
  \[10777] ,
  \[21889] ,
  \[8314] ,
  \[3071] ,
  \[10049] ,
  \[11241] ,
  \[279] ,
  \[611] ,
  \[10774] ,
  \[9176] ,
  \[13632] ,
  \[12439] ,
  \[4603] ,
  \[2215] ,
  \[7851] ,
  \[13294] ,
  \[12433] ,
  \[2946] ,
  \[21891] ,
  \[12440] ,
  \[22359] ,
  \[3411] ,
  \[7126] ,
  \[280] ,
  \[1754] ,
  \[281] ,
  \[282] ,
  \[8320] ,
  \[7859] ,
  \[13634] ,
  \[11976] ,
  \[10058] ,
  \[11250] ,
  \[10057] ,
  \[1759] ,
  \[286] ,
  \[10787] ,
  \[21501] ,
  \[287] ,
  \[22361] ,
  \[3081] ,
  \[9184] ,
  \[10059] ,
  \[288] ,
  \[289] ,
  \[5471] ,
  \[5809] ,
  \[12449] ,
  \[2954] ,
  \[13641] ,
  \[4614] ,
  \[12443] ,
  \[1030] ,
  \[10060] ,
  \[14103] ,
  \[7134] ,
  \[14106] ,
  \[11257] ,
  \[4280] ,
  \[627] ,
  \[3421] ,
  \[1033] ,
  \[13648] ,
  \[1763] ,
  \[290] ,
  \[11259] ,
  \[291] ,
  \[22363] ,
  \[292] ,
  \[7869] ,
  \[293] ,
  \[22365] ,
  \[8331] ,
  \[11986] ,
  \[10068] ,
  \[13646] ,
  \[6675] ,
  \[10797] ,
  \[4288] ,
  \[9194] ,
  \[298] ,
  \[2963] ,
  \[10064] ,
  \[299] ,
  \[3093] ,
  \[14117] ,
  \[10063] ,
  \[13651] ,
  \[12454] ,
  \[634] ,
  \[10795] ,
  \[14114] ,
  \[4625] ,
  \[2237] ,
  \[7143] ,
  \[11600] ,
  \[21519] ,
  \[3430] ,
  \[10072] ,
  \[11602] ,
  \[5488] ,
  \[13657] ,
  \[7877] ,
  \[1776] ,
  \[11993] ,
  \[11266] ,
  \[11608] ,
  \[21521] ,
  \[3438] ,
  \[4298] ,
  \[5827] ,
  \[10079] ,
  \[2973] ,
  \[641] ,
  \[14127] ,
  \[10073] ,
  \[13661] ,
  \[10076] ,
  \[5493] ,
  \[14124] ,
  \[7153] ,
  \[12466] ,
  \[4636] ,
  \[1781] ,
  \[11610] ,
  \[22389] ,
  \[5100] ,
  \[5498] ,
  \[21523] ,
  \[7887] ,
  \[14132] ,
  \[21525] ,
  \[8350] ,
  \[1786] ,
  \[10416] ,
  \[13663] ,
  \[11275] ,
  \[10088] ,
  \[12806] ,
  \[3447] ,
  \[6695] ,
  \[22391] ,
  \[2982] ,
  \[14138] ,
  \[11619] ,
  \[14137] ,
  \[13672] ,
  \[12479] ,
  \[7162] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[4647] ,
  \[2259] ,
  \[22001] ,
  \[7895] ,
  \[19] ,
  \[1063] ,
  \[12817] ,
  \[22393] ,
  \[7501] ,
  \[10426] ,
  \[22395] ,
  \[14141] ,
  \[11285] ,
  \[1798] ,
  \[5845] ,
  \[3457] ,
  \[2990] ,
  \[20] ,
  \[11627] ,
  \[21] ,
  \[13680] ,
  \[11292] ,
  \[10099] ,
  \[22] ,
  \[14148] ,
  \[1404] ,
  \[22003] ,
  \[12822] ,
  \[23] ,
  \[7170] ,
  \[12489] ,
  \[6311] ,
  \[8368] ,
  \[22005] ,
  \[10095] ,
  \[4656] ,
  \[28] ,
  \[21549] ,
  \[29] ,
  \[7176] ,
  \[8707] ,
  \[11294] ,
  \[6319] ,
  \[14152] ,
  \[1076] ,
  \[2605] ,
  \[7511] ,
  \[12824] ,
  \[14151] ,
  \[3465] ,
  \[10435] ,
  \[9569] ,
  \[22017] ,
  \[5855] ,
  \[13686] ,
  \[30] ,
  \[21551] ,
  \[12100] ,
  \[22019] ,
  \[31] ,
  \[10441] ,
  \[32] ,
  \[14158] ,
  \[22013] ,
  \[12832] ,
  \[33] ,
  \[14157] ,
  \[7180] ,
  \[12499] ,
  \[34] ,
  \[672] ,
  \[12494] ,
  \[7519] ,
  \[22015] ,
  \[35] ,
  \[4664] ,
  \[2276] ,
  \[3805] ,
  \[36] ,
  \[11635] ,
  \[37] ,
  \[38] ,
  \[12108] ,
  \[22021] ,
  \[1083] ,
  \[10449] ,
  \[21553] ,
  \[11641] ,
  \[10444] ,
  \[6329] ,
  \[21555] ,
  \[2615] ,
  \[5863] ,
  \[3475] ,
  \[13694] ,
  \[9579] ,
  \[22027] ,
  \[13696] ,
  \[1421] ,
  \[2281] ,
  \[12110] ,
  \[11647] ,
  \[10452] ,
  \[13308] ,
  \[5138] ,
  \[22023] ,
  \[11649] ,
  \[43] ,
  \[8387] ,
  \[44] ,
  \[7529] ,
  \[22025] ,
  \[11643] ,
  \[45] ,
  \[4674] ,
  \[2286] ,
  \[21567] ,
  \[1090] ,
  \[7193] ,
  \[10457] ,
  \[686] ,
  \[14166] ,
  \[21569] ,
  \[3480] ,
  \[12118] ,
  \[12848] ,
  \[6337] ,
  \[10459] ,
  \[21563] ,
  \[2623] ,
  \[10454] ,
  \[21565] ,
  \[3484] ,
  \[13311] ,
  \[5873] ,
  \[12843] ,
  \[9589] ,
  \[12116] ,
  \[22037] ,
  \[21571] ,
  \[21909] ,
  \[22039] ,
  \[11657] ,
  \[13318] ,
  \[1434] ,
  \[7537] ,
  \[14177] ,
  \[4682] ,
  \[8397] ,
  \[3823] ,
  \[12851] ,
  \[54] ,
  \[55] ,
  \[8731] ,
  \[56] ,
  \[21577] ,
  \[11655] ,
  \[57] ,
  \[2298] ,
  \[21911] ,
  \[22041] ,
  \[12127] ,
  \[6347] ,
  \[300] ,
  \[21573] ,
  \[2633] ,
  \[301] ,
  \[10464] ,
  \[5881] ,
  \[12859] ,
  \[302] ,
  \[21575] ,
  \[303] ,
  \[10466] ,
  \[12853] ,
  \[304] ,
  \[305] ,
  \[9202] ,
  \[3497] ,
  \[12125] ,
  \[1441] ,
  \[306] ,
  \[12130] ,
  \[307] ,
  \[61] ,
  \[308] ,
  \[62] ,
  \[10809] ,
  \[21913] ,
  \[7547] ,
  \[63] ,
  \[14187] ,
  \[12861] ,
  \[11664] ,
  \[64] ,
  \[3104] ,
  \[10803] ,
  \[21915] ,
  \[65] ,
  \[4694] ,
  \[8011] ,
  \[11666] ,
  \[66] ,
  \[10805] ,
  \[21587] ,
  \[1448] ,
  \[67] ,
  \[13326] ,
  \[6355] ,
  \[68] ,
  \[21589] ,
  \[2641] ,
  \[5160] ,
  \[12867] ,
  \[11672] ,
  \[8746] ,
  \[5891] ,
  \[12139] ,
  \[10473] ,
  \[313] ,
  \[12133] ,
  \[7552] ,
  \[314] ,
  \[10475] ,
  \[21927] ,
  \[315] ,
  \[4306] ,
  \[9212] ,
  \[10817] ,
  \[5896] ,
  \[21591] ,
  \[21929] ,
  \[22059] ,
  \[3841] ,
  \[10481] ,
  \[14198] ,
  \[21923] ,
  \[7557] ,
  \[12872] ,
  \[73] ,
  \[11674] ,
  \[74] ,
  \[21925] ,
  \[75] ,
  \[10815] ,
  \[10820] ,
  \[6365] ,
  \[13335] ,
  \[21931] ,
  \[2651] ,
  \[8754] ,
  \[22061] ,
  \[12878] ,
  \[13340] ,
  \[10483] ,
  \[12874] ,
  \[9220] ,
  \[8029] ,
  \[21937] ,
  \[12146] ,
  \[4316] ,
  \[10828] ,
  \[11688] ,
  \[6705] ,
  \[21939] ,
  \[2659] ,
  \[13348] ,
  \[21933] ,
  \[9955] ,
  \[1464] ,
  \[22063] ,
  \[11689] ,
  \[5512] ,
  \[84] ,
  \[21935] ,
  \[7569] ,
  \[22065] ,
  \[11683] ,
  \[85] ,
  \[10826] ,
  \[9958] ,
  \[6373] ,
  \[86] ,
  \[3126] ,
  \[22407] ,
  \[87] ,
  \[10830] ,
  \[8763] ,
  \[21941] ,
  \[22409] ,
  \[5517] ,
  \[1803] ,
  \[11692] ,
  \[331] ,
  \[22403] ,
  \[5182] ,
  \[332] ,
  \[10493] ,
  \[12884] ,
  \[333] ,
  \[22405] ,
  \[4324] ,
  \[12153] ,
  \[1807] ,
  \[334] ,
  \[21947] ,
  \[335] ,
  \[6714] ,
  \[1471] ,
  \[7574] ,
  \[11698] ,
  \[336] ,
  \[21949] ,
  \[2669] ,
  \[337] ,
  \[22411] ,
  \[91] ,
  \[3861] ,
  \[338] ,
  \[92] ,
  \[21943] ,
  \[93] ,
  \[12891] ,
  \[94] ,
  \[21945] ,
  \[7579] ,
  \[95] ,
  \[10836] ,
  \[9238] ,
  \[6383] ,
  \[5524] ,
  \[96] ,
  \[13353] ,
  \[1478] ,
  \[10110] ,
  \[7913] ,
  \[22417] ,
  \[97] ,
  \[10840] ,
  \[8773] ,
  \[98] ,
  \[21951] ,
  \[12500] ,
  \[12898] ,
  \[13360] ,
  \[22413] ,
  \[8047] ,
  \[343] ,
  \[6722] ,
  \[22415] ,
  \[4334] ,
  \[12163] ,
  \[12893] ,
  \[344] ,
  \[21957] ,
  \[2677] ,
  \[11305] ,
  \[345] ,
  \[10848] ,
  \[12895] ,
  \[21959] ,
  \[22089] ,
  \[3142] ,
  \[21953] ,
  \[12172] ,
  \[5199] ,
  \[13702] ,
  \[12509] ,
  \[6391] ,
  \[21955] ,
  \[10846] ,
  \[8781] ,
  \[12503] ,
  \[1820] ,
  \[22427] ,
  \[21961] ,
  \[12510] ,
  \[22091] ,
  \[22429] ,
  \[13370] ,
  \[13708] ,
  \[5538] ,
  \[4342] ,
  \[8057] ,
  \[12179] ,
  \[1825] ,
  \[7591] ,
  \[6732] ,
  \[11316] ,
  \[9251] ,
  \[21967] ,
  \[2687] ,
  \[10857] ,
  \[21969] ,
  \[6006] ,
  \[9983] ,
  \[22431] ,
  \[10129] ,
  \[3152] ,
  \[21963] ,
  \[22093] ,
  \[10854] ,
  \[12181] ,
  \[3883] ,
  \[12519] ,
  \[10123] ,
  \[21965] ,
  \[7599] ,
  \[22095] ,
  \[5543] ,
  \[8791] ,
  \[12513] ,
  \[7203] ,
  \[1830] ,
  \[7933] ,
  \[21971] ,
  \[12520] ,
  \[8065] ,
  \[12187] ,
  \[13718] ,
  \[4351] ,
  \[361] ,
  \[6740] ,
  \[1105] ,
  \[12189] ,
  \[362] ,
  \[2695] ,
  \[363] ,
  \[364] ,
  \[21977] ,
  \[9991] ,
  \[11325] ,
  \[365] ,
  \[6015] ,
  \[10137] ,
  \[366] ,
  \[3160] ,
  \[21979] ,
  \[367] ,
  \[13388] ,
  \[8405] ,
  \[11332] ,
  \[368] ,
  \[5550] ,
  \[2303] ,
  \[21973] ,
  \[10134] ,
  \[12529] ,
  \[10133] ,
  \[6749] ,
  \[10863] ,
  \[21975] ,
  \[703] ,
  \[12523] ,
  \[10135] ,
  \[10865] ,
  \[9269] ,
  \[2307] ,
  \[13383] ,
  \[13386] ,
  \[21981] ,
  \[1842] ,
  \[8075] ,
  \[12197] ,
  \[13728] ,
  \[10141] ,
  \[10871] ,
  \[3502] ,
  \[373] ,
  \[1847] ,
  \[374] ,
  \[3506] ,
  \[11335] ,
  \[375] ,
  \[12195] ,
  \[3170] ,
  \[10877] ,
  \[8415] ,
  \[10149] ,
  \[11341] ,
  \[12539] ,
  \[6759] ,
  \[10146] ,
  \[4705] ,
  \[12536] ,
  \[8083] ,
  \[13396] ,
  \[12535] ,
  \[1851] ,
  \[716] ,
  \[3178] ,
  \[1122] ,
  \[7955] ,
  \[13008] ,
  \[5900] ,
  \[7227] ,
  \[13737] ,
  \[12542] ,
  \[6033] ,
  \[10158] ,
  \[2320] ,
  \[8423] ,
  \[13736] ,
  \[21999] ,
  \[4378] ,
  \[3519] ,
  \[14208] ,
  \[11351] ,
  \[10154] ,
  \[10884] ,
  \[13012] ,
  \[5572] ,
  \[2325] ,
  \[723] ,
  \[12543] ,
  \[4716] ,
  \[8093] ,
  \[11358] ,
  \[3188] ,
  \[21609] ,
  \[12550] ,
  \[10892] ,
  \[391] ,
  \[1135] ,
  \[392] ,
  \[6771] ,
  \[393] ,
  \[5913] ,
  \[394] ,
  \[395] ,
  \[2330] ,
  \[8433] ,
  \[13746] ,
  \[1869] ,
  \[396] ,
  \[21611] ,
  \[3528] ,
  \[397] ,
  \[12557] ,
  \[398] ,
  \[10501] ,
  \[730] ,
  \[11361] ,
  \[2335] ,
  \[3196] ,
  \[14213] ,
  \[11368] ,
  \[4727] ,
  \[9633] ,
  \[1142] ,
  \[12560] ,
  \[7975] ,
  \[13028] ,
  \[10509] ,
  \[14220] ,
  \[21613] ,
  \[12561] ,
  \[21615] ,
  \[5923] ,
  \[8441] ,
  \[6053] ,
  \[11366] ,
  \[3536] ,
  \[1149] ,
  \[13756] ,
  \[13025] ,
  \[12900] ,
  \[13030] ,
  \[12567] ,
  \[2343] ,
  \[4002] ,
  \[7250] ,
  \[10176] ,
  \[11703] ,
  \[5594] ,
  \[21627] ,
  \[12566] ,
  \[11705] ,
  \[4007] ,
  \[21629] ,
  \[4738] ,
  \[10181] ,
  \[14230] ,
  \[13037] ,
  \[21623] ,
  \[9645] ,
  \[11711] ,
  \[10514] ,
  \[11374] ,
  \[21625] ,
  \[7259] ,
  \[10516] ,
  \[8451] ,
  \[11376] ,
  \[1887] ,
  \[12903] ,
  \[3546] ,
  \[13763] ,
  \[6794] ,
  \[10520] ,
  \[11380] ,
  \[12905] ,
  \[21631] ,
  \[10522] ,
  \[6401] ,
  \[12911] ,
  \[4013] ,
  \[8458] ,
  \[13771] ,
  \[10186] ,
  \[11713] ,
  \[21637] ,
  \[2357] ,
  \[7993] ,
  \[10528] ,
  \[12575] ,
  \[14236] ,
  \[9653] ,
  \[12917] ,
  \[21633] ,
  \[4749] ,
  \[6070] ,
  \[12582] ,
  \[11389] ,
  \[11721] ,
  \[6409] ,
  \[21635] ,
  \[3554] ,
  \[7269] ,
  \[11383] ,
  \[14241] ,
  \[12913] ,
  \[6074] ,
  \[22107] ,
  \[10530] ,
  \[13046] ,
  \[5216] ,
  \[13775] ,
  \[22109] ,
  \[10199] ,
  \[11391] ,
  \[22103] ,
  \[13782] ,
  \[10193] ,
  \[762] ,
  \[8800] ,
  \[7609] ,
  \[22105] ,
  \[12583] ,
  \[10195] ,
  \[4025] ,
  \[21647] ,
  \[12586] ,
  \[10537] ,
  \[21649] ,
  \[2369] ,
  \[9663] ,
  \[22111] ,
  \[4029] ,
  \[10539] ,
  \[7277] ,
  \[12592] ,
  \[11399] ,
  \[5221] ,
  \[11731] ,
  \[5951] ,
  \[6419] ,
  \[3564] ,
  \[2705] ,
  \[8808] ,
  \[11393] ,
  \[14251] ,
  \[12923] ,
  \[22117] ,
  \[1511] ,
  \[5226] ,
  \[21651] ,
  \[22119] ,
  \[13060] ,
  \[4760] ,
  \[6087] ,
  \[13790] ,
  \[8476] ,
  \[1514] ,
  \[7617] ,
  \[22113] ,
  \[3903] ,
  \[22115] ,
  \[12593] ,
  \[4035] ,
  \[4765] ,
  \[11005] ,
  \[12596] ,
  \[6424] ,
  \[775] ,
  \[11740] ,
  \[10547] ,
  \[14256] ,
  \[9673] ,
  \[1182] ,
  \[12208] ,
  \[22121] ,
  \[13798] ,
  \[3572] ,
  \[7287] ,
  \[2713] ,
  \[12209] ,
  \[6429] ,
  \[12939] ,
  \[14262] ,
  \[8818] ,
  \[12203] ,
  \[12933] ,
  \[10545] ,
  \[13063] ,
  \[22127] ,
  \[11018] ,
  \[6095] ,
  \[13065] ,
  \[22129] ,
  \[4770] ,
  \[2382] ,
  \[7627] ,
  \[22123] ,
  \[782] ,
  \[13409] ,
  \[11013] ,
  \[1526] ,
  \[22125] ,
  \[11746] ,
  \[9681] ,
  \[10558] ,
  \[14263] ,
  \[4047] ,
  \[14266] ,
  \[21669] ,
  \[22131] ,
  \[12948] ,
  \[9684] ,
  \[12217] ,
  \[7296] ,
  \[5240] ,
  \[10559] ,
  \[5970] ,
  \[3582] ,
  \[2723] ,
  \[8826] ,
  \[789] ,
  \[13412] ,
  \[1195] ,
  \[10556] ,
  \[5245] ,
  \[13076] ,
  \[2728] ,
  \[21671] ,
  \[8494] ,
  \[7635] ,
  \[3921] ,
  \[13417] ,
  \[14277] ,
  \[6441] ,
  \[11753] ,
  \[4784] ,
  \[8101] ,
  \[1537] ,
  \[4055] ,
  \[794] ,
  \[11025] ,
  \[11755] ,
  \[10568] ,
  \[10900] ,
  \[14273] ,
  \[14276] ,
  \[3590] ,
  \[13415] ,
  \[12228] ,
  \[6446] ,
  \[12958] ,
  \[11762] ,
  \[13087] ,
  \[21673] ,
  \[4789] ,
  \[2733] ,
  \[8836] ,
  \[11761] ,
  \[2004] ,
  \[5252] ,
  \[10563] ,
  \[21675] ,
  \[403] ,
  \[404] ,
  \[10565] ,
  \[9699] ,
  \[405] ,
  \[10570] ,
  \[7645] ,
  \[22149] ,
  \[3599] ,
  \[10909] ,
  \[5988] ,
  \[6451] ,
  \[12961] ,
  \[9308] ,
  \[8111] ,
  \[4065] ,
  \[3206] ,
  \[14284] ,
  \[21687] ,
  \[13423] ,
  \[11035] ,
  \[1548] ,
  \[11765] ,
  \[10578] ,
  \[10910] ,
  \[14283] ,
  \[4796] ,
  \[21689] ,
  \[13425] ,
  \[8844] ,
  \[22151] ,
  \[21683] ,
  \[11771] ,
  \[12969] ,
  \[14292] ,
  \[2015] ,
  \[21685] ,
  \[13431] ,
  \[12234] ,
  \[2745] ,
  \[10576] ,
  \[8119] ,
  \[12963] ,
  \[414] ,
  \[7653] ,
  \[415] ,
  \[5266] ,
  \[416] ,
  \[21691] ,
  \[3940] ,
  \[12970] ,
  \[417] ,
  \[10919] ,
  \[14298] ,
  \[22153] ,
  \[14297] ,
  \[11044] ,
  \[3214] ,
  \[10913] ,
  \[22155] ,
  \[4074] ,
  \[11773] ,
  \[13434] ,
  \[6463] ,
  \[9319] ,
  \[21697] ,
  \[11775] ,
  \[2750] ,
  \[1559] ,
  \[3948] ,
  \[8854] ,
  \[13440] ,
  \[12247] ,
  \[10921] ,
  \[21693] ,
  \[11051] ,
  \[5271] ,
  \[11781] ,
  \[6800] ,
  \[10584] ,
  \[13442] ,
  \[12979] ,
  \[21695] ,
  \[2755] ,
  \[10586] ,
  \[8129] ,
  \[12243] ,
  \[12973] ,
  \[7663] ,
  \[22167] ,
  \[10927] ,
  \[22169] ,
  \[11787] ,
  \[13448] ,
  \[5278] ,
  \[10929] ,
  \[22163] ,
  \[4082] ,
  \[3223] ,
  \[0] ,
  \[6471] ,
  \[12981] ,
  \[5612] ,
  \[11053] ,
  \[22165] ,
  \[9328] ,
  \[8862] ,
  \[10597] ,
  \[2031] ,
  \[3958] ,
  \[22171] ,
  \[12257] ,
  \[11061] ,
  \[4422] ,
  \[8137] ,
  \[12989] ,
  \[13451] ,
  \[7671] ,
  \[12983] ,
  \[2767] ,
  \[1570] ,
  \[22177] ,
  \[436] ,
  \[22179] ,
  \[437] ,
  \[4091] ,
  \[438] ,
  \[22173] ,
  \[439] ,
  \[9336] ,
  \[6481] ,
  \[10206] ,
  \[22175] ,
  \[13454] ,
  \[8871] ,
  \[11796] ,
  \[10935] ,
  \[3966] ,
  \[11070] ,
  \[11407] ,
  \[22181] ,
  \[13460] ,
  \[12267] ,
  \[10211] ,
  \[5290] ,
  \[440] ,
  \[4431] ,
  \[441] ,
  \[8147] ,
  \[6489] ,
  \[442] ,
  \[13461] ,
  \[2775] ,
  \[7681] ,
  \[443] ,
  \[6822] ,
  \[11405] ,
  \[22187] ,
  \[10948] ,
  \[1581] ,
  \[12995] ,
  \[11077] ,
  \[22189] ,
  \[3241] ,
  \[12607] ,
  \[448] ,
  \[5630] ,
  \[22183] ,
  \[449] ,
  \[9346] ,
  \[12604] ,
  \[7689] ,
  \[22185] ,
  \[13464] ,
  \[3975] ,
  \[8881] ,
  \[12603] ,
  \[10215] ,
  \[8152] ,
  \[11080] ,
  \[22191] ,
  \[10952] ,
  \[13470] ,
  \[11082] ,
  \[450] ,
  \[2053] ,
  \[13807] ,
  \[451] ,
  \[5639] ,
  \[8157] ,
  \[6499] ,
  \[452] ,
  \[2785] ,
  \[11413] ,
  \[1926] ,
  \[453] ,
  \[12273] ,
  \[454] ,
  \[11415] ,
  \[455] ,
  \[11088] ,
  \[6105] ,
  \[456] ,
  \[457] ,
  \[9354] ,
  \[12617] ,
  \[11422] ,
  \[458] ,
  \[10959] ,
  \[12282] ,
  \[6838] ,
  \[13479] ,
  \[13811] ,
  \[12614] ,
  \[7699] ,
  \[3985] ,
  \[1597] ,
  \[12613] ,
  \[13473] ,
  \[7304] ,
  \[11090] ,
  \[8893] ,
  \[1202] ,
  \[12287] ,
  \[5649] ,
  \[12289] ,
  \[2794] ,
  \[11424] ,
  \[13481] ,
  \[463] ,
  \[9360] ,
  \[8169] ,
  \[6113] ,
  \[464] ,
  \[10238] ,
  \[1938] ,
  \[465] ,
  \[1209] ,
  \[11430] ,
  \[12628] ,
  \[4458] ,
  \[3261] ,
  \[13820] ,
  \[11432] ,
  \[10969] ,
  \[13487] ,
  \[11099] ,
  \[2404] ,
  \[3994] ,
  \[10236] ,
  \[11096] ,
  \[10235] ,
  \[7314] ,
  \[2071] ,
  \[8174] ,
  \[10242] ,
  \[5657] ,
  \[12297] ,
  \[6851] ,
  \[8179] ,
  \[6123] ,
  \[474] ,
  \[8512] ,
  \[475] ,
  \[9372] ,
  \[12295] ,
  \[13826] ,
  \[1949] ,
  \[476] ,
  \[4467] ,
  \[12638] ,
  \[477] ,
  \[13100] ,
  \[3609] ,
  \[10979] ,
  \[13497] ,
  \[10976] ,
  \[7322] ,
  \[9379] ,
  \[5667] ,
  \[13838] ,
  \[6131] ,
  \[11443] ,
  \[14301] ,
  \[13103] ,
  \[10987] ,
  \[3618] ,
  \[13835] ,
  \[13110] ,
  \[14308] ,
  \[11451] ,
  \[3283] ,
  \[13112] ,
  \[12649] ,
  \[5672] ,
  \[13841] ,
  \[823] ,
  \[8191] ,
  \[2426] ,
  \[9389] ,
  \[21707] ,
  \[1960] ,
  \[5676] ,
  \[21709] ,
  \[7335] ,
  \[13847] ,
  \[6141] ,
  \[13849] ,
  \[14311] ,
  \[8199] ,
  \[4485] ,
  \[2097] ,
  \[3626] ,
  \[11455] ,
  \[6874] ,
  \[8533] ,
  \[10267] ,
  \[21711] ,
  \[4822] ,
  \[6149] ,
  \[12659] ,
  \[12654] ,
  \[103] ,
  \[10996] ,
  \[104] ,
  \[105] ,
  \[1241] ,
  \[1971] ,
  \[836] ,
  \[14316] ,
  \[13858] ,
  \[5689] ,
  \[9006] ,
  \[13129] ,
  \[11463] ,
  \[14321] ,
  \[10605] ,
  \[9739] ,
  \[13126] ,
  \[3638] ,
  \[13855] ,
  \[11472] ,
  \[4101] ,
  \[6887] ,
  \[14328] ,
  \[13132] ,
  \[2444] ,
  \[6159] ,
  \[11804] ,
  \[12664] ,
  \[843] ,
  \[114] ,
  \[5694] ,
  \[115] ,
  \[9742] ,
  \[116] ,
  \[21729] ,
  \[12670] ,
  \[117] ,
  \[1982] ,
  \[9014] ,
  \[13868] ,
  \[4109] ,
  \[5698] ,
  \[4839] ,
  \[3642] ,
  \[1254] ,
  \[5301] ,
  \[10614] ,
  \[7358] ,
  \[11473] ,
  \[14331] ,
  \[13864] ,
  \[11476] ,
  \[10288] ,
  \[13136] ,
  \[21731] ,
  \[3648] ,
  \[10622] ,
  \[8555] ,
  \[6167] ,
  \[13870] ,
  \[11482] ,
  \[850] ,
  \[121] ,
  \[14337] ,
  \[13142] ,
  \[122] ,
  \[12674] ,
  \[123] ,
  \[11813] ,
  \[14339] ,
  \[12673] ,
  \[124] ,
  \[10285] ,
  \[125] ,
  \[1261] ,
  \[11488] ,
  \[126] ,
  \[11820] ,
  \[127] ,
  \[10292] ,
  \[13878] ,
  \[128] ,
  \[6507] ,
  \[1993] ,
  \[4119] ,
  \[11822] ,
  \[21733] ,
  \[12682] ,
  \[12681] ,
  \[9027] ,
  \[21735] ,
  \[10626] ,
  \[13144] ,
  \[11486] ,
  \[1268] ,
  \[10630] ,
  \[22209] ,
  \[5317] ,
  \[10632] ,
  \[13150] ,
  \[3659] ,
  \[2462] ,
  \[6177] ,
  \[13880] ,
  \[10299] ,
  \[7707] ,
  \[11829] ,
  \[13152] ,
  \[7371] ,
  \[133] ,
  \[10296] ,
  \[134] ,
  \[21747] ,
  \[135] ,
  \[10638] ,
  \[12685] ,
  \[4127] ,
  \[21749] ,
  \[22211] ,
  \[1273] ,
  \[2802] ,
  \[13888] ,
  \[6517] ,
  \[21743] ,
  \[13887] ,
  \[12692] ,
  \[12691] ,
  \[11494] ,
  \[21745] ,
  \[8909] ,
  \[11496] ,
  \[10635] ,
  \[6185] ,
  \[11838] ,
  \[13155] ,
  \[21751] ,
  \[2471] ,
  \[8574] ,
  \[11107] ,
  \[4861] ,
  \[7717] ,
  \[22213] ,
  \[1615] ,
  \[13161] ,
  \[13891] ,
  \[22215] ,
  \[21757] ,
  \[11105] ,
  \[10648] ,
  \[12695] ,
  \[6525] ,
  \[4137] ,
  \[21759] ,
  \[2812] ,
  \[13898] ,
  \[21753] ,
  \[10644] ,
  \[1285] ,
  \[12309] ,
  \[21755] ,
  \[7389] ,
  \[13899] ,
  \[10646] ,
  \[13163] ,
  \[12306] ,
  \[22227] ,
  \[12305] ,
  \[6195] ,
  \[11848] ,
  \[13165] ,
  \[21761] ,
  \[7725] ,
  \[22229] ,
  \[3679] ,
  \[11119] ,
  \[151] ,
  \[22223] ,
  \[5339] ,
  \[152] ,
  \[882] ,
  \[13171] ,
  \[11113] ,
  \[153] ,
  \[22225] ,
  \[9050] ,
  \[11116] ,
  \[154] ,
  \[21767] ,
  \[155] ,
  \[4146] ,
  \[2820] ,
  \[156] ,
  \[6535] ,
  \[21769] ,
  \[2489] ,
  \[13505] ,
  \[157] ,
  \[22231] ,
  \[4878] ,
  \[158] ,
  \[21763] ,
  \[10654] ,
  \[13512] ,
  \[12319] ,
  \[21765] ,
  \[12316] ,
  \[22237] ,
  \[10660] ,
  \[12315] ,
  \[13175] ,
  \[21771] ,
  \[2829] ,
  \[7735] ,
  \[22239] ,
  \[11857] ,
  \[11129] ,
  \[22233] ,
  \[13181] ,
  \[163] ,
  \[22235] ,
  \[4154] ,
  \[11126] ,
  \[8931] ,
  \[164] ,
  \[6543] ,
  \[11125] ,
  \[165] ,
  \[11855] ,
  \[895] ,
  \[22241] ,
  \[13520] ,
  \[4889] ,
  \[12329] ,
  \[13189] ,
  \[8209] ,
  \[9401] ,
  \[13183] ,
  \[7013] ,
  \[7743] ,
  \[22247] ,
  \[3697] ,
  \[11138] ,
  \[11868] ,
  \[2839] ,
  \[22249] ,
  \[10672] ,
  \[22243] ,
  \[3303] ,
  \[13192] ,
  \[4163] ,
  \[13529] ,
  \[22245] ,
  \[6553] ,
  \[11135] ,
  \[2110] ,
  \[21789] ,
  \[13525] ,
  \[22251] ,
  \[13198] ,
  \[5361] ,
  \[8217] ,
  \[4503] ,
  \[13531] ,
  \[7753] ,
  \[7024] ,
  \[2848] ,
  \[9413] ,
  \[21791] ,
  \[13538] ,
  \[10681] ,
  \[1654] ,
  \[181] ,
  \[11879] ,
  \[12341] ,
  \[11144] ,
  \[182] ,
  \[6561] ,
  \[4173] ,
  \[183] ,
  \[11146] ,
  \[184] ,
  \[8952] ,
  \[185] ,
  \[186] ,
  \[187] ,
  \[11152] ,
  \[188] ,
  \[10689] ,
  \[21793] ,
  \[14007] ,
  \[8227] ,
  \[4513] ,
  \[21795] ,
  \[7761] ,
  \[2856] ,
  \[14004] ,
  \[2127] ,
  \[14003] ,
  \[11158] ,
  \[11888] ,
  \[6905] ,
  \[22269] ,
  \[3321] ,
  \[13547] ,
  \[4182] ,
  \[5711] ,
  \[6571] ,
  \[8960] ,
  \[193] ,
  \[194] ,
  \[13543] ,
  \[195] ,
  \[13545] ,
  \[22271] ,
  \[9094] ,
  \[8235] ,
  \[10699] ,
  \[14017] ,
  \[5719] ,
  \[4522] ,
  \[12359] ,
  \[6579] ,
  \[10693] ,
  \[5383] ,
  \[12353] ,
  \[14014] ,
  \[14013] ,
  \[1671] ,
  \[11898] ,
  \[4190] ,
  \[22273] ,
  \[13559] ,
  \[8970] ,
  \[22275] ,
  \[11166] ,
  \[13553] ,
  \[11895] ,
  \[4530] ,
  \[3339] ,
  \[8245] ,
  \[4199] ,
  \[14028] ,
  \[6920] ,
  \[5729] ,
  \[12369] ,
  \[2874] ,
  \[6589] ,
  \[8978] ,
  \[7781] ,
  \[7052] ,
  \[11506] ,
  \[14024] ,
  \[12366] ,
  \[22287] ,
  \[12365] ,
  \[10317] ,
  \[2149] ,
  \[22289] ,
  \[14025] ,
  \[10319] ,
  \[4539] ,
  \[22283] ,
  \[6928] ,
  \[13902] ,
  \[12709] ,
  \[22285] ,
  \[11175] ,
  \[1688] ,
  \[8253] ,
  \[2880] ,
  \[11518] ,
  \[22291] ,
  \[5737] ,
  \[13570] ,
  \[6597] ,
  \[14038] ,
  \[12379] ,
  \[13909] ,
  \[8988] ,
  \[6203] ,
  \[14034] ,
  \[7063] ,
  \[12376] ,
  \[22297] ,
  \[12375] ,
  \[14035] ,
  \[1693] ,
  \[11522] ,
  \[4549] ,
  \[22293] ,
  \[6938] ,
  \[12719] ,
  \[10323] ,
  \[9457] ,
  \[13579] ,
  \[11183] ,
  \[10326] ,
  \[22295] ,
  \[1698] ,
  \[5015] ,
  \[3357] ,
  \[8263] ,
  \[11190] ,
  \[1302] ,
  \[7405] ,
  \[5747] ,
  \[12387] ,
  \[11192] ,
  \[10331] ,
  \[8996] ,
  \[14047] ,
  \[7072] ,
  \[6213] ,
  \[8602] ,
  \[12386] ,
  \[11198] ,
  \[12390] ,
  \[13915] ,
  \[567] ,
  \[6946] ,
  \[4558] ,
  \[9464] ,
  \[13587] ,
  \[11199] ,
  \[902] ,
  \[13921] ,
  \[8271] ,
  \[10335] ,
  \[5755] ,
  \[12725] ,
  \[2171] ,
  \[2509] ,
  \[12730] ,
  \[12397] ,
  \[10341] ,
  \[11539] ,
  \[14057] ,
  \[909] ,
  \[12001] ,
  \[7080] ,
  \[13592] ,
  \[1315] ,
  \[6221] ;
assign
  \[8612]  = ~\[10073]  & (~v15 & ~\[10774] ),
  \[12396]  = ~v1 | (~\[10099]  | (~\[10060]  | ~\[5405] )),
  \[11535]  = ~v11 | (~\[10063]  | ~v12),
  \[10348]  = ~v5 | (~\[10134]  | ~v7),
  \[14053]  = ~v13 | (~\[10088]  | (~v15 | ~\[2097] )),
  \[4566]  = ~\[10059]  & (~v0 & ~v2),
  \[14056]  = ~\[10134]  | (~\[10176]  | (~v0 | ~v2)),
  \[6956]  = ~\[10073]  & (~v15 & (~\[11627]  & ~v13)),
  \[13200]  = ~v1 | (~\[10099]  | ~v3),
  \[4900]  = ~\[10073]  & (~v13 & (~v15 & ~\[12649] )),
  \[12737]  = ~v4 | (~v7 | ~\[10058] ),
  \[13597]  = ~v11 | ~v8,
  \[10344]  = ~v5 | (~\[10134]  | ~v7),
  \[9477]  = ~\[10133]  & (~v12 & (~\[10236]  & ~v4)),
  \[3375]  = ~\[10068]  & (~v9 & ~v12),
  \[8281]  = ~\[10133]  & (~v5 & (~\[10959]  & ~v3)),
  \[4905]  = ~v6 & (~v5 & ~v8),
  \[5765]  = ~v6 & (~v5 & (~\[12217]  & ~v3)),
  \[12005]  = ~v7 | ~\[10236] ,
  \[1322]  = ~\[98]  & (~\[97]  & (~\[96]  & ~\[95] )),
  \[5037]  = ~v6 & (~v5 & ~v8),
  \[12740]  = ~v10 | (~v9 | ~\[10068] ),
  \[10352]  = ~v5 | (~\[10134]  | ~v7),
  \[12012]  = ~v1 | (~\[10099]  | ~v3),
  \[7427]  = ~v9 & (~v7 & ~\[10068] ),
  \[13937]  = ~v10 | (~v9 | ~\[10068] ),
  \[7090]  = ~\[10073]  & (~v15 & (~\[11552]  & ~v13)),
  \[6231]  = ~\[10059]  & (~v0 & (~v2 & ~\[11986] )),
  \[8620]  = ~\[10060]  & (~v1 & ~v3),
  \[8289]  = ~v10 & (~v9 & ~\[10088] ),
  \[3715]  = ~v10 & (~v9 & ~v12),
  \[584]  = ~\[14256]  & (~\[14213]  & ~\[14337] ),
  \[4575]  = ~\[10068]  & (~\[10058]  & ~v12),
  \[11545]  = ~v11 | (~\[10063]  | ~v12),
  \[6964]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[13206]  = ~v15 | (~v13 | ~\[3787] ),
  \[1329]  = ~\[94]  & (~\[93]  & (~\[92]  & ~\[91] )),
  \[14065]  = ~v13 | (~\[10088]  | (~v15 | ~\[2071] )),
  \[9484]  = ~\[10236]  & ~v4,
  \[4910]  = ~\[10060]  & (~v1 & ~v3),
  \[11552]  = ~v11 | ~v8,
  \[7098]  = ~\[10059]  & (~v0 & ~v2),
  \[6239]  = ~\[10068]  & (~v9 & ~v13),
  \[12749]  = ~v4 | (~v7 | ~\[10058] ),
  \[14072]  = ~v10 | ~v9,
  \[14071]  = ~v2 | (~\[10059]  | (~\[10176]  | ~\[2053] )),
  \[5773]  = ~\[10068]  & (~v9 & ~v12),
  \[3385]  = ~\[10133]  & (~v5 & ~\[13388] ),
  \[2526]  = ~\[10072]  & (~v12 & ~v14),
  \[8629]  = ~v10 & (~v9 & ~\[10088] ),
  \[21807]  = ~v13 | (~\[10073]  | (~\[7707]  | ~\[7717] )),
  \[12745]  = ~\[22109]  | (~\[22107]  | (~\[22105]  | ~\[22103] )),
  \[21471]  = ~v9 | (~\[10064]  | ~\[10057] ),
  \[926]  = ~\[299]  & (~\[298]  & (~\[300]  & ~\[12494] )),
  \[21809]  = ~v13 | (~\[10073]  | (~\[7689]  | ~\[7699] )),
  \[12020]  = ~v2 | ~\[10059] ,
  \[13948]  = ~v10 | (~v9 | ~\[10068] ),
  \[2193]  = ~v6 & (~v5 & ~v8),
  \[21803]  = ~v13 | (~\[10073]  | (~\[7743]  | ~\[7753] )),
  \[12752]  = ~v10 | (~v9 | ~\[10068] ),
  \[13219]  = ~v1 | (~\[10099]  | ~v3),
  \[21805]  = ~v13 | (~\[10073]  | (~\[7725]  | ~\[7735] )),
  \[8299]  = ~\[10060]  & (~v1 & (~v3 & ~\[10952] )),
  \[3725]  = ~v6 & (~v5 & (~\[13235]  & ~v3)),
  \[21477]  = ~v15 | (~\[10072]  | (~\[10060]  | ~\[10059] )),
  \[4585]  = ~v6 & (~v5 & ~\[12806] ),
  \[13216]  = ~v15 | ~v13,
  \[21479]  = ~v10 | (~\[10068]  | (~\[10028]  | ~v8)),
  \[21811]  = ~v13 | (~\[10073]  | (~\[7671]  | ~\[7681] )),
  \[12028]  = ~v0 | ~v2,
  \[2531]  = ~\[10058]  & (~v7 & ~v10),
  \[597]  = ~\[464]  & (~\[463]  & (~\[465]  & ~\[14132] )),
  \[10702]  = ~v2 | ~\[10059] ,
  \[14075]  = ~v13 | (~\[10088]  | ~v15),
  \[21473]  = ~v10 | (~\[10068]  | ~\[10049] ),
  \[11561]  = ~v11 | ~v8,
  \[4922]  = ~\[10073]  & (~v13 & (~v15 & ~\[12638] )),
  \[6249]  = ~v6 & (~v5 & ~\[11976] ),
  \[14082]  = ~v10 | ~v9,
  \[21475]  = ~\[10073]  | (~\[10072]  | (~\[10060]  | ~\[10059] )),
  \[3394]  = ~\[10068]  & (~v9 & (~v12 & ~\[13409] )),
  \[14081]  = ~v0 | (~v2 | (~\[10176]  | ~\[2031] )),
  \[5783]  = ~v6 & (~v5 & (~\[12209]  & ~v3)),
  \[933]  = ~\[293]  & (~\[292]  & (~\[291]  & ~\[290] )),
  \[8639]  = ~\[10059]  & (~v0 & (~v2 & ~\[10787] )),
  \[204]  = ~\[11581]  & (~\[11579]  & ~\[11587] ),
  \[21817]  = ~v13 | (~\[10073]  | (~\[7617]  | ~\[7627] )),
  \[5055]  = ~\[10064]  & (~v11 & (~\[10063]  & ~v8)),
  \[205]  = ~\[10073]  & (~v15 & (~\[11593]  & ~\[11591] )),
  \[11568]  = ~v5 | (~\[10134]  | ~v6),
  \[206]  = ~\[10073]  & (~v15 & (~\[11602]  & ~\[11600] )),
  \[3000]  = ~\[10072]  & (~v14 & (~\[13597]  & ~v12)),
  \[21481]  = ~v11 | (~v9 | ~\[10021] ),
  \[21819]  = ~v13 | (~\[10073]  | (~\[7599]  | ~\[7609] )),
  \[4927]  = ~\[10133]  & (~v5 & ~v8),
  \[12760]  = ~v11 | ~v8,
  \[207]  = ~\[10073]  & (~v15 & (~\[11610]  & ~\[11608] )),
  \[13958]  = ~v10 | (~v9 | ~\[10068] ),
  \[13227]  = ~v2 | ~\[10059] ,
  \[21813]  = ~v13 | (~\[10073]  | (~\[7653]  | ~\[7663] )),
  \[1344]  = ~\[87]  & (~\[86]  & (~\[85]  & ~\[84] )),
  \[3733]  = ~v10 & (~v9 & ~v12),
  \[9107]  = ~\[10134]  & ~v6,
  \[4593]  = ~\[10068]  & (~\[10058]  & ~v12),
  \[21815]  = ~v13 | (~\[10073]  | (~\[7635]  | ~\[7645] )),
  \[6982]  = ~\[10059]  & (~v0 & ~v2),
  \[21487]  = ~v12 | (~\[10073]  | (~\[10060]  | ~\[10059] )),
  \[10378]  = ~v1 | (~\[10099]  | ~v2),
  \[3008]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[21489]  = ~v9 | (~\[10064]  | ~\[9991] ),
  \[21821]  = ~\[7574]  | (~\[7579]  | ~\[7591] ),
  \[14085]  = ~v13 | (~\[10088]  | ~v15),
  \[12037]  = ~\[21975]  | (~\[21973]  | (~\[21971]  | ~\[21969] )),
  \[6257]  = ~\[10068]  & (~v9 & ~v13),
  \[10711]  = ~v0 | ~v2,
  \[21483]  = ~v12 | (~v15 | (~\[10060]  | ~\[10059] )),
  \[940]  = ~\[289]  & (~\[288]  & (~\[287]  & ~\[286] )),
  \[4931]  = ~\[10059]  & ~v0,
  \[2543]  = ~\[10060]  & (~v1 & (~v3 & ~\[13811] )),
  \[11571]  = ~v8 | (~\[10133]  | ~v11),
  \[211]  = ~\[10073]  & (~v15 & (~\[11649]  & ~\[11647] )),
  \[5791]  = ~\[10068]  & (~v9 & ~v12),
  \[8647]  = ~\[10058]  & (~v10 & ~\[10088] ),
  \[12769]  = ~v11 | ~v8,
  \[212]  = ~\[10073]  & (~v15 & (~\[11657]  & ~\[11655] )),
  \[11904]  = ~v0 | ~v2,
  \[21485]  = ~v14 | (~v13 | (~\[10076]  | ~\[10007] )),
  \[213]  = ~\[10073]  & (~v15 & (~\[11666]  & ~\[11664] )),
  \[10376]  = ~\[21615]  | (~\[21613]  | (~\[21611]  | ~\[21609] )),
  \[214]  = ~\[10073]  & (~v15 & (~\[11674]  & ~\[11672] )),
  \[21827]  = ~v13 | (~\[10073]  | (~\[7519]  | ~\[7529] )),
  \[9841]  = ~\[10176]  & (~v1 & ~v8),
  \[215]  = ~\[11688]  & ~\[11683] ,
  \[216]  = ~\[11689]  & (~v3 & (~\[11692]  & ~\[11698] )),
  \[21491]  = ~v10 | (~\[10068]  | ~\[9983] ),
  \[21829]  = ~v13 | (~\[10073]  | (~\[7501]  | ~\[7511] )),
  \[7455]  = ~\[10059]  & ~v0,
  \[217]  = ~\[10073]  & (~v15 & (~\[11705]  & ~\[11703] )),
  \[9844]  = ~\[10088]  & ~v14,
  \[13968]  = ~v1 | (~\[10099]  | (~v3 | ~\[2215] )),
  \[218]  = ~\[10073]  & (~v15 & (~\[11713]  & ~\[11711] )),
  \[4209]  = ~v6 & (~v5 & ~\[12995] ),
  \[21823]  = ~\[7552]  | (~\[7557]  | ~\[7569] ),
  \[11579]  = ~v1 | (~\[10099]  | ~v3),
  \[12041]  = ~v5 | (~\[10134]  | ~v6),
  \[3743]  = ~v6 & (~v5 & (~\[13227]  & ~v3)),
  \[21825]  = ~v13 | (~\[10073]  | (~\[7537]  | ~\[7547] )),
  \[13969]  = ~v10 | ~v9,
  \[11576]  = ~\[21877]  | (~\[21875]  | (~\[21873]  | ~\[21871] )),
  \[21497]  = ~v0 | (~\[10060]  | (~v8 | ~\[9958] )),
  \[13963]  = ~\[22365]  | (~\[22363]  | (~\[22361]  | ~\[22359] )),
  \[5405]  = ~\[10133]  & (~v5 & ~v8),
  \[14093]  = ~v4 | (~v7 | ~\[10058] ),
  \[10387]  = ~v1 | (~\[10099]  | ~v2),
  \[3018]  = ~\[10072]  & (~v14 & (~\[13587]  & ~v12)),
  \[6995]  = ~v6 & ~v5,
  \[14096]  = ~v10 | (~v9 | ~\[10068] ),
  \[21499]  = ~v11 | (~v9 | ~\[9955] ),
  \[13235]  = ~v0 | ~v2,
  \[21831]  = ~v13 | (~\[10073]  | (~\[7483]  | ~\[7493] )),
  \[2551]  = ~\[10058]  & (~v10 & ~v12),
  \[6267]  = ~v6 & (~v5 & (~\[11967]  & ~v2)),
  \[21493]  = ~\[10073]  | (~\[10072]  | (~v0 | ~\[10060] )),
  \[11581]  = ~v5 | (~\[10134]  | ~v6),
  \[8657]  = ~\[10133]  & (~v5 & (~\[10777]  & ~v3)),
  \[13972]  = ~v13 | (~\[10088]  | ~v15),
  \[12779]  = ~v8 | (~\[10133]  | ~v11),
  \[10383]  = ~v2 | (~\[10176]  | (~v1 | ~\[10099] )),
  \[11914]  = ~v4 | ~v7,
  \[21495]  = ~v15 | (~\[10072]  | (~v0 | ~\[10060] )),
  \[223]  = ~\[11762]  & (~v2 & (~\[11765]  & ~\[11771] )),
  \[4944]  = ~\[10073]  & (~v13 & (~v15 & ~\[12628] )),
  \[224]  = ~\[11775]  & (~\[11773]  & ~\[11781] ),
  \[954]  = ~\[282]  & (~\[281]  & (~\[280]  & ~\[279] )),
  \[12776]  = ~v5 | (~\[10134]  | ~v6),
  \[225]  = ~v6 & (~v5 & (~\[11755]  & ~\[11761] )),
  \[10728]  = ~\[21697]  | (~\[21695]  | (~\[21693]  | ~\[21691] )),
  \[1361]  = ~\[10449]  & (~\[10416]  & ~\[10514] ),
  \[4217]  = ~\[10058]  & (~v10 & ~v12),
  \[12050]  = ~v4 | ~\[10135] ,
  \[11587]  = ~v8 | (~\[10133]  | (~v11 | ~\[7024] )),
  \[13248]  = ~v5 | (~\[10134]  | ~v6),
  \[3751]  = ~v10 & (~v9 & ~v12),
  \[13978]  = ~v1 | (~\[10099]  | (~v3 | ~\[2259] )),
  \[6607]  = ~\[10059]  & (~v0 & (~v2 & ~\[11796] )),
  \[4949]  = ~\[10133]  & (~v5 & ~v8),
  \[11921]  = ~\[21949]  | (~\[21947]  | ~\[21951] ),
  \[10724]  = ~v8 | (~\[10064]  | ~v12),
  \[6272]  = ~\[10073]  & (~v13 & ~v15),
  \[13979]  = ~v10 | ~v9,
  \[13244]  = ~\[22215]  | (~\[22213]  | (~\[22211]  | ~\[22209] )),
  \[3026]  = ~\[10059]  & (~v0 & ~v2),
  \[7803]  = ~v9 & (~v7 & ~v10),
  \[22307]  = ~v7 | (~\[10236]  | (~\[2856]  | ~\[2848] )),
  \[13245]  = ~v2 | ~\[10059] ,
  \[2561]  = ~\[10134]  & (~v6 & (~\[13826]  & ~v3)),
  \[6276]  = ~v9 & ~v7,
  \[22309]  = ~v13 | (~\[10073]  | (~\[2829]  | ~\[2839] )),
  \[11591]  = ~v1 | (~\[10099]  | (~\[10060]  | ~\[7013] )),
  \v16.0  = \[0] ,
  \[13982]  = ~v13 | (~\[10088]  | ~v15),
  \[12789]  = ~v5 | (~\[10134]  | ~v6),
  \[11924]  = ~\[1083]  | (~\[1090]  | (~\[1076]  | ~\[1063] )),
  \[12784]  = ~\[22117]  | (~\[22115]  | (~\[22113]  | ~\[22111] )),
  \[9130]  = ~\[10060]  & (~v1 & ~v3),
  \[4954]  = ~\[10059]  & (~v0 & ~v2),
  \[12056]  = ~v0 | ~v2,
  \[9861]  = ~v12 & (~v7 & (~\[10135]  & ~\[10134] )),
  \[10738]  = ~v2 | ~\[10059] ,
  \[7474]  = ~\[10059]  & (~v0 & ~v2),
  \[10007]  = ~v2 & (~v1 & ~v12),
  \[6615]  = ~\[10058]  & (~v10 & ~v13),
  \[11930]  = ~v4 | ~v7,
  \[21849]  = ~v7 | (~\[10236]  | (~\[7322]  | ~\[7314] )),
  \[2569]  = ~\[10058]  & (~v10 & ~v12),
  \[22311]  = ~v4 | (~v7 | (~\[2820]  | ~\[2812] )),
  \[3761]  = ~\[10133]  & (~v5 & ~\[13219] ),
  \[11202]  = ~v5 | (~\[10134]  | ~v6),
  \[2902]  = ~\[10072]  & (~v12 & ~v14),
  \[13988]  = ~v1 | (~\[10099]  | (~\[10060]  | ~\[2237] )),
  \[1374]  = ~\[74]  & (~\[73]  & (~\[75]  & ~\[10376] )),
  \[12792]  = ~v8 | (~\[10133]  | ~v11),
  \[10733]  = ~v0 | (~v2 | (~\[10176]  | ~\[8731] )),
  \[13989]  = ~v10 | ~v9,
  \[11593]  = ~v11 | (~v8 | ~\[10072] ),
  \[13254]  = ~v13 | (~\[10088]  | (~v15 | ~\[3659] )),
  \[3036]  = ~\[10072]  & (~v14 & (~\[13579]  & ~v12)),
  \[10735]  = ~v8 | (~\[10064]  | ~v12),
  \[9869]  = ~\[10135]  & (~\[10134]  & ~v7),
  \[1710]  = ~\[10072]  & (~v12 & (~v14 & ~\[14241] )),
  \[22317]  = ~\[2750]  | (~\[2755]  | ~\[2767] ),
  \[13256]  = ~v2 | (~\[10059]  | ~\[10176] ),
  \[11208]  = ~v13 | (~\[10088]  | (~\[10073]  | ~\[7803] )),
  \[11938]  = ~v4 | ~v7,
  \[21851]  = ~v7 | (~\[10236]  | (~\[7304]  | ~\[7296] )),
  \[12068]  = ~v0 | ~v2,
  \[8674]  = ~\[10060]  & (~v1 & ~v3),
  \[12400]  = ~v12 | (~v14 | ~\[10076] ),
  \[22319]  = ~\[2728]  | (~\[2733]  | ~\[2745] ),
  \[5427]  = ~\[10134]  & (~v6 & ~v8),
  \[10741]  = ~v5 | (~\[10134]  | ~v6),
  \[22313]  = ~v4 | (~v7 | (~\[2802]  | ~\[2794] )),
  \[971]  = ~\[12282]  & (~\[12243]  & ~\[12359] ),
  \[13262]  = ~v15 | (~v13 | ~\[3697] ),
  \[6289]  = ~\[10059]  & (~v0 & (~\[10176]  & ~\[11958] )),
  \[13992]  = ~v13 | (~\[10088]  | ~v15),
  \[22315]  = ~v13 | (~\[10073]  | (~\[2775]  | ~\[2785] )),
  \[5094]  = ~v4 & (~v2 & (~\[10059]  & ~v0)),
  \[7483]  = ~v10 & (~v9 & ~v12),
  \[12796]  = ~v1 | ~\[10099] ,
  \[12065]  = ~\[21979]  | (~\[21977]  | ~\[21981] ),
  \[1381]  = ~\[68]  & (~\[67]  & (~\[66]  & ~\[65] )),
  \[11210]  = ~v1 | (~\[10099]  | ~v3),
  \[6625]  = ~v6 & (~v5 & ~\[11787] ),
  \[4237]  = ~\[10058]  & (~v7 & ~v10),
  \[10747]  = ~v12 | (~v14 | (~\[10076]  | ~\[8707] )),
  \[9143]  = ~v6 & ~v5,
  \[3770]  = ~v10 & (~v9 & (~v12 & ~\[13216] )),
  \[2579]  = ~\[10060]  & (~v1 & (~v3 & ~\[13820] )),
  \[12408]  = ~v1 | (~\[10099]  | (~v3 | ~\[5383] )),
  \[22321]  = ~v13 | (~\[10073]  | (~\[2713]  | ~\[2723] )),
  \[11212]  = ~v5 | (~\[10134]  | ~v6),
  \[13998]  = ~\[634]  | (~\[641]  | (~\[627]  | ~\[672] )),
  \[10749]  = ~v0 | ~v2,
  \[21853]  = ~v14 | (~\[10076]  | (~\[7277]  | ~\[7287] )),
  \[12071]  = ~v5 | (~\[10134]  | ~v6),
  \[12409]  = ~v10 | ~v9,
  \[3044]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[21855]  = ~v14 | (~\[10076]  | (~\[7259]  | ~\[7269] )),
  \[13264]  = ~v0 | (~v2 | ~\[10176] ),
  \[1388]  = ~\[64]  & (~\[63]  & (~\[62]  & ~\[61] )),
  \[6294]  = ~\[10073]  & (~v13 & ~v15),
  \[7823]  = ~v10 & (~v9 & ~v12),
  \[22327]  = ~v13 | (~\[10073]  | (~\[2659]  | ~\[2669] )),
  \[11218]  = ~v13 | (~\[10088]  | (~\[10073]  | ~\[7781] )),
  \[2918]  = ~\[10060]  & (~v1 & ~v3),
  \[1721]  = ~v6 & (~v5 & (~v8 & ~\[14236] )),
  \[11948]  = ~v5 | (~\[10134]  | ~v6),
  \[3778]  = ~\[10059]  & (~v0 & ~v2),
  \[22329]  = ~v13 | (~\[10073]  | (~\[2641]  | ~\[2651] )),
  \[10752]  = ~v5 | (~\[10134]  | ~v6),
  \[13270]  = ~v15 | (~v13 | ~\[3679] ),
  \[12077]  = ~v14 | (~\[10072]  | (~\[10076]  | ~\[6053] )),
  \[8685]  = ~\[10058]  & (~v7 & ~v10),
  \[10021]  = ~v2 & (~v1 & ~v8),
  \[4971]  = ~\[10134]  & (~v6 & ~v8),
  \[12412]  = ~v12 | (~v14 | ~\[10076] ),
  \[6298]  = ~v9 & ~v7,
  \[22323]  = ~v13 | (~\[10073]  | (~\[2695]  | ~\[2705] )),
  \[12079]  = ~v2 | (~\[10059]  | ~\[10176] ),
  \[22325]  = ~v13 | (~\[10073]  | (~\[2677]  | ~\[2687] )),
  \[6633]  = ~\[10058]  & (~v10 & ~v13),
  \[21867]  = ~v14 | (~\[10076]  | (~\[7143]  | ~\[7153] )),
  \[2587]  = ~\[10058]  & (~v10 & ~v12),
  \[7493]  = ~\[10099]  & (~\[10060]  & (~v3 & ~\[11335] )),
  \[10028]  = ~v2 & ~v1,
  \[10758]  = ~v12 | (~v14 | (~\[10076]  | ~\[8685] )),
  \[985]  = ~\[269]  & (~\[268]  & (~\[270]  & ~\[12179] )),
  \[256]  = ~\[12068]  & (~v3 & (~\[12071]  & ~\[12077] )),
  \[21869]  = ~v4 | (~v7 | (~\[7134]  | ~\[7126] )),
  \[13605]  = ~v11 | ~v8,
  \[12418]  = ~v2 | (~\[10059]  | (~\[10176]  | ~\[5361] )),
  \[257]  = ~\[10133]  & (~v5 & (~\[12079]  & ~\[12085] )),
  \[22331]  = ~v13 | (~\[10073]  | (~\[2623]  | ~\[2633] )),
  \[13610]  = ~v0 | ~v2,
  \[258]  = ~\[10133]  & (~v5 & (~\[12088]  & ~\[12094] )),
  \[21863]  = ~\[7180]  | (~v11 | (~\[7176]  | ~\[7193] )),
  \[259]  = ~\[10072]  & (~v14 & (~\[12100]  & ~\[12098] )),
  \[12419]  = ~v10 | ~v9,
  \[3054]  = ~\[10072]  & (~v14 & (~\[13570]  & ~v12)),
  \[21865]  = ~v7 | (~\[10236]  | (~\[7170]  | ~\[7162] )),
  \[7833]  = ~\[10059]  & (~v0 & (~\[10176]  & ~\[11183] )),
  \[22337]  = ~v13 | (~\[10073]  | (~\[2569]  | ~\[2579] )),
  \[3787]  = ~v10 & (~v9 & ~v12),
  \[11958]  = ~v5 | (~\[10134]  | ~v6),
  \[21871]  = ~v4 | (~v7 | (~\[7116]  | ~\[7108] )),
  \[12088]  = ~v0 | (~v2 | ~\[10176] ),
  \[1732]  = ~\[10072]  & (~v12 & (~v14 & ~\[14230] )),
  \[22339]  = ~v13 | (~\[10073]  | (~\[2551]  | ~\[2561] )),
  \[10762]  = ~v7 | (~\[10236]  | ~\[8674] ),
  \[260]  = ~\[10073]  & (~v15 & (~\[12110]  & ~\[12108] )),
  \[12422]  = ~v12 | (~v14 | ~\[10076] ),
  \[261]  = ~\[10073]  & (~v15 & (~\[12118]  & ~\[12116] )),
  \[22333]  = ~v13 | (~\[10073]  | (~\[2605]  | ~\[2615] )),
  \[5449]  = ~\[10134]  & (~v6 & ~v8),
  \[7108]  = ~\[10073]  & (~v15 & ~\[11545] ),
  \[11224]  = ~v1 | (~\[10099]  | ~v3),
  \[262]  = ~\[10072]  & (~v14 & (~\[12127]  & ~\[12125] )),
  \[992]  = ~\[263]  & (~\[262]  & (~\[261]  & ~\[260] )),
  \[263]  = ~\[12130]  & (~v2 & (~\[12133]  & ~\[12139] )),
  \[22335]  = ~v13 | (~\[10073]  | (~\[2587]  | ~\[2597] )),
  \[1737]  = ~v6 & (~v5 & ~v8),
  \[9161]  = ~v6 & ~v5,
  \[21877]  = ~\[7052]  | ~\[7063] ,
  \[2597]  = ~v6 & (~v5 & (~\[13798]  & ~v3)),
  \[12085]  = ~v14 | (~\[10076]  | ~\[6033] ),
  \[2931]  = ~\[10134]  & ~v6,
  \[22341]  = ~\[2526]  | (~\[2531]  | ~\[2543] ),
  \[268]  = ~\[10134]  & (~v6 & (~\[12189]  & ~\[12195] )),
  \[4259]  = ~\[10058]  & (~v7 & ~v10),
  \[3062]  = ~\[10059]  & (~v0 & ~v2),
  \[21873]  = ~v4 | (~v7 | (~\[7098]  | ~\[7090] )),
  \[269]  = ~\[10133]  & (~v5 & (~\[12197]  & ~\[12203] )),
  \[10764]  = ~v8 | (~\[10064]  | ~v12),
  \[999]  = ~\[259]  & (~\[258]  & (~\[257]  & ~\[256] )),
  \[13622]  = ~v11 | ~v8,
  \[12429]  = ~v0 | (~v2 | (~\[10176]  | ~\[5339] )),
  \[21875]  = ~v4 | (~v7 | (~\[7080]  | ~\[7072] )),
  \[7841]  = ~v10 & (~v9 & ~v13),
  \[604]  = ~\[458]  & (~\[457]  & (~\[456]  & ~\[455] )),
  \[13283]  = ~v13 | (~\[10088]  | ~v15),
  \[12098]  = ~v4 | (~v7 | ~\[6006] ),
  \[12430]  = ~v10 | ~v9,
  \[1742]  = ~\[10060]  & (~v1 & ~v3),
  \[11967]  = ~v1 | ~\[10099] ,
  \[7116]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[270]  = ~\[10133]  & (~v5 & (~\[12181]  & ~\[12187] )),
  \[3402]  = ~\[10059]  & (~v0 & ~v2),
  \[13627]  = ~\[22297]  | (~\[22295]  | (~\[22293]  | ~\[22291] )),
  \[13291]  = ~v15 | ~v13,
  \[4993]  = ~\[10134]  & (~v6 & ~v8),
  \[8310]  = ~v9 & (~v7 & (~v10 & ~\[10948] )),
  \[12094]  = ~v14 | (~\[10076]  | ~\[6015] ),
  \[11233]  = ~v4 | ~\[10135] ,
  \[6653]  = ~\[10058]  & (~v7 & ~v10),
  \[11966]  = ~\[21959]  | (~\[21957]  | (~\[21955]  | ~\[21953] )),
  \[21887]  = ~v4 | (~\[10135]  | (~\[6964]  | ~\[6956] )),
  \[10777]  = ~v0 | ~v2,
  \[21889]  = ~v7 | (~\[10236]  | (~\[6946]  | ~\[6938] )),
  \[8314]  = ~\[10236]  & ~v4,
  \[3071]  = ~\[10068]  & (~\[10058]  & ~v12),
  \[10049]  = ~v2 & (~v1 & ~v9),
  \[11241]  = ~v1 | (~\[10099]  | ~v3),
  \[279]  = ~\[10072]  & (~v14 & (~\[12289]  & ~\[12287] )),
  \[611]  = ~\[454]  & (~\[453]  & (~\[452]  & ~\[451] )),
  \[10774]  = ~v8 | (~\[10064]  | ~v12),
  \[9176]  = ~\[10073]  & (~v15 & ~\[10493] ),
  \[13632]  = ~v0 | (~v2 | (~\[10176]  | ~\[2931] )),
  \[12439]  = ~v2 | (~\[10059]  | (~\[10176]  | ~\[5317] )),
  \[4603]  = ~v6 & (~v5 & (~\[12796]  & ~v2)),
  \[2215]  = ~\[10133]  & (~v5 & ~v8),
  \[7851]  = ~\[10099]  & (~\[10060]  & (~v3 & ~\[11175] )),
  \[13294]  = ~v0 | ~v2,
  \[12433]  = ~v12 | (~v14 | ~\[10076] ),
  \[2946]  = ~\[10072]  & (~v14 & (~\[13622]  & ~v12)),
  \[21891]  = ~v7 | (~\[10236]  | (~\[6928]  | ~\[6920] )),
  \[12440]  = ~v10 | ~v9,
  \[22359]  = ~\[2335]  | (~v15 | (~\[2343]  | ~\[2357] )),
  \[3411]  = ~\[10068]  & (~v9 & ~v12),
  \[7126]  = ~\[10073]  & (~v15 & ~\[11535] ),
  \[280]  = ~\[10072]  & (~v14 & (~\[12297]  & ~\[12295] )),
  \[1754]  = ~\[10072]  & (~v12 & (~v14 & ~\[14220] )),
  \[281]  = ~\[12306]  & (~v11 & (~\[12309]  & ~\[12305] )),
  \[282]  = ~\[12316]  & (~v11 & (~\[12319]  & ~\[12315] )),
  \[8320]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[7859]  = ~v10 & (~v9 & ~v13),
  \[13634]  = ~v11 | (~v8 | ~\[10088] ),
  \[11976]  = ~v1 | (~\[10099]  | ~v3),
  \[10058]  = ~v8,
  \[11250]  = ~v7 | ~\[10236] ,
  \[10057]  = ~v2 & (~v1 & ~v8),
  \[1759]  = ~\[10133]  & (~v5 & ~v8),
  \[286]  = ~\[12366]  & (~v11 & (~\[12369]  & ~\[12365] )),
  \[10787]  = ~v4 | ~v7,
  \[21501]  = ~v12 | (~v15 | (~v0 | ~\[10060] )),
  \[287]  = ~\[12376]  & (~v11 & (~\[12379]  & ~\[12375] )),
  \[22361]  = ~\[2325]  | (~\[2330]  | ~\[2320] ),
  \[3081]  = ~v6 & (~v5 & ~\[13559] ),
  \[9184]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[10059]  = ~v1,
  \[288]  = ~\[12387]  & (~v11 & (~\[12390]  & ~\[12386] )),
  \[289]  = ~\[12397]  & (~v11 & (~\[12400]  & ~\[12396] )),
  \[5471]  = ~v6 & (~v5 & ~v8),
  \[5809]  = ~\[10068]  & (~v9 & ~v12),
  \[12449]  = ~v0 | (~v2 | ~\[10176] ),
  \[2954]  = ~\[10060]  & (~v1 & ~v3),
  \[13641]  = ~v5 | (~\[10134]  | (~v6 | ~\[2918] )),
  \[4614]  = ~\[10072]  & (~v12 & (~\[10076]  & ~\[12792] )),
  \[12443]  = ~v12 | (~v14 | ~\[10076] ),
  \[1030]  = ~\[12065]  & (~\[12037]  & (~\[12001]  & ~\[11966] )),
  \[10060]  = ~v2,
  \[14103]  = ~v4 | (~v7 | ~\[10058] ),
  \[7134]  = ~\[10060]  & (~v1 & ~v3),
  \[14106]  = ~v10 | (~v9 | ~\[10068] ),
  \[11257]  = ~\[21809]  | (~\[21807]  | (~\[21805]  | ~\[21803] )),
  \[4280]  = ~\[10058]  & (~v10 & (~v12 & ~\[12958] )),
  \[627]  = ~\[449]  & (~\[448]  & (~\[450]  & ~\[13963] )),
  \[3421]  = ~\[10134]  & (~v6 & ~\[13396] ),
  \[1033]  = ~\[13132]  & (~\[12851]  & (~\[12529]  & ~\[12208] )),
  \[13648]  = ~v0 | ~v2,
  \[1763]  = ~\[10059]  & ~v0,
  \[290]  = ~\[12409]  & (~v11 & (~\[12412]  & ~\[12408] )),
  \[11259]  = ~v1 | (~\[10099]  | ~v3),
  \[291]  = ~\[12419]  & (~v11 & (~\[12422]  & ~\[12418] )),
  \[22363]  = ~\[2307]  | (~v3 | (~\[2303]  | ~\[2298] )),
  \[292]  = ~\[12430]  & (~v11 & (~\[12433]  & ~\[12429] )),
  \[7869]  = ~\[10060]  & (~v1 & (~v3 & ~\[11166] )),
  \[293]  = ~\[12440]  & (~v11 & (~\[12443]  & ~\[12439] )),
  \[22365]  = ~\[2281]  | (~\[2286]  | ~\[2276] ),
  \[8331]  = ~v9 & (~v7 & ~v10),
  \[11986]  = ~v4 | ~\[10135] ,
  \[10068]  = ~v11,
  \[13646]  = ~v8 | (~\[10133]  | (~v11 | ~\[2902] )),
  \[6675]  = ~\[10058]  & (~v7 & ~v10),
  \[10797]  = ~\[1322]  | (~\[1329]  | (~\[1315]  | ~\[1302] )),
  \[4288]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[9194]  = ~\[10073]  & (~v15 & ~\[10509] ),
  \[298]  = ~\[12510]  & (~v11 & (~\[12513]  & ~\[12509] )),
  \[2963]  = ~\[10068]  & (~\[10058]  & ~v12),
  \[10064]  = ~v10,
  \[299]  = ~\[12520]  & (~v11 & (~\[12523]  & ~\[12519] )),
  \[3093]  = ~v6 & ~v5,
  \[14117]  = ~v10 | (~v9 | ~\[10068] ),
  \[10063]  = ~v9,
  \[13651]  = ~v5 | (~\[10134]  | ~v6),
  \[12454]  = ~v10 | (~v9 | ~\[10068] ),
  \[634]  = ~\[443]  & (~\[442]  & (~\[441]  & ~\[440] )),
  \[10795]  = ~\[21709]  | (~\[21707]  | (~\[21711]  | ~\[1285] )),
  \[14114]  = ~v4 | (~v7 | ~\[10058] ),
  \[4625]  = ~\[10059]  & (~v0 & (~\[10176]  & ~\[12789] )),
  \[2237]  = ~\[10133]  & (~v5 & ~v8),
  \[7143]  = ~\[10068]  & (~v9 & ~\[10088] ),
  \[11600]  = ~v1 | (~\[10099]  | (~v3 | ~\[6995] )),
  \[21519]  = ~v12 | (~v15 | ~\[9869] ),
  \[3430]  = ~\[10068]  & (~v9 & (~v12 & ~\[13383] )),
  \[10072]  = ~v13,
  \[11602]  = ~v11 | (~v8 | ~\[10072] ),
  \[5488]  = ~\[10088]  & (~\[10073]  & (~v15 & ~\[12329] )),
  \[13657]  = ~v8 | (~\[10133]  | (~v11 | ~\[2880] )),
  \[7877]  = ~v10 & (~v9 & ~v12),
  \[1776]  = ~\[10072]  & (~v12 & (~v14 & ~\[14208] )),
  \[11993]  = ~v1 | (~\[10099]  | ~v3),
  \[11266]  = ~v2 | ~\[10059] ,
  \[11608]  = ~v4 | (~\[10135]  | ~\[6982] ),
  \[21521]  = ~v14 | (~v13 | (~\[10076]  | ~\[9861] )),
  \[3438]  = ~\[10059]  & (~v0 & ~v2),
  \[4298]  = ~\[10076]  & (~\[10072]  & (~\[12948]  & ~v12)),
  \[5827]  = ~\[10068]  & (~v9 & ~v12),
  \[10079]  = ~\[21477]  | (~\[21475]  | (~\[21473]  | ~\[21471] )),
  \[2973]  = ~v6 & (~v5 & (~\[13610]  & ~v3)),
  \[641]  = ~\[439]  & (~\[438]  & (~\[437]  & ~\[436] )),
  \[14127]  = ~v10 | (~v9 | ~\[10068] ),
  \[10073]  = ~v14,
  \[13661]  = ~v7 | (~\[10236]  | ~\[2874] ),
  \[10076]  = ~v15,
  \[5493]  = ~v6 & (~v5 & ~v8),
  \[14124]  = ~v4 | (~v7 | ~\[10058] ),
  \[7153]  = ~\[10133]  & (~v5 & (~\[11522]  & ~v3)),
  \[12466]  = ~v10 | (~\[10068]  | (~v9 | ~\[10058] )),
  \[4636]  = ~\[10072]  & (~v12 & (~\[10076]  & ~\[12779] )),
  \[1781]  = ~\[10133]  & (~v5 & ~v8),
  \[11610]  = ~v11 | (~v8 | ~\[10072] ),
  \[22389]  = ~\[2004]  | ~\[2015] ,
  \[5100]  = ~\[10073]  & (~v13 & ~v15),
  \[5498]  = ~\[10059]  & (~v0 & ~v2),
  \[21523]  = ~v6 | (~v4 | (~\[10133]  | ~\[9844] )),
  \[7887]  = ~\[10059]  & (~v0 & (~v2 & ~\[11158] )),
  \[14132]  = ~\[22395]  | (~\[22393]  | (~\[22391]  | ~\[22389] )),
  \[21525]  = ~v9 | (~\[10064]  | ~\[9841] ),
  \[8350]  = ~v10 & ~v9,
  \[1786]  = ~\[10059]  & (~v0 & ~v2),
  \[10416]  = ~\[21629]  | (~\[21627]  | (~\[21625]  | ~\[21623] )),
  \[13663]  = ~v11 | (~v8 | ~\[10088] ),
  \[11275]  = ~v0 | ~v2,
  \[10088]  = ~v12,
  \[12806]  = ~v1 | (~\[10099]  | ~v3),
  \[3447]  = ~\[10068]  & (~v9 & ~v12),
  \[6695]  = ~\[10058]  & (~v10 & ~v13),
  \[22391]  = ~\[1982]  | ~\[1993] ,
  \[2982]  = ~\[10072]  & (~v14 & (~\[13605]  & ~v12)),
  \[14138]  = ~v10 | ~v9,
  \[11619]  = ~v11 | ~v8,
  \[14137]  = ~v1 | (~\[10099]  | (~\[10060]  | ~\[1869] )),
  \[13672]  = ~v11 | ~v8,
  \[12479]  = ~v10 | (~\[10068]  | (~v9 | ~\[10058] )),
  \[7162]  = ~\[10073]  & (~v15 & ~\[11518] ),
  \[16]  = ~\[10099]  & (~v2 & (~v12 & ~\[10129] )),
  \[17]  = ~\[10088]  & (~v14 & (~\[10099]  & ~v2)),
  \[18]  = ~\[10063]  & (~v8 & (~v10 & ~\[10137] )),
  \[4647]  = ~\[10059]  & (~v0 & (~v2 & ~\[12776] )),
  \[2259]  = ~\[10134]  & (~v6 & ~v8),
  \[22001]  = ~v13 | (~\[10073]  | (~\[5881]  | ~\[5891] )),
  \[7895]  = ~v10 & (~v9 & ~v13),
  \[19]  = ~\[10064]  & (~v9 & (~v11 & ~\[10141] )),
  \[1063]  = ~\[11921]  & (~\[11895]  & (~\[11855]  & ~\[11820] )),
  \[12817]  = ~v11 | ~v8,
  \[22393]  = ~\[1960]  | ~\[1971] ,
  \[7501]  = ~v10 & (~v9 & ~v12),
  \[10426]  = ~v11 | (~v8 | ~v12),
  \[22395]  = ~\[1938]  | ~\[1949] ,
  \[14141]  = ~v13 | (~\[10088]  | ~\[10073] ),
  \[11285]  = ~v4 | ~\[10135] ,
  \[1798]  = ~\[10072]  & (~v12 & (~v14 & ~\[14198] )),
  \[5845]  = ~\[10068]  & (~v9 & ~v12),
  \[3457]  = ~v6 & (~v5 & ~\[13370] ),
  \[2990]  = ~\[10060]  & (~v1 & ~v3),
  \[20]  = ~v14 & (~v13 & (~\[10146]  & ~v7)),
  \[11627]  = ~v11 | ~v8,
  \[21]  = ~\[10076]  & (~v13 & (~\[10149]  & ~v7)),
  \[13680]  = ~v11 | ~v8,
  \[11292]  = ~\[21817]  | (~\[21815]  | (~\[21813]  | ~\[21811] )),
  \[10099]  = ~v0,
  \[22]  = ~\[10064]  & (~\[10058]  & (~v11 & ~\[10154] )),
  \[14148]  = ~v5 | (~v6 | (~\[10133]  | ~\[1926] )),
  \[1404]  = ~\[57]  & (~\[56]  & (~\[55]  & ~\[54] )),
  \[22003]  = ~v13 | (~\[10073]  | (~\[5863]  | ~\[5873] )),
  \[12822]  = ~\[22125]  | (~\[22123]  | (~\[22121]  | ~\[22119] )),
  \[23]  = ~\[10063]  & (~v8 & (~\[10068]  & ~\[10158] )),
  \[7170]  = ~\[10060]  & (~v1 & ~v3),
  \[12489]  = ~v10 | (~v9 | ~\[10068] ),
  \[6311]  = ~\[10059]  & (~v0 & (~v2 & ~\[11948] )),
  \[8368]  = ~v10 & ~v9,
  \[22005]  = ~v13 | (~\[10073]  | (~\[5845]  | ~\[5855] )),
  \[10095]  = ~\[21485]  | (~\[21483]  | (~\[21481]  | ~\[21479] )),
  \[4656]  = ~\[10076]  & (~\[10072]  & (~\[12769]  & ~v12)),
  \[28]  = ~\[10176]  & (~v1 & (~v9 & ~\[10186] )),
  \[21549]  = ~v15 | (~\[10072]  | (~v3 | ~v0)),
  \[29]  = ~v14 & (~v13 & (~\[10176]  & ~v1)),
  \[7176]  = ~\[10088]  & (~\[10073]  & ~v15),
  \[8707]  = ~\[10058]  & (~v7 & ~v10),
  \[11294]  = ~v0 | ~v2,
  \[6319]  = ~\[10068]  & (~v9 & ~v13),
  \[14152]  = ~v13 | ~\[10088] ,
  \[1076]  = ~\[224]  & (~\[223]  & (~\[225]  & ~\[11753] )),
  \[2605]  = ~\[10058]  & (~v10 & ~v12),
  \[7511]  = ~\[10060]  & (~v1 & (~v3 & ~\[11351] )),
  \[12824]  = ~v1 | (~\[10099]  | ~v3),
  \[14151]  = ~v10 | (~\[10068]  | (~v9 | ~\[10058] )),
  \[3465]  = ~\[10068]  & (~v9 & ~v12),
  \[10435]  = ~v11 | (~v8 | ~v12),
  \[9569]  = ~\[10236]  & (~v4 & ~v6),
  \[22017]  = ~v13 | (~\[10073]  | (~\[5737]  | ~\[5747] )),
  \[5855]  = ~\[10059]  & (~v0 & (~v2 & ~\[12172] )),
  \[13686]  = ~v4 | ~v7,
  \[30]  = ~\[10076]  & (~v13 & (~\[10176]  & ~v1)),
  \[21551]  = ~v3 | (~v0 | (~v8 | ~\[9742] )),
  \[12100]  = ~v11 | (~\[10063]  | ~\[10088] ),
  \[22019]  = ~v13 | (~\[10073]  | (~\[5719]  | ~\[5729] )),
  \[31]  = ~\[10064]  & (~v11 & ~\[10195] ),
  \[10441]  = ~v5 | (~\[10134]  | ~v6),
  \[32]  = ~\[10176]  & (~v1 & (~v8 & ~\[10199] )),
  \[14158]  = ~v5 | ~v6,
  \[22013]  = ~v13 | (~\[10073]  | (~\[5773]  | ~\[5783] )),
  \[12832]  = ~v1 | (~\[10099]  | ~v3),
  \[33]  = ~\[10088]  & (~\[10076]  & (~\[10176]  & ~v1)),
  \[14157]  = ~v3 | (~\[10134]  | (~v1 | ~\[10099] )),
  \[7180]  = ~v9 & ~v7,
  \[12499]  = ~v4 | (~v7 | (~\[10058]  | ~\[5160] )),
  \[34]  = ~\[10176]  & (~v1 & (~v12 & ~\[10206] )),
  \[672]  = ~\[13835]  & (~\[13807]  & (~\[13771]  & ~\[13736] )),
  \[12494]  = ~\[22065]  | (~\[22063]  | (~\[22061]  | ~\[22059] )),
  \[7519]  = ~v10 & (~v9 & ~v12),
  \[22015]  = ~v13 | (~\[10073]  | (~\[5755]  | ~\[5765] )),
  \[35]  = ~\[10088]  & (~v14 & (~\[10176]  & ~v1)),
  \[4664]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[2276]  = ~\[10072]  & (~v12 & (~\[10076]  & ~\[13958] )),
  \[3805]  = ~v10 & (~v9 & ~v12),
  \[36]  = ~\[10063]  & (~v10 & (~\[10211]  & ~v8)),
  \[11635]  = ~v11 | ~v8,
  \[37]  = ~\[10064]  & (~v11 & (~\[10215]  & ~v9)),
  \[38]  = ~v14 & (~v13 & (~\[10176]  & ~\[10099] )),
  \[12108]  = ~v4 | (~v7 | ~\[5988] ),
  \[22021]  = ~\[5698]  | (~v11 | (~\[5694]  | ~\[5711] )),
  \[1083]  = ~\[218]  & (~\[217]  & (~\[216]  & ~\[215] )),
  \[10449]  = ~\[21637]  | (~\[21635]  | (~\[21633]  | ~\[21631] )),
  \[21553]  = ~v11 | (~v9 | ~\[9739] ),
  \[11641]  = ~\[21889]  | (~\[21887]  | (~\[21891]  | ~\[1105] )),
  \[10444]  = ~v8 | (~\[10133]  | ~v11),
  \[6329]  = ~\[10059]  & (~v0 & (~\[10176]  & ~\[11938] )),
  \[21555]  = ~v12 | (~v15 | (~v3 | ~v0)),
  \[2615]  = ~v6 & (~v5 & (~\[13790]  & ~v3)),
  \[5863]  = ~\[10068]  & (~v9 & ~v12),
  \[3475]  = ~v6 & (~v5 & (~\[13360]  & ~v2)),
  \[13694]  = ~\[22309]  | (~\[22307]  | (~\[22311]  | ~\[686] )),
  \[9579]  = ~\[10236]  & (~v4 & ~v6),
  \[22027]  = ~v13 | (~\[10073]  | (~\[5639]  | ~\[5649] )),
  \[13696]  = ~\[723]  | (~\[730]  | (~\[716]  | ~\[703] )),
  \[1421]  = ~\[10285]  & (~\[10267]  & ~\[10317] ),
  \[2281]  = ~\[10134]  & (~v6 & ~v8),
  \[12110]  = ~v11 | (~\[10063]  | ~\[10072] ),
  \[11647]  = ~v2 | (~\[10059]  | (~\[10176]  | ~\[6905] )),
  \[10452]  = ~v1 | (~\[10099]  | ~v3),
  \[13308]  = ~v15 | ~v13,
  \[5138]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[22023]  = ~\[5676]  | (~v11 | (~\[5672]  | ~\[5689] )),
  \[11649]  = ~v11 | (~v8 | ~\[10072] ),
  \[43]  = ~\[10073]  & (~\[10072]  & (~v15 & ~\[10242] )),
  \[8387]  = ~v10 & (~v9 & ~\[10088] ),
  \[44]  = ~\[10088]  & (~v14 & (~\[10176]  & ~\[10099] )),
  \[7529]  = ~\[10133]  & (~v5 & (~\[11341]  & ~v3)),
  \[22025]  = ~v13 | (~\[10073]  | (~\[5657]  | ~\[5667] )),
  \[11643]  = ~\[1142]  | (~\[1149]  | (~\[1135]  | ~\[1122] )),
  \[45]  = ~\[10063]  & (~v8 & (~v10 & ~\[10238] )),
  \[4674]  = ~\[10076]  & (~\[10072]  & (~\[12760]  & ~v12)),
  \[2286]  = ~\[10059]  & (~v0 & ~v2),
  \[21567]  = ~v15 | (~\[10072]  | ~\[9681] ),
  \[1090]  = ~\[214]  & (~\[213]  & (~\[212]  & ~\[211] )),
  \[7193]  = ~\[10099]  & (~\[10060]  & (~v3 & ~\[11506] )),
  \[10457]  = ~v8 | (~\[10133]  | ~v11),
  \[686]  = ~\[417]  & (~\[416]  & (~\[415]  & ~\[414] )),
  \[14166]  = ~v13 | (~\[10088]  | (~\[10073]  | ~\[1887] )),
  \[21569]  = ~v10 | (~v8 | (~\[10068]  | ~\[9673] )),
  \[3480]  = ~\[10072]  & (~v12 & ~\[10076] ),
  \[12118]  = ~v11 | (~\[10063]  | ~\[10072] ),
  \[12848]  = ~\[22129]  | (~\[22127]  | ~\[22131] ),
  \[6337]  = ~\[10068]  & (~v9 & ~v13),
  \[10459]  = ~v12 | (~v14 | ~\[10076] ),
  \[21563]  = ~v10 | (~\[10063]  | (~\[10068]  | ~\[9699] )),
  \[2623]  = ~\[10058]  & (~v10 & ~v12),
  \[10454]  = ~v5 | (~\[10134]  | ~v6),
  \[21565]  = ~v6 | (~\[10236]  | (~\[10133]  | ~\[9684] )),
  \[3484]  = ~v9 & ~v7,
  \[13311]  = ~\[22229]  | (~\[22227]  | (~\[22225]  | ~\[22223] )),
  \[5873]  = ~v6 & (~v5 & ~\[12163] ),
  \[12843]  = ~v11 | ~v8,
  \[9589]  = ~\[10236]  & (~v4 & ~v6),
  \[12116]  = ~v4 | (~v7 | ~\[5970] ),
  \[22037]  = ~\[5543]  | (~\[5550]  | ~\[5538] ),
  \[21571]  = ~v9 | (~\[10058]  | (~v11 | ~\[9663] )),
  \[21909]  = ~v14 | (~\[10076]  | (~\[6749]  | ~\[6759] )),
  \[22039]  = ~\[5517]  | (~\[5524]  | ~\[5512] ),
  \[11657]  = ~v11 | (~v8 | ~\[10072] ),
  \[13318]  = ~v15 | ~v13,
  \[1434]  = ~\[44]  & (~\[43]  & (~\[45]  & ~\[10235] )),
  \[7537]  = ~v10 & (~v9 & ~v12),
  \[14177]  = ~v10 | (~v9 | ~\[10068] ),
  \[4682]  = ~\[10059]  & (~v0 & ~v2),
  \[8397]  = ~v6 & (~v5 & (~\[10900]  & ~v3)),
  \[3823]  = ~v10 & (~v9 & ~v12),
  \[12851]  = ~\[902]  | (~\[909]  | (~\[895]  | ~\[882] )),
  \[54]  = ~\[10063]  & (~v8 & (~v10 & ~\[10288] )),
  \[55]  = ~\[10064]  & (~v9 & (~v11 & ~\[10292] )),
  \[8731]  = ~\[10134]  & ~v6,
  \[56]  = ~v14 & (~v13 & (~\[10296]  & ~v6)),
  \[21577]  = ~v12 | (~\[10073]  | ~\[9633] ),
  \[11655]  = ~v0 | (~v2 | (~\[10176]  | ~\[6887] )),
  \[57]  = ~\[10076]  & (~v13 & (~\[10299]  & ~v6)),
  \[2298]  = ~\[10072]  & (~v12 & (~\[10076]  & ~\[13948] )),
  \[21911]  = ~v4 | (~v7 | (~\[6740]  | ~\[6732] )),
  \[22041]  = ~\[5493]  | (~\[5498]  | ~\[5488] ),
  \[12127]  = ~v11 | (~\[10063]  | ~\[10088] ),
  \[6347]  = ~\[10059]  & (~v0 & (~v2 & ~\[11930] )),
  \[300]  = ~\[12500]  & (~v11 & (~\[12503]  & ~\[12499] )),
  \[21573]  = ~v12 | (~v15 | ~\[9653] ),
  \[2633]  = ~\[10133]  & (~v5 & ~\[13782] ),
  \[301]  = ~\[12536]  & (~v11 & (~\[12539]  & ~\[12535] )),
  \[10464]  = ~v1 | (~\[10099]  | (~\[10060]  | ~\[9269] )),
  \[5881]  = ~\[10068]  & (~v9 & ~v12),
  \[12859]  = ~v15 | (~v13 | ~\[4485] ),
  \[302]  = ~\[12543]  & (~v8 & (~\[12542]  & ~\[12550] )),
  \[21575]  = ~v14 | (~v13 | (~\[10076]  | ~\[9645] )),
  \[303]  = ~\[12561]  & (~v15 & (~\[12560]  & ~\[12557] )),
  \[10466]  = ~v11 | (~v8 | ~v12),
  \[12853]  = ~v2 | (~\[10059]  | ~\[10176] ),
  \[304]  = ~\[12567]  & (~v7 & (~\[12566]  & ~\[12575] )),
  \[305]  = ~\[12583]  & (~v11 & (~\[12586]  & ~\[12582] )),
  \[9202]  = ~\[10059]  & (~v0 & ~v2),
  \[3497]  = ~\[10059]  & (~v0 & (~\[10176]  & ~\[13353] )),
  \[12125]  = ~v4 | (~v7 | (~\[5951]  | ~v3)),
  \[1441]  = ~\[38]  & (~\[37]  & (~\[36]  & ~\[35] )),
  \[306]  = ~\[12593]  & (~v11 & (~\[12596]  & ~\[12592] )),
  \[12130]  = ~v1 | ~\[10099] ,
  \[307]  = ~\[12604]  & (~v11 & (~\[12607]  & ~\[12603] )),
  \[61]  = ~\[10073]  & (~\[10072]  & (~v15 & ~\[10323] )),
  \[308]  = ~\[12614]  & (~v11 & (~\[12617]  & ~\[12613] )),
  \[62]  = ~\[10088]  & (~v14 & (~\[10326]  & ~v6)),
  \[10809]  = ~v1 | (~\[10099]  | ~v3),
  \[21913]  = ~v4 | (~v7 | (~\[6722]  | ~\[6714] )),
  \[7547]  = ~\[10060]  & (~v1 & (~v3 & ~\[11325] )),
  \[63]  = ~\[10063]  & (~v8 & (~v10 & ~\[10331] )),
  \[14187]  = ~v10 | (~v9 | ~\[10068] ),
  \[12861]  = ~v0 | (~v2 | ~\[10176] ),
  \[11664]  = ~v4 | (~\[10135]  | ~\[6874] ),
  \[64]  = ~\[10064]  & (~v9 & (~v11 & ~\[10335] )),
  \[3104]  = ~\[10072]  & (~v12 & ~v14),
  \[10803]  = ~v4 | (~v7 | ~\[8602] ),
  \[21915]  = ~v14 | (~\[10076]  | (~\[6695]  | ~\[6705] )),
  \[65]  = ~v14 & (~v13 & ~\[10341] ),
  \[4694]  = ~\[10073]  & (~v13 & (~v15 & ~\[12752] )),
  \[8011]  = ~v10 & (~v9 & ~v13),
  \[11666]  = ~v11 | (~v8 | ~\[10072] ),
  \[66]  = ~\[10076]  & (~v13 & ~\[10344] ),
  \[10805]  = ~v8 | (~\[10064]  | ~v12),
  \[21587]  = ~v10 | (~v8 | (~\[10068]  | ~\[9589] )),
  \[1448]  = ~\[34]  & (~\[33]  & (~\[32]  & ~\[31] )),
  \[67]  = ~\[10064]  & (~\[10058]  & (~v11 & ~\[10348] )),
  \[13326]  = ~v15 | ~v13,
  \[6355]  = ~\[10058]  & (~v10 & ~v13),
  \[68]  = ~\[10063]  & (~v8 & (~\[10068]  & ~\[10352] )),
  \[21589]  = ~v9 | (~\[10058]  | (~v11 | ~\[9579] )),
  \[2641]  = ~\[10058]  & (~v10 & ~v12),
  \[5160]  = ~\[10060]  & (~v1 & ~v3),
  \[12867]  = ~v15 | (~v13 | ~\[4467] ),
  \[11672]  = ~v0 | (~v2 | (~\[10176]  | ~\[6851] )),
  \[8746]  = ~\[10073]  & (~v15 & ~\[10724] ),
  \[5891]  = ~v6 & (~v5 & (~\[12153]  & ~v2)),
  \[12139]  = ~v13 | (~\[10088]  | (~\[10073]  | ~\[5923] )),
  \[10473]  = ~v1 | (~\[10099]  | (~v3 | ~\[9251] )),
  \[313]  = ~\[12682]  & (~v11 & (~\[12685]  & ~\[12681] )),
  \[12133]  = ~v5 | (~\[10134]  | ~v6),
  \[7552]  = ~\[10072]  & (~v12 & ~v14),
  \[314]  = ~\[12692]  & (~v11 & (~\[12695]  & ~\[12691] )),
  \[10475]  = ~v11 | (~v8 | ~v12),
  \[21927]  = ~v14 | (~\[10076]  | (~\[6579]  | ~\[6589] )),
  \[315]  = ~\[12674]  & (~v15 & (~\[12673]  & ~\[12670] )),
  \[4306]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[9212]  = ~\[10073]  & (~v15 & ~\[10501] ),
  \[10817]  = ~v1 | ~\[10099] ,
  \[5896]  = ~\[10072]  & (~v12 & ~v14),
  \[21591]  = ~v12 | (~v15 | ~\[9569] ),
  \[21929]  = ~v14 | (~\[10076]  | (~\[6561]  | ~\[6571] )),
  \[22059]  = ~\[5290]  | ~\[5301] ,
  \[3841]  = ~v10 & (~v9 & ~v12),
  \[10481]  = ~v4 | (~\[10135]  | ~\[9238] ),
  \[14198]  = ~v10 | (~v9 | ~\[10068] ),
  \[21923]  = ~v14 | (~\[10076]  | (~\[6615]  | ~\[6625] )),
  \[7557]  = ~v9 & (~v7 & ~v10),
  \[12872]  = ~v4 | (~\[10135]  | ~\[4458] ),
  \[73]  = ~\[10064]  & (~v9 & (~v11 & ~\[10383] )),
  \[11674]  = ~v11 | (~v8 | ~\[10072] ),
  \[74]  = ~v13 & (~v3 & (~v14 & ~\[10387] )),
  \[21925]  = ~v14 | (~\[10076]  | (~\[6597]  | ~\[6607] )),
  \[75]  = ~v13 & (~v3 & (~\[10076]  & ~\[10378] )),
  \[10815]  = ~v14 | (~\[10076]  | (~\[8574]  | ~v12)),
  \[10820]  = ~v5 | (~\[10134]  | ~v6),
  \[6365]  = ~\[10099]  & (~\[10060]  & (~v3 & ~\[11898] )),
  \[13335]  = ~v15 | ~v13,
  \[21931]  = ~v14 | (~\[10076]  | (~\[6543]  | ~\[6553] )),
  \[2651]  = ~\[10059]  & (~v0 & (~v2 & ~\[13775] )),
  \[8754]  = ~\[10060]  & (~v1 & ~v3),
  \[22061]  = ~\[5271]  | (~\[5278]  | ~\[5266] ),
  \[12878]  = ~v0 | (~v2 | ~\[10176] ),
  \[13340]  = ~v5 | (~\[10134]  | ~v6),
  \[10483]  = ~v11 | (~v8 | ~v12),
  \[12874]  = ~v11 | (~v8 | ~\[10088] ),
  \[9220]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[8029]  = ~v10 & (~v9 & ~v13),
  \[21937]  = ~v14 | (~\[10076]  | (~\[6489]  | ~\[6499] )),
  \[12146]  = ~v5 | (~\[10134]  | ~v6),
  \[4316]  = ~\[10076]  & (~\[10072]  & (~\[12939]  & ~v12)),
  \[10828]  = ~v1 | (~\[10099]  | ~v3),
  \[11688]  = ~v8 | (~\[10133]  | (~v11 | ~\[6822] )),
  \[6705]  = ~\[10059]  & (~v0 & (~\[10176]  & ~\[11746] )),
  \[21939]  = ~v14 | (~\[10076]  | (~\[6471]  | ~\[6481] )),
  \[2659]  = ~\[10058]  & (~v10 & ~v12),
  \[13348]  = ~\[22237]  | (~\[22235]  | (~\[22233]  | ~\[22231] )),
  \[21933]  = ~v14 | (~\[10076]  | (~\[6525]  | ~\[6535] )),
  \[9955]  = ~\[10099]  & (~v2 & ~v8),
  \[1464]  = ~\[29]  & (~\[28]  & (~\[30]  & ~\[10181] )),
  \[22063]  = ~\[5245]  | (~\[5252]  | ~\[5240] ),
  \[11689]  = ~v0 | ~v2,
  \[5512]  = ~\[10088]  & (~\[10073]  & (~v15 & ~\[12353] )),
  \[84]  = ~\[10459]  & (~\[10457]  & (~\[10454]  & ~\[10452] )),
  \[21935]  = ~v14 | (~\[10076]  | (~\[6507]  | ~\[6517] )),
  \[7569]  = ~\[10099]  & (~\[10060]  & (~v3 & ~\[11316] )),
  \[22065]  = ~\[5221]  | (~\[5226]  | ~\[5216] ),
  \[11683]  = ~v5 | (~\[10134]  | (~v6 | ~\[6838] )),
  \[85]  = ~\[10073]  & (~v15 & (~\[10466]  & ~\[10464] )),
  \[10826]  = ~v12 | (~v14 | (~\[10076]  | ~\[8555] )),
  \[9958]  = ~\[10064]  & ~v11,
  \[6373]  = ~\[10058]  & (~v10 & ~v13),
  \[86]  = ~\[10073]  & (~v15 & (~\[10475]  & ~\[10473] )),
  \[3126]  = ~\[10072]  & (~v12 & ~v14),
  \[22407]  = ~\[1807]  | (~v3 | (~\[1803]  | ~\[1798] )),
  \[87]  = ~\[10073]  & (~v15 & (~\[10483]  & ~\[10481] )),
  \[10830]  = ~v5 | (~\[10134]  | ~v6),
  \[8763]  = ~\[10058]  & (~v10 & ~\[10088] ),
  \[21941]  = ~\[6446]  | (~\[6451]  | ~\[6463] ),
  \[22409]  = ~\[1781]  | (~\[1786]  | ~\[1776] ),
  \[5517]  = ~\[10236]  & (~\[10135]  & ~v7),
  \[1803]  = ~\[10134]  & (~v6 & ~v8),
  \[11692]  = ~v5 | (~\[10134]  | ~v6),
  \[331]  = ~v6 & (~v5 & (~\[12853]  & ~\[12859] )),
  \[22403]  = ~\[1851]  | (~v3 | (~\[1847]  | ~\[1842] )),
  \[5182]  = ~\[10059]  & (~v0 & ~v2),
  \[332]  = ~v6 & (~v5 & (~\[12861]  & ~\[12867] )),
  \[10493]  = ~v11 | (~v8 | ~v12),
  \[12884]  = ~v15 | (~v13 | ~\[4431] ),
  \[333]  = ~\[10076]  & (~\[10072]  & (~\[12874]  & ~\[12872] )),
  \[22405]  = ~\[1825]  | (~\[1830]  | ~\[1820] ),
  \[4324]  = ~\[10060]  & (~v1 & ~v3),
  \[12153]  = ~v1 | ~\[10099] ,
  \[1807]  = ~\[10059]  & ~v0,
  \[334]  = ~\[10134]  & (~v6 & (~\[12878]  & ~\[12884] )),
  \[21947]  = ~v14 | (~\[10076]  | (~\[6391]  | ~\[6401] )),
  \[335]  = ~\[12895]  & (~\[12893]  & ~\[12891] ),
  \[6714]  = ~\[10073]  & (~v15 & (~\[11740]  & ~v13)),
  \[1471]  = ~\[23]  & (~\[22]  & (~\[21]  & ~\[20] )),
  \[7574]  = ~\[10072]  & (~v12 & ~v14),
  \[11698]  = ~v8 | (~\[10133]  | (~v11 | ~\[6800] )),
  \[336]  = ~\[12905]  & (~\[12903]  & (~\[12900]  & ~\[12898] )),
  \[21949]  = ~v14 | (~\[10076]  | (~\[6373]  | ~\[6383] )),
  \[2669]  = ~\[10134]  & (~v6 & ~\[13763] ),
  \[337]  = ~\[10076]  & (~\[10072]  & (~\[12913]  & ~\[12911] )),
  \[22411]  = ~\[1763]  | (~v3 | (~\[1759]  | ~\[1754] )),
  \[91]  = ~\[10073]  & (~v15 & (~\[10522]  & ~\[10520] )),
  \[3861]  = ~v9 & (~v7 & ~v10),
  \[338]  = ~\[10133]  & (~v5 & (~\[12917]  & ~\[12923] )),
  \[92]  = ~\[10073]  & (~v15 & (~\[10530]  & ~\[10528] )),
  \[21943]  = ~\[6424]  | (~\[6429]  | ~\[6441] ),
  \[93]  = ~\[10073]  & (~v15 & (~\[10539]  & ~\[10537] )),
  \[12891]  = ~v5 | (~\[10134]  | (~v6 | ~\[4422] )),
  \[94]  = ~\[10073]  & (~v15 & (~\[10547]  & ~\[10545] )),
  \[21945]  = ~v14 | (~\[10076]  | (~\[6409]  | ~\[6419] )),
  \[7579]  = ~v9 & (~v7 & ~v10),
  \[95]  = ~\[10559]  & (~v15 & (~\[10558]  & ~\[10556] )),
  \[10836]  = ~v12 | (~v14 | (~\[10076]  | ~\[8533] )),
  \[9238]  = ~\[10059]  & (~v0 & ~v2),
  \[6383]  = ~\[10060]  & (~v1 & (~v3 & ~\[11914] )),
  \[5524]  = ~\[10176]  & (~v4 & (~\[10059]  & ~v0)),
  \[96]  = ~\[10570]  & (~\[10568]  & (~\[10565]  & ~\[10563] )),
  \[13353]  = ~v5 | (~\[10134]  | ~v6),
  \[1478]  = ~\[19]  & (~\[18]  & (~\[17]  & ~\[16] )),
  \[10110]  = ~\[21493]  | (~\[21491]  | (~\[21489]  | ~\[21487] )),
  \[7913]  = ~v10 & (~v9 & ~v13),
  \[22417]  = ~\[1693]  | (~\[1698]  | ~\[1688] ),
  \[97]  = ~\[10073]  & (~v15 & (~\[10578]  & ~\[10576] )),
  \[10840]  = ~v1 | (~\[10099]  | ~\[10060] ),
  \[8773]  = ~v6 & (~v5 & (~\[10711]  & ~v3)),
  \[98]  = ~\[10073]  & (~v15 & (~\[10586]  & ~\[10584] )),
  \[21951]  = ~v14 | (~\[10076]  | (~\[6355]  | ~\[6365] )),
  \[12500]  = ~v10 | ~v9,
  \[12898]  = ~v0 | (~v2 | ~\[10176] ),
  \[13360]  = ~v1 | ~\[10099] ,
  \[22413]  = ~\[1737]  | (~\[1742]  | ~\[1732] ),
  \[8047]  = ~v10 & (~v9 & ~v13),
  \[343]  = ~\[12970]  & (~v2 & (~\[12973]  & ~\[12979] )),
  \[6722]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[22415]  = ~\[1710]  | ~\[1721] ,
  \[4334]  = ~\[10058]  & (~v10 & (~v12 & ~\[12933] )),
  \[12163]  = ~v1 | (~\[10099]  | ~v3),
  \[12893]  = ~v8 | (~\[10133]  | ~v11),
  \[344]  = ~\[12983]  & (~\[12981]  & ~\[12989] ),
  \[21957]  = ~\[6298]  | (~v11 | (~\[6294]  | ~\[6311] )),
  \[2677]  = ~\[10058]  & (~v10 & ~v12),
  \[11305]  = ~v5 | (~\[10134]  | ~v6),
  \[345]  = ~v6 & (~v5 & (~\[12963]  & ~\[12969] )),
  \[10848]  = ~v1 | (~\[10099]  | ~v3),
  \[12895]  = ~v13 | (~\[10088]  | ~v15),
  \[21959]  = ~\[6276]  | (~v11 | (~\[6272]  | ~\[6289] )),
  \[22089]  = ~\[4949]  | (~\[4954]  | ~\[4944] ),
  \[3142]  = ~\[10059]  & (~v0 & ~v2),
  \[21953]  = ~v14 | (~\[10076]  | (~\[6337]  | ~\[6347] )),
  \[12172]  = ~v4 | ~\[10135] ,
  \[5199]  = ~\[10133]  & (~v5 & ~v8),
  \[13702]  = ~v11 | ~v8,
  \[12509]  = ~v0 | (~v2 | (~\[10176]  | ~\[5199] )),
  \[6391]  = ~\[10058]  & (~v10 & ~v13),
  \[21955]  = ~v14 | (~\[10076]  | (~\[6319]  | ~\[6329] )),
  \[10846]  = ~v14 | (~\[10076]  | (~\[8512]  | ~v12)),
  \[8781]  = ~\[10058]  & (~v10 & ~\[10088] ),
  \[12503]  = ~v12 | (~v14 | ~\[10076] ),
  \[1820]  = ~\[10072]  & (~v12 & (~v14 & ~\[14187] )),
  \[22427]  = ~\[1570]  | ~\[1581] ,
  \[21961]  = ~v14 | (~\[10076]  | (~\[6257]  | ~\[6267] )),
  \[12510]  = ~v10 | ~v9,
  \[22091]  = ~\[4931]  | (~v3 | (~\[4927]  | ~\[4922] )),
  \[22429]  = ~\[1548]  | ~\[1559] ,
  \[13370]  = ~v1 | (~\[10099]  | ~v3),
  \[13708]  = ~v4 | ~v7,
  \[5538]  = ~\[10088]  & (~\[10073]  & (~v15 & ~\[12341] )),
  \[4342]  = ~\[10059]  & (~v0 & ~v2),
  \[8057]  = ~\[10133]  & (~v5 & ~\[11053] ),
  \[12179]  = ~\[22005]  | (~\[22003]  | (~\[22001]  | ~\[21999] )),
  \[1825]  = ~\[10134]  & (~v6 & ~v8),
  \[7591]  = ~\[10060]  & (~v1 & (~v3 & ~\[11305] )),
  \[6732]  = ~\[10073]  & (~v15 & (~\[11731]  & ~v13)),
  \[11316]  = ~v5 | (~\[10134]  | ~v6),
  \[9251]  = ~v6 & ~v5,
  \[21967]  = ~v14 | (~\[10076]  | (~\[6203]  | ~\[6213] )),
  \[2687]  = ~\[10059]  & (~v0 & (~v2 & ~\[13756] )),
  \[10857]  = ~v1 | (~\[10099]  | ~\[10060] ),
  \[21969]  = ~v14 | (~\[10076]  | (~\[6185]  | ~\[6195] )),
  \[6006]  = ~\[10059]  & (~v0 & ~v2),
  \[9983]  = ~\[10099]  & (~v2 & ~v9),
  \[22431]  = ~\[1526]  | ~\[1537] ,
  \[10129]  = ~v14 | (~v13 | ~\[10076] ),
  \[3152]  = ~\[10072]  & (~v14 & (~\[13520]  & ~v12)),
  \[21963]  = ~v14 | (~\[10076]  | (~\[6239]  | ~\[6249] )),
  \[22093]  = ~\[4905]  | (~\[4910]  | ~\[4900] ),
  \[10854]  = ~v14 | (~\[10076]  | (~\[8494]  | ~v12)),
  \[12181]  = ~v1 | (~\[10099]  | ~v3),
  \[3883]  = ~v9 & (~v7 & ~v10),
  \[12519]  = ~v4 | (~v7 | (~\[10058]  | ~\[5182] )),
  \[10123]  = ~\[21501]  | (~\[21499]  | (~\[21497]  | ~\[21495] )),
  \[21965]  = ~v14 | (~\[10076]  | (~\[6221]  | ~\[6231] )),
  \[7599]  = ~v10 & (~v9 & ~v12),
  \[22095]  = ~\[4878]  | ~\[4889] ,
  \[5543]  = ~\[10236]  & (~\[10135]  & ~v7),
  \[8791]  = ~v6 & (~v5 & (~\[10702]  & ~v3)),
  \[12513]  = ~v12 | (~v14 | ~\[10076] ),
  \[7203]  = ~v9 & (~v7 & ~\[10068] ),
  \[1830]  = ~\[10059]  & (~v0 & ~v2),
  \[7933]  = ~v9 & (~v7 & ~v10),
  \[21971]  = ~v14 | (~\[10076]  | (~\[6167]  | ~\[6177] )),
  \[12520]  = ~v10 | ~v9,
  \[8065]  = ~v10 & (~v9 & ~v13),
  \[12187]  = ~v13 | (~\[10073]  | ~\[5791] ),
  \[13718]  = ~v5 | (~\[10134]  | ~v6),
  \[4351]  = ~\[10068]  & (~\[10058]  & ~v12),
  \[361]  = ~\[10134]  & (~\[10133]  & (~\[13136]  & ~\[13142] )),
  \[6740]  = ~\[10060]  & (~v1 & ~v3),
  \[1105]  = ~\[207]  & (~\[206]  & (~\[205]  & ~\[204] )),
  \[12189]  = ~v1 | (~\[10099]  | ~v3),
  \[362]  = ~\[10134]  & (~\[10133]  & (~\[13144]  & ~\[13150] )),
  \[2695]  = ~\[10058]  & (~v10 & ~v12),
  \[363]  = ~\[13152]  & (~v2 & (~\[13155]  & ~\[13161] )),
  \[364]  = ~\[13165]  & (~\[13163]  & ~\[13171] ),
  \[21977]  = ~v14 | (~\[10076]  | (~\[6113]  | ~\[6123] )),
  \[9991]  = ~\[10099]  & (~v2 & ~v8),
  \[11325]  = ~v7 | ~\[10236] ,
  \[365]  = ~v6 & (~v5 & (~\[13175]  & ~\[13181] )),
  \[6015]  = ~\[10068]  & (~v9 & ~v13),
  \[10137]  = ~v6 | (~v4 | ~\[10133] ),
  \[366]  = ~v6 & (~v5 & (~\[13183]  & ~\[13189] )),
  \[3160]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[21979]  = ~v14 | (~\[10076]  | (~\[6095]  | ~\[6105] )),
  \[367]  = ~\[10134]  & (~v6 & (~\[13192]  & ~\[13198] )),
  \[13388]  = ~v1 | (~\[10099]  | ~v3),
  \[8405]  = ~v10 & (~v9 & ~\[10088] ),
  \[11332]  = ~\[21825]  | (~\[21823]  | (~\[21821]  | ~\[21819] )),
  \[368]  = ~\[10134]  & (~v6 & (~\[13200]  & ~\[13206] )),
  \[5550]  = ~v4 & (~v2 & (~\[10059]  & ~v0)),
  \[2303]  = ~v6 & (~v5 & ~v8),
  \[21973]  = ~v14 | (~\[10076]  | (~\[6149]  | ~\[6159] )),
  \[10134]  = ~v4,
  \[12529]  = ~\[933]  | (~\[940]  | (~\[926]  | ~\[971] )),
  \[10133]  = ~v7,
  \[6749]  = ~\[10058]  & (~v10 & ~v13),
  \[10863]  = ~v14 | (~\[10076]  | (~\[8476]  | ~v12)),
  \[21975]  = ~v14 | (~\[10076]  | (~\[6131]  | ~\[6141] )),
  \[703]  = ~\[13627]  & (~\[13592]  & ~\[13694] ),
  \[12523]  = ~v14 | (~\[10072]  | ~\[10076] ),
  \[10135]  = ~v6,
  \[10865]  = ~v1 | (~\[10099]  | ~v3),
  \[9269]  = ~v6 & ~v5,
  \[2307]  = ~\[10059]  & ~v0,
  \[13383]  = ~v15 | ~v13,
  \[13386]  = ~\[22245]  | (~\[22243]  | (~\[22241]  | ~\[22239] )),
  \[21981]  = ~\[6074]  | (~v11 | (~\[6070]  | ~\[6087] )),
  \[1842]  = ~\[10072]  & (~v12 & (~v14 & ~\[14177] )),
  \[8075]  = ~\[10059]  & (~v0 & (~v2 & ~\[11070] )),
  \[12197]  = ~v1 | (~\[10099]  | ~\[10060] ),
  \[13728]  = ~v5 | (~\[10134]  | ~v6),
  \[10141]  = ~v6 | (~v4 | ~\[10133] ),
  \[10871]  = ~v14 | (~\[10076]  | (~\[8458]  | ~v12)),
  \[3502]  = ~\[10072]  & (~v12 & ~\[10076] ),
  \[373]  = ~\[10134]  & (~v6 & (~\[13256]  & ~\[13262] )),
  \[1847]  = ~v6 & (~v5 & ~v8),
  \[374]  = ~\[10134]  & (~v6 & (~\[13264]  & ~\[13270] )),
  \[3506]  = ~v9 & ~v7,
  \[11335]  = ~v4 | ~v7,
  \[375]  = ~\[13245]  & (~v3 & (~\[13248]  & ~\[13254] )),
  \[12195]  = ~v13 | (~\[10073]  | ~\[5827] ),
  \[3170]  = ~\[10072]  & (~v14 & (~\[13512]  & ~v12)),
  \[10877]  = ~v7 | ~\[10236] ,
  \[8415]  = ~v6 & (~v5 & (~\[10892]  & ~v3)),
  \[10149]  = ~v6 | ~v4,
  \[11341]  = ~v0 | ~v2,
  \[12539]  = ~v12 | (~v14 | ~\[10076] ),
  \[6759]  = ~\[10059]  & (~v0 & (~v2 & ~\[11721] )),
  \[10146]  = ~v6 | ~v4,
  \[4705]  = ~\[10099]  & (~\[10060]  & (~v3 & ~\[12749] )),
  \[12536]  = ~v10 | ~v9,
  \[8083]  = ~v10 & (~v9 & ~v13),
  \[13396]  = ~v1 | (~\[10099]  | ~v3),
  \[12535]  = ~v4 | (~v7 | (~\[10058]  | ~\[5138] )),
  \[1851]  = ~\[10059]  & ~v0,
  \[716]  = ~\[404]  & (~\[403]  & (~\[405]  & ~\[13525] )),
  \[3178]  = ~\[10059]  & (~v0 & ~v2),
  \[1122]  = ~\[11576]  & (~\[11539]  & ~\[11641] ),
  \[7955]  = ~v9 & (~v7 & ~v10),
  \[13008]  = ~v15 | ~v13,
  \[5900]  = ~v9 & ~v7,
  \[7227]  = ~\[10134]  & ~v6,
  \[13737]  = ~v1 | ~\[10099] ,
  \[12542]  = ~v1 | (~\[10099]  | ~v3),
  \[6033]  = ~\[10068]  & (~v9 & ~v13),
  \[10158]  = ~v6 | (~v4 | ~\[10133] ),
  \[2320]  = ~\[10072]  & (~v12 & (~\[10076]  & ~\[13937] )),
  \[8423]  = ~v10 & (~v9 & ~\[10088] ),
  \[13736]  = ~\[22319]  | (~\[22317]  | (~\[22315]  | ~\[22313] )),
  \[21999]  = ~\[5900]  | (~v11 | (~\[5896]  | ~\[5913] )),
  \[4378]  = ~\[10060]  & (~v1 & ~v3),
  \[3519]  = ~\[10059]  & (~v0 & (~v2 & ~\[13340] )),
  \[14208]  = ~v10 | (~v9 | ~\[10068] ),
  \[11351]  = ~v4 | ~v7,
  \[10154]  = ~v6 | (~v4 | ~\[10133] ),
  \[10884]  = ~v1 | (~\[10099]  | ~v3),
  \[13012]  = ~v1 | (~\[10099]  | ~v3),
  \[5572]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[2325]  = ~v6 & (~v5 & ~v8),
  \[723]  = ~\[398]  & (~\[397]  & (~\[396]  & ~\[395] )),
  \[12543]  = ~v4 | ~v7,
  \[4716]  = ~\[10073]  & (~v13 & (~v15 & ~\[12740] )),
  \[8093]  = ~\[10134]  & (~v6 & ~\[11061] ),
  \[11358]  = ~\[21829]  | (~\[21827]  | ~\[21831] ),
  \[3188]  = ~\[10068]  & (~v9 & (~v12 & ~\[13505] )),
  \[21609]  = ~v12 | (~v15 | (~\[9484]  | ~v7)),
  \[12550]  = ~v10 | (~v9 | (~\[10068]  | ~\[5100] )),
  \[10892]  = ~v2 | ~\[10059] ,
  \[391]  = ~v6 & (~v5 & (~\[13417]  & ~\[13423] )),
  \[1135]  = ~\[194]  & (~\[193]  & (~\[195]  & ~\[11472] )),
  \[392]  = ~v6 & (~v5 & (~\[13425]  & ~\[13431] )),
  \[6771]  = ~\[10133]  & ~v5,
  \[393]  = ~\[10134]  & (~v6 & (~\[13434]  & ~\[13440] )),
  \[5913]  = ~\[10059]  & (~v0 & (~\[10176]  & ~\[12146] )),
  \[394]  = ~\[10134]  & (~v6 & (~\[13442]  & ~\[13448] )),
  \[395]  = ~\[13451]  & (~v3 & (~\[13454]  & ~\[13460] )),
  \[2330]  = ~\[10059]  & (~v0 & ~v2),
  \[8433]  = ~\[10133]  & (~v5 & ~\[10884] ),
  \[13746]  = ~v1 | (~\[10099]  | ~v3),
  \[1869]  = ~v6 & (~v5 & ~v8),
  \[396]  = ~\[13461]  & (~v3 & (~\[13464]  & ~\[13470] )),
  \[21611]  = ~v14 | (~v13 | (~\[10076]  | ~\[9477] )),
  \[3528]  = ~\[10068]  & (~v9 & (~v12 & ~\[13335] )),
  \[397]  = ~\[10133]  & (~v5 & (~\[13473]  & ~\[13479] )),
  \[12557]  = ~v5 | (~v6 | (~\[10133]  | ~\[5094] )),
  \[398]  = ~\[10133]  & (~v5 & (~\[13481]  & ~\[13487] )),
  \[10501]  = ~v11 | (~v8 | ~v12),
  \[730]  = ~\[394]  & (~\[393]  & (~\[392]  & ~\[391] )),
  \[11361]  = ~\[1202]  | (~\[1209]  | (~\[1195]  | ~\[1182] )),
  \[2335]  = ~\[10072]  & ~v12,
  \[3196]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[14213]  = ~\[22409]  | (~\[22407]  | (~\[22405]  | ~\[22403] )),
  \[11368]  = ~v11 | (~\[10063]  | ~v12),
  \[4727]  = ~\[10060]  & (~v1 & (~v3 & ~\[12737] )),
  \[9633]  = ~\[10135]  & (~v5 & ~v7),
  \[1142]  = ~\[188]  & (~\[187]  & (~\[186]  & ~\[185] )),
  \[12560]  = ~v10 | (~\[10068]  | (~v9 | ~\[10058] )),
  \[7975]  = ~v10 & (~v9 & ~v13),
  \[13028]  = ~\[22169]  | (~\[22167]  | (~\[22165]  | ~\[22163] )),
  \[10509]  = ~v11 | (~v8 | ~v12),
  \[14220]  = ~v10 | (~v9 | ~\[10068] ),
  \[21613]  = ~v12 | (~\[10073]  | (~\[9464]  | ~v7)),
  \[12561]  = ~v14 | ~\[10072] ,
  \[21615]  = ~v9 | (~\[10058]  | (~\[10064]  | ~\[9457] )),
  \[5923]  = ~v9 & (~v7 & ~\[10068] ),
  \[8441]  = ~v10 & (~v9 & ~\[10088] ),
  \[6053]  = ~v9 & (~v7 & ~\[10068] ),
  \[11366]  = ~v4 | (~v7 | ~\[7474] ),
  \[3536]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[1149]  = ~\[184]  & (~\[183]  & (~\[182]  & ~\[181] )),
  \[13756]  = ~v4 | ~\[10135] ,
  \[13025]  = ~v15 | ~v13,
  \[12900]  = ~v5 | (~\[10134]  | ~v6),
  \[13030]  = ~v1 | (~\[10099]  | ~v3),
  \[12567]  = ~v5 | ~v6,
  \[2343]  = ~\[10064]  & (~v11 & (~\[10063]  & ~v8)),
  \[4002]  = ~\[10060]  & (~v1 & ~v3),
  \[7250]  = ~\[10060]  & (~v1 & ~v3),
  \[10176]  = ~v3,
  \[11703]  = ~v7 | (~\[10236]  | ~\[6794] ),
  \[5594]  = ~\[10059]  & (~v0 & ~v2),
  \[21627]  = ~v12 | (~\[10176]  | (~v15 | ~\[9389] )),
  \[12566]  = ~v3 | (~\[10134]  | (~v1 | ~\[10099] )),
  \[11705]  = ~v11 | (~v8 | ~\[10072] ),
  \[4007]  = ~\[10072]  & ~v12,
  \[21629]  = ~\[9372]  | ~\[9379] ,
  \[4738]  = ~\[10073]  & (~v13 & (~v15 & ~\[12730] )),
  \[10181]  = ~\[21525]  | (~\[21523]  | (~\[21521]  | ~\[21519] )),
  \[14230]  = ~v10 | (~v9 | ~\[10068] ),
  \[13037]  = ~v2 | ~\[10059] ,
  \[21623]  = ~v10 | (~v8 | (~\[10068]  | ~\[9413] )),
  \[9645]  = ~v12 & (~v7 & (~\[10135]  & ~v5)),
  \[11711]  = ~v0 | (~v2 | (~\[10176]  | ~\[6771] )),
  \[10514]  = ~\[21649]  | (~\[21647]  | (~\[21651]  | ~\[1344] )),
  \[11374]  = ~v4 | (~v7 | (~\[7455]  | ~v3)),
  \[21625]  = ~v9 | (~\[10058]  | (~v11 | ~\[9401] )),
  \[7259]  = ~\[10068]  & (~v9 & ~\[10088] ),
  \[10516]  = ~\[1381]  | (~\[1388]  | (~\[1374]  | ~\[1361] )),
  \[8451]  = ~\[10059]  & (~v0 & (~v2 & ~\[10877] )),
  \[11376]  = ~v11 | (~\[10063]  | ~v12),
  \[1887]  = ~\[10064]  & (~v11 & (~\[10063]  & ~v8)),
  \[12903]  = ~v8 | (~\[10133]  | ~v11),
  \[3546]  = ~\[10068]  & (~v9 & (~v12 & ~\[13326] )),
  \[13763]  = ~v1 | (~\[10099]  | ~v3),
  \[6794]  = ~\[10060]  & (~v1 & ~v3),
  \[10520]  = ~v2 | (~\[10059]  | (~\[10176]  | ~\[9161] )),
  \[11380]  = ~v1 | ~\[10099] ,
  \[12905]  = ~v13 | (~\[10088]  | ~v15),
  \[21631]  = ~v1 | (~\[10099]  | (~v2 | ~\[9360] )),
  \[10522]  = ~v11 | (~v8 | ~v12),
  \[6401]  = ~\[10133]  & (~v5 & (~\[11904]  & ~v3)),
  \[12911]  = ~v7 | (~\[10236]  | ~\[4378] ),
  \[4013]  = ~\[10058]  & (~v7 & ~v10),
  \[8458]  = ~v10 & ~v9,
  \[13771]  = ~\[22327]  | (~\[22325]  | (~\[22323]  | ~\[22321] )),
  \[10186]  = ~v10 | ~\[10068] ,
  \[11713]  = ~v11 | (~v8 | ~\[10072] ),
  \[21637]  = ~\[9308]  | ~\[9319] ,
  \[2357]  = ~\[10236]  & (~\[10135]  & (~v7 & ~\[13921] )),
  \[7993]  = ~v10 & (~v9 & ~v13),
  \[10528]  = ~v0 | (~v2 | (~\[10176]  | ~\[9143] )),
  \[12575]  = ~v14 | (~\[10072]  | (~\[10076]  | ~\[5055] )),
  \[14236]  = ~v0 | (~v2 | ~\[10176] ),
  \[9653]  = ~\[10135]  & (~v5 & ~v7),
  \[12917]  = ~v0 | (~v2 | ~\[10176] ),
  \[21633]  = ~v4 | (~v7 | (~\[9354]  | ~\[9346] )),
  \[4749]  = ~\[10133]  & (~v5 & (~v8 & ~\[12725] )),
  \[6070]  = ~\[10073]  & (~v13 & ~v15),
  \[12582]  = ~v1 | (~\[10099]  | (~\[10060]  | ~\[5037] )),
  \[11389]  = ~v12 | (~v14 | (~\[10076]  | ~\[7427] )),
  \[11721]  = ~v4 | ~v7,
  \[6409]  = ~\[10058]  & (~v10 & ~v13),
  \[21635]  = ~v4 | (~v7 | (~\[9336]  | ~\[9328] )),
  \[3554]  = ~\[10059]  & (~v0 & ~v2),
  \[7269]  = ~v6 & (~v5 & (~\[11463]  & ~v3)),
  \[11383]  = ~v5 | (~\[10134]  | ~v6),
  \[14241]  = ~v10 | (~v9 | ~\[10068] ),
  \[12913]  = ~v11 | (~v8 | ~\[10088] ),
  \[6074]  = ~v9 & ~v7,
  \[22107]  = ~\[4738]  | ~\[4749] ,
  \[10530]  = ~v11 | (~v8 | ~v12),
  \[13046]  = ~v0 | ~v2,
  \[5216]  = ~\[10088]  & (~\[10073]  & (~v15 & ~\[12489] )),
  \[13775]  = ~v7 | ~\[10236] ,
  \[22109]  = ~\[4716]  | ~\[4727] ,
  \[10199]  = ~v11 | ~v9,
  \[11391]  = ~v1 | (~\[10099]  | ~v3),
  \[22103]  = ~\[4789]  | (~\[4796]  | ~\[4784] ),
  \[13782]  = ~v1 | (~\[10099]  | ~v3),
  \[10193]  = ~\[1471]  | (~\[1478]  | (~\[1464]  | ~\[1511] )),
  \[762]  = ~\[13412]  & (~\[13386]  & (~\[13348]  & ~\[13311] )),
  \[8800]  = ~\[10073]  & (~v15 & ~\[10699] ),
  \[7609]  = ~\[10134]  & (~v6 & (~\[11294]  & ~v3)),
  \[22105]  = ~\[4765]  | (~\[4770]  | ~\[4760] ),
  \[12583]  = ~v10 | ~v9,
  \[10195]  = ~v3 | (~\[10059]  | ~v8),
  \[4025]  = ~\[10099]  & (~\[10060]  & (~v3 & ~\[13087] )),
  \[21647]  = ~v4 | (~\[10135]  | (~\[9220]  | ~\[9212] )),
  \[12586]  = ~v14 | (~\[10072]  | ~\[10076] ),
  \[10537]  = ~v4 | (~\[10135]  | ~\[9130] ),
  \[21649]  = ~v7 | (~\[10236]  | (~\[9202]  | ~\[9194] )),
  \[2369]  = ~\[10064]  & (~v11 & (~\[10063]  & ~v8)),
  \[9663]  = ~\[10135]  & (~v5 & ~v7),
  \[22111]  = ~\[4694]  | ~\[4705] ,
  \[4029]  = ~\[10072]  & ~v12,
  \[10539]  = ~v11 | (~v8 | ~v12),
  \[7277]  = ~\[10068]  & (~v9 & ~\[10088] ),
  \[12592]  = ~v1 | (~\[10099]  | (~v3 | ~\[5015] )),
  \[11399]  = ~v12 | (~v14 | (~\[10076]  | ~\[7405] )),
  \[5221]  = ~\[10133]  & (~v5 & ~v8),
  \[11731]  = ~v11 | ~v8,
  \[5951]  = ~\[10059]  & ~v0,
  \[6419]  = ~\[10060]  & (~v1 & (~v3 & ~\[11888] )),
  \[3564]  = ~v10 & (~v9 & (~v12 & ~\[13318] )),
  \[2705]  = ~v6 & (~v5 & ~\[13746] ),
  \[8808]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[11393]  = ~v5 | (~\[10134]  | ~v6),
  \[14251]  = ~v10 | (~v9 | ~\[10068] ),
  \[12923]  = ~v15 | (~v13 | ~\[4351] ),
  \[22117]  = ~\[4636]  | ~\[4647] ,
  \[1511]  = ~\[10123]  & (~\[10110]  & (~\[10095]  & ~\[10079] )),
  \[5226]  = ~\[10060]  & (~v1 & ~v3),
  \[21651]  = ~v7 | (~\[10236]  | (~\[9184]  | ~\[9176] )),
  \[22119]  = ~\[4614]  | ~\[4625] ,
  \[13060]  = ~v15 | ~v13,
  \[4760]  = ~\[10073]  & (~v13 & (~v15 & ~\[12719] )),
  \[6087]  = ~\[10060]  & (~v1 & (~v3 & ~\[12041] )),
  \[13790]  = ~v2 | ~\[10059] ,
  \[8476]  = ~v10 & ~v9,
  \[1514]  = ~\[10797]  & (~\[10516]  & (~\[10319]  & ~\[10193] )),
  \[7617]  = ~v10 & (~v9 & ~v12),
  \[22113]  = ~v4 | (~v7 | (~\[4682]  | ~\[4674] )),
  \[3903]  = ~v10 & (~v9 & ~v12),
  \[22115]  = ~v4 | (~v7 | (~\[4664]  | ~\[4656] )),
  \[12593]  = ~v10 | ~v9,
  \[4035]  = ~\[10058]  & (~v7 & ~v10),
  \[4765]  = ~\[10133]  & (~v5 & ~v8),
  \[11005]  = ~v5 | (~\[10134]  | ~v6),
  \[12596]  = ~v14 | (~\[10072]  | ~\[10076] ),
  \[6424]  = ~\[10073]  & (~v13 & ~v15),
  \[775]  = ~\[374]  & (~\[373]  & (~\[375]  & ~\[13244] )),
  \[11740]  = ~v11 | ~v8,
  \[10547]  = ~v11 | (~v8 | ~v12),
  \[14256]  = ~\[22417]  | (~\[22415]  | (~\[22413]  | ~\[22411] )),
  \[9673]  = ~\[10135]  & (~v5 & ~v7),
  \[1182]  = ~\[11358]  & (~\[11332]  & (~\[11292]  & ~\[11257] )),
  \[12208]  = ~\[992]  | (~\[999]  | (~\[985]  | ~\[1030] )),
  \[22121]  = ~v15 | (~v13 | (~\[4593]  | ~\[4603] )),
  \[13798]  = ~v0 | ~v2,
  \[3572]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[7287]  = ~v6 & (~v5 & (~\[11455]  & ~v3)),
  \[2713]  = ~\[10058]  & (~v10 & ~v12),
  \[12209]  = ~v2 | ~\[10059] ,
  \[6429]  = ~\[10058]  & (~v7 & ~v10),
  \[12939]  = ~v11 | ~v8,
  \[14262]  = ~v0 | (~v2 | (~\[10176]  | ~\[1671] )),
  \[8818]  = ~\[10073]  & (~v15 & ~\[10689] ),
  \[12203]  = ~v13 | (~\[10073]  | ~\[5809] ),
  \[12933]  = ~v15 | ~v13,
  \[10545]  = ~v0 | (~v2 | (~\[10176]  | ~\[9107] )),
  \[13063]  = ~\[22177]  | (~\[22175]  | (~\[22173]  | ~\[22171] )),
  \[22127]  = ~v15 | (~v13 | (~\[4539]  | ~\[4549] )),
  \[11018]  = ~v5 | (~\[10134]  | ~v6),
  \[6095]  = ~\[10068]  & (~v9 & ~v13),
  \[13065]  = ~v0 | ~v2,
  \[22129]  = ~v7 | (~\[10236]  | (~\[4530]  | ~\[4522] )),
  \[4770]  = ~\[10060]  & (~v1 & ~v3),
  \[2382]  = ~v4 & (~v2 & (~\[10059]  & ~v0)),
  \[7627]  = ~\[10060]  & (~v1 & (~v3 & ~\[11285] )),
  \[22123]  = ~v15 | (~v13 | (~\[4575]  | ~\[4585] )),
  \[782]  = ~\[368]  & (~\[367]  & (~\[366]  & ~\[365] )),
  \[13409]  = ~v15 | ~v13,
  \[11013]  = ~\[21757]  | (~\[21755]  | (~\[21753]  | ~\[21751] )),
  \[1526]  = ~\[10072]  & (~v12 & (~v14 & ~\[14311] )),
  \[22125]  = ~v4 | (~\[10135]  | (~\[4566]  | ~\[4558] )),
  \[11746]  = ~v4 | ~v7,
  \[9681]  = ~\[10135]  & (~v5 & ~v7),
  \[10558]  = ~v8 | (~\[10133]  | ~v11),
  \[14263]  = ~v10 | ~v9,
  \[4047]  = ~\[10060]  & (~v1 & (~v3 & ~\[13076] )),
  \[14266]  = ~v13 | (~\[10088]  | ~\[10073] ),
  \[21669]  = ~v4 | (~v7 | (~\[9014]  | ~\[9006] )),
  \[22131]  = ~v15 | (~v13 | (~\[4503]  | ~\[4513] )),
  \[12948]  = ~v11 | ~v8,
  \[9684]  = ~v14 & ~v13,
  \[12217]  = ~v0 | ~v2,
  \[7296]  = ~\[10073]  & (~v15 & ~\[11451] ),
  \[5240]  = ~\[10088]  & (~\[10073]  & (~v15 & ~\[12479] )),
  \[10559]  = ~v12 | ~v14,
  \[5970]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[3582]  = ~v10 & (~v9 & (~v12 & ~\[13308] )),
  \[2723]  = ~v6 & (~v5 & (~\[13737]  & ~v2)),
  \[8826]  = ~\[10059]  & (~v0 & ~v2),
  \[789]  = ~\[364]  & (~\[363]  & (~\[362]  & ~\[361] )),
  \[13412]  = ~\[22249]  | (~\[22247]  | ~\[22251] ),
  \[1195]  = ~\[164]  & (~\[163]  & (~\[165]  & ~\[11190] )),
  \[10556]  = ~v5 | (~\[10134]  | (~v6 | ~\[9094] )),
  \[5245]  = ~\[10236]  & (~\[10135]  & ~v7),
  \[13076]  = ~v5 | (~\[10134]  | ~v6),
  \[2728]  = ~\[10072]  & (~v12 & ~v14),
  \[21671]  = ~v4 | (~v7 | (~\[8996]  | ~\[8988] )),
  \[8494]  = ~v10 & ~v9,
  \[7635]  = ~v10 & (~v9 & ~v12),
  \[3921]  = ~\[10058]  & (~v10 & ~v12),
  \[13417]  = ~v2 | (~\[10059]  | ~\[10176] ),
  \[14277]  = ~v13 | ~\[10088] ,
  \[6441]  = ~\[10099]  & (~\[10060]  & (~v3 & ~\[11879] )),
  \[11753]  = ~\[21915]  | (~\[21913]  | (~\[21911]  | ~\[21909] )),
  \[4784]  = ~\[10073]  & (~v13 & (~v15 & ~\[12709] )),
  \[8101]  = ~v10 & (~v9 & ~v13),
  \[1537]  = ~\[10099]  & (~\[10060]  & (~v3 & ~\[14308] )),
  \[4055]  = ~\[10058]  & (~v10 & ~v12),
  \[794]  = ~\[14339]  & (~\[13998]  & (~\[13696]  & ~\[13415] )),
  \[11025]  = ~v1 | ~\[10099] ,
  \[11755]  = ~v1 | (~\[10099]  | ~\[10060] ),
  \[10568]  = ~v8 | (~\[10133]  | ~v11),
  \[10900]  = ~v0 | ~v2,
  \[14273]  = ~v5 | (~v6 | (~\[10133]  | ~\[1654] )),
  \[14276]  = ~v10 | (~\[10068]  | (~v9 | ~\[10058] )),
  \[3590]  = ~\[10060]  & (~v1 & ~v3),
  \[13415]  = ~\[782]  | (~\[789]  | (~\[775]  | ~\[762] )),
  \[12228]  = ~v4 | ~\[10135] ,
  \[6446]  = ~\[10073]  & (~v13 & ~v15),
  \[12958]  = ~v15 | ~v13,
  \[11762]  = ~v1 | ~\[10099] ,
  \[13087]  = ~v5 | (~\[10134]  | ~v6),
  \[21673]  = ~v4 | (~v7 | (~\[8978]  | ~\[8970] )),
  \[4789]  = ~\[10236]  & (~\[10135]  & ~v7),
  \[2733]  = ~\[10058]  & (~v7 & ~v10),
  \[8836]  = ~\[10073]  & (~v15 & ~\[10681] ),
  \[11761]  = ~v14 | (~\[10076]  | ~\[6633] ),
  \[2004]  = ~\[10072]  & (~v12 & (~v14 & ~\[14096] )),
  \[5252]  = ~v4 & (~v3 & (~\[10099]  & ~\[10060] )),
  \[10563]  = ~v0 | (~v2 | ~\[10176] ),
  \[21675]  = ~v4 | (~v7 | (~\[8960]  | ~\[8952] )),
  \[403]  = ~\[13543]  & ~\[13538] ,
  \[404]  = ~\[13547]  & (~\[13545]  & ~\[13553] ),
  \[10565]  = ~v5 | (~\[10134]  | ~v6),
  \[9699]  = ~\[10135]  & (~v5 & ~v7),
  \[405]  = ~\[10072]  & (~v14 & (~\[13531]  & ~\[13529] )),
  \[10570]  = ~v12 | (~v14 | ~\[10076] ),
  \[7645]  = ~v6 & (~v5 & (~\[11275]  & ~v3)),
  \[22149]  = ~v4 | (~v7 | (~\[4342]  | ~\[4334] )),
  \[3599]  = ~v10 & (~v9 & ~v12),
  \[10909]  = ~\[21735]  | (~\[21733]  | (~\[21731]  | ~\[21729] )),
  \[5988]  = ~\[10060]  & (~v1 & ~v3),
  \[6451]  = ~\[10058]  & (~v7 & ~v10),
  \[12961]  = ~\[22155]  | (~\[22153]  | (~\[22151]  | ~\[22149] )),
  \[9308]  = ~\[10088]  & (~\[10073]  & (~v15 & ~\[10444] )),
  \[8111]  = ~\[10059]  & (~v0 & (~v2 & ~\[11044] )),
  \[4065]  = ~\[10134]  & (~v6 & (~\[13065]  & ~v3)),
  \[3206]  = ~\[10068]  & (~v9 & (~v12 & ~\[13497] )),
  \[14284]  = ~v5 | ~v6,
  \[21687]  = ~v4 | (~\[10135]  | (~\[8844]  | ~\[8836] )),
  \[13423]  = ~v15 | (~v13 | ~\[3357] ),
  \[11035]  = ~v1 | (~\[10099]  | ~v3),
  \[1548]  = ~\[10072]  & (~v12 & (~v14 & ~\[14331] )),
  \[11765]  = ~v5 | (~\[10134]  | ~v6),
  \[10578]  = ~v11 | (~v8 | ~v12),
  \[10910]  = ~v2 | ~\[10059] ,
  \[14283]  = ~\[10134]  | (~\[10176]  | (~v0 | ~v2)),
  \[4796]  = ~v4 & (~v3 & (~\[10099]  & ~\[10060] )),
  \[21689]  = ~v7 | (~\[10236]  | (~\[8826]  | ~\[8818] )),
  \[13425]  = ~v0 | (~v2 | ~\[10176] ),
  \[8844]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[22151]  = ~v4 | (~v7 | (~\[4324]  | ~\[4316] )),
  \[21683]  = ~v14 | (~\[10076]  | (~\[8871]  | ~\[8881] )),
  \[11771]  = ~v14 | (~\[10072]  | (~\[10076]  | ~\[6675] )),
  \[12969]  = ~v15 | (~v13 | ~\[4217] ),
  \[14292]  = ~v13 | (~\[10088]  | (~\[10073]  | ~\[1615] )),
  \[2015]  = ~\[10059]  & (~v0 & (~v2 & ~\[14093] )),
  \[21685]  = ~v4 | (~\[10135]  | (~\[8862]  | ~\[8854] )),
  \[13431]  = ~v15 | (~v13 | ~\[3339] ),
  \[12234]  = ~v0 | ~v2,
  \[2745]  = ~\[10059]  & (~v0 & (~\[10176]  & ~\[13728] )),
  \[10576]  = ~v7 | (~\[10236]  | ~\[9050] ),
  \[8119]  = ~v10 & (~v9 & ~v13),
  \[12963]  = ~v1 | (~\[10099]  | ~\[10060] ),
  \[414]  = ~\[10072]  & (~v14 & (~\[13634]  & ~\[13632] )),
  \[7653]  = ~v10 & (~v9 & ~v12),
  \[415]  = ~\[13646]  & ~\[13641] ,
  \[5266]  = ~\[10088]  & (~\[10073]  & (~v15 & ~\[12466] )),
  \[416]  = ~\[13648]  & (~v3 & (~\[13651]  & ~\[13657] )),
  \[21691]  = ~v7 | (~\[10236]  | (~\[8808]  | ~\[8800] )),
  \[3940]  = ~\[10058]  & (~v10 & (~v12 & ~\[13110] )),
  \[12970]  = ~v1 | ~\[10099] ,
  \[417]  = ~\[10072]  & (~v14 & (~\[13663]  & ~\[13661] )),
  \[10919]  = ~v12 | (~v14 | (~\[10076]  | ~\[8331] )),
  \[14298]  = ~v10 | ~v9,
  \[22153]  = ~v4 | (~v7 | (~\[4306]  | ~\[4298] )),
  \[14297]  = ~v2 | (~\[10059]  | (~\[10176]  | ~\[1597] )),
  \[11044]  = ~v4 | ~\[10135] ,
  \[3214]  = ~\[10060]  & (~v1 & ~v3),
  \[10913]  = ~v5 | (~\[10134]  | ~v6),
  \[22155]  = ~v4 | (~v7 | (~\[4288]  | ~\[4280] )),
  \[4074]  = ~\[10058]  & (~v10 & (~v12 & ~\[13060] )),
  \[11773]  = ~v1 | (~\[10099]  | ~v3),
  \[13434]  = ~v2 | (~\[10059]  | ~\[10176] ),
  \[6463]  = ~\[10060]  & (~v1 & (~v3 & ~\[11868] )),
  \[9319]  = ~\[10059]  & (~v0 & (~v2 & ~\[10441] )),
  \[21697]  = ~v4 | (~\[10135]  | (~\[8754]  | ~\[8746] )),
  \[11775]  = ~v5 | (~\[10134]  | ~v6),
  \[2750]  = ~\[10072]  & (~v12 & ~v14),
  \[1559]  = ~\[10060]  & (~v1 & (~v3 & ~\[14328] )),
  \[3948]  = ~\[10060]  & (~v1 & ~v3),
  \[8854]  = ~\[10073]  & (~v15 & ~\[10672] ),
  \[13440]  = ~v15 | (~v13 | ~\[3321] ),
  \[12247]  = ~v5 | (~\[10134]  | ~v6),
  \[10921]  = ~v2 | (~\[10059]  | ~\[10176] ),
  \[21693]  = ~v14 | (~\[10076]  | (~\[8781]  | ~\[8791] )),
  \[11051]  = ~\[21765]  | (~\[21763]  | (~\[21761]  | ~\[21759] )),
  \[5271]  = ~\[10236]  & (~\[10135]  & ~v7),
  \[11781]  = ~v14 | (~\[10072]  | (~\[10076]  | ~\[6653] )),
  \[6800]  = ~\[10073]  & (~v13 & ~v15),
  \[10584]  = ~v0 | (~v2 | (~\[10176]  | ~\[9027] )),
  \[13442]  = ~v0 | (~v2 | ~\[10176] ),
  \[12979]  = ~v13 | (~\[10088]  | (~v15 | ~\[4259] )),
  \[21695]  = ~v14 | (~\[10076]  | (~\[8763]  | ~\[8773] )),
  \[2755]  = ~\[10058]  & (~v7 & ~v10),
  \[10586]  = ~v11 | (~v8 | ~v12),
  \[8129]  = ~v6 & (~v5 & ~\[11035] ),
  \[12243]  = ~\[22019]  | (~\[22017]  | (~\[22015]  | ~\[22013] )),
  \[12973]  = ~v5 | (~\[10134]  | ~v6),
  \[7663]  = ~v6 & (~v5 & (~\[11266]  & ~v3)),
  \[22167]  = ~v15 | (~v13 | (~\[4163]  | ~\[4173] )),
  \[10927]  = ~v14 | (~\[10076]  | (~\[8368]  | ~v12)),
  \[22169]  = ~v7 | (~\[10236]  | (~\[4154]  | ~\[4146] )),
  \[11787]  = ~v1 | (~\[10099]  | ~v3),
  \[13448]  = ~v15 | (~v13 | ~\[3303] ),
  \[5278]  = ~v4 & (~v3 & (~\[10060]  & ~v1)),
  \[10929]  = ~v0 | (~v2 | ~\[10176] ),
  \[22163]  = ~v15 | (~v13 | (~\[4199]  | ~\[4209] )),
  \[4082]  = ~\[10060]  & (~v1 & ~v3),
  \[3223]  = ~\[10068]  & (~v9 & ~v12),
  \[0]  = ~\[794]  | (~\[1033]  | (~\[1273]  | ~\[1514] )),
  \[6471]  = ~\[10058]  & (~v10 & ~v13),
  \[12981]  = ~v1 | (~\[10099]  | ~v3),
  \[5612]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[11053]  = ~v1 | (~\[10099]  | ~v3),
  \[22165]  = ~v4 | (~\[10135]  | (~\[4190]  | ~\[4182] )),
  \[9328]  = ~\[10073]  & (~v15 & ~\[10435] ),
  \[8862]  = ~\[10059]  & (~v0 & ~v2),
  \[10597]  = ~v8 | (~\[10064]  | ~v12),
  \[2031]  = ~\[10133]  & (~v5 & ~v8),
  \[3958]  = ~v10 & (~v9 & (~v12 & ~\[13126] )),
  \[22171]  = ~v15 | (~v13 | (~\[4127]  | ~\[4137] )),
  \[12257]  = ~v5 | (~\[10134]  | ~v6),
  \[11061]  = ~v1 | (~\[10099]  | ~v3),
  \[4422]  = ~\[10060]  & (~v1 & ~v3),
  \[8137]  = ~v10 & (~v9 & ~v13),
  \[12989]  = ~v13 | (~\[10088]  | (~v15 | ~\[4237] )),
  \[13451]  = ~v2 | ~\[10059] ,
  \[7671]  = ~v10 & (~v9 & ~v12),
  \[12983]  = ~v5 | (~\[10134]  | ~v6),
  \[2767]  = ~\[10059]  & (~v0 & (~v2 & ~\[13718] )),
  \[1570]  = ~\[10072]  & (~v12 & (~v14 & ~\[14321] )),
  \[22177]  = ~v4 | (~\[10135]  | (~\[4082]  | ~\[4074] )),
  \[436]  = ~\[13838]  & (~v3 & (~\[13841]  & ~\[13847] )),
  \[22179]  = ~v15 | (~v13 | (~\[4055]  | ~\[4065] )),
  \[437]  = ~\[10133]  & (~v5 & (~\[13849]  & ~\[13855] )),
  \[4091]  = ~\[10058]  & (~v10 & ~v12),
  \[438]  = ~\[10133]  & (~v5 & (~\[13858]  & ~\[13864] )),
  \[22173]  = ~v15 | (~v13 | (~\[4109]  | ~\[4119] )),
  \[439]  = ~\[10072]  & (~v14 & (~\[13870]  & ~\[13868] )),
  \[9336]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[6481]  = ~\[10134]  & (~v6 & (~\[11857]  & ~v3)),
  \[10206]  = ~v14 | (~v13 | ~\[10076] ),
  \[22175]  = ~v15 | (~v13 | (~\[4091]  | ~\[4101] )),
  \[13454]  = ~v5 | (~\[10134]  | ~v6),
  \[8871]  = ~\[10058]  & (~v10 & ~\[10088] ),
  \[11796]  = ~v4 | ~\[10135] ,
  \[10935]  = ~v14 | (~\[10076]  | (~\[8350]  | ~v12)),
  \[3966]  = ~\[10059]  & (~v0 & ~v2),
  \[11070]  = ~v7 | ~\[10236] ,
  \[11407]  = ~v11 | (~\[10063]  | ~v12),
  \[22181]  = ~\[4029]  | (~v15 | (~\[4035]  | ~\[4047] )),
  \[13460]  = ~v13 | (~\[10088]  | (~v15 | ~\[3283] )),
  \[12267]  = ~v7 | ~\[10236] ,
  \[10211]  = ~v3 | ~v0,
  \[5290]  = ~\[10088]  & (~\[10073]  & (~v15 & ~\[12454] )),
  \[440]  = ~\[10072]  & (~v14 & (~\[13880]  & ~\[13878] )),
  \[4431]  = ~\[10068]  & (~\[10058]  & ~v12),
  \[441]  = ~\[13888]  & (~v11 & (~\[13891]  & ~\[13887] )),
  \[8147]  = ~v6 & (~v5 & (~\[11025]  & ~v2)),
  \[6489]  = ~\[10058]  & (~v10 & ~v13),
  \[442]  = ~\[13899]  & (~v11 & (~\[13902]  & ~\[13898] )),
  \[13461]  = ~v0 | ~v2,
  \[2775]  = ~\[10058]  & (~v10 & ~v12),
  \[7681]  = ~\[10133]  & (~v5 & ~\[11259] ),
  \[443]  = ~\[13915]  & ~\[13909] ,
  \[6822]  = ~\[10073]  & (~v13 & ~v15),
  \[11405]  = ~v1 | (~\[10099]  | (~\[10060]  | ~\[7389] )),
  \[22187]  = ~v15 | (~v13 | (~\[3975]  | ~\[3985] )),
  \[10948]  = ~v12 | (~v14 | ~\[10076] ),
  \[1581]  = ~\[10133]  & (~v5 & (~v8 & ~\[14316] )),
  \[12995]  = ~v1 | (~\[10099]  | ~v3),
  \[11077]  = ~\[21769]  | (~\[21767]  | ~\[21771] ),
  \[22189]  = ~v4 | (~v7 | (~\[3966]  | ~\[3958] )),
  \[3241]  = ~\[10068]  & (~v9 & ~v12),
  \[12607]  = ~v14 | (~\[10072]  | ~\[10076] ),
  \[448]  = ~\[13979]  & (~v11 & (~\[13982]  & ~\[13978] )),
  \[5630]  = ~\[10060]  & (~v1 & ~v3),
  \[22183]  = ~\[4007]  | (~v15 | (~\[4013]  | ~\[4025] )),
  \[449]  = ~\[13989]  & (~v11 & (~\[13992]  & ~\[13988] )),
  \[9346]  = ~\[10073]  & (~v15 & ~\[10426] ),
  \[12604]  = ~v10 | ~v9,
  \[7689]  = ~v10 & (~v9 & ~v12),
  \[22185]  = ~v7 | (~\[10236]  | (~\[4002]  | ~\[3994] )),
  \[13464]  = ~v5 | (~\[10134]  | ~v6),
  \[3975]  = ~\[10058]  & (~v10 & ~v12),
  \[8881]  = ~v6 & (~v5 & ~\[10660] ),
  \[12603]  = ~v1 | (~\[10099]  | (~\[10060]  | ~\[4993] )),
  \[10215]  = ~v3 | ~v0,
  \[8152]  = ~\[10073]  & (~v13 & ~v15),
  \[11080]  = ~\[1261]  | (~\[1268]  | (~\[1254]  | ~\[1241] )),
  \[22191]  = ~v4 | (~v7 | (~\[3948]  | ~\[3940] )),
  \[10952]  = ~v7 | ~\[10236] ,
  \[13470]  = ~v13 | (~\[10088]  | (~v15 | ~\[3261] )),
  \[11082]  = ~v2 | (~\[10059]  | ~\[10176] ),
  \[450]  = ~\[13969]  & (~v11 & (~\[13972]  & ~\[13968] )),
  \[2053]  = ~\[10133]  & (~v5 & ~v8),
  \[13807]  = ~\[22335]  | (~\[22333]  | (~\[22331]  | ~\[22329] )),
  \[451]  = ~\[14004]  & (~v11 & (~\[14007]  & ~\[14003] )),
  \[5639]  = ~\[10068]  & (~v9 & ~v12),
  \[8157]  = ~v9 & (~v7 & ~v10),
  \[6499]  = ~\[10060]  & (~v1 & (~v3 & ~\[11848] )),
  \[452]  = ~\[14014]  & (~v11 & (~\[14017]  & ~\[14013] )),
  \[2785]  = ~\[10059]  & (~v0 & (~\[10176]  & ~\[13708] )),
  \[11413]  = ~v1 | (~\[10099]  | (~v3 | ~\[7371] )),
  \[1926]  = ~v4 & (~v2 & (~\[10059]  & ~v0)),
  \[453]  = ~\[14025]  & (~v11 & (~\[14028]  & ~\[14024] )),
  \[12273]  = ~v0 | ~v2,
  \[454]  = ~\[14035]  & (~v11 & (~\[14038]  & ~\[14034] )),
  \[11415]  = ~v11 | (~\[10063]  | ~v12),
  \[455]  = ~\[14053]  & ~\[14047] ,
  \[11088]  = ~v14 | (~\[10076]  | ~\[8029] ),
  \[6105]  = ~\[10134]  & (~v6 & (~\[12056]  & ~v3)),
  \[456]  = ~\[14057]  & (~v7 & (~\[14056]  & ~\[14065] )),
  \[457]  = ~\[14072]  & (~v11 & (~\[14075]  & ~\[14071] )),
  \[9354]  = ~\[10059]  & (~v0 & ~v2),
  \[12617]  = ~v14 | (~\[10072]  | ~\[10076] ),
  \[11422]  = ~v4 | (~\[10135]  | ~\[7358] ),
  \[458]  = ~\[14082]  & (~v11 & (~\[14085]  & ~\[14081] )),
  \[10959]  = ~v0 | ~v2,
  \[12282]  = ~\[22027]  | (~\[22025]  | (~\[22023]  | ~\[22021] )),
  \[6838]  = ~\[10060]  & (~v1 & ~v3),
  \[13479]  = ~v15 | (~v13 | ~\[3241] ),
  \[13811]  = ~v5 | (~\[10134]  | ~v6),
  \[12614]  = ~v10 | ~v9,
  \[7699]  = ~\[10059]  & (~v0 & (~v2 & ~\[11250] )),
  \[3985]  = ~\[10133]  & (~v5 & (~\[13112]  & ~v3)),
  \[1597]  = ~\[10133]  & (~v5 & ~v8),
  \[12613]  = ~v1 | (~\[10099]  | (~v3 | ~\[4971] )),
  \[13473]  = ~v2 | (~\[10059]  | ~\[10176] ),
  \[7304]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[11090]  = ~v0 | (~v2 | ~\[10176] ),
  \[8893]  = ~v6 & ~v5,
  \[1202]  = ~\[158]  & (~\[157]  & (~\[156]  & ~\[155] )),
  \[12287]  = ~v4 | (~v7 | ~\[5630] ),
  \[5649]  = ~\[10133]  & (~v5 & (~\[12273]  & ~v3)),
  \[12289]  = ~v11 | (~\[10063]  | ~\[10088] ),
  \[2794]  = ~\[10072]  & (~v14 & (~\[13702]  & ~v12)),
  \[11424]  = ~v11 | (~\[10063]  | ~v12),
  \[13481]  = ~v0 | (~v2 | ~\[10176] ),
  \[463]  = ~\[14152]  & (~v14 & (~\[14151]  & ~\[14148] )),
  \[9360]  = ~\[10088]  & (~v3 & ~v14),
  \[8169]  = ~\[10059]  & (~v0 & (~\[10176]  & ~\[11018] )),
  \[6113]  = ~\[10068]  & (~v9 & ~v13),
  \[464]  = ~\[14158]  & (~v7 & (~\[14157]  & ~\[14166] )),
  \[10238]  = ~v6 | (~\[10236]  | ~\[10133] ),
  \[1938]  = ~\[10072]  & (~v12 & (~v14 & ~\[14127] )),
  \[465]  = ~\[14138]  & (~v11 & (~\[14141]  & ~\[14137] )),
  \[1209]  = ~\[154]  & (~\[153]  & (~\[152]  & ~\[151] )),
  \[11430]  = ~v1 | (~\[10099]  | (~v3 | ~\[7335] )),
  \[12628]  = ~v10 | (~v9 | ~\[10068] ),
  \[4458]  = ~\[10060]  & (~v1 & ~v3),
  \[3261]  = ~v9 & (~v7 & ~\[10068] ),
  \[13820]  = ~v4 | ~\[10135] ,
  \[11432]  = ~v11 | (~\[10063]  | ~v12),
  \[10969]  = ~v4 | ~v7,
  \[13487]  = ~v15 | (~v13 | ~\[3223] ),
  \[11099]  = ~v2 | (~\[10059]  | ~\[10176] ),
  \[2404]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[3994]  = ~\[10058]  & (~v10 & (~v12 & ~\[13100] )),
  \[10236]  = ~v5,
  \[11096]  = ~v14 | (~\[10076]  | ~\[8011] ),
  \[10235]  = ~\[21555]  | (~\[21553]  | (~\[21551]  | ~\[21549] )),
  \[7314]  = ~\[10073]  & (~v15 & ~\[11443] ),
  \[2071]  = ~\[10064]  & (~v11 & (~\[10063]  & ~v8)),
  \[8174]  = ~\[10073]  & (~v13 & ~v15),
  \[10242]  = ~v3 | (~v0 | ~\[10088] ),
  \[5657]  = ~\[10068]  & (~v9 & ~v12),
  \[12297]  = ~v11 | (~\[10063]  | ~\[10088] ),
  \[6851]  = ~\[10134]  & ~v6,
  \[8179]  = ~v9 & (~v7 & ~v10),
  \[6123]  = ~\[10060]  & (~v1 & (~v3 & ~\[12050] )),
  \[474]  = ~\[14263]  & (~v11 & (~\[14266]  & ~\[14262] )),
  \[8512]  = ~v10 & ~v9,
  \[475]  = ~\[14277]  & (~v14 & (~\[14276]  & ~\[14273] )),
  \[9372]  = ~\[10073]  & (~v15 & (~\[10072]  & ~v12)),
  \[12295]  = ~v4 | (~v7 | ~\[5612] ),
  \[13826]  = ~v0 | ~v2,
  \[1949]  = ~\[10059]  & (~v0 & (~\[10176]  & ~\[14124] )),
  \[476]  = ~\[14284]  & (~v7 & (~\[14283]  & ~\[14292] )),
  \[4467]  = ~\[10068]  & (~\[10058]  & ~v12),
  \[12638]  = ~v10 | (~v9 | ~\[10068] ),
  \[477]  = ~\[14298]  & (~v11 & (~\[14301]  & ~\[14297] )),
  \[13100]  = ~v15 | ~v13,
  \[3609]  = ~\[10133]  & (~v5 & (~\[13294]  & ~v3)),
  \[10979]  = ~v4 | ~v7,
  \[13497]  = ~v15 | ~v13,
  \[10976]  = ~\[21749]  | (~\[21747]  | (~\[21745]  | ~\[21743] )),
  \[7322]  = ~\[10059]  & (~v0 & ~v2),
  \[9379]  = ~\[10060]  & (~v3 & (~\[10059]  & ~v0)),
  \[5667]  = ~\[10060]  & (~v1 & (~v3 & ~\[12267] )),
  \[13838]  = ~v0 | ~v2,
  \[6131]  = ~\[10068]  & (~v9 & ~v13),
  \[11443]  = ~v11 | (~\[10063]  | ~v12),
  \[14301]  = ~v13 | (~\[10088]  | ~\[10073] ),
  \[13103]  = ~\[22185]  | (~\[22183]  | (~\[22181]  | ~\[22179] )),
  \[10987]  = ~v4 | ~v7,
  \[3618]  = ~v10 & (~v9 & (~v12 & ~\[13291] )),
  \[13835]  = ~\[22339]  | (~\[22337]  | ~\[22341] ),
  \[13110]  = ~v15 | ~v13,
  \[14308]  = ~v4 | (~v7 | ~\[10058] ),
  \[11451]  = ~v11 | (~\[10063]  | ~v12),
  \[3283]  = ~v9 & (~v7 & ~\[10068] ),
  \[13112]  = ~v0 | ~v2,
  \[12649]  = ~v10 | (~v9 | ~\[10068] ),
  \[5672]  = ~\[10072]  & (~v12 & ~v14),
  \[13841]  = ~v5 | (~\[10134]  | ~v6),
  \[823]  = ~\[13129]  & (~\[13103]  & (~\[13063]  & ~\[13028] )),
  \[8191]  = ~\[10059]  & (~v0 & (~v2 & ~\[11005] )),
  \[2426]  = ~\[10059]  & (~v0 & ~v2),
  \[9389]  = ~\[10059]  & (~v0 & ~\[10060] ),
  \[21707]  = ~v14 | (~\[10076]  | (~\[8647]  | ~\[8657] )),
  \[1960]  = ~\[10072]  & (~v12 & (~\[10076]  & ~\[14117] )),
  \[5676]  = ~v9 & ~v7,
  \[21709]  = ~v14 | (~\[10076]  | (~\[8629]  | ~\[8639] )),
  \[7335]  = ~\[10134]  & ~v6,
  \[13847]  = ~v13 | (~\[10088]  | (~\[10073]  | ~\[2509] )),
  \[6141]  = ~v6 & (~v5 & (~\[12028]  & ~v3)),
  \[13849]  = ~v2 | (~\[10059]  | ~\[10176] ),
  \[14311]  = ~v10 | (~v9 | ~\[10068] ),
  \[8199]  = ~v10 & (~v9 & ~v13),
  \[4485]  = ~\[10068]  & (~\[10058]  & ~v12),
  \[2097]  = ~\[10064]  & (~v11 & (~\[10063]  & ~v8)),
  \[3626]  = ~\[10060]  & (~v1 & ~v3),
  \[11455]  = ~v2 | ~\[10059] ,
  \[6874]  = ~\[10060]  & (~v1 & ~v3),
  \[8533]  = ~v9 & (~v7 & ~v10),
  \[10267]  = ~\[21569]  | (~\[21567]  | (~\[21565]  | ~\[21563] )),
  \[21711]  = ~v4 | (~v7 | (~\[8620]  | ~\[8612] )),
  \[4822]  = ~v4 & (~v3 & (~\[10060]  & ~v1)),
  \[6149]  = ~\[10068]  & (~v9 & ~v13),
  \[12659]  = ~v10 | (~v9 | ~\[10068] ),
  \[12654]  = ~v0 | (~v2 | ~\[10176] ),
  \[103]  = ~\[10635]  & (~v2 & (~\[10638]  & ~\[10644] )),
  \[10996]  = ~v4 | ~v7,
  \[104]  = ~\[10648]  & (~\[10646]  & ~\[10654] ),
  \[105]  = ~\[10073]  & (~v15 & (~\[10632]  & ~\[10630] )),
  \[1241]  = ~\[11077]  & (~\[11051]  & (~\[11013]  & ~\[10976] )),
  \[1971]  = ~\[10099]  & (~\[10060]  & (~v3 & ~\[14114] )),
  \[836]  = ~\[344]  & (~\[343]  & (~\[345]  & ~\[12961] )),
  \[14316]  = ~v0 | (~v2 | ~\[10176] ),
  \[13858]  = ~v0 | (~v2 | ~\[10176] ),
  \[5689]  = ~\[10099]  & (~\[10060]  & (~v3 & ~\[12257] )),
  \[9006]  = ~\[10073]  & (~v15 & ~\[10597] ),
  \[13129]  = ~\[22189]  | (~\[22187]  | ~\[22191] ),
  \[11463]  = ~v0 | ~v2,
  \[14321]  = ~v10 | (~v9 | ~\[10068] ),
  \[10605]  = ~v11 | (~v8 | ~v12),
  \[9739]  = ~\[10176]  & (~\[10099]  & ~v8),
  \[13126]  = ~v15 | ~v13,
  \[3638]  = ~v9 & (~v7 & (~v10 & ~\[13283] )),
  \[13855]  = ~v13 | (~\[10073]  | ~\[2489] ),
  \[11472]  = ~\[21855]  | (~\[21853]  | (~\[21851]  | ~\[21849] )),
  \[4101]  = ~v6 & (~v5 & (~\[13046]  & ~v3)),
  \[6887]  = ~v6 & ~v5,
  \[14328]  = ~v4 | (~v7 | ~\[10058] ),
  \[13132]  = ~\[843]  | (~\[850]  | (~\[836]  | ~\[823] )),
  \[2444]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[6159]  = ~v6 & (~v5 & (~\[12020]  & ~v3)),
  \[11804]  = ~v1 | (~\[10099]  | ~v3),
  \[12664]  = ~\[22095]  | (~\[22093]  | (~\[22091]  | ~\[22089] )),
  \[843]  = ~\[338]  & (~\[337]  & (~\[336]  & ~\[335] )),
  \[114]  = ~\[10073]  & (~v15 & (~\[10735]  & ~\[10733] )),
  \[5694]  = ~\[10072]  & (~v12 & ~v14),
  \[115]  = ~\[10738]  & (~v3 & (~\[10741]  & ~\[10747] )),
  \[9742]  = ~\[10064]  & ~v11,
  \[116]  = ~\[10749]  & (~v3 & (~\[10752]  & ~\[10758] )),
  \[21729]  = ~v14 | (~\[10076]  | (~\[8441]  | ~\[8451] )),
  \[12670]  = ~v5 | (~v6 | (~\[10133]  | ~\[4822] )),
  \[117]  = ~\[10073]  & (~v15 & (~\[10764]  & ~\[10762] )),
  \[1982]  = ~\[10072]  & (~v12 & (~\[10076]  & ~\[14106] )),
  \[9014]  = ~\[10059]  & (~v0 & ~v2),
  \[13868]  = ~v4 | (~v7 | ~\[2462] ),
  \[4109]  = ~\[10058]  & (~v10 & ~v12),
  \[5698]  = ~v9 & ~v7,
  \[4839]  = ~\[10134]  & (~v6 & ~v8),
  \[3642]  = ~\[10236]  & ~v4,
  \[1254]  = ~\[134]  & (~\[133]  & (~\[135]  & ~\[10909] )),
  \[5301]  = ~\[10134]  & (~v6 & (~v8 & ~\[12449] )),
  \[10614]  = ~v11 | (~v8 | ~v12),
  \[7358]  = ~\[10059]  & (~v0 & ~v2),
  \[11473]  = ~v2 | ~\[10059] ,
  \[14331]  = ~v10 | (~v9 | ~\[10068] ),
  \[13864]  = ~v13 | (~\[10073]  | ~\[2471] ),
  \[11476]  = ~v5 | (~\[10134]  | ~v6),
  \[10288]  = ~v5 | (~\[10134]  | ~\[10135] ),
  \[13136]  = ~v0 | (~v2 | ~\[10176] ),
  \[21731]  = ~v14 | (~\[10076]  | (~\[8423]  | ~\[8433] )),
  \[3648]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[10622]  = ~v8 | (~\[10064]  | ~v12),
  \[8555]  = ~v9 & (~v7 & ~v10),
  \[6167]  = ~\[10068]  & (~v9 & ~v13),
  \[13870]  = ~v8 | (~\[10064]  | ~\[10088] ),
  \[11482]  = ~v12 | (~v14 | (~\[10076]  | ~\[7203] )),
  \[850]  = ~\[334]  & (~\[333]  & (~\[332]  & ~\[331] )),
  \[121]  = ~\[10073]  & (~v15 & (~\[10805]  & ~\[10803] )),
  \[14337]  = ~\[22429]  | (~\[22427]  | (~\[22431]  | ~\[567] )),
  \[13142]  = ~v15 | (~v13 | ~\[3921] ),
  \[122]  = ~\[10134]  & (~\[10133]  & (~\[10809]  & ~\[10815] )),
  \[12674]  = ~v14 | ~\[10072] ,
  \[123]  = ~\[10817]  & (~v2 & (~\[10820]  & ~\[10826] )),
  \[11813]  = ~v7 | ~\[10236] ,
  \[14339]  = ~\[604]  | (~\[611]  | (~\[597]  | ~\[584] )),
  \[12673]  = ~v10 | (~\[10068]  | (~v9 | ~\[10058] )),
  \[124]  = ~\[10830]  & (~\[10828]  & ~\[10836] ),
  \[10285]  = ~\[21577]  | (~\[21575]  | (~\[21573]  | ~\[21571] )),
  \[125]  = ~v6 & (~v5 & (~\[10840]  & ~\[10846] )),
  \[1261]  = ~\[128]  & (~\[127]  & (~\[126]  & ~\[125] )),
  \[11488]  = ~v11 | (~\[10063]  | ~v12),
  \[126]  = ~v6 & (~v5 & (~\[10848]  & ~\[10854] )),
  \[11820]  = ~\[21929]  | (~\[21927]  | (~\[21925]  | ~\[21923] )),
  \[127]  = ~\[10134]  & (~v6 & (~\[10857]  & ~\[10863] )),
  \[10292]  = ~v5 | (~\[10134]  | ~\[10135] ),
  \[13878]  = ~v4 | (~v7 | ~\[2444] ),
  \[128]  = ~\[10134]  & (~v6 & (~\[10865]  & ~\[10871] )),
  \[6507]  = ~\[10058]  & (~v10 & ~v13),
  \[1993]  = ~\[10060]  & (~v1 & (~v3 & ~\[14103] )),
  \[4119]  = ~v6 & (~v5 & (~\[13037]  & ~v3)),
  \[11822]  = ~v1 | (~\[10099]  | ~v3),
  \[21733]  = ~v14 | (~\[10076]  | (~\[8405]  | ~\[8415] )),
  \[12682]  = ~v10 | ~v9,
  \[12681]  = ~v2 | (~\[10059]  | (~\[10176]  | ~\[4861] )),
  \[9027]  = ~\[10133]  & ~v5,
  \[21735]  = ~v14 | (~\[10076]  | (~\[8387]  | ~\[8397] )),
  \[10626]  = ~\[21675]  | (~\[21673]  | (~\[21671]  | ~\[21669] )),
  \[13144]  = ~v1 | (~\[10099]  | ~v3),
  \[11486]  = ~v4 | (~\[10135]  | ~\[7250] ),
  \[1268]  = ~\[124]  & (~\[123]  & (~\[122]  & ~\[121] )),
  \[10630]  = ~v1 | (~\[10099]  | (~\[10060]  | ~\[8893] )),
  \[22209]  = ~v7 | (~\[10236]  | (~\[3778]  | ~\[3770] )),
  \[5317]  = ~\[10134]  & (~v6 & ~v8),
  \[10632]  = ~v8 | (~\[10064]  | ~v12),
  \[13150]  = ~v15 | (~v13 | ~\[3903] ),
  \[3659]  = ~v9 & (~v7 & ~v10),
  \[2462]  = ~\[10060]  & (~v1 & ~v3),
  \[6177]  = ~\[10133]  & (~v5 & ~\[12012] ),
  \[13880]  = ~v8 | (~\[10064]  | ~\[10088] ),
  \[10299]  = ~v5 | ~\[10134] ,
  \[7707]  = ~v10 & (~v9 & ~v12),
  \[11829]  = ~v2 | ~\[10059] ,
  \[13152]  = ~v1 | ~\[10099] ,
  \[7371]  = ~v6 & ~v5,
  \[133]  = ~\[10134]  & (~v6 & (~\[10921]  & ~\[10927] )),
  \[10296]  = ~v5 | ~\[10134] ,
  \[134]  = ~\[10134]  & (~v6 & (~\[10929]  & ~\[10935] )),
  \[21747]  = ~v14 | (~\[10076]  | (~\[8271]  | ~\[8281] )),
  \[135]  = ~\[10910]  & (~v3 & (~\[10913]  & ~\[10919] )),
  \[10638]  = ~v5 | (~\[10134]  | ~v6),
  \[12685]  = ~v14 | (~\[10072]  | ~\[10076] ),
  \[4127]  = ~\[10058]  & (~v10 & ~v12),
  \[21749]  = ~v14 | (~\[10076]  | (~\[8253]  | ~\[8263] )),
  \[22211]  = ~v15 | (~v13 | (~\[3751]  | ~\[3761] )),
  \[1273]  = ~\[11924]  & (~\[11643]  & (~\[11361]  & ~\[11080] )),
  \[2802]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[13888]  = ~v10 | ~v9,
  \[6517]  = ~v6 & (~v5 & (~\[11838]  & ~v3)),
  \[21743]  = ~\[8314]  | (~v6 | (~\[8320]  | ~\[8310] )),
  \[13887]  = ~v4 | (~v7 | (~\[10058]  | ~\[2426] )),
  \[12692]  = ~v10 | ~v9,
  \[12691]  = ~v0 | (~v2 | (~\[10176]  | ~\[4839] )),
  \[11494]  = ~v0 | (~v2 | (~\[10176]  | ~\[7227] )),
  \[21745]  = ~v14 | (~\[10076]  | (~\[8289]  | ~\[8299] )),
  \[8909]  = ~\[10058]  & (~v7 & ~v10),
  \[11496]  = ~v11 | (~\[10063]  | ~v12),
  \[10635]  = ~v1 | ~\[10099] ,
  \[6185]  = ~\[10068]  & (~v9 & ~v13),
  \[11838]  = ~v0 | ~v2,
  \[13155]  = ~v5 | (~\[10134]  | ~v6),
  \[21751]  = ~v14 | (~\[10076]  | (~\[8235]  | ~\[8245] )),
  \[2471]  = ~\[10058]  & (~v10 & ~v12),
  \[8574]  = ~v10 & ~v9,
  \[11107]  = ~v0 | (~v2 | ~\[10176] ),
  \[4861]  = ~\[10134]  & (~v6 & ~v8),
  \[7717]  = ~\[10134]  & (~v6 & ~\[11241] ),
  \[22213]  = ~v15 | (~v13 | (~\[3733]  | ~\[3743] )),
  \[1615]  = ~\[10064]  & (~v11 & (~\[10063]  & ~v8)),
  \[13161]  = ~v13 | (~\[10088]  | (~v15 | ~\[3883] )),
  \[13891]  = ~v13 | (~\[10088]  | ~v15),
  \[22215]  = ~v15 | (~v13 | (~\[3715]  | ~\[3725] )),
  \[21757]  = ~\[8174]  | (~\[8179]  | ~\[8191] ),
  \[11105]  = ~v14 | (~\[10076]  | ~\[7993] ),
  \[10648]  = ~v5 | (~\[10134]  | ~v6),
  \[12695]  = ~v14 | (~\[10072]  | ~\[10076] ),
  \[6525]  = ~\[10058]  & (~v10 & ~v13),
  \[4137]  = ~\[10133]  & (~v5 & ~\[13030] ),
  \[21759]  = ~\[8152]  | (~\[8157]  | ~\[8169] ),
  \[2812]  = ~\[10072]  & (~v14 & (~\[13672]  & ~v12)),
  \[13898]  = ~v4 | (~v7 | (~\[10058]  | ~\[2404] )),
  \[21753]  = ~v14 | (~\[10076]  | (~\[8217]  | ~\[8227] )),
  \[10644]  = ~v12 | (~v14 | (~\[10076]  | ~\[8931] )),
  \[1285]  = ~\[117]  & (~\[116]  & (~\[115]  & ~\[114] )),
  \[12309]  = ~v12 | (~v14 | ~\[10076] ),
  \[21755]  = ~v14 | (~\[10076]  | (~\[8199]  | ~\[8209] )),
  \[7389]  = ~v6 & ~v5,
  \[13899]  = ~v10 | ~v9,
  \[10646]  = ~v1 | (~\[10099]  | ~v3),
  \[13163]  = ~v1 | (~\[10099]  | ~v3),
  \[12306]  = ~v10 | ~v9,
  \[22227]  = ~v15 | (~v13 | (~\[3599]  | ~\[3609] )),
  \[12305]  = ~v4 | (~v7 | (~\[10058]  | ~\[5594] )),
  \[6195]  = ~\[10059]  & (~v0 & (~v2 & ~\[12005] )),
  \[11848]  = ~v4 | ~\[10135] ,
  \[13165]  = ~v5 | (~\[10134]  | ~v6),
  \[21761]  = ~v14 | (~\[10076]  | (~\[8137]  | ~\[8147] )),
  \[7725]  = ~v10 & (~v9 & ~v12),
  \[22229]  = ~v4 | (~v7 | (~\[3590]  | ~\[3582] )),
  \[3679]  = ~v10 & (~v9 & ~v12),
  \[11119]  = ~v5 | (~\[10134]  | ~v6),
  \[151]  = ~v6 & (~v5 & (~\[11082]  & ~\[11088] )),
  \[22223]  = ~\[3642]  | (~v6 | (~\[3648]  | ~\[3638] )),
  \[5339]  = ~v6 & (~v5 & ~v8),
  \[152]  = ~v6 & (~v5 & (~\[11090]  & ~\[11096] )),
  \[882]  = ~\[12848]  & (~\[12822]  & (~\[12784]  & ~\[12745] )),
  \[13171]  = ~v13 | (~\[10088]  | (~v15 | ~\[3861] )),
  \[11113]  = ~v14 | (~\[10076]  | ~\[7975] ),
  \[153]  = ~\[10134]  & (~v6 & (~\[11099]  & ~\[11105] )),
  \[22225]  = ~v7 | (~\[10236]  | (~\[3626]  | ~\[3618] )),
  \[9050]  = ~\[10060]  & (~v1 & ~v3),
  \[11116]  = ~v2 | ~\[10059] ,
  \[154]  = ~\[10134]  & (~v6 & (~\[11107]  & ~\[11113] )),
  \[21767]  = ~v14 | (~\[10076]  | (~\[8083]  | ~\[8093] )),
  \[155]  = ~\[11116]  & (~v3 & (~\[11119]  & ~\[11125] )),
  \[4146]  = ~\[10058]  & (~v10 & (~v12 & ~\[13025] )),
  \[2820]  = ~\[10060]  & (~v1 & ~v3),
  \[156]  = ~\[11126]  & (~v3 & (~\[11129]  & ~\[11135] )),
  \[6535]  = ~v6 & (~v5 & (~\[11829]  & ~v3)),
  \[21769]  = ~v14 | (~\[10076]  | (~\[8065]  | ~\[8075] )),
  \[2489]  = ~\[10058]  & (~v10 & ~v12),
  \[13505]  = ~v15 | ~v13,
  \[157]  = ~\[10133]  & (~v5 & (~\[11138]  & ~\[11144] )),
  \[22231]  = ~v4 | (~v7 | (~\[3572]  | ~\[3564] )),
  \[4878]  = ~\[10073]  & (~v13 & (~v15 & ~\[12659] )),
  \[158]  = ~\[10133]  & (~v5 & (~\[11146]  & ~\[11152] )),
  \[21763]  = ~v14 | (~\[10076]  | (~\[8119]  | ~\[8129] )),
  \[10654]  = ~v12 | (~v14 | (~\[10076]  | ~\[8909] )),
  \[13512]  = ~v11 | ~v8,
  \[12319]  = ~v12 | (~v14 | ~\[10076] ),
  \[21765]  = ~v14 | (~\[10076]  | (~\[8101]  | ~\[8111] )),
  \[12316]  = ~v10 | ~v9,
  \[22237]  = ~\[3506]  | (~v11 | (~\[3502]  | ~\[3519] )),
  \[10660]  = ~v1 | (~\[10099]  | ~v3),
  \[12315]  = ~v4 | (~v7 | (~\[10058]  | ~\[5572] )),
  \[13175]  = ~v1 | (~\[10099]  | ~\[10060] ),
  \[21771]  = ~v14 | (~\[10076]  | (~\[8047]  | ~\[8057] )),
  \[2829]  = ~\[10058]  & (~v10 & ~v12),
  \[7735]  = ~\[10059]  & (~v0 & (~v2 & ~\[11233] )),
  \[22239]  = ~\[3484]  | (~v11 | (~\[3480]  | ~\[3497] )),
  \[11857]  = ~v0 | ~v2,
  \[11129]  = ~v5 | (~\[10134]  | ~v6),
  \[22233]  = ~v4 | (~v7 | (~\[3554]  | ~\[3546] )),
  \[13181]  = ~v15 | (~v13 | ~\[3841] ),
  \[163]  = ~\[11199]  & (~v2 & (~\[11202]  & ~\[11208] )),
  \[22235]  = ~v4 | (~v7 | (~\[3536]  | ~\[3528] )),
  \[4154]  = ~\[10059]  & (~v0 & ~v2),
  \[11126]  = ~v0 | ~v2,
  \[8931]  = ~\[10058]  & (~v7 & ~v10),
  \[164]  = ~\[11212]  & (~\[11210]  & ~\[11218] ),
  \[6543]  = ~\[10058]  & (~v10 & ~v13),
  \[11125]  = ~v14 | (~\[10072]  | (~\[10076]  | ~\[7955] )),
  \[165]  = ~v6 & (~v5 & (~\[11192]  & ~\[11198] )),
  \[11855]  = ~\[21937]  | (~\[21935]  | (~\[21933]  | ~\[21931] )),
  \[895]  = ~\[314]  & (~\[313]  & (~\[315]  & ~\[12664] )),
  \[22241]  = ~v15 | (~v13 | (~\[3465]  | ~\[3475] )),
  \[13520]  = ~v11 | ~v8,
  \[4889]  = ~v6 & (~v5 & (~v8 & ~\[12654] )),
  \[12329]  = ~v10 | (~v9 | ~\[10068] ),
  \[13189]  = ~v15 | (~v13 | ~\[3823] ),
  \[8209]  = ~\[10059]  & (~v0 & (~\[10176]  & ~\[10996] )),
  \[9401]  = ~\[10060]  & (~v3 & (~\[10059]  & ~v0)),
  \[13183]  = ~v1 | (~\[10099]  | ~v3),
  \[7013]  = ~v6 & ~v5,
  \[7743]  = ~v10 & (~v9 & ~v12),
  \[22247]  = ~v15 | (~v13 | (~\[3411]  | ~\[3421] )),
  \[3697]  = ~v10 & (~v9 & ~v12),
  \[11138]  = ~v2 | (~\[10059]  | ~\[10176] ),
  \[11868]  = ~v5 | (~\[10134]  | ~v6),
  \[2839]  = ~\[10059]  & (~v0 & (~v2 & ~\[13686] )),
  \[22249]  = ~v7 | (~\[10236]  | (~\[3402]  | ~\[3394] )),
  \[10672]  = ~v8 | (~\[10064]  | ~v12),
  \[22243]  = ~v15 | (~v13 | (~\[3447]  | ~\[3457] )),
  \[3303]  = ~\[10068]  & (~v9 & ~v12),
  \[13192]  = ~v1 | (~\[10099]  | ~\[10060] ),
  \[4163]  = ~\[10058]  & (~v10 & ~v12),
  \[13529]  = ~v1 | (~\[10099]  | (~\[10060]  | ~\[3093] )),
  \[22245]  = ~v4 | (~\[10135]  | (~\[3438]  | ~\[3430] )),
  \[6553]  = ~\[10133]  & (~v5 & ~\[11822] ),
  \[11135]  = ~v14 | (~\[10072]  | (~\[10076]  | ~\[7933] )),
  \[2110]  = ~v4 & (~v3 & (~\[10060]  & ~v1)),
  \[21789]  = ~v13 | (~\[10073]  | (~\[7877]  | ~\[7887] )),
  \[13525]  = ~\[22275]  | (~\[22273]  | (~\[22271]  | ~\[22269] )),
  \[22251]  = ~v15 | (~v13 | (~\[3375]  | ~\[3385] )),
  \[13198]  = ~v15 | (~v13 | ~\[3805] ),
  \[5361]  = ~v6 & (~v5 & ~v8),
  \[8217]  = ~v10 & (~v9 & ~\[10088] ),
  \[4503]  = ~\[10068]  & (~\[10058]  & ~v12),
  \[13531]  = ~v11 | (~v8 | ~\[10088] ),
  \[7753]  = ~v6 & (~v5 & ~\[11224] ),
  \[7024]  = ~\[10073]  & (~v13 & ~v15),
  \[2848]  = ~\[10072]  & (~v14 & (~\[13680]  & ~v12)),
  \[9413]  = ~\[10060]  & (~v3 & (~\[10059]  & ~v0)),
  \[21791]  = ~v14 | (~\[10076]  | (~\[7859]  | ~\[7869] )),
  \[13538]  = ~v5 | (~\[10134]  | (~v6 | ~\[3142] )),
  \[10681]  = ~v8 | (~\[10064]  | ~v12),
  \[1654]  = ~v4 & (~v3 & (~\[10060]  & ~v1)),
  \[181]  = ~\[10073]  & (~v15 & (~\[11368]  & ~\[11366] )),
  \[11879]  = ~v5 | (~\[10134]  | ~v6),
  \[12341]  = ~v10 | (~\[10068]  | (~v9 | ~\[10058] )),
  \[11144]  = ~v14 | (~\[10076]  | ~\[7913] ),
  \[182]  = ~\[10073]  & (~v15 & (~\[11376]  & ~\[11374] )),
  \[6561]  = ~\[10058]  & (~v10 & ~v13),
  \[4173]  = ~\[10134]  & (~v6 & ~\[13012] ),
  \[183]  = ~\[11380]  & (~v2 & (~\[11383]  & ~\[11389] )),
  \[11146]  = ~v0 | (~v2 | ~\[10176] ),
  \[184]  = ~\[11393]  & (~\[11391]  & ~\[11399] ),
  \[8952]  = ~\[10073]  & (~v15 & ~\[10622] ),
  \[185]  = ~\[10073]  & (~v15 & (~\[11407]  & ~\[11405] )),
  \[186]  = ~\[10073]  & (~v15 & (~\[11415]  & ~\[11413] )),
  \[187]  = ~\[10073]  & (~v15 & (~\[11424]  & ~\[11422] )),
  \[11152]  = ~v14 | (~\[10076]  | ~\[7895] ),
  \[188]  = ~\[10073]  & (~v15 & (~\[11432]  & ~\[11430] )),
  \[10689]  = ~v8 | (~\[10064]  | ~v12),
  \[21793]  = ~v14 | (~\[10076]  | (~\[7841]  | ~\[7851] )),
  \[14007]  = ~v13 | (~\[10088]  | ~v15),
  \[8227]  = ~\[10099]  & (~\[10060]  & (~v3 & ~\[10987] )),
  \[4513]  = ~\[10133]  & (~v5 & ~\[12824] ),
  \[21795]  = ~v13 | (~\[10073]  | (~\[7823]  | ~\[7833] )),
  \[7761]  = ~v10 & (~v9 & ~v12),
  \[2856]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[14004]  = ~v10 | ~v9,
  \[2127]  = ~\[10134]  & (~v6 & ~v8),
  \[14003]  = ~v2 | (~\[10059]  | (~\[10176]  | ~\[2193] )),
  \[11158]  = ~v4 | ~v7,
  \[11888]  = ~v7 | ~\[10236] ,
  \[6905]  = ~v6 & ~v5,
  \[22269]  = ~v4 | (~v7 | (~\[3214]  | ~\[3206] )),
  \[3321]  = ~\[10068]  & (~v9 & ~v12),
  \[13547]  = ~v5 | (~\[10134]  | ~v6),
  \[4182]  = ~\[10058]  & (~v10 & (~v12 & ~\[13008] )),
  \[5711]  = ~\[10060]  & (~v1 & (~v3 & ~\[12247] )),
  \[6571]  = ~\[10059]  & (~v0 & (~v2 & ~\[11813] )),
  \[8960]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[193]  = ~\[10073]  & (~v15 & (~\[11488]  & ~\[11486] )),
  \[194]  = ~\[10073]  & (~v15 & (~\[11496]  & ~\[11494] )),
  \[13543]  = ~v8 | (~\[10133]  | (~v11 | ~\[3126] )),
  \[195]  = ~\[11473]  & (~v3 & (~\[11476]  & ~\[11482] )),
  \[13545]  = ~v1 | (~\[10099]  | ~v3),
  \[22271]  = ~v4 | (~v7 | (~\[3196]  | ~\[3188] )),
  \[9094]  = ~\[10060]  & (~v1 & ~v3),
  \[8235]  = ~v10 & (~v9 & ~\[10088] ),
  \[10699]  = ~v8 | (~\[10064]  | ~v12),
  \[14017]  = ~v13 | (~\[10088]  | ~v15),
  \[5719]  = ~\[10068]  & (~v9 & ~v12),
  \[4522]  = ~\[10076]  & (~\[10072]  & (~\[12843]  & ~v12)),
  \[12359]  = ~\[22039]  | (~\[22037]  | (~\[22041]  | ~\[954] )),
  \[6579]  = ~\[10058]  & (~v10 & ~v13),
  \[10693]  = ~\[21689]  | (~\[21687]  | (~\[21685]  | ~\[21683] )),
  \[5383]  = ~\[10133]  & (~v5 & ~v8),
  \[12353]  = ~v10 | (~\[10068]  | (~v9 | ~\[10058] )),
  \[14014]  = ~v10 | ~v9,
  \[14013]  = ~v0 | (~v2 | (~\[10176]  | ~\[2171] )),
  \[1671]  = ~\[10134]  & (~v6 & ~v8),
  \[11898]  = ~v4 | ~v7,
  \[4190]  = ~\[10059]  & (~v0 & ~v2),
  \[22273]  = ~v4 | (~v7 | (~\[3178]  | ~\[3170] )),
  \[13559]  = ~v1 | (~\[10099]  | ~v3),
  \[8970]  = ~\[10073]  & (~v15 & ~\[10614] ),
  \[22275]  = ~v4 | (~v7 | (~\[3160]  | ~\[3152] )),
  \[11166]  = ~v4 | ~v7,
  \[13553]  = ~v8 | (~\[10133]  | (~v11 | ~\[3104] )),
  \[11895]  = ~\[21945]  | (~\[21943]  | (~\[21941]  | ~\[21939] )),
  \[4530]  = ~\[10059]  & (~v0 & ~v2),
  \[3339]  = ~\[10068]  & (~v9 & ~v12),
  \[8245]  = ~\[10060]  & (~v1 & (~v3 & ~\[10979] )),
  \[4199]  = ~\[10058]  & (~v10 & ~v12),
  \[14028]  = ~v13 | (~\[10088]  | ~v15),
  \[6920]  = ~\[10073]  & (~v15 & (~\[11619]  & ~v13)),
  \[5729]  = ~\[10134]  & (~v6 & (~\[12234]  & ~v3)),
  \[12369]  = ~v12 | (~v14 | ~\[10076] ),
  \[2874]  = ~\[10060]  & (~v1 & ~v3),
  \[6589]  = ~\[10134]  & (~v6 & ~\[11804] ),
  \[8978]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[7781]  = ~v9 & (~v7 & ~v10),
  \[7052]  = ~\[10073]  & (~v13 & (~v15 & ~\[11571] )),
  \[11506]  = ~v5 | (~\[10134]  | ~v6),
  \[14024]  = ~v2 | (~\[10059]  | (~\[10176]  | ~\[2149] )),
  \[12366]  = ~v10 | ~v9,
  \[22287]  = ~v4 | (~\[10135]  | (~\[3044]  | ~\[3036] )),
  \[12365]  = ~v1 | (~\[10099]  | (~v3 | ~\[5471] )),
  \[10317]  = ~\[21589]  | (~\[21587]  | (~\[21591]  | ~\[1404] )),
  \[2149]  = ~\[10134]  & (~v6 & ~v8),
  \[22289]  = ~v7 | (~\[10236]  | (~\[3026]  | ~\[3018] )),
  \[14025]  = ~v10 | ~v9,
  \[10319]  = ~\[1441]  | (~\[1448]  | (~\[1434]  | ~\[1421] )),
  \[4539]  = ~\[10068]  & (~\[10058]  & ~v12),
  \[22283]  = ~v13 | (~\[10073]  | (~\[3071]  | ~\[3081] )),
  \[6928]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[13902]  = ~v13 | (~\[10088]  | ~v15),
  \[12709]  = ~v10 | (~\[10068]  | (~v9 | ~\[10058] )),
  \[22285]  = ~v4 | (~\[10135]  | (~\[3062]  | ~\[3054] )),
  \[11175]  = ~v4 | ~v7,
  \[1688]  = ~\[10072]  & (~v12 & (~v14 & ~\[14251] )),
  \[8253]  = ~v10 & (~v9 & ~v13),
  \[2880]  = ~\[10072]  & (~v12 & ~v14),
  \[11518]  = ~v11 | (~\[10063]  | ~v12),
  \[22291]  = ~v7 | (~\[10236]  | (~\[3008]  | ~\[3000] )),
  \[5737]  = ~\[10068]  & (~v9 & ~v12),
  \[13570]  = ~v11 | ~v8,
  \[6597]  = ~\[10058]  & (~v10 & ~v13),
  \[14038]  = ~v13 | (~\[10088]  | ~v15),
  \[12379]  = ~v12 | (~v14 | ~\[10076] ),
  \[13909]  = ~v5 | (~v6 | (~\[10133]  | ~\[2382] )),
  \[8988]  = ~\[10073]  & (~v15 & ~\[10605] ),
  \[6203]  = ~\[10068]  & (~v9 & ~v13),
  \[14034]  = ~v0 | (~v2 | (~\[10176]  | ~\[2127] )),
  \[7063]  = ~\[10059]  & (~v0 & (~v2 & ~\[11568] )),
  \[12376]  = ~v10 | ~v9,
  \[22297]  = ~v4 | (~\[10135]  | (~\[2954]  | ~\[2946] )),
  \[12375]  = ~v1 | (~\[10099]  | (~\[10060]  | ~\[5449] )),
  \[14035]  = ~v10 | ~v9,
  \[1693]  = ~\[10134]  & (~v6 & ~v8),
  \[11522]  = ~v0 | ~v2,
  \[4549]  = ~\[10134]  & (~v6 & ~\[12832] ),
  \[22293]  = ~\[10135]  | (~\[10236]  | (~\[2990]  | ~\[2982] )),
  \[6938]  = ~\[10073]  & (~v15 & (~\[11635]  & ~v13)),
  \[12719]  = ~v10 | (~v9 | ~\[10068] ),
  \[10323]  = ~\[10088]  | (~\[10135]  | (~v5 | ~\[10134] )),
  \[9457]  = ~\[10060]  & (~v3 & (~\[10059]  & ~v0)),
  \[13579]  = ~v11 | ~v8,
  \[11183]  = ~v4 | ~v7,
  \[10326]  = ~v5 | ~\[10134] ,
  \[22295]  = ~v13 | (~\[10073]  | (~\[2963]  | ~\[2973] )),
  \[1698]  = ~\[10060]  & (~v1 & ~v3),
  \[5015]  = ~v6 & (~v5 & ~v8),
  \[3357]  = ~\[10068]  & (~v9 & ~v12),
  \[8263]  = ~\[10059]  & (~v0 & (~v2 & ~\[10969] )),
  \[11190]  = ~\[21795]  | (~\[21793]  | (~\[21791]  | ~\[21789] )),
  \[1302]  = ~\[10728]  & (~\[10693]  & ~\[10795] ),
  \[7405]  = ~v9 & (~v7 & ~\[10068] ),
  \[5747]  = ~\[10060]  & (~v1 & (~v3 & ~\[12228] )),
  \[12387]  = ~v10 | ~v9,
  \[11192]  = ~v1 | (~\[10099]  | ~\[10060] ),
  \[10331]  = ~v5 | (~\[10134]  | ~v7),
  \[8996]  = ~\[10060]  & (~v1 & ~v3),
  \[14047]  = ~v5 | (~v6 | (~\[10133]  | ~\[2110] )),
  \[7072]  = ~\[10073]  & (~v15 & (~\[11561]  & ~v13)),
  \[6213]  = ~\[10134]  & (~v6 & ~\[11993] ),
  \[8602]  = ~\[10099]  & (~\[10060]  & ~v3),
  \[12386]  = ~v1 | (~\[10099]  | (~v3 | ~\[5427] )),
  \[11198]  = ~v13 | (~\[10073]  | ~\[7761] ),
  \[12390]  = ~v12 | (~v14 | ~\[10076] ),
  \[13915]  = ~v13 | (~\[10088]  | (~v15 | ~\[2369] )),
  \[567]  = ~\[477]  & (~\[476]  & (~\[475]  & ~\[474] )),
  \[6946]  = ~\[10059]  & (~v0 & ~v2),
  \[4558]  = ~\[10076]  & (~\[10072]  & (~\[12817]  & ~v12)),
  \[9464]  = ~\[10236]  & ~v4,
  \[13587]  = ~v11 | ~v8,
  \[11199]  = ~v1 | ~\[10099] ,
  \[902]  = ~\[308]  & (~\[307]  & (~\[306]  & ~\[305] )),
  \[13921]  = ~v3 | (~\[10134]  | (~v1 | ~\[10099] )),
  \[8271]  = ~v10 & (~v9 & ~\[10088] ),
  \[10335]  = ~v5 | (~\[10134]  | ~v7),
  \[5755]  = ~\[10068]  & (~v9 & ~v12),
  \[12725]  = ~v0 | (~v2 | ~\[10176] ),
  \[2171]  = ~v6 & (~v5 & ~v8),
  \[2509]  = ~\[10058]  & (~v7 & ~v10),
  \[12730]  = ~v10 | (~v9 | ~\[10068] ),
  \[12397]  = ~v10 | ~v9,
  \[10341]  = ~v5 | (~\[10134]  | ~v7),
  \[11539]  = ~\[21869]  | (~\[21867]  | (~\[21865]  | ~\[21863] )),
  \[14057]  = ~v5 | ~v6,
  \[909]  = ~\[304]  & (~\[303]  & (~\[302]  & ~\[301] )),
  \[12001]  = ~\[21967]  | (~\[21965]  | (~\[21963]  | ~\[21961] )),
  \[7080]  = ~\[10059]  & (~v0 & ~\[10176] ),
  \[13592]  = ~\[22289]  | (~\[22287]  | (~\[22285]  | ~\[22283] )),
  \[1315]  = ~\[104]  & (~\[103]  & (~\[105]  & ~\[10626] )),
  \[6221]  = ~\[10068]  & (~v9 & ~v13);
endmodule

