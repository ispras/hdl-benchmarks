module s38584_bench(
  blif_clk_net,
  blif_reset_net,
  g35,
  g36,
  g6744,
  g6745,
  g6746,
  g6747,
  g6748,
  g6749,
  g6750,
  g6751,
  g6752,
  g6753,
  g7243,
  g7245,
  g7257,
  g7260,
  g7540,
  g7916,
  g7946,
  g8132,
  g8178,
  g8215,
  g8235,
  g8277,
  g8279,
  g8283,
  g8291,
  g8342,
  g8344,
  g8353,
  g8358,
  g8398,
  g8403,
  g8416,
  g8475,
  g8719,
  g8783,
  g8784,
  g8785,
  g8786,
  g8787,
  g8788,
  g8789,
  g8839,
  g8870,
  g8915,
  g8916,
  g8917,
  g8918,
  g8919,
  g8920,
  g9019,
  g9048,
  g9251,
  g9497,
  g9553,
  g9555,
  g9615,
  g9617,
  g9680,
  g9682,
  g9741,
  g9743,
  g9817,
  g10122,
  g10306,
  g10500,
  g10527,
  g11349,
  g11388,
  g11418,
  g11447,
  g11678,
  g11770,
  g12184,
  g12238,
  g12300,
  g12350,
  g12368,
  g12422,
  g12470,
  g12832,
  g12919,
  g12923,
  g13039,
  g13049,
  g13068,
  g13085,
  g13099,
  g13259,
  g13272,
  g13865,
  g13881,
  g13895,
  g13906,
  g13926,
  g13966,
  g14096,
  g14125,
  g14147,
  g14167,
  g14189,
  g14201,
  g14217,
  g14421,
  g14451,
  g14518,
  g14597,
  g14635,
  g14662,
  g14673,
  g14694,
  g14705,
  g14738,
  g14749,
  g14779,
  g14828,
  g16603,
  g16624,
  g16627,
  g16656,
  g16659,
  g16686,
  g16693,
  g16718,
  g16722,
  g16744,
  g16748,
  g16775,
  g16874,
  g16924,
  g16955,
  g17291,
  g17316,
  g17320,
  g17400,
  g17404,
  g17423,
  g17519,
  g17577,
  g17580,
  g17604,
  g17607,
  g17639,
  g17646,
  g17649,
  g17674,
  g17678,
  g17685,
  g17688,
  g17711,
  g17715,
  g17722,
  g17739,
  g17743,
  g17760,
  g17764,
  g17778,
  g17787,
  g17813,
  g17819,
  g17845,
  g17871,
  g18092,
  g18094,
  g18095,
  g18096,
  g18097,
  g18098,
  g18099,
  g18100,
  g18101,
  g18881,
  g19334,
  g19357,
  g20049,
  g20557,
  g20652,
  g20654,
  g20763,
  g20899,
  g20901,
  g21176,
  g21245,
  g21270,
  g21292,
  g21698,
  g21727,
  g23002,
  g23190,
  g23612,
  g23652,
  g23683,
  g23759,
  g24151,
  g25114,
  g25167,
  g25219,
  g25259,
  g25582,
  g25583,
  g25584,
  g25585,
  g25586,
  g25587,
  g25588,
  g25589,
  g25590,
  g26801,
  g26875,
  g26876,
  g26877,
  g27831,
  g28030,
  g28041,
  g28042,
  g28753,
  g29210,
  g29211,
  g29212,
  g29213,
  g29214,
  g29215,
  g29216,
  g29217,
  g29218,
  g29219,
  g29220,
  g29221,
  g30327,
  g30329,
  g30330,
  g30331,
  g30332,
  g31521,
  g31656,
  g31665,
  g31793,
  g31860,
  g31861,
  g31862,
  g31863,
  g32185,
  g32429,
  g32454,
  g32975,
  g33079,
  g33435,
  g33533,
  g33636,
  g33659,
  g33874,
  g33894,
  g33935,
  g33945,
  g33946,
  g33947,
  g33948,
  g33949,
  g33950,
  g33959,
  g34201,
  g34221,
  g34232,
  g34233,
  g34234,
  g34235,
  g34236,
  g34237,
  g34238,
  g34239,
  g34240,
  g34383,
  g34425,
  g34435,
  g34436,
  g34437,
  g34597,
  g34788,
  g34839,
  g34913,
  g34915,
  g34917,
  g34919,
  g34921,
  g34923,
  g34925,
  g34927,
  g34956,
  g34972);
input blif_clk_net;
input blif_reset_net;
input g35;
input g36;
input g6744;
input g6745;
input g6746;
input g6747;
input g6748;
input g6749;
input g6750;
input g6751;
input g6752;
input g6753;
output g7243;
output g7245;
output g7257;
output g7260;
output g7540;
output g7916;
output g7946;
output g8132;
output g8178;
output g8215;
output g8235;
output g8277;
output g8279;
output g8283;
output g8291;
output g8342;
output g8344;
output g8353;
output g8358;
output g8398;
output g8403;
output g8416;
output g8475;
output g8719;
output g8783;
output g8784;
output g8785;
output g8786;
output g8787;
output g8788;
output g8789;
output g8839;
output g8870;
output g8915;
output g8916;
output g8917;
output g8918;
output g8919;
output g8920;
output g9019;
output g9048;
output g9251;
output g9497;
output g9553;
output g9555;
output g9615;
output g9617;
output g9680;
output g9682;
output g9741;
output g9743;
output g9817;
output g10122;
output g10306;
output g10500;
output g10527;
output g11349;
output g11388;
output g11418;
output g11447;
output g11678;
output g11770;
output g12184;
output g12238;
output g12300;
output g12350;
output g12368;
output g12422;
output g12470;
output g12832;
output g12919;
output g12923;
output g13039;
output g13049;
output g13068;
output g13085;
output g13099;
output g13259;
output g13272;
output g13865;
output g13881;
output g13895;
output g13906;
output g13926;
output g13966;
output g14096;
output g14125;
output g14147;
output g14167;
output g14189;
output g14201;
output g14217;
output g14421;
output g14451;
output g14518;
output g14597;
output g14635;
output g14662;
output g14673;
output g14694;
output g14705;
output g14738;
output g14749;
output g14779;
output g14828;
output g16603;
output g16624;
output g16627;
output g16656;
output g16659;
output g16686;
output g16693;
output g16718;
output g16722;
output g16744;
output g16748;
output g16775;
output g16874;
output g16924;
output g16955;
output g17291;
output g17316;
output g17320;
output g17400;
output g17404;
output g17423;
output g17519;
output g17577;
output g17580;
output g17604;
output g17607;
output g17639;
output g17646;
output g17649;
output g17674;
output g17678;
output g17685;
output g17688;
output g17711;
output g17715;
output g17722;
output g17739;
output g17743;
output g17760;
output g17764;
output g17778;
output g17787;
output g17813;
output g17819;
output g17845;
output g17871;
output g18092;
output g18094;
output g18095;
output g18096;
output g18097;
output g18098;
output g18099;
output g18100;
output g18101;
output g18881;
output g19334;
output g19357;
output g20049;
output g20557;
output g20652;
output g20654;
output g20763;
output g20899;
output g20901;
output g21176;
output g21245;
output g21270;
output g21292;
output g21698;
output g21727;
output g23002;
output g23190;
output g23612;
output g23652;
output g23683;
output g23759;
output g24151;
output g25114;
output g25167;
output g25219;
output g25259;
output g25582;
output g25583;
output g25584;
output g25585;
output g25586;
output g25587;
output g25588;
output g25589;
output g25590;
output g26801;
output g26875;
output g26876;
output g26877;
output g27831;
output g28030;
output g28041;
output g28042;
output g28753;
output g29210;
output g29211;
output g29212;
output g29213;
output g29214;
output g29215;
output g29216;
output g29217;
output g29218;
output g29219;
output g29220;
output g29221;
output g30327;
output g30329;
output g30330;
output g30331;
output g30332;
output g31521;
output g31656;
output g31665;
output g31793;
output g31860;
output g31861;
output g31862;
output g31863;
output g32185;
output g32429;
output g32454;
output g32975;
output g33079;
output g33435;
output g33533;
output g33636;
output g33659;
output g33874;
output g33894;
output g33935;
output g33945;
output g33946;
output g33947;
output g33948;
output g33949;
output g33950;
output g33959;
output g34201;
output g34221;
output g34232;
output g34233;
output g34234;
output g34235;
output g34236;
output g34237;
output g34238;
output g34239;
output g34240;
output g34383;
output g34425;
output g34435;
output g34436;
output g34437;
output g34597;
output g34788;
output g34839;
output g34913;
output g34915;
output g34917;
output g34919;
output g34921;
output g34923;
output g34925;
output g34927;
output g34956;
output g34972;
reg g72;
reg g73;
reg g84;
reg g90;
reg g91;
reg g92;
reg g99;
reg g100;
reg g110;
reg g112;
reg g113;
reg g114;
reg g115;
reg g116;
reg g120;
reg g124;
reg g125;
reg g126;
reg g127;
reg g134;
reg g135;
reg g44;
reg g45;
reg g46;
reg g47;
reg g48;
reg g49;
reg g50;
reg g51;
reg g52;
reg g53;
reg g54;
reg g55;
reg g56;
reg g57;
reg g58;
reg g63;
reg g71;
reg g85;
reg g93;
reg g101;
reg g111;
reg g43;
reg g64;
reg g65;
reg g70;
reg g4507;
reg g4459;
reg g4369;
reg g4473;
reg g4462;
reg g4581;
reg g4467;
reg g4474;
reg g4477;
reg g4480;
reg g4495;
reg g4498;
reg g4501;
reg g4504;
reg g4512;
reg g4521;
reg g4527;
reg g4515;
reg g4519;
reg g4520;
reg g4483;
reg g4486;
reg g4489;
reg g4492;
reg g4537;
reg g4423;
reg g4540;
reg g4543;
reg g4567;
reg g4546;
reg g4549;
reg g4552;
reg g4570;
reg g4571;
reg g4555;
reg g4558;
reg g4561;
reg g4564;
reg g4534;
reg g4420;
reg g4438;
reg g4449;
reg g4443;
reg g4446;
reg g4452;
reg g4434;
reg g4430;
reg g4427;
reg g4375;
reg g4414;
reg g4411;
reg g4408;
reg g4405;
reg g4401;
reg g4388;
reg g4382;
reg g4417;
reg g4392;
reg g4456;
reg g4455;
reg g1;
reg g4304;
reg g4308;
reg g2932;
reg g4639;
reg g4621;
reg g4628;
reg g4633;
reg g4643;
reg g4340;
reg g4349;
reg g4358;
reg g66;
reg g4531;
reg g4311;
reg g4322;
reg g4332;
reg g4584;
reg g4593;
reg g4601;
reg g4608;
reg g4616;
reg g4366;
reg g4372;
reg g4836;
reg g4864;
reg g4871;
reg g4878;
reg g4843;
reg g4849;
reg g4854;
reg g4859;
reg g4917;
reg g4922;
reg g4907;
reg g4912;
reg g4927;
reg g4931;
reg g4932;
reg g4572;
reg g4578;
reg g4999;
reg g5002;
reg g5005;
reg g5008;
reg g4983;
reg g4991;
reg g4966;
reg g4975;
reg g4899;
reg g4894;
reg g4888;
reg g4939;
reg g4933;
reg g4950;
reg g4944;
reg g4961;
reg g4955;
reg g4646;
reg g4674;
reg g4681;
reg g4688;
reg g4653;
reg g4659;
reg g4664;
reg g4669;
reg g4727;
reg g4732;
reg g4717;
reg g4722;
reg g4737;
reg g4741;
reg g4742;
reg g59;
reg g4575;
reg g4809;
reg g4812;
reg g4815;
reg g4818;
reg g4793;
reg g4801;
reg g4776;
reg g4785;
reg g4709;
reg g4704;
reg g4698;
reg g4749;
reg g4743;
reg g4760;
reg g4754;
reg g4771;
reg g4765;
reg g5313;
reg g5290;
reg g5320;
reg g5276;
reg g5283;
reg g5308;
reg g5327;
reg g5331;
reg g5335;
reg g5339;
reg g5343;
reg g5348;
reg g5352;
reg g5357;
reg g5297;
reg g5101;
reg g5109;
reg g5062;
reg g5105;
reg g5112;
reg g5022;
reg g5016;
reg g5029;
reg g5033;
reg g5037;
reg g5041;
reg g5046;
reg g5052;
reg g5057;
reg g5069;
reg g5073;
reg g5077;
reg g5080;
reg g5084;
reg g5092;
reg g5097;
reg g86;
reg g5164;
reg g5170;
reg g5176;
reg g5180;
reg g5188;
reg g5196;
reg g5224;
reg g5240;
reg g5256;
reg g5204;
reg g5200;
reg g5228;
reg g5244;
reg g5260;
reg g5212;
reg g5208;
reg g5232;
reg g5248;
reg g5264;
reg g5220;
reg g5216;
reg g5236;
reg g5252;
reg g5268;
reg g5272;
reg g128;
reg g5156;
reg g5120;
reg g5115;
reg g5124;
reg g5128;
reg g5134;
reg g5138;
reg g5142;
reg g5148;
reg g5152;
reg g5160;
reg g5659;
reg g5637;
reg g5666;
reg g5623;
reg g5630;
reg g5654;
reg g5673;
reg g5677;
reg g5681;
reg g5685;
reg g5689;
reg g5694;
reg g5698;
reg g5703;
reg g5644;
reg g5448;
reg g5456;
reg g5406;
reg g5452;
reg g5459;
reg g5366;
reg g5360;
reg g5373;
reg g5377;
reg g5381;
reg g5385;
reg g5390;
reg g5396;
reg g5401;
reg g5413;
reg g5417;
reg g5421;
reg g5424;
reg g5428;
reg g5436;
reg g5441;
reg g5445;
reg g5511;
reg g5517;
reg g5523;
reg g5527;
reg g5535;
reg g5543;
reg g5571;
reg g5587;
reg g5603;
reg g5551;
reg g5547;
reg g5575;
reg g5591;
reg g5607;
reg g5559;
reg g5555;
reg g5579;
reg g5595;
reg g5611;
reg g5567;
reg g5563;
reg g5583;
reg g5599;
reg g5615;
reg g5619;
reg g4821;
reg g5503;
reg g5467;
reg g5462;
reg g5471;
reg g5475;
reg g5481;
reg g5485;
reg g5489;
reg g5495;
reg g5499;
reg g5507;
reg g6005;
reg g5983;
reg g6012;
reg g5969;
reg g5976;
reg g6000;
reg g6019;
reg g6023;
reg g6027;
reg g6031;
reg g6035;
reg g6040;
reg g6044;
reg g6049;
reg g5990;
reg g5794;
reg g5802;
reg g5752;
reg g5798;
reg g5805;
reg g5712;
reg g5706;
reg g5719;
reg g5723;
reg g5727;
reg g5731;
reg g5736;
reg g5742;
reg g5747;
reg g5759;
reg g5763;
reg g5767;
reg g5770;
reg g5774;
reg g5782;
reg g5787;
reg g5791;
reg g5857;
reg g5863;
reg g5869;
reg g5873;
reg g5881;
reg g5889;
reg g5917;
reg g5933;
reg g5949;
reg g5897;
reg g5893;
reg g5921;
reg g5937;
reg g5953;
reg g5905;
reg g5901;
reg g5925;
reg g5941;
reg g5957;
reg g5913;
reg g5909;
reg g5929;
reg g5945;
reg g5961;
reg g5965;
reg g4831;
reg g5849;
reg g5813;
reg g5808;
reg g5817;
reg g5821;
reg g5827;
reg g5831;
reg g5835;
reg g5841;
reg g5845;
reg g5853;
reg g6351;
reg g6329;
reg g6358;
reg g6315;
reg g6322;
reg g6346;
reg g6365;
reg g6369;
reg g6373;
reg g6377;
reg g6381;
reg g6386;
reg g6390;
reg g6395;
reg g6336;
reg g6140;
reg g6148;
reg g6098;
reg g6144;
reg g6151;
reg g6058;
reg g6052;
reg g6065;
reg g6069;
reg g6073;
reg g6077;
reg g6082;
reg g6088;
reg g6093;
reg g6105;
reg g6109;
reg g6113;
reg g6116;
reg g6120;
reg g6128;
reg g6133;
reg g6137;
reg g6203;
reg g6209;
reg g6215;
reg g6219;
reg g6227;
reg g6235;
reg g6263;
reg g6279;
reg g6295;
reg g6243;
reg g6239;
reg g6267;
reg g6283;
reg g6299;
reg g6251;
reg g6247;
reg g6271;
reg g6287;
reg g6303;
reg g6259;
reg g6255;
reg g6275;
reg g6291;
reg g6307;
reg g6311;
reg g4826;
reg g6195;
reg g6159;
reg g6154;
reg g6163;
reg g6167;
reg g6173;
reg g6177;
reg g6181;
reg g6187;
reg g6191;
reg g6199;
reg g6697;
reg g6675;
reg g6704;
reg g6661;
reg g6668;
reg g6692;
reg g6711;
reg g6715;
reg g6719;
reg g6723;
reg g6727;
reg g6732;
reg g6736;
reg g6741;
reg g6682;
reg g6486;
reg g6494;
reg g6444;
reg g6490;
reg g6497;
reg g6404;
reg g6398;
reg g6411;
reg g6415;
reg g6419;
reg g6423;
reg g6428;
reg g6434;
reg g6439;
reg g6451;
reg g6455;
reg g6459;
reg g6462;
reg g6466;
reg g6474;
reg g6479;
reg g6483;
reg g6549;
reg g6555;
reg g6561;
reg g6565;
reg g6573;
reg g6581;
reg g6609;
reg g6625;
reg g6641;
reg g6589;
reg g6585;
reg g6613;
reg g6629;
reg g6645;
reg g6597;
reg g6593;
reg g6617;
reg g6633;
reg g6649;
reg g6605;
reg g6601;
reg g6621;
reg g6637;
reg g6653;
reg g6657;
reg g5011;
reg g6541;
reg g6505;
reg g6500;
reg g6509;
reg g6513;
reg g6519;
reg g6523;
reg g6527;
reg g6533;
reg g6537;
reg g6545;
reg g3303;
reg g3281;
reg g3310;
reg g3267;
reg g3274;
reg g3298;
reg g3317;
reg g3321;
reg g3325;
reg g3329;
reg g3338;
reg g3343;
reg g3347;
reg g3352;
reg g3288;
reg g3092;
reg g3100;
reg g3050;
reg g3096;
reg g3103;
reg g3010;
reg g3004;
reg g3017;
reg g3021;
reg g3025;
reg g3029;
reg g3034;
reg g3040;
reg g3045;
reg g3057;
reg g3061;
reg g3065;
reg g3068;
reg g3072;
reg g3080;
reg g3085;
reg g3089;
reg g3155;
reg g3161;
reg g3167;
reg g3171;
reg g3179;
reg g3187;
reg g3215;
reg g3231;
reg g3247;
reg g3195;
reg g3191;
reg g3219;
reg g3235;
reg g3251;
reg g3203;
reg g3199;
reg g3223;
reg g3239;
reg g3255;
reg g3211;
reg g3207;
reg g3227;
reg g3243;
reg g3259;
reg g3263;
reg g3333;
reg g3147;
reg g3111;
reg g3106;
reg g3115;
reg g3119;
reg g3125;
reg g3129;
reg g3133;
reg g3139;
reg g3143;
reg g3151;
reg g3654;
reg g3632;
reg g3661;
reg g3618;
reg g3625;
reg g3649;
reg g3668;
reg g3672;
reg g3676;
reg g3680;
reg g3689;
reg g3694;
reg g3698;
reg g3703;
reg g3639;
reg g3443;
reg g3451;
reg g3401;
reg g3447;
reg g3454;
reg g3361;
reg g3355;
reg g3368;
reg g3372;
reg g3376;
reg g3380;
reg g3385;
reg g3391;
reg g3396;
reg g3408;
reg g3412;
reg g3416;
reg g3419;
reg g3423;
reg g3431;
reg g3436;
reg g3440;
reg g3506;
reg g3512;
reg g3518;
reg g3522;
reg g3530;
reg g3538;
reg g3566;
reg g3582;
reg g3598;
reg g3546;
reg g3542;
reg g3570;
reg g3586;
reg g3602;
reg g3554;
reg g3550;
reg g3574;
reg g3590;
reg g3606;
reg g3562;
reg g3558;
reg g3578;
reg g3594;
reg g3610;
reg g3614;
reg g3684;
reg g3498;
reg g3462;
reg g3457;
reg g3466;
reg g3470;
reg g3476;
reg g3480;
reg g3484;
reg g3490;
reg g3494;
reg g3502;
reg g4005;
reg g3983;
reg g4012;
reg g3969;
reg g3976;
reg g4000;
reg g4019;
reg g4023;
reg g4027;
reg g4031;
reg g4040;
reg g4045;
reg g4049;
reg g4054;
reg g3990;
reg g3794;
reg g3802;
reg g3752;
reg g3798;
reg g3805;
reg g3712;
reg g3706;
reg g3719;
reg g3723;
reg g3727;
reg g3731;
reg g3736;
reg g3742;
reg g3747;
reg g3759;
reg g3763;
reg g3767;
reg g3770;
reg g3774;
reg g3782;
reg g3787;
reg g3791;
reg g3857;
reg g3863;
reg g3869;
reg g3873;
reg g3881;
reg g3889;
reg g3917;
reg g3933;
reg g3949;
reg g3897;
reg g3893;
reg g3921;
reg g3937;
reg g3953;
reg g3905;
reg g3901;
reg g3925;
reg g3941;
reg g3957;
reg g3913;
reg g3909;
reg g3929;
reg g3945;
reg g3961;
reg g3965;
reg g4035;
reg g3849;
reg g3813;
reg g3808;
reg g3817;
reg g3821;
reg g3827;
reg g3831;
reg g3835;
reg g3841;
reg g3845;
reg g3853;
reg g4165;
reg g4169;
reg g4125;
reg g4072;
reg g4064;
reg g4057;
reg g4141;
reg g4082;
reg g4076;
reg g4087;
reg g4093;
reg g4098;
reg g4108;
reg g4104;
reg g4145;
reg g4112;
reg g4116;
reg g4119;
reg g4122;
reg g4153;
reg g4164;
reg g4129;
reg g4132;
reg g4135;
reg g4138;
reg g4172;
reg g4176;
reg g4146;
reg g4157;
reg g4258;
reg g4264;
reg g4269;
reg g4273;
reg g4239;
reg g4294;
reg g4297;
reg g4300;
reg g4253;
reg g4249;
reg g4245;
reg g4277;
reg g4281;
reg g4284;
reg g4287;
reg g4291;
reg g2946;
reg g4191;
reg g4188;
reg g4194;
reg g4197;
reg g4200;
reg g4204;
reg g4207;
reg g4210;
reg g4180;
reg g4185;
reg g4213;
reg g4216;
reg g4219;
reg g4222;
reg g4226;
reg g4229;
reg g4232;
reg g4235;
reg g4242;
reg g305;
reg g311;
reg g336;
reg g324;
reg g316;
reg g319;
reg g329;
reg g333;
reg g344;
reg g347;
reg g351;
reg g355;
reg g74;
reg g106;
reg g341;
reg g637;
reg g640;
reg g559;
reg g562;
reg g568;
reg g572;
reg g586;
reg g577;
reg g582;
reg g590;
reg g595;
reg g599;
reg g604;
reg g608;
reg g613;
reg g617;
reg g622;
reg g626;
reg g632;
reg g859;
reg g869;
reg g875;
reg g878;
reg g881;
reg g884;
reg g887;
reg g872;
reg g225;
reg g255;
reg g232;
reg g262;
reg g239;
reg g269;
reg g246;
reg g446;
reg g890;
reg g862;
reg g896;
reg g901;
reg g391;
reg g365;
reg g358;
reg g370;
reg g376;
reg g385;
reg g203;
reg g854;
reg g847;
reg g703;
reg g837;
reg g843;
reg g812;
reg g817;
reg g832;
reg g822;
reg g827;
reg g723;
reg g645;
reg g681;
reg g699;
reg g650;
reg g655;
reg g718;
reg g661;
reg g728;
reg g79;
reg g691;
reg g686;
reg g667;
reg g671;
reg g676;
reg g714;
reg g499;
reg g504;
reg g513;
reg g518;
reg g528;
reg g482;
reg g490;
reg g417;
reg g411;
reg g424;
reg g475;
reg g441;
reg g437;
reg g433;
reg g429;
reg g401;
reg g392;
reg g405;
reg g182;
reg g174;
reg g168;
reg g460;
reg g452;
reg g457;
reg g471;
reg g464;
reg g468;
reg g479;
reg g102;
reg g496;
reg g732;
reg g753;
reg g799;
reg g802;
reg g736;
reg g739;
reg g744;
reg g749;
reg g758;
reg g763;
reg g767;
reg g772;
reg g776;
reg g781;
reg g785;
reg g790;
reg g794;
reg g807;
reg g554;
reg g538;
reg g546;
reg g542;
reg g534;
reg g550;
reg g136;
reg g199;
reg g278;
reg g283;
reg g287;
reg g291;
reg g294;
reg g298;
reg g142;
reg g146;
reg g164;
reg g150;
reg g153;
reg g157;
reg g160;
reg g301;
reg g222;
reg g194;
reg g191;
reg g209;
reg g215;
reg g218;
reg g1249;
reg g1266;
reg g1280;
reg g1252;
reg g1256;
reg g1259;
reg g1263;
reg g1270;
reg g1274;
reg g1277;
reg g1418;
reg g1422;
reg g1426;
reg g1430;
reg g1548;
reg g1564;
reg g1559;
reg g1554;
reg g1570;
reg g1585;
reg g1589;
reg g1576;
reg g1579;
reg g1339;
reg g1500;
reg g1582;
reg g1333;
reg g1399;
reg g1459;
reg g1322;
reg g1514;
reg g1526;
reg g1521;
reg g1306;
reg g1532;
reg g1536;
reg g1542;
reg g1413;
reg g1395;
reg g1404;
reg g1319;
reg g1312;
reg g1351;
reg g1345;
reg g1361;
reg g1367;
reg g1373;
reg g1379;
reg g1384;
reg g1389;
reg g1489;
reg g1495;
reg g1442;
reg g1437;
reg g1478;
reg g1454;
reg g1448;
reg g1467;
reg g1472;
reg g1484;
reg g1300;
reg g1291;
reg g1296;
reg g1283;
reg g1287;
reg g1311;
reg g929;
reg g904;
reg g921;
reg g936;
reg g907;
reg g911;
reg g914;
reg g918;
reg g925;
reg g930;
reg g933;
reg g1075;
reg g1079;
reg g1083;
reg g1087;
reg g1205;
reg g1221;
reg g1216;
reg g1211;
reg g1227;
reg g1242;
reg g1246;
reg g1233;
reg g1236;
reg g996;
reg g1157;
reg g1239;
reg g990;
reg g1056;
reg g1116;
reg g979;
reg g1171;
reg g1183;
reg g1178;
reg g962;
reg g1189;
reg g1193;
reg g1199;
reg g1070;
reg g1052;
reg g1061;
reg g976;
reg g969;
reg g1008;
reg g1002;
reg g1018;
reg g1024;
reg g1030;
reg g1036;
reg g1041;
reg g1046;
reg g1146;
reg g1152;
reg g1099;
reg g1094;
reg g1135;
reg g1111;
reg g1105;
reg g1124;
reg g1129;
reg g1141;
reg g956;
reg g947;
reg g952;
reg g939;
reg g943;
reg g967;
reg g968;
reg g1592;
reg g1644;
reg g1636;
reg g1668;
reg g1682;
reg g1687;
reg g1604;
reg g1600;
reg g1608;
reg g1620;
reg g1616;
reg g1612;
reg g1632;
reg g1624;
reg g1648;
reg g1664;
reg g1657;
reg g1677;
reg g1691;
reg g1696;
reg g1700;
reg g1706;
reg g1710;
reg g1714;
reg g1720;
reg g1724;
reg g1728;
reg g1779;
reg g1772;
reg g1802;
reg g1816;
reg g1821;
reg g1740;
reg g1736;
reg g1744;
reg g1756;
reg g1752;
reg g1748;
reg g1768;
reg g1760;
reg g1783;
reg g1798;
reg g1792;
reg g1811;
reg g1825;
reg g1830;
reg g1834;
reg g1840;
reg g1844;
reg g1848;
reg g1854;
reg g1858;
reg g1862;
reg g1913;
reg g1906;
reg g1936;
reg g1950;
reg g1955;
reg g1874;
reg g1870;
reg g1878;
reg g1890;
reg g1886;
reg g1882;
reg g1902;
reg g1894;
reg g1917;
reg g1932;
reg g1926;
reg g1945;
reg g1959;
reg g1964;
reg g1968;
reg g1974;
reg g1978;
reg g1982;
reg g1988;
reg g1992;
reg g1996;
reg g2047;
reg g2040;
reg g2070;
reg g2084;
reg g2089;
reg g2008;
reg g2004;
reg g2012;
reg g2024;
reg g2020;
reg g2016;
reg g2036;
reg g2028;
reg g2051;
reg g2066;
reg g2060;
reg g2079;
reg g2093;
reg g2098;
reg g2102;
reg g2108;
reg g2112;
reg g2116;
reg g2122;
reg g2126;
reg g2130;
reg g2138;
reg g2145;
reg g2151;
reg g2152;
reg g2153;
reg g2204;
reg g2197;
reg g2227;
reg g2241;
reg g2246;
reg g2165;
reg g2161;
reg g2169;
reg g2181;
reg g2177;
reg g2173;
reg g2193;
reg g2185;
reg g2208;
reg g2223;
reg g2217;
reg g2236;
reg g2250;
reg g2255;
reg g2259;
reg g2265;
reg g2269;
reg g2273;
reg g2279;
reg g2283;
reg g2287;
reg g2338;
reg g2331;
reg g2361;
reg g2375;
reg g2380;
reg g2299;
reg g2295;
reg g2303;
reg g2315;
reg g2311;
reg g2307;
reg g2327;
reg g2319;
reg g2342;
reg g2357;
reg g2351;
reg g2370;
reg g2384;
reg g2389;
reg g2393;
reg g2399;
reg g2403;
reg g2407;
reg g2413;
reg g2417;
reg g2421;
reg g2472;
reg g2465;
reg g2495;
reg g2509;
reg g2514;
reg g2433;
reg g2429;
reg g2437;
reg g2449;
reg g2445;
reg g2441;
reg g2461;
reg g2453;
reg g2476;
reg g2491;
reg g2485;
reg g2504;
reg g2518;
reg g2523;
reg g2527;
reg g2533;
reg g2537;
reg g2541;
reg g2547;
reg g2551;
reg g2555;
reg g2606;
reg g2599;
reg g2629;
reg g2643;
reg g2648;
reg g2567;
reg g2563;
reg g2571;
reg g2583;
reg g2579;
reg g2575;
reg g2595;
reg g2587;
reg g2610;
reg g2625;
reg g2619;
reg g2638;
reg g2652;
reg g2657;
reg g2661;
reg g2667;
reg g2671;
reg g2675;
reg g2681;
reg g2685;
reg g2689;
reg g2697;
reg g2704;
reg g2710;
reg g2711;
reg g2837;
reg g2841;
reg g2712;
reg g2715;
reg g2719;
reg g2724;
reg g2729;
reg g2735;
reg g2741;
reg g2748;
reg g2756;
reg g2759;
reg g2763;
reg g2767;
reg g2779;
reg g2791;
reg g2795;
reg g2787;
reg g2783;
reg g2775;
reg g2771;
reg g2831;
reg g121;
reg g2799;
reg g2811;
reg g2823;
reg g2827;
reg g2819;
reg g2815;
reg g2807;
reg g2803;
reg g2834;
reg g117;
reg g2999;
reg g2994;
reg g2988;
reg g2868;
reg g2873;
reg g2890;
reg g2844;
reg g2852;
reg g2860;
reg g2894;
reg g37;
reg g94;
reg g2848;
reg g2856;
reg g2864;
reg g2898;
reg g2882;
reg g2878;
reg g2886;
reg g2980;
reg g2984;
reg g2907;
reg g2912;
reg g2922;
reg g2936;
reg g2950;
reg g2960;
reg g2970;
reg g2902;
reg g2917;
reg g2927;
reg g2941;
reg g2955;
reg g2965;
reg g2975;
reg g3003;
reg g5;
reg g6;
reg g7;
reg g8;
reg g9;
reg g16;
reg g19;
reg g28;
reg g31;
reg g34;
reg g12;
reg g22;
reg g25;
wire II28897;
wire g20592;
wire g18281;
wire II26071;
wire g24124;
wire g31542;
wire g31799;
wire II13463;
wire g30503;
wire g22225;
wire g24850;
wire g32057;
wire g13491;
wire g28911;
wire g14745;
wire II15363;
wire II15147;
wire g30086;
wire g24362;
wire g21718;
wire g8508;
wire II14712;
wire g30484;
wire g32453;
wire g33602;
wire g29928;
wire g20549;
wire g34089;
wire g9977;
wire g27059;
wire g20649;
wire g21930;
wire g9700;
wire g17417;
wire g32491;
wire II32535;
wire g30384;
wire g24396;
wire g32767;
wire g21693;
wire g19524;
wire g31471;
wire g34351;
wire g34132;
wire II18509;
wire g16508;
wire g24600;
wire g22712;
wire g13626;
wire g22527;
wire g28160;
wire II12994;
wire g27547;
wire g24903;
wire g21458;
wire g16530;
wire g26632;
wire g7252;
wire g22719;
wire II20203;
wire g32879;
wire g34370;
wire g32226;
wire II21802;
wire g8938;
wire g32852;
wire g23609;
wire g18644;
wire g24985;
wire g25907;
wire II13240;
wire g34643;
wire g15647;
wire g14394;
wire g28840;
wire II20542;
wire g33470;
wire II12041;
wire g7521;
wire g29308;
wire g33097;
wire II18307;
wire g32274;
wire g17296;
wire g29740;
wire g12855;
wire g32910;
wire g33592;
wire g31239;
wire g15348;
wire g21780;
wire g31883;
wire g12193;
wire g25200;
wire II16526;
wire g22036;
wire g19765;
wire g32438;
wire II21047;
wire g17694;
wire g22220;
wire g29295;
wire g28186;
wire gbuf3;
wire g23276;
wire g28773;
wire g28619;
wire g8106;
wire g10230;
wire g29301;
wire g19449;
wire g32943;
wire g11232;
wire g6847;
wire g33669;
wire g31772;
wire g10882;
wire g27481;
wire g19638;
wire g29873;
wire g22625;
wire g25317;
wire g20573;
wire g15809;
wire g23984;
wire g15053;
wire II32225;
wire II12070;
wire g18334;
wire g6827;
wire g29846;
wire g34706;
wire g14764;
wire g8130;
wire II13509;
wire g20240;
wire g23183;
wire g32772;
wire g24196;
wire g24906;
wire g29336;
wire g25544;
wire g30376;
wire g8123;
wire g25630;
wire g12868;
wire g34249;
wire g30608;
wire g32803;
wire g16066;
wire g11907;
wire g8032;
wire g18465;
wire g23297;
wire g25564;
wire g17652;
wire g11584;
wire g23313;
wire g13413;
wire g32663;
wire g32510;
wire II26880;
wire g19432;
wire g32343;
wire II23321;
wire g34544;
wire g21876;
wire g33694;
wire II17919;
wire g18250;
wire g30219;
wire g31762;
wire g30423;
wire g32131;
wire II11682;
wire g21657;
wire g25639;
wire g28052;
wire g34193;
wire g19903;
wire g14489;
wire g29575;
wire g34833;
wire g12921;
wire g33675;
wire g17821;
wire g32914;
wire g31278;
wire g27523;
wire g32312;
wire g34334;
wire g11900;
wire g29151;
wire g17136;
wire g10217;
wire g23051;
wire g34112;
wire g32557;
wire II29218;
wire g25232;
wire g10117;
wire g8804;
wire g33088;
wire g20273;
wire g22142;
wire g29246;
wire g28361;
wire g34272;
wire g23994;
wire II14332;
wire g27479;
wire g32830;
wire g15148;
wire g28059;
wire g33729;
wire g7297;
wire II11753;
wire II17207;
wire g11811;
wire g32211;
wire II16460;
wire g18994;
wire g23337;
wire g32987;
wire g16701;
wire g30469;
wire g24796;
wire g7132;
wire g33233;
wire g24189;
wire g30333;
wire g32933;
wire g26277;
wire g32895;
wire g18389;
wire g27138;
wire g30302;
wire g9360;
wire g34406;
wire g17790;
wire g30150;
wire g10400;
wire g26301;
wire g24946;
wire g22638;
wire g27184;
wire g18349;
wire g8678;
wire g9011;
wire g18391;
wire g12804;
wire g20496;
wire g8137;
wire g10405;
wire g22855;
wire II14893;
wire g28151;
wire g12179;
wire II22845;
wire g24565;
wire g29362;
wire g7537;
wire g28344;
wire g32283;
wire g16661;
wire g10099;
wire g9582;
wire g22086;
wire g24149;
wire g30491;
wire g13656;
wire g15720;
wire g26606;
wire g33888;
wire g24069;
wire g31301;
wire g33109;
wire g17637;
wire II29720;
wire g9914;
wire g33090;
wire g13047;
wire g15867;
wire g34880;
wire g24427;
wire g32356;
wire g16179;
wire g25740;
wire g12126;
wire g11169;
wire g12041;
wire g33128;
wire g13138;
wire g25781;
wire g29948;
wire g12122;
wire II26004;
wire g20614;
wire g16795;
wire II22900;
wire g6900;
wire g22117;
wire g18803;
wire g30228;
wire g18531;
wire g33881;
wire g11344;
wire g30245;
wire g24300;
wire g23917;
wire g17954;
wire g27575;
wire g26357;
wire g16767;
wire g34728;
wire g17740;
wire g27693;
wire g30998;
wire g26667;
wire g34252;
wire g25106;
wire g29485;
wire g16766;
wire g34152;
wire II26440;
wire g9825;
wire g13477;
wire g27401;
wire g27635;
wire g14376;
wire g8373;
wire g18263;
wire g12217;
wire g34242;
wire g32609;
wire g11045;
wire g16800;
wire g24003;
wire II13054;
wire g18954;
wire g25032;
wire g24088;
wire g25946;
wire g30265;
wire g25131;
wire g15911;
wire g14443;
wire II15702;
wire II12314;
wire g29996;
wire g18286;
wire g34566;
wire g33625;
wire g31803;
wire g33974;
wire g21248;
wire g10373;
wire g24045;
wire g11924;
wire g18917;
wire g26161;
wire g30550;
wire II29447;
wire II23971;
wire g23215;
wire g23563;
wire g9200;
wire g14785;
wire g29973;
wire g10762;
wire g30568;
wire g24359;
wire g16752;
wire g29257;
wire g12233;
wire II18143;
wire g18268;
wire g30344;
wire II18285;
wire g34001;
wire II20167;
wire II16679;
wire g27133;
wire g30010;
wire g26145;
wire g17809;
wire II28594;
wire g17608;
wire g15966;
wire g33287;
wire g31797;
wire g33778;
wire g16886;
wire g18427;
wire g30526;
wire g32441;
wire II26960;
wire g26614;
wire II13374;
wire II31256;
wire g27508;
wire g30296;
wire g18884;
wire g24034;
wire II11992;
wire g30403;
wire g26206;
wire g18791;
wire g13098;
wire g20133;
wire g30288;
wire g10616;
wire g32085;
wire g25788;
wire g12340;
wire g10543;
wire g25977;
wire g7495;
wire g29175;
wire g27317;
wire g29943;
wire g25627;
wire g18656;
wire g12505;
wire g24257;
wire g34311;
wire g28211;
wire g20526;
wire g23489;
wire g10165;
wire II25606;
wire g17793;
wire g26872;
wire g16708;
wire g32742;
wire g33131;
wire g26826;
wire g14309;
wire II13889;
wire g7049;
wire g19861;
wire g34462;
wire II27492;
wire g33056;
wire g25261;
wire g25994;
wire g18811;
wire g27298;
wire g30159;
wire g8844;
wire g33322;
wire g34593;
wire g34980;
wire g17157;
wire g13022;
wire g33823;
wire g18373;
wire g29288;
wire g18653;
wire II19759;
wire g33102;
wire gbuf130;
wire g16733;
wire II29973;
wire g29641;
wire g17248;
wire g6977;
wire II15088;
wire g25165;
wire g27590;
wire g31839;
wire II18373;
wire g21939;
wire g16484;
wire II15052;
wire II15782;
wire g26902;
wire g32498;
wire g29478;
wire II14427;
wire II12278;
wire g24237;
wire g25596;
wire g11324;
wire g10140;
wire II15213;
wire g14616;
wire g6804;
wire gbuf35;
wire g34769;
wire g31658;
wire g7908;
wire g28220;
wire g23781;
wire g32483;
wire II23587;
wire g33492;
wire g19782;
wire g33868;
wire g24846;
wire g21913;
wire II32840;
wire g27310;
wire g28612;
wire II19487;
wire g24673;
wire II27927;
wire g23863;
wire g23476;
wire g18188;
wire g28918;
wire g23289;
wire g19686;
wire II32815;
wire g15562;
wire g13251;
wire g28761;
wire II16855;
wire II31056;
wire II22894;
wire g10043;
wire g28524;
wire g10653;
wire g28903;
wire g23941;
wire II17140;
wire g28977;
wire g18402;
wire g28108;
wire II15334;
wire g27252;
wire g19720;
wire g8026;
wire g25833;
wire g23234;
wire g33796;
wire g34314;
wire g17597;
wire II14455;
wire g25924;
wire g9305;
wire g20385;
wire g24725;
wire g17491;
wire g17578;
wire g34124;
wire g27772;
wire g23433;
wire g22980;
wire II27429;
wire II16613;
wire g25517;
wire II18120;
wire g29181;
wire g17177;
wire g33809;
wire g24973;
wire g32575;
wire g29093;
wire g31926;
wire g8131;
wire g18439;
wire g15118;
wire g17844;
wire g16646;
wire g8426;
wire g19710;
wire g15747;
wire g29267;
wire g25533;
wire g19371;
wire g33619;
wire g30200;
wire g24411;
wire g34672;
wire g34288;
wire g23352;
wire g13909;
wire g13498;
wire g26610;
wire g18777;
wire g31850;
wire II13723;
wire II33152;
wire g21609;
wire g21755;
wire g22045;
wire g29591;
wire g13540;
wire g20004;
wire g26572;
wire g32600;
wire II32074;
wire g23410;
wire g8434;
wire g18719;
wire g18939;
wire g34295;
wire g23252;
wire g21993;
wire g23436;
wire g14993;
wire g14516;
wire g25067;
wire gbuf121;
wire II16629;
wire g34497;
wire g15843;
wire g18726;
wire g21306;
wire g27692;
wire g25057;
wire g24014;
wire g28693;
wire g20265;
wire II17750;
wire g33553;
wire II31500;
wire g34793;
wire g14094;
wire II23118;
wire g20516;
wire g19397;
wire g21746;
wire g16670;
wire II32096;
wire g32182;
wire g14173;
wire g29005;
wire gbuf23;
wire g32336;
wire g22869;
wire g25715;
wire g28255;
wire g30521;
wire g33511;
wire g22147;
wire g12847;
wire g7869;
wire g10102;
wire g22179;
wire II23378;
wire g16524;
wire gbuf76;
wire g19421;
wire II30537;
wire g34738;
wire g10175;
wire II12141;
wire g18541;
wire g15121;
wire g31374;
wire g18203;
wire g30026;
wire g25667;
wire g30123;
wire g34069;
wire g30593;
wire g32013;
wire g31527;
wire g8531;
wire g27653;
wire g26154;
wire g22862;
wire g32651;
wire g27675;
wire g19490;
wire g32054;
wire g16688;
wire g15810;
wire g21751;
wire g31248;
wire g14192;
wire g7095;
wire g26124;
wire g16839;
wire g34922;
wire g11884;
wire g17687;
wire II15340;
wire g27086;
wire g25967;
wire g14014;
wire g13972;
wire g34850;
wire II22419;
wire g6995;
wire g29638;
wire g30382;
wire g27570;
wire II31307;
wire g10918;
wire g11989;
wire g29911;
wire g13432;
wire g34971;
wire II18634;
wire g9040;
wire g22660;
wire g29515;
wire g10204;
wire g21268;
wire g11834;
wire g21970;
wire g17416;
wire g33385;
wire g32523;
wire g8620;
wire g18735;
wire g21812;
wire g34444;
wire II22965;
wire g32750;
wire g16225;
wire g33267;
wire II13391;
wire g21823;
wire g11237;
wire g30061;
wire g24009;
wire g11248;
wire g21977;
wire g33984;
wire g30205;
wire g12978;
wire g7926;
wire g28518;
wire g15723;
wire II12773;
wire g31207;
wire g8069;
wire g27907;
wire II20130;
wire g13853;
wire g14782;
wire g15799;
wire g18228;
wire g23459;
wire g24160;
wire g25758;
wire g34514;
wire g14521;
wire g29661;
wire g20199;
wire g33051;
wire g15073;
wire g8187;
wire g33357;
wire g16930;
wire II12770;
wire g28242;
wire g20053;
wire g28938;
wire g27119;
wire g21846;
wire g33500;
wire II26195;
wire g14573;
wire g30670;
wire g14933;
wire g27435;
wire g14680;
wire g10902;
wire g20639;
wire g11033;
wire g20209;
wire g26753;
wire g33138;
wire g33066;
wire g16479;
wire g13075;
wire g32252;
wire g25706;
wire g33424;
wire II12841;
wire g23009;
wire g12796;
wire g23854;
wire g10365;
wire g28102;
wire g31623;
wire g25526;
wire g31505;
wire g32208;
wire g30042;
wire II33182;
wire g18714;
wire g34851;
wire II22316;
wire II11865;
wire II31701;
wire g16193;
wire g13518;
wire g12884;
wire g32348;
wire g17122;
wire g6986;
wire II15105;
wire g25451;
wire g28466;
wire g16681;
wire II27738;
wire II32947;
wire g33002;
wire g26835;
wire II12583;
wire g22154;
wire g34789;
wire g18303;
wire g26957;
wire II33034;
wire g9214;
wire g26330;
wire g33827;
wire g10607;
wire II29961;
wire g33992;
wire g34986;
wire g30229;
wire g24998;
wire g24078;
wire g29761;
wire g32925;
wire g28997;
wire g26882;
wire g15124;
wire g32711;
wire g9630;
wire g12337;
wire g25110;
wire g26821;
wire g28381;
wire g21673;
wire g21335;
wire g18183;
wire g24172;
wire II31142;
wire g25022;
wire g30598;
wire II15474;
wire II19707;
wire g21275;
wire II31002;
wire g12645;
wire g6941;
wire g20720;
wire g19613;
wire g24714;
wire II30741;
wire g14882;
wire g29510;
wire g32932;
wire g33715;
wire g13280;
wire g32260;
wire g32581;
wire g9766;
wire II15533;
wire g24337;
wire g15091;
wire g21298;
wire g16579;
wire g25019;
wire g32174;
wire g27236;
wire g25922;
wire g10586;
wire II27232;
wire g25239;
wire g19597;
wire g34196;
wire II26531;
wire g12197;
wire g10475;
wire g23052;
wire g20157;
wire g31868;
wire g31832;
wire g25655;
wire g9257;
wire g33375;
wire g24180;
wire g16635;
wire g26390;
wire g33341;
wire g19932;
wire II21930;
wire g23452;
wire g24726;
wire g26920;
wire g31121;
wire g32116;
wire gbuf55;
wire g32622;
wire g24098;
wire g18607;
wire g32229;
wire g13805;
wire g27697;
wire II21849;
wire g33501;
wire g31014;
wire g34947;
wire g22834;
wire g12819;
wire g13621;
wire g26487;
wire g25600;
wire g10935;
wire g22923;
wire g9442;
wire g33877;
wire g33121;
wire g27315;
wire g17529;
wire g29226;
wire g10019;
wire g14002;
wire g24536;
wire g30937;
wire g24022;
wire g22973;
wire g8341;
wire g27032;
wire g21354;
wire g17188;
wire g10515;
wire g10427;
wire g23746;
wire g10649;
wire g11669;
wire g24154;
wire II33155;
wire g21330;
wire g26686;
wire g25642;
wire g12947;
wire II22711;
wire II21776;
wire g7201;
wire g29192;
wire II12344;
wire g24588;
wire g29508;
wire g19206;
wire g20663;
wire II15167;
wire g31128;
wire g26948;
wire g26022;
wire g28316;
wire g10396;
wire g17431;
wire II24474;
wire II31337;
wire g12024;
wire g33240;
wire g30371;
wire g29888;
wire g34457;
wire g23512;
wire g33899;
wire g13896;
wire g28249;
wire g11316;
wire II24705;
wire g8005;
wire II14647;
wire g15873;
wire g24572;
wire g32537;
wire g22685;
wire g26323;
wire g26083;
wire g27369;
wire g29494;
wire g29018;
wire II12189;
wire g16986;
wire g17755;
wire g19736;
wire g13297;
wire g8354;
wire g34768;
wire g24083;
wire II31477;
wire g27279;
wire g29639;
wire II12735;
wire g27251;
wire g13469;
wire g32793;
wire g34488;
wire g18741;
wire g33966;
wire g15935;
wire g31931;
wire g14744;
wire g18177;
wire g31295;
wire II26687;
wire g25151;
wire g26927;
wire g28631;
wire g29049;
wire g13939;
wire g33231;
wire g8690;
wire II31267;
wire g28141;
wire g19542;
wire g30242;
wire II31724;
wire g21859;
wire g28421;
wire g31230;
wire g17682;
wire g25770;
wire g24037;
wire II31187;
wire II22380;
wire g9672;
wire g31320;
wire g21356;
wire g27544;
wire g28439;
wire g23245;
wire gbuf124;
wire g13969;
wire g16672;
wire g22858;
wire g13738;
wire g8238;
wire g25448;
wire g29556;
wire g34481;
wire g24267;
wire g14740;
wire II17114;
wire II21922;
wire g32637;
wire g19369;
wire g18409;
wire g22092;
wire g34011;
wire g27408;
wire g19351;
wire II25907;
wire g13638;
wire II29269;
wire gbuf92;
wire g30239;
wire g33140;
wire II27543;
wire g18710;
wire g32982;
wire g20779;
wire g28078;
wire g10675;
wire g31751;
wire g28359;
wire g19874;
wire II33173;
wire II12463;
wire g16533;
wire II11737;
wire g32744;
wire g29628;
wire g19535;
wire g23964;
wire II18865;
wire g9100;
wire g20733;
wire II13078;
wire g18160;
wire g12078;
wire g29791;
wire g7161;
wire g19699;
wire II12545;
wire II33041;
wire II22571;
wire g13134;
wire II14896;
wire g17647;
wire g22885;
wire g27582;
wire g33806;
wire g9496;
wire g21205;
wire g18773;
wire g22588;
wire g31814;
wire g24243;
wire g30019;
wire g7002;
wire g18515;
wire II24051;
wire g28552;
wire g31975;
wire g14861;
wire g29283;
wire g9369;
wire g25837;
wire g11707;
wire g12108;
wire II20165;
wire II17324;
wire g11762;
wire g33115;
wire g23812;
wire g28069;
wire g11207;
wire g18898;
wire II28540;
wire g27271;
wire g19560;
wire g14234;
wire g22120;
wire II30971;
wire g11336;
wire g19476;
wire g18008;
wire g23499;
wire g34811;
wire g31254;
wire g34762;
wire g33788;
wire g32370;
wire g29908;
wire g32795;
wire g21819;
wire g24897;
wire II21074;
wire g24310;
wire g30030;
wire g17568;
wire gbuf43;
wire g28598;
wire g19518;
wire g21946;
wire g8526;
wire g18506;
wire g14817;
wire g34173;
wire g25983;
wire g13065;
wire g20436;
wire g20175;
wire g19277;
wire II12415;
wire g24199;
wire g34307;
wire g34693;
wire g16096;
wire g32008;
wire g24581;
wire g31993;
wire g34381;
wire II28434;
wire g8301;
wire g25699;
wire g27228;
wire g10415;
wire g32219;
wire II17436;
wire g32049;
wire g25010;
wire g7174;
wire g10420;
wire g26958;
wire g11216;
wire g25086;
wire g7423;
wire g29749;
wire II14924;
wire g12904;
wire g29270;
wire g10036;
wire g21180;
wire g16658;
wire g27973;
wire g31671;
wire g22929;
wire g13033;
wire g28656;
wire g22645;
wire g34628;
wire g13835;
wire g33164;
wire g33842;
wire g28513;
wire II15647;
wire g12540;
wire g32837;
wire g28281;
wire g34697;
wire g10147;
wire g34399;
wire g22875;
wire g10378;
wire II11743;
wire II15130;
wire II27777;
wire g18788;
wire II16555;
wire g11537;
wire g32425;
wire II13511;
wire g30392;
wire g14082;
wire II26367;
wire g13008;
wire g24378;
wire g29736;
wire g31125;
wire g22754;
wire g32108;
wire g18649;
wire II21234;
wire g34363;
wire g22848;
wire II22801;
wire II13335;
wire g9274;
wire g24386;
wire g18193;
wire g28678;
wire g18790;
wire g16601;
wire g20920;
wire g27820;
wire g28349;
wire g12932;
wire g12111;
wire g20185;
wire g34758;
wire g33011;
wire g30058;
wire g24208;
wire g15711;
wire g34993;
wire g26815;
wire g28600;
wire g28581;
wire II12437;
wire g10027;
wire g23443;
wire g29965;
wire g21433;
wire II33218;
wire g26869;
wire II23372;
wire g15757;
wire g34808;
wire g29143;
wire g23301;
wire g30361;
wire g25289;
wire g14924;
wire g9963;
wire g33275;
wire g22650;
wire g8944;
wire g24782;
wire II32516;
wire g24841;
wire g22908;
wire g26951;
wire g25316;
wire g29872;
wire II11620;
wire g14895;
wire II12987;
wire g24223;
wire g17486;
wire g20508;
wire g20644;
wire II18740;
wire g20232;
wire g18259;
wire g34962;
wire g27958;
wire g27414;
wire g18991;
wire g32924;
wire II11635;
wire g26609;
wire g16198;
wire g21012;
wire g26976;
wire g11956;
wire g34687;
wire g34714;
wire g14794;
wire g19408;
wire g13460;
wire II21486;
wire II20819;
wire g7528;
wire g24999;
wire g25147;
wire g25123;
wire g23182;
wire g32396;
wire g24475;
wire g13486;
wire g26019;
wire g12708;
wire g17663;
wire g29347;
wire g25124;
wire g7985;
wire g25215;
wire g12186;
wire g33599;
wire g27540;
wire g24778;
wire g27288;
wire g33575;
wire g20234;
wire g29563;
wire g22841;
wire g17785;
wire g34526;
wire g25388;
wire g30235;
wire g17531;
wire g8171;
wire g29685;
wire g33861;
wire g23129;
wire g25688;
wire g34417;
wire g21362;
wire g31767;
wire g11631;
wire g17148;
wire g15718;
wire g9311;
wire g34635;
wire g14386;
wire g24431;
wire g28923;
wire g22192;
wire II31016;
wire g24053;
wire g24406;
wire II32222;
wire g26232;
wire g20780;
wire g10319;
wire g8647;
wire g31818;
wire g27455;
wire II12112;
wire g27207;
wire g9536;
wire g7549;
wire g9818;
wire g33988;
wire g34105;
wire g31186;
wire g11200;
wire g25555;
wire g21903;
wire g28661;
wire II32752;
wire II17405;
wire g7442;
wire g21405;
wire g14222;
wire g16024;
wire II21199;
wire g28192;
wire g33828;
wire g23952;
wire g17769;
wire g23408;
wire g32125;
wire II16181;
wire g17810;
wire g13026;
wire g21998;
wire g25664;
wire g10754;
wire g9839;
wire g28073;
wire g11736;
wire II22111;
wire g33830;
wire g29316;
wire g24930;
wire g7634;
wire II32881;
wire g27661;
wire g29866;
wire g24913;
wire g15114;
wire g30478;
wire g24367;
wire g19795;
wire g21850;
wire g25681;
wire g28816;
wire g30073;
wire g18356;
wire g17606;
wire g30326;
wire g32466;
wire g32777;
wire II20562;
wire g18368;
wire g26165;
wire II11896;
wire g28237;
wire g14182;
wire g24763;
wire g31515;
wire g23351;
wire g10741;
wire g32759;
wire g7178;
wire g28477;
wire g17586;
wire g24730;
wire g17643;
wire g34805;
wire g34262;
wire g27303;
wire g16022;
wire g9832;
wire g32762;
wire g33463;
wire g21965;
wire g34039;
wire g33766;
wire g11029;
wire g31268;
wire g18613;
wire II15705;
wire g17717;
wire g10154;
wire II29182;
wire g32032;
wire g32546;
wire II24579;
wire g26120;
wire g32671;
wire g30105;
wire g9903;
wire g21709;
wire g27266;
wire g21468;
wire g34022;
wire II26100;
wire II30980;
wire g24921;
wire II31282;
wire II12758;
wire g25227;
wire g23170;
wire g8086;
wire g27937;
wire g24522;
wire g18398;
wire g27281;
wire g22077;
wire g32309;
wire g8011;
wire g27683;
wire g28110;
wire g28680;
wire g31770;
wire g30460;
wire g16660;
wire g14950;
wire II27576;
wire g26158;
wire g9174;
wire g26855;
wire g21870;
wire g33482;
wire g11796;
wire g27105;
wire g18909;
wire g20853;
wire g26127;
wire g21665;
wire g12112;
wire g26860;
wire g24342;
wire g7244;
wire g34663;
wire g9186;
wire g11190;
wire g13303;
wire g18745;
wire g11998;
wire g18493;
wire g11933;
wire g11470;
wire g20715;
wire g25194;
wire g29118;
wire g27345;
wire II20650;
wire g9223;
wire g14018;
wire g12785;
wire g34259;
wire g10737;
wire g29771;
wire g18187;
wire g25603;
wire g19437;
wire g33610;
wire g27980;
wire g21387;
wire g25738;
wire g29565;
wire g21717;
wire g24187;
wire g33900;
wire g21894;
wire g32489;
wire g30563;
wire g32814;
wire II12205;
wire g13887;
wire g24119;
wire g8720;
wire g25062;
wire g34599;
wire g27535;
wire g24182;
wire g32842;
wire g28687;
wire g30525;
wire g34916;
wire g31491;
wire g17737;
wire II12046;
wire g21222;
wire g14205;
wire g8400;
wire g11194;
wire II15915;
wire g25072;
wire g21411;
wire g32401;
wire g33677;
wire g32302;
wire II18555;
wire II17111;
wire g30119;
wire g18458;
wire g34281;
wire g28498;
wire g13346;
wire g14752;
wire g12852;
wire g29776;
wire g28537;
wire g20768;
wire g10106;
wire II14480;
wire g31210;
wire g10857;
wire g28259;
wire g33907;
wire g28607;
wire g29734;
wire g11411;
wire g24804;
wire g34008;
wire g12051;
wire g20433;
wire g16875;
wire g17150;
wire g29756;
wire g20919;
wire II26581;
wire II22864;
wire g34518;
wire g32780;
wire g13273;
wire g29666;
wire g8967;
wire g7512;
wire g27024;
wire g8631;
wire g29601;
wire g24147;
wire II23986;
wire g14335;
wire g24444;
wire g20539;
wire g17128;
wire g14776;
wire g28212;
wire g25832;
wire g21983;
wire g11971;
wire g29164;
wire g10501;
wire g22143;
wire g18596;
wire g24807;
wire g32633;
wire g34331;
wire g17571;
wire g20084;
wire g25819;
wire g18827;
wire g30253;
wire II29582;
wire g26783;
wire g24233;
wire g8795;
wire g18897;
wire II31878;
wire g14317;
wire g33403;
wire g31847;
wire g23610;
wire g20586;
wire g14011;
wire g13976;
wire g7841;
wire g34826;
wire g31001;
wire g23011;
wire g19912;
wire g16583;
wire g18570;
wire g18415;
wire II13851;
wire g11855;
wire g6870;
wire g15578;
wire g11979;
wire g29353;
wire g27504;
wire g9920;
wire g10897;
wire g18558;
wire g23524;
wire g10061;
wire g7285;
wire g16612;
wire g34581;
wire II17276;
wire gbuf84;
wire II32782;
wire g11048;
wire g26814;
wire g28569;
wire g28982;
wire g33026;
wire g33426;
wire g14104;
wire g23507;
wire g19592;
wire g15701;
wire g23012;
wire g30512;
wire g24276;
wire g33970;
wire g28199;
wire g22110;
wire II12608;
wire g14378;
wire g32700;
wire g25158;
wire g34410;
wire g16275;
wire g22546;
wire g25098;
wire II13718;
wire g13290;
wire g20379;
wire g27595;
wire g30004;
wire g10356;
wire g21836;
wire g33705;
wire g14503;
wire II31296;
wire g25775;
wire g31482;
wire g18578;
wire g25753;
wire g9450;
wire g15065;
wire II18667;
wire g11366;
wire II29139;
wire g30051;
wire g27246;
wire g11030;
wire g18797;
wire g15880;
wire g23389;
wire g8997;
wire g34212;
wire g10970;
wire II23671;
wire g18136;
wire II20937;
wire g20210;
wire g24620;
wire II18248;
wire II14258;
wire g27039;
wire g34050;
wire g26055;
wire II33197;
wire II31022;
wire g23770;
wire II17491;
wire g34075;
wire g7661;
wire g22591;
wire II18762;
wire II17475;
wire g14563;
wire g29807;
wire g11543;
wire II15765;
wire g30915;
wire II12402;
wire g9194;
wire g32579;
wire g12983;
wire g29234;
wire g32688;
wire g31871;
wire g10896;
wire II18114;
wire II21483;
wire g16804;
wire g33064;
wire g10386;
wire g31489;
wire g32709;
wire g14029;
wire g12346;
wire g26097;
wire II32757;
wire g25510;
wire g21343;
wire g21056;
wire g28935;
wire g16309;
wire g22176;
wire g32293;
wire g18906;
wire g20625;
wire g15874;
wire II17741;
wire g17511;
wire g30337;
wire g29130;
wire g22065;
wire g24305;
wire g31281;
wire g32178;
wire g10000;
wire g10960;
wire g28099;
wire II22830;
wire g11383;
wire g28230;
wire g14732;
wire g18290;
wire g14674;
wire g13947;
wire g31942;
wire g30604;
wire g19617;
wire g10776;
wire II18588;
wire g24112;
wire g7598;
wire g23570;
wire g16846;
wire g33007;
wire g11171;
wire g11403;
wire g30448;
wire g7591;
wire g33818;
wire g16176;
wire g23656;
wire g16472;
wire g12752;
wire g21288;
wire g33528;
wire g16076;
wire g30279;
wire g34168;
wire g16323;
wire g14600;
wire g25183;
wire g14538;
wire g7809;
wire g19489;
wire g18748;
wire g14031;
wire g19674;
wire II33067;
wire g25956;
wire g12998;
wire g22010;
wire g21805;
wire g34328;
wire g15506;
wire g30008;
wire II33050;
wire II12848;
wire g24812;
wire g25036;
wire g16261;
wire g10626;
wire g34782;
wire g24179;
wire g24669;
wire g34550;
wire g22123;
wire g14364;
wire g14708;
wire g32267;
wire g19384;
wire g24165;
wire g31935;
wire g25007;
wire g8765;
wire g16619;
wire g27687;
wire g21705;
wire II17416;
wire g13324;
wire g26264;
wire II31176;
wire g18975;
wire g27256;
wire g19695;
wire g32591;
wire g27558;
wire II32827;
wire g8542;
wire g26078;
wire g9753;
wire g18761;
wire g34719;
wire g32618;
wire g22635;
wire II18879;
wire g9690;
wire g34600;
wire g20495;
wire g20551;
wire g30249;
wire g29045;
wire g6988;
wire g30262;
wire g20619;
wire g18523;
wire g34618;
wire g33684;
wire g34392;
wire g26848;
wire g33248;
wire g12419;
wire g12255;
wire g10808;
wire g25671;
wire g10079;
wire II11879;
wire g30544;
wire g31147;
wire g11916;
wire g32668;
wire g34056;
wire II22871;
wire g29496;
wire g30166;
wire g14415;
wire g22131;
wire g13564;
wire g23196;
wire g25135;
wire g24356;
wire g32514;
wire g30269;
wire g33505;
wire g28720;
wire g9269;
wire g21881;
wire II26584;
wire g24451;
wire g8666;
wire gbuf50;
wire II22729;
wire g12970;
wire II12654;
wire g26929;
wire g21656;
wire II14800;
wire g33436;
wire g26854;
wire g32198;
wire g34996;
wire g7939;
wire g20602;
wire g32920;
wire II22989;
wire g20673;
wire g26932;
wire g10136;
wire gbuf118;
wire g25000;
wire g18320;
wire g13737;
wire g22105;
wire g12925;
wire g26213;
wire g33318;
wire II22824;
wire II13403;
wire g22002;
wire g25366;
wire g21768;
wire II14789;
wire g8102;
wire g33334;
wire g20034;
wire g12306;
wire II23354;
wire g31167;
wire g34476;
wire g26919;
wire g29282;
wire g30733;
wire g27214;
wire II12345;
wire g25581;
wire g15033;
wire II31066;
wire g28896;
wire g21889;
wire g33392;
wire g16736;
wire g16513;
wire g14665;
wire g8364;
wire g12915;
wire g15786;
wire g19964;
wire g28716;
wire g27516;
wire g19070;
wire g31243;
wire g25249;
wire g27363;
wire g32543;
wire g18243;
wire g9821;
wire g7418;
wire g9883;
wire g24951;
wire g12491;
wire g34107;
wire II31171;
wire g25349;
wire g28695;
wire g28545;
wire g25856;
wire g13574;
wire g34572;
wire g24681;
wire g10123;
wire g20011;
wire g26514;
wire g16725;
wire g18141;
wire g27099;
wire g13989;
wire g24218;
wire g28954;
wire II18117;
wire g32644;
wire g16694;
wire g13661;
wire II19238;
wire g27115;
wire g24091;
wire g20322;
wire g25374;
wire g16810;
wire g14542;
wire g16208;
wire g24920;
wire g10039;
wire g31310;
wire g19338;
wire g27090;
wire g7601;
wire gbuf74;
wire II13390;
wire g28500;
wire g9714;
wire II30962;
wire g18406;
wire II21294;
wire g30358;
wire g26100;
wire g12463;
wire g15847;
wire g20556;
wire g23347;
wire g28267;
wire g26944;
wire g34140;
wire g33259;
wire g20522;
wire II17606;
wire g24219;
wire II29228;
wire g31654;
wire g24654;
wire g34554;
wire II32391;
wire g30223;
wire g34965;
wire g33438;
wire g28131;
wire g32726;
wire g13287;
wire g16518;
wire II17679;
wire g18239;
wire g13851;
wire g30087;
wire g18983;
wire g34347;
wire g24984;
wire g25814;
wire g12476;
wire II21792;
wire g8097;
wire g20998;
wire g23022;
wire g18218;
wire g14767;
wire g7779;
wire g28068;
wire II14563;
wire g16926;
wire g19682;
wire g19778;
wire g18661;
wire g12016;
wire II14290;
wire g18234;
wire g30140;
wire g11559;
wire g19769;
wire g11213;
wire g16771;
wire g26866;
wire g34467;
wire g23197;
wire g17582;
wire g16812;
wire g28298;
wire g14614;
wire g28508;
wire g7802;
wire g30074;
wire g11842;
wire g19487;
wire g28301;
wire g18731;
wire g21453;
wire II15194;
wire g24093;
wire g13797;
wire g17085;
wire g28597;
wire g18316;
wire II24064;
wire g21986;
wire g26970;
wire g30029;
wire g22309;
wire g16893;
wire g19345;
wire g24678;
wire II22561;
wire g8241;
wire g8575;
wire g24546;
wire g27007;
wire g17616;
wire g8478;
wire g19555;
wire II15987;
wire gbuf119;
wire g25550;
wire g15373;
wire g18115;
wire g15852;
wire g23383;
wire g24139;
wire g25275;
wire II15650;
wire g32658;
wire g8443;
wire g18152;
wire g25282;
wire g9559;
wire g12662;
wire g17058;
wire g8595;
wire g26308;
wire g30174;
wire g20169;
wire g18171;
wire g30480;
wire g27389;
wire II14663;
wire g11702;
wire g26256;
wire g25820;
wire g21281;
wire g30232;
wire g32887;
wire II15243;
wire g15785;
wire g34679;
wire g20911;
wire g27269;
wire g23684;
wire g29291;
wire g29528;
wire g18418;
wire g30342;
wire gbuf33;
wire g14055;
wire g13061;
wire g20136;
wire g32222;
wire g21175;
wire g32446;
wire g34644;
wire g19661;
wire g15084;
wire g12099;
wire g34879;
wire g27881;
wire g18270;
wire II13149;
wire II17494;
wire g16642;
wire g33541;
wire II21036;
wire g27018;
wire g11721;
wire g34149;
wire g23883;
wire g25209;
wire g6809;
wire g24642;
wire II32089;
wire g15830;
wire g24777;
wire g20777;
wire gbuf17;
wire g23761;
wire g12833;
wire g23429;
wire g10725;
wire g32232;
wire g13118;
wire g30168;
wire g33305;
wire g30364;
wire g25692;
wire g29538;
wire g8803;
wire g34897;
wire g29072;
wire II14967;
wire g22407;
wire g27046;
wire g29924;
wire g25608;
wire g10583;
wire g23875;
wire g16282;
wire g29597;
wire II32482;
wire g26800;
wire g18496;
wire g25432;
wire g19602;
wire g29522;
wire g34755;
wire g25599;
wire g19470;
wire g8249;
wire g30576;
wire g11890;
wire g20610;
wire II12083;
wire g34340;
wire g29206;
wire g8712;
wire g34143;
wire g17301;
wire g24315;
wire g27015;
wire g27154;
wire g12440;
wire g18385;
wire g32528;
wire g23992;
wire g8477;
wire g16652;
wire g20658;
wire II21934;
wire g8046;
wire g12412;
wire g24698;
wire g34503;
wire g12146;
wire g28640;
wire g29581;
wire g20567;
wire II14326;
wire g10183;
wire g11370;
wire g29266;
wire g27360;
wire g15158;
wire g22987;
wire g13014;
wire g23602;
wire g14654;
wire g17710;
wire g19678;
wire g12729;
wire g12101;
wire g16868;
wire g26943;
wire g7395;
wire g25950;
wire II33079;
wire g22008;
wire g20063;
wire g11692;
wire g30930;
wire g22715;
wire g31893;
wire g10715;
wire g31749;
wire g25143;
wire g23715;
wire g12245;
wire g21731;
wire g31828;
wire g17590;
wire g13763;
wire g18279;
wire g25439;
wire g13377;
wire II31848;
wire g34218;
wire g33581;
wire II27528;
wire g18708;
wire g7750;
wire g17758;
wire g23768;
wire g16289;
wire g34030;
wire g13876;
wire g23920;
wire g8165;
wire g18327;
wire g13525;
wire g14876;
wire g13980;
wire g22033;
wire g28555;
wire g18580;
wire g32189;
wire g28336;
wire g17642;
wire g10072;
wire g11995;
wire g25990;
wire g10498;
wire g28705;
wire g6789;
wire g26683;
wire g31132;
wire g29502;
wire g33350;
wire II27495;
wire g14810;
wire g12632;
wire g24463;
wire g23264;
wire g10619;
wire II18360;
wire II24685;
wire g31475;
wire g32682;
wire g12292;
wire g25768;
wire g11965;
wire II14169;
wire g22022;
wire g12223;
wire g17365;
wire g32962;
wire g26364;
wire g11714;
wire g28746;
wire g15938;
wire g22165;
wire II31332;
wire g32376;
wire g33916;
wire g34650;
wire g18224;
wire g18524;
wire g33363;
wire g25157;
wire g20128;
wire g15480;
wire g23422;
wire g28080;
wire g28701;
wire g24959;
wire g28273;
wire g27323;
wire g26961;
wire g32956;
wire g32535;
wire g22070;
wire g33071;
wire g16749;
wire g19571;
wire g24106;
wire g23956;
wire g25978;
wire g21775;
wire g20100;
wire g29604;
wire II20870;
wire II31261;
wire II18709;
wire g25745;
wire g14713;
wire g7785;
wire g28081;
wire g18755;
wire g27235;
wire g18158;
wire g31950;
wire g18120;
wire g18475;
wire g34449;
wire II17925;
wire g32690;
wire g22472;
wire g9155;
wire g22939;
wire g7685;
wire g12054;
wire g12952;
wire g18876;
wire g23377;
wire g28036;
wire g21826;
wire g32158;
wire g25140;
wire g25092;
wire g23417;
wire II31868;
wire g14714;
wire g15851;
wire gbuf65;
wire g14202;
wire g28305;
wire g27571;
wire g11409;
wire g18552;
wire g33922;
wire g8350;
wire g20785;
wire g8659;
wire g20389;
wire g24176;
wire II23163;
wire II22718;
wire g21605;
wire g10939;
wire g7470;
wire g30204;
wire g13473;
wire g18213;
wire II20781;
wire g6888;
wire g18480;
wire II12541;
wire g14425;
wire II31853;
wire g27615;
wire g23698;
wire g30120;
wire g24328;
wire g11928;
wire g12459;
wire g34875;
wire g23112;
wire g28203;
wire g29008;
wire g27467;
wire g13665;
wire g20904;
wire g29784;
wire g31272;
wire g34657;
wire g30109;
wire g19146;
wire g27593;
wire g25274;
wire g15568;
wire g13495;
wire g12524;
wire g20638;
wire gbuf26;
wire g29660;
wire g21339;
wire g34157;
wire g19730;
wire g16956;
wire II18579;
wire g14253;
wire g23214;
wire g13139;
wire g10519;
wire g32564;
wire g31864;
wire g18950;
wire g34466;
wire g29313;
wire II12483;
wire II31252;
wire g29952;
wire g31509;
wire g28734;
wire g18469;
wire g34015;
wire g15567;
wire g24623;
wire g13175;
wire g15133;
wire g25485;
wire g19749;
wire g16183;
wire II24363;
wire g25423;
wire g29571;
wire g27295;
wire g15742;
wire g15727;
wire g30982;
wire g14185;
wire g18282;
wire g28571;
wire g27392;
wire g14291;
wire g23272;
wire g13011;
wire g27028;
wire II14991;
wire g33419;
wire g27439;
wire g18880;
wire II25243;
wire g18652;
wire II13454;
wire II32651;
wire g30407;
wire g23485;
wire g29550;
wire g30283;
wire g10003;
wire g30187;
wire g24926;
wire g34830;
wire g14120;
wire g26693;
wire g32861;
wire II12096;
wire g19654;
wire g8859;
wire g22994;
wire g17153;
wire g24062;
wire g24286;
wire g31219;
wire g33944;
wire g12937;
wire g11385;
wire g27314;
wire g28970;
wire g31794;
wire g33458;
wire g14433;
wire g23105;
wire g29148;
wire g24609;
wire g25265;
wire g15048;
wire g8737;
wire g15077;
wire g9300;
wire g24253;
wire II12172;
wire g33389;
wire II25351;
wire g23970;
wire g18648;
wire g25577;
wire g31250;
wire g31817;
wire g26840;
wire g19375;
wire g32846;
wire II22793;
wire g10274;
wire g28065;
wire g25730;
wire g27927;
wire g24144;
wire g24173;
wire g24365;
wire g24842;
wire g32785;
wire g22896;
wire g33841;
wire g18206;
wire g10657;
wire g30442;
wire g34323;
wire g6973;
wire g30132;
wire II32204;
wire g26209;
wire g34453;
wire g13554;
wire g32525;
wire II11809;
wire g24559;
wire g34299;
wire g17221;
wire g18435;
wire g8583;
wire g7184;
wire g24041;
wire g28098;
wire g24388;
wire g24605;
wire g12289;
wire g24497;
wire g28137;
wire g25216;
wire g19529;
wire II17302;
wire g26731;
wire g32807;
wire g29253;
wire II21058;
wire g18264;
wire g31907;
wire g12252;
wire g29305;
wire II16117;
wire g18361;
wire g22041;
wire g19451;
wire g14965;
wire g28171;
wire g11320;
wire g23871;
wire g16488;
wire g33410;
wire g24552;
wire g17593;
wire g29082;
wire g14130;
wire II17008;
wire g33326;
wire II13452;
wire g32284;
wire g9698;
wire II21013;
wire g29260;
wire g20269;
wire g33304;
wire g27527;
wire g25721;
wire g14038;
wire g23788;
wire g33096;
wire g15672;
wire g23284;
wire II31052;
wire II32675;
wire II26664;
wire g9407;
wire II32982;
wire g26576;
wire II28062;
wire II12056;
wire g26260;
wire g20732;
wire g28990;
wire g10799;
wire g23413;
wire II32812;
wire g20195;
wire g25611;
wire II30399;
wire II13110;
wire g14781;
wire g34114;
wire g23978;
wire g18679;
wire g25949;
wire g18441;
wire g29992;
wire g20766;
wire g25676;
wire g26178;
wire g23238;
wire II13597;
wire g24747;
wire g22851;
wire II15623;
wire g20172;
wire II18370;
wire g12975;
wire g28224;
wire g32476;
wire g23945;
wire g28907;
wire g30193;
wire g29709;
wire II16676;
wire g23567;
wire g12369;
wire g12861;
wire g12428;
wire g28652;
wire g26832;
wire g10980;
wire g32290;
wire g19793;
wire g24478;
wire g20088;
wire II29245;
wire g16763;
wire g10169;
wire g23135;
wire g31876;
wire II12850;
wire g33967;
wire g28966;
wire g8451;
wire g18744;
wire g20857;
wire g13190;
wire g34065;
wire g16209;
wire g22200;
wire II30760;
wire g6904;
wire g30322;
wire g16720;
wire g34137;
wire g30022;
wire g9284;
wire g21797;
wire g15631;
wire g19658;
wire g30488;
wire g12589;
wire g26702;
wire II20864;
wire II16417;
wire g27779;
wire g25537;
wire g30238;
wire g30055;
wire II26710;
wire II14761;
wire II12793;
wire g26712;
wire II14531;
wire g15017;
wire g31775;
wire g10658;
wire g23989;
wire gbuf150;
wire II14970;
wire II13990;
wire g19753;
wire g20542;
wire g22300;
wire g32947;
wire g10397;
wire g17734;
wire g31153;
wire g7239;
wire g34533;
wire g10219;
wire II16969;
wire g30428;
wire g18674;
wire g33836;
wire g22983;
wire II14619;
wire g8514;
wire g32245;
wire g34530;
wire g24561;
wire g28778;
wire g24392;
wire g27454;
wire II25190;
wire II18310;
wire g19681;
wire g33596;
wire g13832;
wire g23654;
wire II13037;
wire II23099;
wire g32332;
wire g33835;
wire g27427;
wire g25082;
wire II17885;
wire g29900;
wire g25128;
wire g12843;
wire g25727;
wire g33106;
wire g14549;
wire g17677;
wire II18417;
wire g23473;
wire g10096;
wire g32315;
wire g10676;
wire g9321;
wire g32604;
wire g29624;
wire g20650;
wire gbuf114;
wire g27705;
wire g26679;
wire g33878;
wire g27562;
wire g8284;
wire g25591;
wire g18394;
wire g32103;
wire g22360;
wire g32464;
wire g9973;
wire g21784;
wire g26517;
wire g32278;
wire g28480;
wire g15164;
wire g32070;
wire g6816;
wire g32977;
wire g28615;
wire g22310;
wire II17639;
wire g18519;
wire g10087;
wire g32856;
wire g28164;
wire g32024;
wire g22998;
wire g18323;
wire g34810;
wire g25909;
wire g32970;
wire g33811;
wire g13093;
wire II15800;
wire g24993;
wire g14927;
wire g34291;
wire g7118;
wire g26345;
wire II29285;
wire II22640;
wire g30154;
wire II31076;
wire g32855;
wire g14892;
wire g14142;
wire g27181;
wire g7411;
wire g25712;
wire g24705;
wire g31824;
wire g30209;
wire g25942;
wire g29117;
wire g24525;
wire II22488;
wire g17724;
wire g9613;
wire II20957;
wire g6832;
wire g16704;
wire g23018;
wire II20569;
wire g32166;
wire g19552;
wire g32495;
wire g19718;
wire g28406;
wire II27449;
wire g28055;
wire g7519;
wire g27567;
wire g18352;
wire g26306;
wire g25228;
wire g9397;
wire II14733;
wire g17465;
wire g25119;
wire g25635;
wire II17733;
wire g32418;
wire g24533;
wire g33871;
wire II31287;
wire g24192;
wire g14588;
wire g19605;
wire g27485;
wire g24891;
wire g29249;
wire g9681;
wire II33189;
wire g10401;
wire g17464;
wire g20576;
wire g18377;
wire g28117;
wire g10540;
wire g15144;
wire g7846;
wire g30334;
wire g26819;
wire g14254;
wire g17133;
wire g11028;
wire II14833;
wire g17670;
wire g28870;
wire g18683;
wire g6846;
wire g24281;
wire g24074;
wire g23394;
wire g23292;
wire g28367;
wire g9828;
wire II31111;
wire g32677;
wire g10080;
wire g33237;
wire g34785;
wire II14611;
wire II15929;
wire g10564;
wire g27737;
wire g27150;
wire g28877;
wire g33417;
wire g25231;
wire g34374;
wire II14818;
wire g29327;
wire g11496;
wire g19761;
wire II28336;
wire g29242;
wire g13942;
wire g21181;
wire g9911;
wire II15824;
wire g32121;
wire g34151;
wire g34144;
wire g7581;
wire II32648;
wire g19952;
wire g15057;
wire g23553;
wire g29332;
wire g19907;
wire II20205;
wire g30427;
wire g7443;
wire g34933;
wire g30096;
wire g29577;
wire II33146;
wire g27083;
wire II31873;
wire g28294;
wire g32940;
wire g33977;
wire g16841;
wire g18254;
wire g31309;
wire g18699;
wire II32855;
wire g10078;
wire g21793;
wire g28348;
wire g33903;
wire g12321;
wire g22517;
wire g26765;
wire g23999;
wire g23776;
wire g11107;
wire g18453;
wire g20247;
wire g8267;
wire g31305;
wire g8297;
wire g7631;
wire g25616;
wire g18337;
wire II13065;
wire g21863;
wire g21653;
wire g19748;
wire g12083;
wire g27733;
wire g19559;
wire g31840;
wire g21452;
wire g15863;
wire g11741;
wire g32352;
wire g13334;
wire g9586;
wire g9015;
wire g23265;
wire g21720;
wire g30537;
wire g18997;
wire g33327;
wire II13749;
wire g30479;
wire g8697;
wire g8150;
wire g29370;
wire g25382;
wire g7886;
wire g17708;
wire g29687;
wire g18346;
wire g32437;
wire II17876;
wire g26079;
wire g23534;
wire g7293;
wire g14879;
wire g13913;
wire II33030;
wire g23382;
wire g28181;
wire II31528;
wire II26479;
wire g33567;
wire g29552;
wire g13018;
wire g26087;
wire g25031;
wire g14262;
wire g34064;
wire g30341;
wire II32665;
wire g19637;
wire g10392;
wire g30156;
wire II30983;
wire g11443;
wire II18476;
wire g18889;
wire g13625;
wire g20094;
wire g26423;
wire g6826;
wire g24158;
wire II32479;
wire g19731;
wire II18627;
wire g20599;
wire g28467;
wire g17779;
wire g7690;
wire g7697;
wire g34386;
wire g26743;
wire g9856;
wire II12991;
wire g30495;
wire g29014;
wire g34623;
wire g11203;
wire g23335;
wire g8635;
wire g28228;
wire g25749;
wire g23582;
wire g21736;
wire g33609;
wire g8234;
wire g24584;
wire II33109;
wire g21779;
wire g24027;
wire g7050;
wire g22689;
wire g10032;
wire g33124;
wire g27679;
wire g21463;
wire g11183;
wire g14630;
wire g14940;
wire g34700;
wire g8180;
wire g31990;
wire g25717;
wire II18906;
wire g25132;
wire g11244;
wire g32748;
wire g30579;
wire g32204;
wire g23716;
wire g21353;
wire g14064;
wire g31914;
wire g33761;
wire g27500;
wire g19365;
wire g14902;
wire g14444;
wire g16632;
wire g17523;
wire g33646;
wire g9055;
wire g28981;
wire g21010;
wire g15160;
wire g23754;
wire g21049;
wire g30268;
wire g24631;
wire g7909;
wire g26080;
wire g34664;
wire g28178;
wire g31708;
wire II29013;
wire g19479;
wire g24323;
wire g32615;
wire g23042;
wire g24125;
wire II21477;
wire g29923;
wire g25607;
wire g7121;
wire g33687;
wire g17569;
wire II16538;
wire g33346;
wire g32792;
wire g31968;
wire g32164;
wire g32918;
wire g24407;
wire II28582;
wire g23742;
wire g28425;
wire g28215;
wire g25702;
wire gbuf95;
wire g13104;
wire g20562;
wire g31324;
wire g27372;
wire gbuf136;
wire g28358;
wire g18610;
wire g22053;
wire g24261;
wire g27990;
wire g33456;
wire g34350;
wire g29795;
wire g34580;
wire g16675;
wire g19410;
wire g19530;
wire g13084;
wire g26286;
wire g19061;
wire g32799;
wire g28285;
wire g33119;
wire g11415;
wire g30083;
wire II18367;
wire g25709;
wire g10710;
wire g30452;
wire g17096;
wire II27518;
wire g12885;
wire g27012;
wire g29171;
wire II29002;
wire g12908;
wire g12028;
wire II32696;
wire g18988;
wire g15814;
wire g19394;
wire II14046;
wire g27147;
wire gbuf128;
wire g24018;
wire g28900;
wire g29081;
wire g8873;
wire g32965;
wire g28312;
wire II23684;
wire g18715;
wire g11372;
wire g23249;
wire g34492;
wire g13298;
wire g10290;
wire g14001;
wire II12826;
wire g30052;
wire g11279;
wire g28727;
wire II32062;
wire g18382;
wire g13042;
wire II14499;
wire g33895;
wire II21787;
wire II29204;
wire g9402;
wire g32570;
wire g24989;
wire g29915;
wire g33864;
wire g13311;
wire g17014;
wire g11867;
wire g31667;
wire g14277;
wire g24011;
wire g29594;
wire g14212;
wire II15308;
wire II29296;
wire g33112;
wire g29369;
wire g18230;
wire g13069;
wire g27586;
wire g34862;
wire g32833;
wire g25015;
wire g14342;
wire g23849;
wire g10207;
wire g16290;
wire g30374;
wire g8345;
wire g8745;
wire g10554;
wire g18766;
wire g34707;
wire g24304;
wire g34338;
wire g30729;
wire g12222;
wire g28280;
wire II13473;
wire g25240;
wire g19128;
wire g24881;
wire II33161;
wire g30387;
wire g16605;
wire g7927;
wire g30179;
wire g33657;
wire g33244;
wire II13548;
wire II18492;
wire II15195;
wire g32325;
wire g12020;
wire g27328;
wire g16536;
wire g26274;
wire g26252;
wire II12719;
wire g19785;
wire g25647;
wire g13264;
wire g28455;
wire g32141;
wire g26327;
wire g34428;
wire g27342;
wire g33958;
wire g25695;
wire g33360;
wire g21427;
wire g9390;
wire g29970;
wire II32994;
wire g31997;
wire g18342;
wire g22096;
wire g32693;
wire II32997;
wire g13993;
wire g25541;
wire II18304;
wire II24582;
wire g32672;
wire g33367;
wire g18629;
wire II16610;
wire g25762;
wire g24357;
wire g14228;
wire g31245;
wire g12824;
wire g26968;
wire II14644;
wire g28517;
wire II18320;
wire g26244;
wire g34371;
wire g33504;
wire g34981;
wire g29129;
wire g18979;
wire g7087;
wire g11012;
wire g26346;
wire g24033;
wire II15593;
wire g33620;
wire g14511;
wire g24893;
wire g34975;
wire g34721;
wire g31523;
wire g28601;
wire g16528;
wire II33214;
wire g13597;
wire g28730;
wire g34046;
wire g20450;
wire g8740;
wire g24234;
wire g34059;
wire g10822;
wire g32520;
wire g12478;
wire g23893;
wire II22619;
wire g20978;
wire II19235;
wire g20697;
wire g32736;
wire II16770;
wire g10367;
wire g24756;
wire g24700;
wire g33516;
wire g24950;
wire g15823;
wire g8057;
wire II24365;
wire g13727;
wire g24489;
wire g14098;
wire II13044;
wire g18816;
wire g11677;
wire g18624;
wire g22641;
wire II17834;
wire g28739;
wire g32367;
wire g26393;
wire g26770;
wire g20682;
wire g7349;
wire g23059;
wire g25046;
wire g17634;
wire g21678;
wire g26777;
wire g26936;
wire II24445;
wire g27121;
wire g33934;
wire II20399;
wire g16243;
wire II11864;
wire g14520;
wire g33250;
wire g23835;
wire g25041;
wire II25221;
wire g27696;
wire g27265;
wire g20648;
wire g29110;
wire g32458;
wire g16777;
wire g18430;
wire g15655;
wire g16684;
wire II24505;
wire g32017;
wire g14643;
wire g27559;
wire g21974;
wire II16660;
wire II14764;
wire g16423;
wire II32185;
wire g32569;
wire g20057;
wire g13857;
wire g16965;
wire g24650;
wire g17683;
wire g28299;
wire gbuf79;
wire g12460;
wire g30127;
wire g23165;
wire g25937;
wire g11428;
wire g17198;
wire g21843;
wire g30352;
wire g33260;
wire g12198;
wire g34954;
wire g25101;
wire g32387;
wire g34510;
wire II18845;
wire g28251;
wire g27670;
wire g12656;
wire g34612;
wire g33380;
wire g23356;
wire g25529;
wire gbuf145;
wire g20093;
wire g24245;
wire g33143;
wire g31887;
wire g19335;
wire g18727;
wire g15736;
wire g9992;
wire gbuf51;
wire g30215;
wire g9691;
wire II13539;
wire g19541;
wire g34751;
wire g21807;
wire g28064;
wire g34860;
wire g32871;
wire g24577;
wire g10362;
wire g27128;
wire g18686;
wire g27829;
wire g15159;
wire g32937;
wire g9749;
wire g34440;
wire g16867;
wire g14999;
wire II14899;
wire g34733;
wire g20025;
wire g17309;
wire g22108;
wire g13798;
wire g34111;
wire g19951;
wire II18716;
wire g13697;
wire gbuf8;
wire II29965;
wire g27647;
wire g28324;
wire g15120;
wire II31107;
wire g16760;
wire g34943;
wire g24772;
wire g18313;
wire g28106;
wire g25988;
wire II32051;
wire g29518;
wire g32172;
wire g12898;
wire g18169;
wire g31296;
wire g34935;
wire g33288;
wire g32921;
wire g28156;
wire g22216;
wire g33371;
wire g21402;
wire g33534;
wire II31782;
wire gbuf27;
wire II13510;
wire g6955;
wire g21936;
wire g10379;
wire II12372;
wire g30541;
wire g30082;
wire g29765;
wire g25409;
wire g33376;
wire g32508;
wire g29489;
wire gbuf20;
wire g32040;
wire g23967;
wire g9576;
wire II26578;
wire g30047;
wire II21029;
wire g33420;
wire g16700;
wire g18947;
wire g13409;
wire g22153;
wire g11293;
wire g20153;
wire gbuf42;
wire II12382;
wire g27484;
wire g33885;
wire g27035;
wire g13252;
wire g13544;
wire g22830;
wire g15794;
wire II31006;
wire g33046;
wire g33858;
wire g24722;
wire g34858;
wire g14160;
wire g34310;
wire g18603;
wire g32585;
wire g33083;
wire g7301;
wire II15051;
wire g22682;
wire g18722;
wire g29744;
wire g34797;
wire g33702;
wire g28560;
wire g21865;
wire g18545;
wire g29057;
wire g33443;
wire g20770;
wire II12963;
wire II12530;
wire g34182;
wire II18538;
wire g30594;
wire II27364;
wire g23850;
wire g26886;
wire g22158;
wire g28374;
wire II32935;
wire g32150;
wire g11178;
wire g29168;
wire g15856;
wire g12846;
wire g19566;
wire g30481;
wire g29616;
wire g31070;
wire g22104;
wire g11302;
wire g22083;
wire g21156;
wire g16431;
wire g14272;
wire g21271;
wire g20005;
wire g22048;
wire g25071;
wire g27349;
wire g33282;
wire g26352;
wire g6756;
wire g32719;
wire g23947;
wire g33802;
wire g15732;
wire g30436;
wire g14163;
wire II25366;
wire II27564;
wire II11878;
wire g29032;
wire g14209;
wire g29186;
wire g31148;
wire g29968;
wire g32811;
wire g29276;
wire g10568;
wire g25095;
wire g21399;
wire g20164;
wire g29861;
wire g25750;
wire g27600;
wire g34773;
wire II12026;
wire g21302;
wire g11511;
wire g18365;
wire II15262;
wire g17242;
wire g18696;
wire g12259;
wire g25573;
wire II27730;
wire g26905;
wire g17745;
wire g25198;
wire g31285;
wire g15800;
wire g23547;
wire g23932;
wire g33299;
wire II25786;
wire g23611;
wire g14279;
wire g34568;
wire g7392;
wire g34160;
wire II12611;
wire g28559;
wire g12779;
wire g21743;
wire g21854;
wire II19917;
wire g18987;
wire g8791;
wire g21890;
wire g17817;
wire g13144;
wire g7643;
wire g26267;
wire g16260;
wire g33927;
wire g20371;
wire g27930;
wire g29028;
wire g21193;
wire g28521;
wire g34255;
wire g10312;
wire g28684;
wire g29774;
wire g25370;
wire g10157;
wire g6800;
wire g24639;
wire g34989;
wire g27555;
wire g31300;
wire g26363;
wire g27255;
wire g22114;
wire II12728;
wire g16969;
wire II31292;
wire g31220;
wire g19483;
wire g31240;
wire g14330;
wire g26792;
wire g16582;
wire II31535;
wire g8964;
wire g15070;
wire g20659;
wire g16523;
wire g16099;
wire g11666;
wire g29669;
wire g12869;
wire g22171;
wire g18823;
wire g32999;
wire g21991;
wire g28430;
wire g6917;
wire g32596;
wire g24672;
wire II31196;
wire g26248;
wire g23085;
wire g23822;
wire g29344;
wire II17989;
wire II14241;
wire g29717;
wire g29286;
wire g34608;
wire g31496;
wire g28492;
wire g16587;
wire II13937;
wire g24657;
wire g30508;
wire g18308;
wire gbuf141;
wire g30102;
wire g7673;
wire g14406;
wire g7436;
wire g33996;
wire g34189;
wire g29237;
wire II32929;
wire g27239;
wire g24047;
wire g21410;
wire g32866;
wire g28132;
wire g18411;
wire II32904;
wire II17098;
wire II27524;
wire g28142;
wire g34269;
wire g34214;
wire II30469;
wire g25193;
wire II32967;
wire g17249;
wire g29646;
wire g22654;
wire g20132;
wire g7594;
wire g24977;
wire g8928;
wire g25848;
wire II31137;
wire g23929;
wire g33572;
wire g27177;
wire g19879;
wire g10531;
wire II12544;
wire g24272;
wire g28428;
wire g23446;
wire g28556;
wire g34563;
wire g9372;
wire II23961;
wire g12894;
wire g25881;
wire g14946;
wire g20113;
wire g23751;
wire g25929;
wire g15741;
wire g18635;
wire g16735;
wire II21976;
wire g15978;
wire g29230;
wire g9645;
wire g14697;
wire g24808;
wire g27405;
wire g30188;
wire g21249;
wire g8906;
wire g18574;
wire g32380;
wire g33709;
wire g32817;
wire g22524;
wire g32392;
wire g21051;
wire g22594;
wire g18317;
wire g18478;
wire II22604;
wire g25974;
wire g17515;
wire II29254;
wire gbuf131;
wire g21764;
wire g12721;
wire g30243;
wire g28390;
wire g28300;
wire g25623;
wire g28389;
wire g29203;
wire g27241;
wire g14678;
wire II31121;
wire g24963;
wire g25875;
wire g22168;
wire g25211;
wire g26670;
wire g29854;
wire g30400;
wire g25450;
wire g16713;
wire g30275;
wire g34624;
wire g6855;
wire g9924;
wire g17953;
wire g23574;
wire g25997;
wire g14357;
wire g20214;
wire g28586;
wire g15608;
wire g34121;
wire g18784;
wire g16172;
wire g17396;
wire g21369;
wire II15821;
wire g22871;
wire g17518;
wire g34710;
wire g32705;
wire II14687;
wire II13634;
wire gbuf81;
wire II20486;
wire II15176;
wire II26409;
wire g24070;
wire g29069;
wire g32903;
wire II20867;
wire g23540;
wire g28830;
wire g19356;
wire g33614;
wire II32591;
wire g9003;
wire g10382;
wire g34208;
wire g16228;
wire g19866;
wire II32775;
wire g26093;
wire g18294;
wire g32030;
wire g28494;
wire g29620;
wire g26547;
wire g7479;
wire II31336;
wire g11119;
wire g12837;
wire g34079;
wire II17873;
wire g21291;
wire g25684;
wire g17144;
wire g16621;
wire g12115;
wire g33073;
wire g34918;
wire II14346;
wire g26397;
wire g22068;
wire g30443;
wire II32843;
wire g9601;
wire g19574;
wire g31259;
wire II15298;
wire g32039;
wire g7765;
wire g27985;
wire g29961;
wire g28564;
wire g22866;
wire g25323;
wire II12064;
wire g33691;
wire g34754;
wire g9967;
wire g25223;
wire g22651;
wire II18574;
wire II19799;
wire g29746;
wire g23840;
wire g30258;
wire g19799;
wire g33537;
wire II17932;
wire g12227;
wire g9631;
wire g9983;
wire g23902;
wire g22358;
wire g11936;
wire g27665;
wire g32045;
wire g33730;
wire g15837;
wire g8480;
wire g22128;
wire g30397;
wire II17924;
wire g29339;
wire g34396;
wire II18180;
wire g23518;
wire g33726;
wire g33588;
wire g12680;
wire g21070;
wire g14258;
wire g18194;
wire g23299;
wire g13046;
wire g21160;
wire II26438;
wire g23000;
wire g22845;
wire g25545;
wire g14845;
wire II31227;
wire g14867;
wire g17773;
wire g30112;
wire II22331;
wire g19442;
wire g32986;
wire g34229;
wire g23386;
wire II31087;
wire g18148;
wire g23541;
wire g18893;
wire g15714;
wire g17482;
wire II16452;
wire g26781;
wire g21611;
wire g26313;
wire g31764;
wire g26236;
wire g27433;
wire g7995;
wire g25551;
wire g14119;
wire g11618;
wire g6983;
wire g32696;
wire g20231;
wire g12194;
wire g33530;
wire g25285;
wire g27480;
wire g12153;
wire g22494;
wire gbuf103;
wire g30556;
wire g34881;
wire II14883;
wire g21935;
wire g25900;
wire g17476;
wire g16196;
wire g25127;
wire g15903;
wire g9694;
wire g24402;
wire g13257;
wire g34414;
wire g21251;
wire g21942;
wire gbuf115;
wire g20660;
wire g12553;
wire g23907;
wire g26648;
wire g20072;
wire II26643;
wire g19789;
wire g20196;
wire g30991;
wire g30438;
wire g27101;
wire g31226;
wire g24916;
wire g12183;
wire II31201;
wire g14226;
wire g28417;
wire II18341;
wire g23520;
wire g24855;
wire II13852;
wire g11951;
wire g34819;
wire g9626;
wire g33085;
wire g27204;
wire g24712;
wire g23681;
wire g28218;
wire g34939;
wire II31607;
wire II32868;
wire g23361;
wire g29041;
wire g14110;
wire II20468;
wire g15595;
wire g31903;
wire g21830;
wire g31291;
wire g14151;
wire g18630;
wire g25735;
wire g16127;
wire g23404;
wire g30474;
wire g34366;
wire g16540;
wire II15837;
wire g27993;
wire g28034;
wire II31262;
wire g28667;
wire g34222;
wire g9685;
wire g16923;
wire g22708;
wire g32340;
wire g18808;
wire g19587;
wire g34101;
wire g31478;
wire g24094;
wire g26342;
wire g32994;
wire g19633;
wire g28530;
wire g34575;
wire g17315;
wire g20238;
wire g24307;
wire II16217;
wire II27539;
wire g20595;
wire g34346;
wire g16757;
wire g34607;
wire g23124;
wire g28476;
wire g30036;
wire g32479;
wire g30530;
wire g26296;
wire g24750;
wire g7558;
wire g26973;
wire g20189;
wire g29999;
wire g34274;
wire g15104;
wire g23318;
wire II32231;
wire g11534;
wire g8948;
wire g21388;
wire g27306;
wire g11136;
wire g7557;
wire g23620;
wire g14385;
wire g24352;
wire g25660;
wire g12587;
wire g30091;
wire II22745;
wire g32755;
wire g32236;
wire g22940;
wire g21669;
wire g8571;
wire g25042;
wire g25299;
wire g26281;
wire g24934;
wire g32129;
wire g11561;
wire g22758;
wire g18330;
wire g33276;
wire g11975;
wire g26839;
wire g30379;
wire II16289;
wire II13236;
wire g30410;
wire II28913;
wire g30416;
wire g22073;
wire g23887;
wire g26865;
wire g24227;
wire g27284;
wire g34026;
wire g32876;
wire g13306;
wire g18536;
wire g29568;
wire g8530;
wire g24374;
wire g30419;
wire g32404;
wire g21961;
wire g34423;
wire g28370;
wire gbuf6;
wire g19505;
wire II16606;
wire g33408;
wire g31827;
wire g22905;
wire g22716;
wire g33032;
wire g23462;
wire g10200;
wire g32240;
wire g24346;
wire g27137;
wire g28360;
wire g34035;
wire g34086;
wire g32321;
wire g26278;
wire g6874;
wire g24786;
wire II16401;
wire g20923;
wire g19773;
wire II16468;
wire g12738;
wire g14124;
wire g26915;
wire g28623;
wire II15590;
wire g9640;
wire g34911;
wire g28401;
wire II23363;
wire II31206;
wire g25778;
wire II25555;
wire g9467;
wire g20583;
wire g8125;
wire g32223;
wire g23608;
wire g27723;
wire g29843;
wire g22639;
wire g32385;
wire g26912;
wire g31519;
wire g29598;
wire g32764;
wire g10874;
wire g7617;
wire g10665;
wire g29365;
wire g25659;
wire g33059;
wire g14953;
wire g10733;
wire II21230;
wire g10759;
wire g16897;
wire g17759;
wire g11473;
wire II31167;
wire g29800;
wire g25189;
wire g32936;
wire g32306;
wire g33698;
wire g9815;
wire g24030;
wire g31182;
wire g27379;
wire g24636;
wire II11617;
wire g29903;
wire g12207;
wire g19265;
wire g27587;
wire II32837;
wire g29585;
wire g24423;
wire g33912;
wire gbuf16;
wire g24087;
wire g18061;
wire g27041;
wire II30717;
wire II18526;
wire II14079;
wire g27274;
wire g20915;
wire g27552;
wire g18584;
wire II17476;
wire g14411;
wire g14723;
wire g21923;
wire g27440;
wire g30613;
wire g10934;
wire g6836;
wire g32654;
wire g8591;
wire II12878;
wire II22938;
wire g24866;
wire g24686;
wire g34303;
wire II24689;
wire g32503;
wire g17509;
wire g12591;
wire g18105;
wire g34090;
wire g26965;
wire g25851;
wire g25982;
wire II18682;
wire g23590;
wire g30307;
wire g30170;
wire g29600;
wire g21424;
wire g20274;
wire g29506;
wire g19276;
wire g23321;
wire g12413;
wire g30139;
wire g12066;
wire II22754;
wire g32718;
wire g9380;
wire g29384;
wire g12762;
wire g29752;
wire g31287;
wire g10820;
wire g29977;
wire g11223;
wire II17447;
wire g27019;
wire g25206;
wire g29271;
wire g31745;
wire g34847;
wire g20916;
wire g18488;
wire g22020;
wire g11705;
wire g24202;
wire g21185;
wire g23067;
wire g33160;
wire g28489;
wire g27350;
wire II30992;
wire g12333;
wire g9778;
wire g28914;
wire g24311;
wire g9568;
wire g30368;
wire II31097;
wire II32431;
wire g17611;
wire g11772;
wire g27877;
wire g33187;
wire g24417;
wire g25973;
wire g30116;
wire g20709;
wire II24461;
wire g15572;
wire g20203;
wire g20773;
wire II30959;
wire g24197;
wire II12749;
wire g32823;
wire g32147;
wire g34992;
wire g26273;
wire g27767;
wire g24709;
wire g29231;
wire g34570;
wire g23493;
wire g30522;
wire II32203;
wire II12811;
wire g29208;
wire II28419;
wire g7717;
wire II11623;
wire II26309;
wire II24839;
wire g32155;
wire II25105;
wire g10487;
wire g29533;
wire g32518;
wire g33433;
wire g25961;
wire g14832;
wire g22059;
wire g23302;
wire g16161;
wire g18274;
wire g13057;
wire g34203;
wire g15705;
wire g24291;
wire II24038;
wire g10143;
wire g29194;
wire II14213;
wire g10707;
wire g11165;
wire II17814;
wire g18702;
wire g18359;
wire g29750;
wire g23397;
wire g34097;
wire g23924;
wire g28085;
wire g25764;
wire II32243;
wire II31047;
wire g27223;
wire g28246;
wire g15110;
wire g24792;
wire g15483;
wire g30573;
wire g29988;
wire g18883;
wire g28084;
wire II18485;
wire g18554;
wire g22536;
wire g32069;
wire g19610;
wire g9239;
wire g16745;
wire g27353;
wire g11969;
wire g17768;
wire g35000;
wire g28931;
wire II15306;
wire g12317;
wire g9461;
wire g17420;
wire g24467;
wire g24268;
wire g20008;
wire g20499;
wire g23764;
wire g21139;
wire g12968;
wire g23426;
wire g20504;
wire g20147;
wire g20067;
wire g21815;
wire g25548;
wire g16286;
wire g17326;
wire g28708;
wire g33652;
wire g30173;
wire II15448;
wire g28638;
wire g21853;
wire gbuf88;
wire g27087;
wire II14955;
wire g21885;
wire g26299;
wire g24318;
wire II16391;
wire g9483;
wire gbuf69;
wire g28576;
wire g25507;
wire g29374;
wire g7880;
wire g21756;
wire gbuf90;
wire g25435;
wire II31864;
wire gbuf13;
wire g34840;
wire II18460;
wire g15154;
wire g10084;
wire g32890;
wire II26466;
wire II24018;
wire g34654;
wire g30567;
wire g32486;
wire g18156;
wire g31115;
wire g14448;
wire g30313;
wire g28127;
wire g24116;
wire II18785;
wire g16206;
wire g34874;
wire g22007;
wire g7322;
wire g21771;
wire g13060;
wire g10572;
wire g25741;
wire g26052;
wire g7564;
wire g30516;
wire g23937;
wire g29323;
wire II11655;
wire g30218;
wire g18591;
wire g22369;
wire g20104;
wire g32531;
wire g26512;
wire g22667;
wire g18627;
wire g33039;
wire II15166;
wire g8608;
wire g24161;
wire g34791;
wire g14314;
wire II13094;
wire g18751;
wire g23606;
wire g21706;
wire g9744;
wire g20702;
wire g23390;
wire g24102;
wire g25652;
wire g15753;
wire g25917;
wire g23576;
wire g29524;
wire g34431;
wire g32625;
wire g29878;
wire g15884;
wire g18933;
wire g11468;
wire g34585;
wire g19714;
wire g32875;
wire g21400;
wire g31910;
wire g16303;
wire g10803;
wire II31504;
wire g23255;
wire g7805;
wire g9663;
wire II31322;
wire g12087;
wire g23599;
wire g8769;
wire g16615;
wire g21801;
wire g24339;
wire g34009;
wire II15287;
wire g29647;
wire g16591;
wire g26843;
wire g34732;
wire II18293;
wire g34317;
wire g24995;
wire g24203;
wire g12640;
wire II26522;
wire g28673;
wire g21958;
wire g30920;
wire II18875;
wire II31172;
wire g14637;
wire g9761;
wire g30145;
wire g6990;
wire II13497;
wire II29969;
wire g19068;
wire g13580;
wire g10622;
wire g26181;
wire g7933;
wire g18130;
wire II31555;
wire II32103;
wire g12118;
wire g27954;
wire g23374;
wire g17504;
wire g13522;
wire g7267;
wire g13283;
wire g8733;
wire g13288;
wire g16729;
wire g27210;
wire II24393;
wire g28504;
wire g34715;
wire g20634;
wire g20432;
wire g17789;
wire g29981;
wire g34181;
wire II24546;
wire g28604;
wire g25025;
wire II11824;
wire g9960;
wire g14583;
wire II12176;
wire g27224;
wire g31009;
wire II31463;
wire g27563;
wire g34559;
wire g33548;
wire g10411;
wire g28780;
wire g20037;
wire g8218;
wire g15612;
wire g13036;
wire g32194;
wire g20714;
wire II17128;
wire g28329;
wire g22760;
wire II12092;
wire II18700;
wire g34096;
wire II19818;
wire g15805;
wire g22849;
wire g13932;
wire g33509;
wire II24228;
wire g10352;
wire g32263;
wire II27349;
wire g18561;
wire g33014;
wire g18145;
wire g24383;
wire II17425;
wire g29893;
wire g21379;
wire g7624;
wire g23305;
wire g18460;
wire II12074;
wire g30162;
wire g33354;
wire g22357;
wire g15717;
wire g26148;
wire g24646;
wire g12036;
wire g28852;
wire g24134;
wire g21278;
wire g29001;
wire II18518;
wire g23188;
wire g30318;
wire II24022;
wire g17602;
wire g26336;
wire g20606;
wire g30548;
wire g14419;
wire g32800;
wire II23351;
wire g25867;
wire g34742;
wire g22101;
wire g28593;
wire g22136;
wire II16626;
wire g34335;
wire g32560;
wire g28645;
wire g34590;
wire g33313;
wire g24549;
wire g8229;
wire g22014;
wire g24668;
wire g14176;
wire g31835;
wire g24077;
wire g12358;
wire g22305;
wire g31143;
wire g32647;
wire g6999;
wire g17191;
wire g30917;
wire II31001;
wire g16699;
wire g28093;
wire g31638;
wire g21682;
wire g17086;
wire g10387;
wire g23250;
wire II31622;
wire g13634;
wire II22946;
wire g20014;
wire g21787;
wire II13520;
wire II23969;
wire g20443;
wire II33258;
wire g27494;
wire g15589;
wire g11355;
wire g11679;
wire g32687;
wire g22854;
wire g14912;
wire g28233;
wire g13527;
wire g12467;
wire g18446;
wire g33466;
wire g15080;
wire g31882;
wire g14677;
wire g11450;
wire g33338;
wire g20552;
wire g21409;
wire g31068;
wire g34558;
wire g34118;
wire g15087;
wire g7516;
wire II18238;
wire g33255;
wire g16000;
wire g22207;
wire g16598;
wire g24215;
wire g18705;
wire g27658;
wire g25186;
wire g10795;
wire g23191;
wire II17612;
wire g8725;
wire g29787;
wire g16691;
wire g14610;
wire g13570;
wire II15893;
wire g14566;
wire g23897;
wire g28549;
wire g26360;
wire g34801;
wire g32179;
wire g9792;
wire g33135;
wire II22760;
wire g18609;
wire g25367;
wire g20010;
wire g12911;
wire g25466;
wire g8070;
wire g17124;
wire g24348;
wire g13349;
wire g8404;
wire g26898;
wire g15782;
wire g32733;
wire g9688;
wire g24214;
wire g30199;
wire g9729;
wire gbuf153;
wire g25888;
wire g22409;
wire g23015;
wire II24075;
wire II29214;
wire g14987;
wire g10150;
wire g33720;
wire g19962;
wire g21295;
wire g33061;
wire g16234;
wire g24680;
wire g24452;
wire g21430;
wire g8841;
wire g13883;
wire g8848;
wire g27262;
wire g18905;
wire g14719;
wire g25078;
wire g22035;
wire g34562;
wire g11990;
wire g26851;
wire g33557;
wire g15818;
wire g17121;
wire g21994;
wire II23756;
wire g14035;
wire g14248;
wire g20513;
wire g34969;
wire g20326;
wire g18248;
wire g28263;
wire g22146;
wire g16231;
wire g31856;
wire g16514;
wire g24505;
wire g32255;
wire g28541;
wire g12296;
wire g12462;
wire gbuf70;
wire g27217;
wire g13342;
wire II12227;
wire g23355;
wire g18513;
wire g21701;
wire g31988;
wire g30003;
wire g30078;
wire g30066;
wire g30457;
wire g32898;
wire g29379;
wire g29839;
wire g24679;
wire g27463;
wire g17325;
wire g23439;
wire g28386;
wire g34051;
wire g28710;
wire g33963;
wire g25245;
wire II24527;
wire g32880;
wire g10357;
wire g32362;
wire g10179;
wire g28666;
wire II28002;
wire g30183;
wire g20451;
wire g9907;
wire g25170;
wire g34948;
wire g28130;
wire g22897;
wire g15651;
wire g13794;
wire g21985;
wire g33057;
wire g24651;
wire g18315;
wire g23341;
wire g10917;
wire g13793;
wire g33519;
wire g26155;
wire II17658;
wire g32012;
wire g19948;
wire g27510;
wire g17676;
wire g18062;
wire g30590;
wire g17415;
wire g25759;
wire g10042;
wire g24517;
wire g34511;
wire g14555;
wire II18221;
wire g27116;
wire g13431;
wire g12772;
wire g14089;
wire g19585;
wire g32576;
wire g7763;
wire g14851;
wire g27773;
wire g15072;
wire g19781;
wire g15722;
wire g30357;
wire g28519;
wire g11249;
wire g34375;
wire g33031;
wire g29810;
wire g30141;
wire g28010;
wire g28871;
wire g34426;
wire II31317;
wire g18235;
wire g25716;
wire g7352;
wire g18980;
wire g24884;
wire g7314;
wire g13971;
wire g16869;
wire g12811;
wire g10571;
wire II33020;
wire g18219;
wire g34859;
wire II23366;
wire g33358;
wire g34506;
wire g25966;
wire g29477;
wire g7867;
wire g31242;
wire g10666;
wire g33981;
wire g18567;
wire g26123;
wire g33847;
wire g7696;
wire g16427;
wire g10561;
wire g11325;
wire g31829;
wire g16774;
wire g8728;
wire g17585;
wire g10998;
wire g33256;
wire g15693;
wire g9715;
wire g20696;
wire g24587;
wire g28261;
wire g17473;
wire g16724;
wire g13101;
wire g19398;
wire g13593;
wire g18747;
wire g28510;
wire II32297;
wire g13140;
wire g33448;
wire gbuf71;
wire g13604;
wire g28256;
wire g31879;
wire g19337;
wire II15106;
wire g33525;
wire g20083;
wire g28077;
wire II18832;
wire II14862;
wire g7073;
wire g11424;
wire g21804;
wire II22929;
wire II16829;
wire g20776;
wire g34983;
wire II12144;
wire g12085;
wire II27271;
wire g7192;
wire g13928;
wire g28266;
wire g29844;
wire g13662;
wire g29762;
wire II12954;
wire g22839;
wire g10176;
wire g19491;
wire II12907;
wire g34887;
wire g24944;
wire g26381;
wire g13700;
wire g31526;
wire g29611;
wire g34617;
wire II12109;
wire g12256;
wire g28523;
wire g22213;
wire g8112;
wire g28721;
wire g29225;
wire g31120;
wire g31964;
wire g32723;
wire g19498;
wire g34007;
wire g34348;
wire g12173;
wire g16200;
wire g13846;
wire g19979;
wire g33716;
wire g7626;
wire g30599;
wire g16424;
wire g30369;
wire g33508;
wire II17704;
wire g19947;
wire g34964;
wire g22132;
wire g26324;
wire g33693;
wire g20616;
wire g31798;
wire II14291;
wire g19744;
wire g18760;
wire g30543;
wire g7523;
wire g31127;
wire g23882;
wire g18220;
wire II15250;
wire g32109;
wire g26916;
wire g18792;
wire g28671;
wire II27192;
wire II21734;
wire g28039;
wire g26947;
wire g34319;
wire g17776;
wire g31015;
wire g34995;
wire g28327;
wire II17653;
wire II17839;
wire g18677;
wire II22973;
wire g28284;
wire g17748;
wire g13709;
wire g13946;
wire II32645;
wire g27503;
wire g28735;
wire g28060;
wire g33249;
wire g27488;
wire g26853;
wire g13736;
wire g28290;
wire g27127;
wire g24390;
wire g23675;
wire g32266;
wire g11034;
wire g17405;
wire g25389;
wire g25470;
wire g24490;
wire g19554;
wire g10625;
wire g31706;
wire g34243;
wire g25705;
wire II31032;
wire g28939;
wire II31849;
wire g27222;
wire g13074;
wire g32372;
wire g18520;
wire II15033;
wire g27259;
wire g20382;
wire g25800;
wire g29484;
wire g17681;
wire g12797;
wire g27515;
wire g23733;
wire g24002;
wire II26679;
wire g34325;
wire g32111;
wire g25117;
wire g24168;
wire g16680;
wire g7023;
wire g31189;
wire II18048;
wire g12883;
wire g13517;
wire g6989;
wire g33001;
wire g28817;
wire g24997;
wire g33340;
wire g24484;
wire g32095;
wire g8680;
wire g10374;
wire g19510;
wire g29514;
wire g10366;
wire g25150;
wire g18687;
wire II15869;
wire g12979;
wire g15123;
wire g18501;
wire g32347;
wire g11913;
wire II27481;
wire g26311;
wire g18549;
wire g9750;
wire g18713;
wire g23231;
wire g26845;
wire g27400;
wire g11706;
wire g10320;
wire II25579;
wire g19981;
wire g18974;
wire g32186;
wire g8558;
wire g10410;
wire g28594;
wire g26050;
wire g33013;
wire g29284;
wire g13315;
wire g12293;
wire g24983;
wire g12893;
wire g20507;
wire g28665;
wire g10618;
wire g21334;
wire g27407;
wire g29631;
wire g22091;
wire g13176;
wire g9951;
wire g34044;
wire II14370;
wire gbuf60;
wire g33898;
wire II14964;
wire g16671;
wire II14230;
wire g16668;
wire g29042;
wire g22157;
wire g9678;
wire g29322;
wire g19735;
wire II32809;
wire g28274;
wire g23027;
wire g33038;
wire g17756;
wire g12226;
wire g12163;
wire g13080;
wire g8186;
wire g13108;
wire g21357;
wire g33114;
wire g24580;
wire g14180;
wire g21355;
wire II29261;
wire gbuf64;
wire gbuf139;
wire g8673;
wire II13287;
wire g27335;
wire g27104;
wire g25018;
wire g29596;
wire g17820;
wire II31191;
wire II24440;
wire g14825;
wire g34012;
wire g25790;
wire g16626;
wire g31321;
wire g34126;
wire g17521;
wire g34759;
wire II12709;
wire g14513;
wire II21250;
wire g30241;
wire g32339;
wire g24316;
wire g14339;
wire II30193;
wire II15906;
wire g10499;
wire g33043;
wire g24645;
wire g8340;
wire g30305;
wire g29144;
wire g33122;
wire g19687;
wire g18161;
wire g32154;
wire g24952;
wire g27031;
wire g24153;
wire g22921;
wire II16077;
wire g32743;
wire II12086;
wire II14305;
wire g33563;
wire g23384;
wire g32773;
wire II24787;
wire g24023;
wire g8033;
wire g32132;
wire g28579;
wire g19579;
wire g33146;
wire g26545;
wire g14875;
wire g21732;
wire II12546;
wire g31971;
wire g29792;
wire g25080;
wire II12132;
wire II19837;
wire g9644;
wire g14101;
wire g31500;
wire g27237;
wire g23331;
wire g8876;
wire g19734;
wire g7202;
wire g12946;
wire g31133;
wire g30146;
wire II12469;
wire g8456;
wire g28150;
wire g8064;
wire g32704;
wire g10395;
wire g34458;
wire g31748;
wire g17641;
wire g34389;
wire g22541;
wire g25481;
wire g12023;
wire g26085;
wire g32534;
wire g26084;
wire g22399;
wire g12437;
wire g29622;
wire g25821;
wire g24619;
wire g28032;
wire g20523;
wire g33999;
wire g32342;
wire g25641;
wire g21408;
wire g16215;
wire g15758;
wire g11273;
wire g31670;
wire g12980;
wire g20046;
wire g18477;
wire g11441;
wire g12145;
wire g10726;
wire g16531;
wire g21849;
wire g32582;
wire g27263;
wire g26162;
wire g11419;
wire II14331;
wire II31132;
wire II32446;
wire g9638;
wire g21694;
wire g17093;
wire g10881;
wire g25568;
wire g16155;
wire g25633;
wire g12848;
wire g22751;
wire g14015;
wire g18408;
wire g9808;
wire g34692;
wire g13241;
wire g28289;
wire g25939;
wire g24601;
wire g27014;
wire g19473;
wire g6767;
wire g33280;
wire g33366;
wire g32009;
wire g29228;
wire II15636;
wire g23586;
wire g26962;
wire g34863;
wire gbuf123;
wire g15734;
wire g12515;
wire g30169;
wire g13064;
wire g29887;
wire g27646;
wire g28641;
wire g11609;
wire g34696;
wire g10231;
wire g22193;
wire g19395;
wire g20162;
wire g11185;
wire g26378;
wire g13385;
wire g10158;
wire g23246;
wire g15479;
wire g26350;
wire g25984;
wire g11786;
wire g18948;
wire g24428;
wire g8068;
wire g26950;
wire g34384;
wire g12077;
wire g23819;
wire II13079;
wire II12217;
wire g7069;
wire g20386;
wire g9619;
wire g30214;
wire g29627;
wire g15680;
wire g14091;
wire g14688;
wire g28888;
wire g25969;
wire II24497;
wire g12037;
wire g33600;
wire g34302;
wire g21423;
wire g18423;
wire g19691;
wire g33952;
wire g19614;
wire g20910;
wire g32794;
wire g13877;
wire g18247;
wire g34802;
wire g28603;
wire g31996;
wire II20840;
wire II12262;
wire g16653;
wire g14237;
wire g19268;
wire g23338;
wire g18172;
wire g7003;
wire g26844;
wire g23645;
wire g10878;
wire g26309;
wire g32796;
wire g33891;
wire g25199;
wire g23226;
wire g22085;
wire g13670;
wire g29503;
wire g23373;
wire g9708;
wire II32991;
wire II20929;
wire g26899;
wire g32289;
wire g33070;
wire g34676;
wire g27957;
wire g14190;
wire g24242;
wire g25414;
wire g26255;
wire g24905;
wire g29309;
wire g33471;
wire g25011;
wire g30039;
wire g32973;
wire g30059;
wire g12432;
wire g23281;
wire g32467;
wire g11658;
wire g11810;
wire g26633;
wire g15969;
wire g29296;
wire g31855;
wire g9909;
wire g32460;
wire II23309;
wire g22064;
wire g25904;
wire g7635;
wire g33815;
wire g13997;
wire g24031;
wire g29104;
wire g22979;
wire g24368;
wire g32126;
wire g25543;
wire g18931;
wire g9728;
wire g14535;
wire g6828;
wire g18625;
wire g24186;
wire g28920;
wire g11231;
wire g10518;
wire g26611;
wire g15632;
wire g18812;
wire g21562;
wire g14797;
wire g29610;
wire g14545;
wire g18190;
wire g20582;
wire g6817;
wire g34023;
wire g21708;
wire II14429;
wire g19207;
wire g34509;
wire g11016;
wire II13875;
wire g27520;
wire gbuf142;
wire g30377;
wire II12487;
wire g14399;
wire g34377;
wire g7943;
wire g24403;
wire g34246;
wire g23555;
wire g32545;
wire g16044;
wire g31495;
wire g26654;
wire g34294;
wire g13092;
wire II30330;
wire g12558;
wire g12929;
wire II29891;
wire g17673;
wire g28051;
wire II13740;
wire g24353;
wire g16485;
wire g34537;
wire g25734;
wire g27995;
wire g34133;
wire II26394;
wire g24858;
wire g31768;
wire II17633;
wire g18616;
wire g8703;
wire g31255;
wire g28125;
wire g26349;
wire II26378;
wire g30502;
wire g22027;
wire g32698;
wire g7804;
wire g24249;
wire g9337;
wire g21432;
wire g11215;
wire g18636;
wire g25789;
wire g32768;
wire g8651;
wire II13672;
wire g34102;
wire g22332;
wire II30751;
wire g30090;
wire g34477;
wire g26710;
wire g21820;
wire g33857;
wire g32225;
wire g25932;
wire gbuf4;
wire g16509;
wire g28295;
wire g28091;
wire II33047;
wire g32490;
wire g19766;
wire g9970;
wire g16100;
wire g14033;
wire II15364;
wire g22856;
wire g32257;
wire g33485;
wire g32878;
wire g14221;
wire g31801;
wire g33742;
wire g34924;
wire g14437;
wire g33274;
wire g18367;
wire II17462;
wire g30475;
wire g18798;
wire II13462;
wire g8287;
wire g12486;
wire g23965;
wire g25958;
wire g11923;
wire g30931;
wire g18260;
wire g28161;
wire g20546;
wire g17478;
wire g15169;
wire g18357;
wire g20453;
wire g10951;
wire g32433;
wire g32556;
wire g8497;
wire g27185;
wire g22637;
wire g12123;
wire g25224;
wire g33889;
wire g10406;
wire g26302;
wire g30295;
wire g29939;
wire g20497;
wire g16192;
wire g20515;
wire II12855;
wire g11031;
wire g33162;
wire g29363;
wire g18695;
wire g23842;
wire g24089;
wire g23908;
wire g20615;
wire II20433;
wire g27564;
wire g27272;
wire g13256;
wire g31754;
wire g20192;
wire g29348;
wire g21795;
wire g28874;
wire g33478;
wire g31231;
wire g23859;
wire g7228;
wire II20529;
wire g23475;
wire g30317;
wire g22686;
wire g30559;
wire g12000;
wire g8010;
wire g19745;
wire II14369;
wire g26303;
wire g10180;
wire g20182;
wire g12692;
wire g12933;
wire g30211;
wire g23496;
wire g28565;
wire g13048;
wire g31765;
wire g7857;
wire g26818;
wire g19696;
wire g10216;
wire g28846;
wire g25927;
wire g8172;
wire g32913;
wire g8138;
wire g32397;
wire II32517;
wire g25214;
wire g33862;
wire g7536;
wire g16801;
wire g31317;
wire g27368;
wire g31902;
wire g19798;
wire g23001;
wire g21060;
wire g33413;
wire g12345;
wire g17139;
wire g29033;
wire g14529;
wire g23519;
wire g16727;
wire g17468;
wire g15579;
wire g19441;
wire g9739;
wire g32662;
wire g21725;
wire g32778;
wire g21069;
wire g18758;
wire g28319;
wire II32071;
wire g32867;
wire g25638;
wire g20781;
wire g8087;
wire II16541;
wire g24226;
wire g31791;
wire g12922;
wire g24131;
wire g34192;
wire g8500;
wire g15857;
wire g22902;
wire g22874;
wire g23490;
wire g33801;
wire g27456;
wire g32313;
wire g10114;
wire g21269;
wire g31277;
wire g24377;
wire g18280;
wire g23267;
wire g21719;
wire g32944;
wire g10490;
wire g16808;
wire g25558;
wire g33087;
wire g27524;
wire g30151;
wire g8679;
wire g30422;
wire g14146;
wire II23396;
wire g11906;
wire g34545;
wire g24058;
wire g18225;
wire g10334;
wire g31229;
wire g20641;
wire g33232;
wire g9913;
wire II29909;
wire g34689;
wire g22000;
wire g28113;
wire g15912;
wire g21412;
wire g10026;
wire g23451;
wire g8211;
wire g32802;
wire g27903;
wire g29245;
wire g16987;
wire g16031;
wire g26398;
wire g32028;
wire g17847;
wire g18258;
wire g18165;
wire g21891;
wire II14289;
wire g24510;
wire g21869;
wire g15155;
wire II28866;
wire g33269;
wire g13960;
wire g11492;
wire g31467;
wire g18426;
wire g32781;
wire g13478;
wire g27598;
wire g16326;
wire g33930;
wire II14352;
wire g30160;
wire g27178;
wire g28185;
wire II15335;
wire g17408;
wire g25035;
wire g34074;
wire g26207;
wire g13097;
wire II15550;
wire g31898;
wire g32868;
wire g26166;
wire g20445;
wire g11116;
wire g33759;
wire g30601;
wire g14695;
wire g33321;
wire g7017;
wire g33006;
wire II14475;
wire g17657;
wire g18555;
wire g26053;
wire g31275;
wire g20589;
wire g16927;
wire g13416;
wire g32552;
wire g33103;
wire g32386;
wire g33605;
wire g29165;
wire g30527;
wire g22535;
wire g15129;
wire g33391;
wire g23912;
wire g10278;
wire g27299;
wire g28611;
wire g19389;
wire g7462;
wire g24662;
wire g34629;
wire g21767;
wire g23032;
wire II31357;
wire g26146;
wire g23789;
wire g33653;
wire g31134;
wire g16173;
wire g8890;
wire g26200;
wire II18482;
wire g15932;
wire g23398;
wire g10223;
wire g33713;
wire g27064;
wire g19935;
wire g17794;
wire g23013;
wire g11350;
wire II32788;
wire g32667;
wire g7701;
wire II30734;
wire g28803;
wire g9686;
wire g34662;
wire g33027;
wire II12644;
wire g14204;
wire g8363;
wire g7850;
wire g21914;
wire g9824;
wire g32173;
wire g34727;
wire g18659;
wire g31504;
wire g14045;
wire II17507;
wire g32294;
wire g23218;
wire g28754;
wire g22592;
wire g18896;
wire g25602;
wire g24256;
wire g30338;
wire g18291;
wire g16319;
wire II16671;
wire g28917;
wire g29940;
wire g25624;
wire g32434;
wire g12739;
wire g11345;
wire g28209;
wire g34036;
wire g18916;
wire g19650;
wire g15979;
wire g18459;
wire g32608;
wire g8616;
wire g11483;
wire II23586;
wire g15563;
wire g18911;
wire g30351;
wire g18289;
wire g29200;
wire g11761;
wire g12527;
wire II18443;
wire g30569;
wire g33611;
wire g13551;
wire II32963;
wire g12450;
wire II26070;
wire g18155;
wire g34584;
wire g24080;
wire g17180;
wire g12423;
wire g32993;
wire g25136;
wire g18537;
wire g10082;
wire g21740;
wire g23564;
wire g27817;
wire II31497;
wire g14947;
wire II32985;
wire II16795;
wire g34282;
wire g9326;
wire g15137;
wire g14126;
wire g23270;
wire II18758;
wire g29319;
wire g7167;
wire g18180;
wire g23825;
wire g34125;
wire g33906;
wire g32086;
wire g23353;
wire g30208;
wire g20527;
wire g23763;
wire g30383;
wire g23257;
wire g13715;
wire II16695;
wire g25532;
wire g23732;
wire g20708;
wire g21754;
wire g17791;
wire g9567;
wire g31870;
wire g13497;
wire II17783;
wire g18412;
wire g29189;
wire g24148;
wire g24474;
wire g23275;
wire g25168;
wire g34673;
wire II15626;
wire g23481;
wire II26516;
wire g23862;
wire g18938;
wire g18778;
wire g32601;
wire g26573;
wire g22106;
wire II22923;
wire g17570;
wire g24289;
wire g30287;
wire g10587;
wire g28402;
wire II16663;
wire II14579;
wire g29350;
wire g27709;
wire g19458;
wire g34258;
wire g26838;
wire g34138;
wire g19630;
wire g32335;
wire g34744;
wire g24556;
wire g17575;
wire II18635;
wire g16310;
wire g23458;
wire II24400;
wire g12067;
wire g6976;
wire g24385;
wire g19361;
wire g23692;
wire g30990;
wire g12860;
wire g13938;
wire II16709;
wire g25818;
wire g32151;
wire g14753;
wire II33103;
wire II18028;
wire g23391;
wire g10141;
wire g21300;
wire g27025;
wire g19379;
wire g24238;
wire g10652;
wire g33795;
wire g33476;
wire g27038;
wire g33882;
wire g34866;
wire g14295;
wire g28088;
wire g30220;
wire g28976;
wire g16185;
wire g25834;
wire g15570;
wire g26615;
wire II29255;
wire g26901;
wire g15092;
wire II22893;
wire g32697;
wire II27235;
wire g16805;
wire g29883;
wire g31842;
wire g8566;
wire g18269;
wire g31923;
wire g25357;
wire g23509;
wire g24230;
wire g17492;
wire g25159;
wire g14504;
wire g8921;
wire g34339;
wire g6940;
wire g31820;
wire g30167;
wire g32884;
wire g14414;
wire II13139;
wire g34332;
wire g19210;
wire g27674;
wire g34553;
wire g32559;
wire g34601;
wire g30375;
wire II22966;
wire g21274;
wire g21280;
wire II18647;
wire g21880;
wire g15858;
wire II25567;
wire g33544;
wire g25087;
wire g30925;
wire g34445;
wire II14398;
wire g17194;
wire g34195;
wire g20550;
wire g19446;
wire II18614;
wire g9417;
wire g19330;
wire g16638;
wire g12614;
wire g13246;
wire g21299;
wire gbuf44;
wire g7781;
wire g20559;
wire g20603;
wire g18486;
wire II13402;
wire g32870;
wire g14615;
wire g19965;
wire g32197;
wire g25744;
wire g24727;
wire g28655;
wire g11512;
wire g33082;
wire II13066;
wire g20033;
wire II13202;
wire g31846;
wire g24113;
wire II25683;
wire g15824;
wire g24279;
wire g31146;
wire g29789;
wire g29733;
wire g23794;
wire g16696;
wire g25921;
wire g21888;
wire g29984;
wire g10353;
wire g26190;
wire g33076;
wire g30580;
wire g25476;
wire II24191;
wire II12840;
wire g13078;
wire g20674;
wire II12123;
wire g25334;
wire g14589;
wire g20568;
wire II32824;
wire gbuf36;
wire g16473;
wire g26754;
wire g22498;
wire g29490;
wire g22835;
wire g8357;
wire g7854;
wire g12999;
wire g32758;
wire g8139;
wire g22303;
wire g22119;
wire II15954;
wire g14030;
wire g22078;
wire g34794;
wire g12190;
wire g31853;
wire g15507;
wire g17472;
wire gbuf111;
wire II17772;
wire II24619;
wire g27578;
wire g22011;
wire g9755;
wire g20144;
wire g16090;
wire g20734;
wire g34080;
wire g32482;
wire g25006;
wire g18828;
wire g25957;
wire g34067;
wire g29757;
wire g17617;
wire g14365;
wire II13360;
wire g26049;
wire g15713;
wire g25331;
wire g18137;
wire g32326;
wire g14509;
wire g18174;
wire g27201;
wire g19620;
wire g18189;
wire g18669;
wire II16898;
wire g22882;
wire g23063;
wire g23975;
wire g21834;
wire g30005;
wire g30027;
wire g8541;
wire g12644;
wire g20329;
wire g14800;
wire g21655;
wire g23086;
wire g9527;
wire g9509;
wire II30750;
wire II13352;
wire gbuf56;
wire g32389;
wire g25670;
wire g32957;
wire g18113;
wire gbuf9;
wire g17200;
wire g30501;
wire g27714;
wire g13524;
wire g32788;
wire g18231;
wire II18333;
wire g24282;
wire g32390;
wire g31206;
wire g34683;
wire g32827;
wire g16069;
wire g15107;
wire g7778;
wire g31786;
wire g16519;
wire g21686;
wire g25462;
wire g15100;
wire g29836;
wire g23198;
wire g30075;
wire II14823;
wire II25552;
wire g29912;
wire g34047;
wire g9889;
wire g21187;
wire g30409;
wire g24509;
wire g27213;
wire g16235;
wire g24502;
wire II18825;
wire g29006;
wire g28509;
wire g15840;
wire g20670;
wire g15779;
wire g18738;
wire II20412;
wire g33957;
wire g22003;
wire g21845;
wire g33333;
wire II31067;
wire II25594;
wire g30464;
wire g16258;
wire II22580;
wire g13155;
wire g34952;
wire g18151;
wire g9820;
wire g15817;
wire g28544;
wire g28692;
wire g23253;
wire g34461;
wire II15564;
wire g20321;
wire g9933;
wire g18242;
wire g16510;
wire g18091;
wire g24682;
wire g34820;
wire g7212;
wire g13573;
wire g27394;
wire g14700;
wire g25527;
wire g29564;
wire g26310;
wire g10172;
wire g19763;
wire II20187;
wire g30009;
wire g16288;
wire g34571;
wire g12901;
wire g27627;
wire g27560;
wire g34053;
wire g11944;
wire g26515;
wire g33510;
wire g34767;
wire g24217;
wire gbuf77;
wire g31874;
wire g23346;
wire g34611;
wire g21704;
wire g22649;
wire g25174;
wire g11729;
wire g18571;
wire g27381;
wire g25328;
wire g18407;
wire g26881;
wire g16207;
wire g31802;
wire g19996;
wire g9339;
wire g33794;
wire g14193;
wire g10031;
wire g6830;
wire g13854;
wire g13886;
wire g12479;
wire g23767;
wire g10805;
wire g15146;
wire g33462;
wire g9086;
wire g6839;
wire g12336;
wire g26101;
wire g34647;
wire g8821;
wire g24677;
wire g11964;
wire g23428;
wire g34148;
wire g33251;
wire g27511;
wire g18304;
wire g27388;
wire g13494;
wire g23760;
wire g33866;
wire g32140;
wire g7197;
wire g27720;
wire g10869;
wire g12834;
wire g22644;
wire g24397;
wire g27010;
wire g25693;
wire g29684;
wire g26251;
wire g15795;
wire II13252;
wire g27357;
wire II18205;
wire g18662;
wire g7670;
wire g33965;
wire g27250;
wire II24684;
wire g13296;
wire II31122;
wire II18379;
wire g26822;
wire II18894;
wire g29580;
wire g9551;
wire g14816;
wire g34017;
wire II13744;
wire g22852;
wire g28706;
wire g34306;
wire g20579;
wire g34298;
wire g13266;
wire g19475;
wire g32908;
wire g15838;
wire g23874;
wire g11626;
wire g8718;
wire II31838;
wire g24699;
wire g10275;
wire g32233;
wire g28906;
wire g32628;
wire II28147;
wire II17154;
wire II17819;
wire g9310;
wire g18492;
wire g17493;
wire g20101;
wire g11720;
wire g24649;
wire g15345;
wire g10414;
wire g14168;
wire g15060;
wire g33010;
wire g22406;
wire II24482;
wire g15585;
wire g29299;
wire g27584;
wire g9091;
wire g11961;
wire g24121;
wire g12443;
wire II17448;
wire g16821;
wire g27684;
wire g28173;
wire g23815;
wire g15030;
wire g8764;
wire g27581;
wire II24384;
wire g23745;
wire g34170;
wire g18516;
wire g25185;
wire g7566;
wire g19750;
wire II15242;
wire g13131;
wire g31483;
wire g32592;
wire g30432;
wire g8240;
wire II12902;
wire g23666;
wire g32963;
wire II17181;
wire g29265;
wire g19904;
wire II26461;
wire g31185;
wire g26023;
wire g33295;
wire g31117;
wire g32950;
wire g16594;
wire g8449;
wire g17591;
wire II15284;
wire g32160;
wire g33296;
wire g23263;
wire g32894;
wire g10611;
wire g14915;
wire II33235;
wire g25283;
wire g19887;
wire g18935;
wire g32683;
wire g29725;
wire g18128;
wire g14636;
wire II14033;
wire II17695;
wire g14181;
wire g29656;
wire g15737;
wire g18335;
wire II12899;
wire g20993;
wire g33421;
wire II26049;
wire II16486;
wire g18419;
wire g24988;
wire g27880;
wire g12109;
wire g18271;
wire g26486;
wire g17216;
wire g32981;
wire g18740;
wire g34489;
wire g34665;
wire g17503;
wire g31932;
wire g12563;
wire II29279;
wire g24625;
wire II25736;
wire g27085;
wire g18474;
wire g27276;
wire g21811;
wire g32507;
wire g22663;
wire II21722;
wire g28702;
wire g34186;
wire g26924;
wire g24084;
wire g31915;
wire g30046;
wire g6956;
wire g7224;
wire g23357;
wire g23799;
wire g7753;
wire g7835;
wire II20385;
wire g17189;
wire g24105;
wire II12003;
wire g28745;
wire g15853;
wire g21929;
wire g29530;
wire g24035;
wire g23041;
wire g23379;
wire g25970;
wire g21906;
wire g21824;
wire g18544;
wire g34482;
wire g20026;
wire gbuf18;
wire g10307;
wire g22859;
wire II30986;
wire g19350;
wire g24260;
wire g26285;
wire g24295;
wire g12053;
wire g24547;
wire g34470;
wire g14712;
wire g31969;
wire g20563;
wire g27972;
wire g18210;
wire g12411;
wire g22023;
wire g34961;
wire g24399;
wire g20009;
wire g31865;
wire g21950;
wire g25243;
wire g12436;
wire g31894;
wire g19675;
wire g33582;
wire II22502;
wire g32399;
wire II25790;
wire g18121;
wire g26969;
wire g22009;
wire g13620;
wire g20593;
wire g27091;
wire g22976;
wire g14608;
wire g18978;
wire g32205;
wire g19679;
wire g24333;
wire g31138;
wire g24220;
wire II12782;
wire g25951;
wire g15372;
wire g25142;
wire g24054;
wire g13584;
wire g25182;
wire g9234;
wire g31812;
wire II32659;
wire II23694;
wire g16746;
wire g18114;
wire g21287;
wire g10347;
wire g8790;
wire g15745;
wire g34844;
wire g11852;
wire g23020;
wire g23208;
wire II32452;
wire g19532;
wire g16281;
wire g31974;
wire g11996;
wire g23921;
wire g25979;
wire g22032;
wire II18626;
wire g21338;
wire g13474;
wire g17062;
wire g23372;
wire g18276;
wire II31331;
wire g16221;
wire g13897;
wire g7327;
wire g28159;
wire g34403;
wire g9649;
wire II20216;
wire g31282;
wire g20135;
wire II33158;
wire g34320;
wire g18328;
wire g18550;
wire g15166;
wire g28599;
wire II33053;
wire g29380;
wire II14277;
wire II13166;
wire g34761;
wire gbuf110;
wire g21347;
wire g28049;
wire g25784;
wire II20750;
wire g20233;
wire g12187;
wire g33978;
wire g32563;
wire g29653;
wire g32273;
wire g27662;
wire g32170;
wire g7520;
wire g24945;
wire g26802;
wire g12301;
wire g9546;
wire g27043;
wire II33064;
wire II32770;
wire g24195;
wire g19431;
wire g18569;
wire g33915;
wire g28774;
wire g24439;
wire g16197;
wire II15843;
wire g18127;
wire g11708;
wire g21947;
wire g11955;
wire g25559;
wire g24974;
wire g33869;
wire g28534;
wire g23312;
wire g22900;
wire g25084;
wire g21404;
wire g22152;
wire g17500;
wire g11972;
wire g17485;
wire g32475;
wire g20235;
wire g30227;
wire g18532;
wire g12539;
wire g30301;
wire g24914;
wire g19603;
wire II16590;
wire II31082;
wire II21254;
wire g30494;
wire g34185;
wire g12044;
wire g10124;
wire II12253;
wire g33593;
wire g32105;
wire g34523;
wire g32923;
wire g20052;
wire g20536;
wire g21509;
wire g16602;
wire g25645;
wire g27309;
wire g34686;
wire g18386;
wire g11038;
wire II27677;
wire II18852;
wire g18787;
wire g24387;
wire g33129;
wire g32346;
wire g23523;
wire g29176;
wire g29642;
wire g9299;
wire g24306;
wire II26366;
wire g29354;
wire g32691;
wire g34364;
wire g23626;
wire g26231;
wire g12735;
wire II13336;
wire g17782;
wire g32048;
wire g17510;
wire g34642;
wire g7235;
wire g24138;
wire II15981;
wire II16564;
wire g24762;
wire g28620;
wire g27208;
wire g15870;
wire g24073;
wire g19502;
wire g34827;
wire g28090;
wire g15710;
wire g7640;
wire g23955;
wire II28572;
wire g8124;
wire g27858;
wire g30547;
wire g33362;
wire g29964;
wire II12730;
wire g32806;
wire g18583;
wire g34809;
wire g25610;
wire g30348;
wire g32329;
wire g12180;
wire II31983;
wire g33706;
wire g32212;
wire II32973;
wire g27538;
wire g30385;
wire g27247;
wire g20218;
wire g29184;
wire g32909;
wire g14157;
wire g18641;
wire g24379;
wire g26934;
wire II12470;
wire g28953;
wire g29539;
wire g13051;
wire g28435;
wire g27489;
wire g27326;
wire g25563;
wire g8107;
wire g9777;
wire g13304;
wire g23870;
wire g34638;
wire gbuf53;
wire g28270;
wire g33787;
wire g12113;
wire g20270;
wire g7170;
wire g23400;
wire g8903;
wire g24566;
wire g28528;
wire g21955;
wire g24320;
wire g14397;
wire g25878;
wire g23571;
wire g18390;
wire g22513;
wire g32033;
wire g29152;
wire II19661;
wire II31237;
wire g29847;
wire II12030;
wire g27963;
wire g9000;
wire g27304;
wire g26977;
wire g15050;
wire g27267;
wire g33721;
wire g34029;
wire g9012;
wire g10502;
wire g32859;
wire g26177;
wire g21858;
wire g34632;
wire g25040;
wire g16882;
wire g26949;
wire g25201;
wire g9904;
wire g31773;
wire g16845;
wire g14150;
wire g33805;
wire g7577;
wire g23407;
wire g20572;
wire II31266;
wire g17321;
wire g26650;
wire II29248;
wire g28660;
wire g12875;
wire g21973;
wire g18690;
wire g11017;
wire g23019;
wire g18908;
wire g9833;
wire g11930;
wire II32687;
wire II14450;
wire g26861;
wire g33369;
wire g13030;
wire g17691;
wire II13280;
wire g20090;
wire II18469;
wire g18804;
wire g27280;
wire II17879;
wire g20064;
wire g12244;
wire g20076;
wire g30393;
wire g21666;
wire g32308;
wire g27931;
wire g7410;
wire g29735;
wire g18251;
wire II13857;
wire g34167;
wire g25021;
wire g10738;
wire g33497;
wire g19570;
wire II32681;
wire g34587;
wire g9037;
wire g18709;
wire g29865;
wire g25309;
wire g30236;
wire g24965;
wire g28910;
wire g33834;
wire gbuf143;
wire g30033;
wire g26666;
wire II17404;
wire g32407;
wire g32243;
wire II12837;
wire g20664;
wire g26709;
wire g21326;
wire g31909;
wire g8509;
wire g29927;
wire g28193;
wire g28627;
wire g12073;
wire g20530;
wire g34454;
wire g13009;
wire g22312;
wire g29193;
wire g16655;
wire g32087;
wire g31886;
wire g8644;
wire g26048;
wire g17707;
wire g30485;
wire g23056;
wire II15872;
wire g28714;
wire g7553;
wire g24496;
wire II25530;
wire II31017;
wire g10755;
wire g16027;
wire g17811;
wire g22089;
wire g25049;
wire II32884;
wire g7175;
wire g12588;
wire g18360;
wire g31474;
wire g7834;
wire g34369;
wire g22039;
wire g34031;
wire g15113;
wire g25195;
wire g21419;
wire g14687;
wire g12700;
wire g17489;
wire g11819;
wire II21067;
wire II17916;
wire g34273;
wire g25562;
wire g34739;
wire g34321;
wire g20111;
wire II16231;
wire II23985;
wire g23449;
wire g22493;
wire g10155;
wire g29705;
wire g12872;
wire g16739;
wire g18438;
wire g26276;
wire g32992;
wire g18429;
wire g29858;
wire g29864;
wire g25308;
wire g33550;
wire g21365;
wire g32634;
wire g21982;
wire g21221;
wire g15045;
wire g28213;
wire g25356;
wire g19469;
wire g27711;
wire g33399;
wire g22658;
wire g20655;
wire g7396;
wire g25267;
wire g32287;
wire g20391;
wire g31000;
wire g23651;
wire g15746;
wire g23121;
wire II18897;
wire g30254;
wire g18579;
wire g30190;
wire g21989;
wire g15796;
wire g21909;
wire g28969;
wire g7963;
wire g9946;
wire g14332;
wire g30732;
wire g22308;
wire II28883;
wire g12546;
wire II16688;
wire g19333;
wire g21190;
wire g25518;
wire g25068;
wire II13552;
wire II18900;
wire g13541;
wire g11615;
wire g34289;
wire g32753;
wire g7511;
wire g31927;
wire g22118;
wire II19813;
wire g17784;
wire II18587;
wire g16600;
wire II17763;
wire g25911;
wire g21460;
wire g16586;
wire g15277;
wire g8431;
wire g21384;
wire g17870;
wire g25054;
wire g32542;
wire g16607;
wire g15709;
wire g34781;
wire g23639;
wire g29777;
wire II31829;
wire II23300;
wire g7647;
wire g29772;
wire II12497;
wire g33641;
wire g34604;
wire g21055;
wire g30250;
wire g24849;
wire g12711;
wire g23128;
wire g12013;
wire g22044;
wire g31776;
wire g27926;
wire g30128;
wire II22794;
wire g17391;
wire g10224;
wire g11744;
wire II24089;
wire g9875;
wire g13250;
wire g27453;
wire g18764;
wire g13345;
wire g12288;
wire II23979;
wire g23855;
wire g20211;
wire g28717;
wire g34000;
wire g15066;
wire g28497;
wire g24366;
wire g29995;
wire g25679;
wire g19777;
wire g31490;
wire g32301;
wire g32529;
wire g29079;
wire II26925;
wire II18092;
wire g9332;
wire g23293;
wire g34806;
wire g29013;
wire g17587;
wire g19873;
wire g28688;
wire g33786;
wire g34251;
wire g11193;
wire gbuf109;
wire II23333;
wire g29713;
wire II32079;
wire II12346;
wire g28238;
wire g12234;
wire II20166;
wire g26098;
wire g7518;
wire g28139;
wire g19862;
wire II20910;
wire g29149;
wire g14306;
wire g17178;
wire g25885;
wire g24042;
wire g11544;
wire g7885;
wire g31002;
wire g10598;
wire g28813;
wire g30553;
wire g21381;
wire g23755;
wire g34592;
wire g33920;
wire g30278;
wire g7142;
wire g30914;
wire g9007;
wire g19504;
wire II13334;
wire g32708;
wire g10385;
wire g27438;
wire g31960;
wire g29806;
wire g18298;
wire g25663;
wire g30404;
wire g20626;
wire g27404;
wire g17777;
wire g17424;
wire g34265;
wire g19717;
wire g22679;
wire g10961;
wire g18466;
wire g28089;
wire g30449;
wire g16971;
wire g29944;
wire g25628;
wire g11170;
wire g16620;
wire II22889;
wire g28796;
wire g31267;
wire g12343;
wire g28231;
wire g17653;
wire gbuf102;
wire g30435;
wire g18374;
wire g13023;
wire II28597;
wire g23618;
wire g32714;
wire g14452;
wire g8836;
wire g10604;
wire g9740;
wire g16180;
wire II29286;
wire II18034;
wire II31182;
wire g13485;
wire g24618;
wire g32113;
wire g27346;
wire II13519;
wire g11020;
wire g24277;
wire g26784;
wire g25260;
wire g13504;
wire gbuf138;
wire g33577;
wire g16126;
wire g18215;
wire g18353;
wire g13321;
wire g16768;
wire g32090;
wire g18450;
wire g19525;
wire g9379;
wire g25871;
wire g14218;
wire g28698;
wire g22842;
wire g28304;
wire g22626;
wire g22545;
wire g7345;
wire II20982;
wire g33622;
wire g30122;
wire g21837;
wire II17101;
wire g11261;
wire g29256;
wire g24157;
wire g29198;
wire g23914;
wire g9030;
wire g22861;
wire g21857;
wire II11843;
wire g7472;
wire II31341;
wire g8224;
wire II31141;
wire g29333;
wire g24177;
wire g11135;
wire g11639;
wire g10370;
wire g11917;
wire g28341;
wire g32820;
wire g14962;
wire g33975;
wire g24717;
wire g13119;
wire g34315;
wire g12716;
wire II22422;
wire g25063;
wire II32059;
wire g9414;
wire II16755;
wire II13708;
wire g32747;
wire g25504;
wire II17883;
wire g31325;
wire g28980;
wire g30578;
wire g13603;
wire g24628;
wire II22816;
wire g24702;
wire g18795;
wire g34393;
wire g32053;
wire g34653;
wire g19549;
wire g28635;
wire g31807;
wire g32350;
wire g16578;
wire g32929;
wire g17522;
wire g30261;
wire g22145;
wire g29481;
wire g20503;
wire g30426;
wire gbuf68;
wire g22028;
wire g25718;
wire g12897;
wire g23533;
wire g25701;
wire II18486;
wire g28245;
wire g32966;
wire g26518;
wire g33345;
wire g19538;
wire g21350;
wire g23962;
wire g24324;
wire II32432;
wire g14833;
wire II23387;
wire II24128;
wire g22052;
wire g23023;
wire g24571;
wire g28895;
wire g22709;
wire g18754;
wire g14626;
wire g30523;
wire g14438;
wire g25014;
wire g16160;
wire g30088;
wire g9154;
wire g14683;
wire gbuf135;
wire g18200;
wire g34430;
wire g18895;
wire g12892;
wire II31181;
wire g30340;
wire g12082;
wire g33317;
wire g34407;
wire g20095;
wire g27960;
wire g14505;
wire g11184;
wire II29295;
wire g9679;
wire II30904;
wire g8872;
wire g15754;
wire g11396;
wire g13081;
wire II14708;
wire g11128;
wire g19355;
wire g33733;
wire II18083;
wire g25248;
wire g17645;
wire II16492;
wire g29922;
wire g25606;
wire g29987;
wire g31943;
wire II17692;
wire g9556;
wire g10391;
wire g27275;
wire II16917;
wire g33292;
wire g26422;
wire g6869;
wire g15062;
wire g18689;
wire g26088;
wire g32874;
wire g30053;
wire g14786;
wire g13319;
wire g27362;
wire II27549;
wire II14248;
wire g32530;
wire II26417;
wire g24292;
wire g26223;
wire g9492;
wire g17496;
wire g24992;
wire g24771;
wire g31780;
wire g33562;
wire g29229;
wire g9892;
wire II13043;
wire g26744;
wire g18684;
wire g15083;
wire II24030;
wire g16520;
wire g22986;
wire g32375;
wire g27352;
wire II32240;
wire g33186;
wire g22920;
wire g13830;
wire g33018;
wire g31116;
wire g15806;
wire g34485;
wire g34385;
wire g25767;
wire g15151;
wire g19953;
wire g27311;
wire g24026;
wire g19739;
wire g28333;
wire g33111;
wire g31899;
wire g30564;
wire g17147;
wire II33044;
wire g31655;
wire g25899;
wire g31744;
wire g21464;
wire g17367;
wire g12149;
wire g20275;
wire g19366;
wire g13265;
wire g29976;
wire g15163;
wire g27678;
wire g29623;
wire g23542;
wire g26680;
wire g34620;
wire g14315;
wire g32905;
wire g31787;
wire g28575;
wire g34228;
wire g31318;
wire g17594;
wire g18207;
wire g18383;
wire g23961;
wire g20202;
wire g10584;
wire g32513;
wire g19618;
wire g7451;
wire g21184;
wire g13872;
wire II32550;
wire g13056;
wire g32494;
wire II23393;
wire g28463;
wire g23472;
wire II11626;
wire g25058;
wire g8607;
wire g26894;
wire g26328;
wire II22009;
wire g29745;
wire g23506;
wire g28851;
wire g9523;
wire g18888;
wire g32519;
wire g18932;
wire g22102;
wire g23549;
wire g30136;
wire g27975;
wire g19738;
wire II13383;
wire g28616;
wire g11448;
wire g20914;
wire g16537;
wire g15654;
wire g18343;
wire g21722;
wire g28646;
wire g13764;
wire g19411;
wire g18106;
wire g13910;
wire g32571;
wire II15241;
wire g19913;
wire g33551;
wire g27998;
wire g23898;
wire II27758;
wire g26966;
wire g12027;
wire g33053;
wire II14623;
wire g29383;
wire g23494;
wire g27008;
wire g23775;
wire g16534;
wire g23256;
wire g21818;
wire g31554;
wire g23227;
wire g19367;
wire g8592;
wire g12399;
wire g30451;
wire g25936;
wire II22211;
wire g33142;
wire g24637;
wire g34040;
wire g15095;
wire g29796;
wire g22127;
wire g8438;
wire g9804;
wire g23220;
wire g31755;
wire g17243;
wire g21908;
wire g11204;
wire g23968;
wire g34848;
wire g23320;
wire g28468;
wire II14498;
wire gbuf127;
wire g32549;
wire g23154;
wire g29904;
wire g11562;
wire g31299;
wire g12844;
wire g19429;
wire g19264;
wire g30210;
wire g19713;
wire g12201;
wire g27378;
wire g30673;
wire g24424;
wire g29676;
wire g34134;
wire g33865;
wire g16606;
wire g14829;
wire g9616;
wire II15620;
wire II15123;
wire II33252;
wire g31578;
wire g32775;
wire g34502;
wire g32016;
wire g24210;
wire g20645;
wire II22458;
wire g10565;
wire g27112;
wire g18431;
wire g9166;
wire g34685;
wire g13282;
wire g24038;
wire g32734;
wire II12950;
wire II26395;
wire g10191;
wire g18734;
wire g28126;
wire g14889;
wire g31292;
wire g34740;
wire II31011;
wire II14765;
wire g21964;
wire g26195;
wire g32897;
wire g28514;
wire g30049;
wire g34625;
wire g9044;
wire g34498;
wire g6972;
wire II13141;
wire g33985;
wire gbuf152;
wire g20512;
wire II26334;
wire g25171;
wire g21827;
wire g13037;
wire g21774;
wire g29121;
wire g21873;
wire II32284;
wire g13633;
wire g14864;
wire g22622;
wire g18309;
wire g16630;
wire g15885;
wire g9499;
wire g21036;
wire g23166;
wire g34422;
wire II27381;
wire g18628;
wire g30462;
wire g24244;
wire g21677;
wire g26126;
wire gbuf146;
wire g6840;
wire g32502;
wire g11189;
wire g18319;
wire g32938;
wire g32161;
wire g26942;
wire g25547;
wire g34117;
wire g29852;
wire g28225;
wire g16529;
wire g33062;
wire g33378;
wire g30196;
wire g14512;
wire g12482;
wire g12823;
wire g33791;
wire g25680;
wire g8407;
wire g11663;
wire g11201;
wire II31823;
wire g28728;
wire g34329;
wire II12519;
wire II25391;
wire g32862;
wire II17754;
wire g31021;
wire g30934;
wire g26831;
wire g34427;
wire g33442;
wire g24481;
wire g31522;
wire g9704;
wire g28861;
wire g20448;
wire g32412;
wire g15844;
wire g8056;
wire g17401;
wire g32673;
wire g7565;
wire g20887;
wire g16641;
wire g24528;
wire g31514;
wire g18525;
wire g24755;
wire g17514;
wire g25178;
wire g11986;
wire g32262;
wire g16249;
wire g27227;
wire II14589;
wire g17624;
wire g33252;
wire g26159;
wire g11590;
wire g28945;
wire g16489;
wire g24140;
wire g25371;
wire g16928;
wire g24010;
wire g29766;
wire g29980;
wire g31067;
wire g18510;
wire g24940;
wire II20913;
wire g31836;
wire g28315;
wire g12297;
wire g32041;
wire g16428;
wire g20152;
wire g30117;
wire II14006;
wire g11245;
wire II12277;
wire g20713;
wire g13221;
wire g33962;
wire g33645;
wire g7992;
wire g16244;
wire g32717;
wire g21303;
wire II17801;
wire gbuf34;
wire g27462;
wire g24821;
wire g25696;
wire g18285;
wire g28326;
wire g26871;
wire g34741;
wire II31217;
wire g29488;
wire g16474;
wire g6991;
wire g7863;
wire g24285;
wire g32727;
wire g10603;
wire g23066;
wire g33475;
wire II27573;
wire g18505;
wire g8685;
wire II25220;
wire g29743;
wire II12098;
wire g15726;
wire g28262;
wire g16590;
wire g27034;
wire g16685;
wire II26741;
wire g28426;
wire g21800;
wire g9541;
wire g14090;
wire g29378;
wire g28731;
wire g33457;
wire g22126;
wire g9908;
wire g6895;
wire g23167;
wire g33388;
wire g21024;
wire g30595;
wire g25830;
wire g21204;
wire g25064;
wire g9931;
wire g28590;
wire g34955;
wire g25763;
wire g33459;
wire g25687;
wire g11948;
wire g24312;
wire g33312;
wire II18537;
wire g9664;
wire g18718;
wire II13109;
wire g31124;
wire g24017;
wire gbuf120;
wire g7356;
wire g19067;
wire g25325;
wire g18481;
wire g9692;
wire g10113;
wire g20170;
wire g32171;
wire g15076;
wire g18728;
wire g19692;
wire g8201;
wire g15508;
wire g10205;
wire g28035;
wire g22137;
wire g21253;
wire g22634;
wire g29517;
wire g9732;
wire II16724;
wire II15697;
wire II13566;
wire g31845;
wire g10621;
wire g19445;
wire II16143;
wire g12088;
wire g32568;
wire g18445;
wire g31936;
wire g34991;
wire g10489;
wire g32976;
wire g34200;
wire II18449;
wire g32127;
wire g24506;
wire g31018;
wire g31911;
wire g9760;
wire g34968;
wire g9860;
wire g24164;
wire II14275;
wire g33118;
wire g26750;
wire g28072;
wire g15128;
wire II22267;
wire g10555;
wire g24145;
wire g27142;
wire II15102;
wire g16873;
wire II11708;
wire g18951;
wire g18984;
wire g12793;
wire g25987;
wire g13512;
wire g10368;
wire g27528;
wire II14660;
wire g29853;
wire g24553;
wire g16322;
wire g25876;
wire g15002;
wire g25102;
wire g10109;
wire g12953;
wire g11042;
wire g28414;
wire II17136;
wire g26380;
wire g18364;
wire g21744;
wire g17605;
wire g19416;
wire g32381;
wire g30282;
wire g26297;
wire g24922;
wire g18657;
wire g31508;
wire gbuf85;
wire g22870;
wire g31790;
wire g30292;
wire g30189;
wire g27339;
wire g12639;
wire g22111;
wire g13012;
wire II27970;
wire g17497;
wire g23926;
wire g21910;
wire g29169;
wire g10337;
wire g28991;
wire II17108;
wire g18770;
wire II16090;
wire g25887;
wire g34078;
wire g15936;
wire g23513;
wire g27232;
wire g24252;
wire g33873;
wire g15628;
wire g7499;
wire II18835;
wire II24215;
wire g24532;
wire g25424;
wire g29668;
wire g14691;
wire g25429;
wire II33170;
wire g33998;
wire g28570;
wire II21246;
wire g24658;
wire g14731;
wire g15875;
wire g12571;
wire g14541;
wire g18564;
wire g22993;
wire g20166;
wire g27981;
wire II19778;
wire g33615;
wire II24709;
wire g24048;
wire g20114;
wire gbuf61;
wire g13096;
wire g22838;
wire g25941;
wire g21864;
wire g24159;
wire g19741;
wire II13453;
wire g19461;
wire g11142;
wire g17873;
wire g32969;
wire g31130;
wire g24576;
wire g18295;
wire g28689;
wire g26813;
wire II16160;
wire II23978;
wire g32137;
wire g28205;
wire g21155;
wire II33137;
wire g33971;
wire g32393;
wire g24798;
wire II16618;
wire II20861;
wire g28750;
wire g27332;
wire g31477;
wire g25774;
wire g20667;
wire g7627;
wire g21763;
wire g14078;
wire II13699;
wire II16780;
wire g22082;
wire g18214;
wire g14424;
wire g23416;
wire g26987;
wire g21608;
wire II23162;
wire g14517;
wire g16705;
wire II31854;
wire g25620;
wire II17529;
wire g12523;
wire g17183;
wire g18300;
wire g7183;
wire II31972;
wire II25115;
wire gbuf147;
wire g10041;
wire g34656;
wire g18473;
wire II19734;
wire g30531;
wire g14450;
wire g21917;
wire g28429;
wire g13666;
wire g23971;
wire g33598;
wire g20109;
wire g24624;
wire g11367;
wire g13412;
wire g30203;
wire gbuf134;
wire g21999;
wire g17686;
wire g15569;
wire g31470;
wire g32953;
wire g29643;
wire gbuf25;
wire g25210;
wire g30482;
wire g23395;
wire g34156;
wire g30142;
wire g27616;
wire g34465;
wire g28375;
wire g32011;
wire g32082;
wire g17264;
wire g7335;
wire g30401;
wire g34254;
wire g33095;
wire II14481;
wire g33303;
wire g7231;
wire g33418;
wire g17574;
wire g32331;
wire g13222;
wire g32586;
wire g10529;
wire g20737;
wire g14208;
wire II31291;
wire g31920;
wire g20704;
wire II20221;
wire g8330;
wire g25722;
wire g33926;
wire g29578;
wire g6801;
wire g26776;
wire II13444;
wire g24606;
wire g32605;
wire g12361;
wire g33886;
wire g23948;
wire II26512;
wire g23271;
wire g29615;
wire g25948;
wire II21918;
wire g23130;
wire g20769;
wire g24746;
wire g12850;
wire II29352;
wire g18817;
wire g23412;
wire g16957;
wire g34159;
wire II14054;
wire g29204;
wire g23162;
wire g30065;
wire II31197;
wire g33612;
wire g9639;
wire g33034;
wire g10213;
wire g20449;
wire g9187;
wire g32998;
wire g22047;
wire g23787;
wire II17787;
wire II12563;
wire g29248;
wire g8113;
wire g32098;
wire g23568;
wire g22099;
wire g26203;
wire II14684;
wire g11755;
wire II32170;
wire g34776;
wire g34722;
wire g19376;
wire g7548;
wire II32106;
wire g16761;
wire II24558;
wire g19659;
wire II18376;
wire g28674;
wire g22755;
wire g16826;
wire g9340;
wire g15078;
wire g19655;
wire g19454;
wire II24463;
wire g9501;
wire g25572;
wire g9443;
wire g20900;
wire g25536;
wire II15253;
wire g17736;
wire g29838;
wire g10656;
wire II18160;
wire g27828;
wire g22997;
wire g29901;
wire g32526;
wire g25094;
wire g9974;
wire g18440;
wire g27393;
wire g31616;
wire g11292;
wire g7666;
wire g12835;
wire g13027;
wire g17581;
wire g18676;
wire g31211;
wire g25791;
wire g9689;
wire g31608;
wire II26448;
wire g17744;
wire g28149;
wire g28136;
wire g24358;
wire g29277;
wire g16734;
wire g12730;
wire g32841;
wire II12333;
wire g13350;
wire g13902;
wire g30441;
wire g18265;
wire g30133;
wire g21284;
wire g7393;
wire II23600;
wire II19345;
wire g14095;
wire g23885;
wire g8519;
wire g19629;
wire g11812;
wire g30224;
wire g34027;
wire g29634;
wire g28889;
wire g11412;
wire II18868;
wire g24343;
wire g19740;
wire g29665;
wire g27617;
wire g29614;
wire g20524;
wire g8387;
wire g22717;
wire g8002;
wire g21610;
wire g33819;
wire g28711;
wire g28659;
wire g18612;
wire II18523;
wire II30755;
wire g27428;
wire II29315;
wire g18397;
wire II11685;
wire g14539;
wire g30824;
wire g14085;
wire g12581;
wire g33134;
wire g30106;
wire g34380;
wire g18404;
wire II15736;
wire II31136;
wire g30388;
wire g27073;
wire g25118;
wire g28165;
wire II11665;
wire g29572;
wire g18502;
wire g34290;
wire II20469;
wire g26858;
wire g16815;
wire g25805;
wire g33279;
wire g28033;
wire g34539;
wire II12033;
wire g29178;
wire II15921;
wire g31825;
wire g25658;
wire g27334;
wire g22067;
wire g12838;
wire g22318;
wire II32476;
wire g7437;
wire II18795;
wire II14742;
wire g10706;
wire g22518;
wire g32253;
wire II24699;
wire g31152;
wire II20882;
wire g33481;
wire g33870;
wire g9724;
wire g26713;
wire II14530;
wire g15018;
wire II15834;
wire g28973;
wire g28066;
wire g26703;
wire g23560;
wire g21749;
wire g15143;
wire g14121;
wire g33498;
wire g31251;
wire g23988;
wire g17271;
wire g30094;
wire g33679;
wire g33589;
wire g34890;
wire g21796;
wire g8183;
wire g8504;
wire g16268;
wire g25250;
wire g23559;
wire g18632;
wire II32874;
wire g8088;
wire g28779;
wire II30727;
wire g27292;
wire g30471;
wire g10491;
wire g25083;
wire g24745;
wire g9281;
wire g33670;
wire g23430;
wire g32246;
wire g11533;
wire g28440;
wire g34493;
wire g20543;
wire g17636;
wire g30325;
wire g19609;
wire g19762;
wire g34278;
wire g34225;
wire g33107;
wire II16010;
wire g30023;
wire g14154;
wire g7764;
wire g7247;
wire g23479;
wire g24430;
wire g32478;
wire g31256;
wire g22341;
wire g32316;
wire g22489;
wire g11027;
wire g19634;
wire II27538;
wire g24181;
wire g25728;
wire g18743;
wire g30097;
wire II29242;
wire g17700;
wire g31304;
wire g11139;
wire g20186;
wire g27732;
wire g18990;
wire g32146;
wire g31769;
wire II12401;
wire g32917;
wire g19908;
wire g31709;
wire g31225;
wire g22224;
wire g30270;
wire g21250;
wire g21451;
wire g28675;
wire g21557;
wire g18892;
wire g21978;
wire g17119;
wire g23998;
wire g32928;
wire II21959;
wire g21934;
wire g12154;
wire g22981;
wire g27432;
wire g24720;
wire g13019;
wire g27459;
wire g14873;
wire g22906;
wire g23235;
wire g26732;
wire II18003;
wire g26636;
wire II31494;
wire g23997;
wire g21799;
wire g23515;
wire g7117;
wire g25619;
wire g10077;
wire II22799;
wire g18691;
wire g31959;
wire g34150;
wire g19558;
wire g8880;
wire g15702;
wire g20611;
wire g21792;
wire g26362;
wire g25122;
wire g10407;
wire g32192;
wire g24373;
wire II17395;
wire g29116;
wire g16214;
wire g24854;
wire g13333;
wire g14855;
wire g15862;
wire g29679;
wire g11236;
wire g28101;
wire g24941;
wire g7876;
wire g12307;
wire g16613;
wire g12048;
wire g24063;
wire II13726;
wire g24663;
wire g24711;
wire g34061;
wire g31313;
wire g21952;
wire g29241;
wire g29345;
wire II25750;
wire g32948;
wire g33236;
wire g25893;
wire II24530;
wire g30155;
wire g23055;
wire g11444;
wire g25554;
wire g32419;
wire g23657;
wire II21815;
wire g32626;
wire g19436;
wire g34906;
wire g34540;
wire g32270;
wire g25220;
wire g13070;
wire g33576;
wire g14261;
wire g34549;
wire g28180;
wire g23005;
wire g34532;
wire g27736;
wire g14772;
wire g27956;
wire g18673;
wire g24569;
wire g20071;
wire g14255;
wire g20838;
wire g8879;
wire g12888;
wire g33416;
wire g18195;
wire g13941;
wire g12659;
wire g26616;
wire g20632;
wire II31177;
wire g30035;
wire g25286;
wire g9912;
wire g27134;
wire g30511;
wire II27519;
wire II22512;
wire g16840;
wire g25651;
wire g25754;
wire g28582;
wire II12799;
wire g29553;
wire g25865;
wire g26953;
wire g16201;
wire g32652;
wire g34784;
wire g28058;
wire g25634;
wire g10218;
wire g32110;
wire g23317;
wire g27568;
wire g30555;
wire g31308;
wire g23079;
wire g34790;
wire g21926;
wire g33351;
wire g22941;
wire g32067;
wire g33919;
wire g9898;
wire II22880;
wire g14051;
wire g30178;
wire g8744;
wire g31262;
wire g31978;
wire g32144;
wire g29916;
wire g33432;
wire g8840;
wire g13870;
wire g12332;
wire g25646;
wire g17612;
wire g22338;
wire g33991;
wire g23905;
wire g34344;
wire II24680;
wire g11894;
wire g30306;
wire g24634;
wire g18589;
wire g23501;
wire g27724;
wire g12768;
wire g32643;
wire II31650;
wire g27876;
wire II32607;
wire g11868;
wire g15117;
wire g29209;
wire II31327;
wire g11779;
wire g16709;
wire II17471;
wire g20922;
wire g24968;
wire g27011;
wire II33164;
wire II17699;
wire g26513;
wire II21181;
wire g13173;
wire g14572;
wire g18666;
wire g11771;
wire g30735;
wire g27327;
wire g26272;
wire II13321;
wire g17733;
wire g16136;
wire g34110;
wire g8822;
wire II32202;
wire g33045;
wire g11394;
wire g29799;
wire g25566;
wire g28229;
wire g26799;
wire II31779;
wire g23662;
wire g25540;
wire g21711;
wire g26180;
wire g28456;
wire g18701;
wire g28647;
wire g32524;
wire g31833;
wire g32083;
wire g29534;
wire g9600;
wire g27216;
wire g15069;
wire g7749;
wire g14911;
wire II15078;
wire II22601;
wire g17389;
wire II23330;
wire g10615;
wire g33953;
wire g30355;
wire g11432;
wire g9071;
wire g25801;
wire g13637;
wire g27042;
wire g20266;
wire g12416;
wire g23811;
wire g27146;
wire g23647;
wire g23839;
wire g28083;
wire II25847;
wire g10551;
wire g26289;
wire g25039;
wire g29549;
wire g28155;
wire g11724;
wire g8146;
wire II18270;
wire g16776;
wire g26341;
wire g35001;
wire g27358;
wire g13279;
wire g26956;
wire g22522;
wire g20435;
wire g6782;
wire g14822;
wire II26654;
wire g19916;
wire g29593;
wire g12159;
wire g23202;
wire g29896;
wire g29366;
wire g18437;
wire g13043;
wire g18124;
wire g34823;
wire g32720;
wire g25465;
wire g24129;
wire g29272;
wire II17381;
wire g27585;
wire g24453;
wire g23425;
wire g32242;
wire g12418;
wire g30260;
wire II18364;
wire g33521;
wire II17842;
wire g18144;
wire g16728;
wire g33212;
wire II31086;
wire g21699;
wire g18878;
wire g8179;
wire g13105;
wire g16732;
wire g30312;
wire g10719;
wire g33933;
wire g14449;
wire g23881;
wire g11024;
wire g11547;
wire g16954;
wire g13679;
wire II18680;
wire g24126;
wire g34708;
wire g24464;
wire g28387;
wire g7689;
wire gbuf98;
wire g7831;
wire g20105;
wire g12050;
wire g30000;
wire g24701;
wire g16205;
wire II31863;
wire g11897;
wire g19531;
wire g20701;
wire g31965;
wire g18943;
wire g21461;
wire g16853;
wire g27287;
wire II30998;
wire g19536;
wire g30015;
wire g8847;
wire g23936;
wire g24301;
wire g33547;
wire II13518;
wire g27410;
wire g21604;
wire g22109;
wire II12000;
wire II12360;
wire g24101;
wire gbuf14;
wire g26921;
wire g10083;
wire g32701;
wire g25438;
wire g23262;
wire g8993;
wire g29722;
wire g33554;
wire g25492;
wire g21048;
wire g34946;
wire g29694;
wire II28872;
wire g29375;
wire II25908;
wire II28585;
wire g10419;
wire II33056;
wire g33911;
wire g18275;
wire g11841;
wire g28345;
wire g8632;
wire g16210;
wire g11166;
wire g23925;
wire g23204;
wire g7704;
wire g26911;
wire g8715;
wire II18138;
wire g20383;
wire II25695;
wire g19611;
wire g14197;
wire g24685;
wire g24793;
wire g8259;
wire g12761;
wire g25521;
wire g18882;
wire g22432;
wire g25601;
wire g22938;
wire g12150;
wire g13624;
wire g15992;
wire g18750;
wire g23332;
wire g33568;
wire g18425;
wire g22846;
wire g28758;
wire g30612;
wire g12969;
wire g29094;
wire g10074;
wire g32201;
wire g19478;
wire g8080;
wire g24020;
wire g25772;
wire g13831;
wire g19754;
wire g18324;
wire g19882;
wire g21378;
wire g23209;
wire g34578;
wire g15573;
wire g33515;
wire g10819;
wire g16742;
wire g19671;
wire g16285;
wire g14656;
wire II18031;
wire g9484;
wire g25666;
wire g29584;
wire g27149;
wire g32237;
wire g27163;
wire II22725;
wire g24050;
wire g24235;
wire g13015;
wire g27371;
wire II18728;
wire g25501;
wire II20690;
wire g24213;
wire g30561;
wire g14584;
wire g28724;
wire g8217;
wire g11968;
wire g9051;
wire II16646;
wire g24723;
wire g32193;
wire g24774;
wire g24336;
wire g18560;
wire g29358;
wire g28061;
wire g30148;
wire g33372;
wire g22169;
wire g13569;
wire g20633;
wire g32421;
wire g13141;
wire g18765;
wire g18461;
wire g7623;
wire g34569;
wire II16803;
wire g25868;
wire g15613;
wire g24109;
wire g20596;
wire II23312;
wire g27592;
wire g24076;
wire g28252;
wire g30217;
wire g27553;
wire g24621;
wire g27534;
wire g23082;
wire g20607;
wire g18587;
wire g24514;
wire g23187;
wire g34336;
wire g30163;
wire g23342;
wire g29786;
wire II14630;
wire g12487;
wire II15316;
wire g34095;
wire g28561;
wire g22831;
wire g26885;
wire g13808;
wire II29363;
wire g21660;
wire g19071;
wire g17599;
wire g24817;
wire g34084;
wire g34473;
wire g32836;
wire g13130;
wire g27824;
wire g29877;
wire g19999;
wire g29589;
wire g28094;
wire g10358;
wire g31631;
wire g10476;
wire g34441;
wire g18989;
wire g30070;
wire g20612;
wire g34637;
wire g10804;
wire g18606;
wire g17308;
wire g20903;
wire g22217;
wire g34798;
wire g28105;
wire II28349;
wire g9759;
wire g32555;
wire II18060;
wire gbuf91;
wire g28589;
wire gbuf52;
wire g21959;
wire g30921;
wire g10371;
wire g34752;
wire g33503;
wire II31321;
wire g29753;
wire g34324;
wire g20640;
wire II16150;
wire g31142;
wire g22074;
wire g8440;
wire g14063;
wire g28783;
wire g24117;
wire g20148;
wire g32094;
wire g32710;
wire g20875;
wire g17506;
wire g27667;
wire II29239;
wire g21995;
wire g18774;
wire g9462;
wire g16616;
wire g28321;
wire g34318;
wire g23605;
wire g34557;
wire g13698;
wire g21361;
wire g30589;
wire g32272;
wire g24418;
wire g34019;
wire g9479;
wire II12805;
wire g15820;
wire g28391;
wire II15341;
wire g8734;
wire g32597;
wire g14366;
wire g11147;
wire g18229;
wire g22640;
wire g27120;
wire g11991;
wire g10118;
wire g34641;
wire g16663;
wire g9220;
wire II18313;
wire g26937;
wire g28520;
wire g22202;
wire II26093;
wire II27509;
wire g17057;
wire g14034;
wire g34876;
wire g32256;
wire g30928;
wire g30540;
wire g27230;
wire g19517;
wire g25133;
wire g30267;
wire g28709;
wire g22623;
wire g26394;
wire g24135;
wire g21842;
wire g25368;
wire g7216;
wire g27652;
wire g17412;
wire g21457;
wire g7490;
wire g34772;
wire g30470;
wire g33264;
wire g22408;
wire g33384;
wire II23755;
wire g28540;
wire g30079;
wire g14418;
wire g33674;
wire g32888;
wire g21700;
wire g16515;
wire g24962;
wire g27768;
wire g30456;
wire g13882;
wire g17601;
wire g20127;
wire g31918;
wire g30126;
wire g24110;
wire g16224;
wire g34871;
wire g22034;
wire g22015;
wire g28431;
wire g21786;
wire g8686;
wire g27095;
wire g30299;
wire II12271;
wire II31186;
wire II12241;
wire g19480;
wire II31012;
wire g18877;
wire g26542;
wire g33241;
wire g28558;
wire g6887;
wire g13858;
wire g32646;
wire II22974;
wire g18621;
wire g7405;
wire g20068;
wire g25003;
wire g21778;
wire g7970;
wire g21393;
wire g29525;
wire g28965;
wire II21769;
wire g18499;
wire g25030;
wire g30468;
wire g18321;
wire g29648;
wire g25838;
wire g12076;
wire II32093;
wire g13920;
wire g34734;
wire g24066;
wire g33848;
wire II22280;
wire g20555;
wire g31881;
wire g27491;
wire g13799;
wire g23304;
wire g34668;
wire g29876;
wire g7116;
wire g32428;
wire g18831;
wire g33467;
wire II32621;
wire g30538;
wire g27254;
wire II21994;
wire g30515;
wire g23192;
wire g31168;
wire g20979;
wire g30194;
wire g19385;
wire g25756;
wire g12995;
wire g11676;
wire g32493;
wire g28548;
wire g23193;
wire g22304;
wire g16631;
wire g22021;
wire g13242;
wire g10184;
wire g19963;
wire g18706;
wire g10823;
wire g19755;
wire g27634;
wire g24349;
wire g13521;
wire g14611;
wire g25880;
wire g16692;
wire g18312;
wire g29312;
wire g22763;
wire g28339;
wire g33558;
wire g11976;
wire g28651;
wire g32881;
wire g20325;
wire g14331;
wire g34016;
wire g16449;
wire g14868;
wire g20651;
wire g33409;
wire g24447;
wire gbuf37;
wire g34211;
wire g10509;
wire g22497;
wire g21418;
wire g34884;
wire g7674;
wire g29991;
wire g25675;
wire g26358;
wire g10266;
wire g9439;
wire g22713;
wire g23619;
wire g14676;
wire g19388;
wire g21960;
wire g26607;
wire g34615;
wire II27504;
wire II25534;
wire g30398;
wire g24803;
wire g9510;
wire g13967;
wire g15147;
wire II21911;
wire g32099;
wire II24920;
wire g8237;
wire g13005;
wire II31251;
wire II24416;
wire g32904;
wire g33995;
wire g29551;
wire g15142;
wire g34609;
wire g12017;
wire g24477;
wire g20444;
wire g28491;
wire g30259;
wire g29238;
wire g34893;
wire II20793;
wire g29801;
wire g9699;
wire g23650;
wire g25091;
wire g15749;
wire g18305;
wire g26095;
wire g6918;
wire II15494;
wire II16129;
wire g21898;
wire g8411;
wire g31499;
wire g22752;
wire g28551;
wire g31906;
wire g25595;
wire g17197;
wire g20165;
wire g33283;
wire II15087;
wire g28234;
wire g18168;
wire II14905;
wire g33840;
wire g25229;
wire g28679;
wire II31356;
wire g25166;
wire g27966;
wire g34670;
wire g9518;
wire g8805;
wire g33486;
wire g27539;
wire g19452;
wire g32810;
wire II21162;
wire g33969;
wire g13215;
wire II12493;
wire g24141;
wire g21681;
wire g14164;
wire g22160;
wire g13341;
wire g17480;
wire g33921;
wire II16246;
wire g34268;
wire g15733;
wire g27469;
wire g22040;
wire g34161;
wire II16778;
wire g30362;
wire II18842;
wire g21054;
wire g32818;
wire II29225;
wire g29732;
wire g18575;
wire g32845;
wire g26904;
wire g20215;
wire g16597;
wire g21398;
wire g29605;
wire II24695;
wire g24174;
wire g33022;
wire g24761;
wire II29585;
wire g24797;
wire g7515;
wire g28143;
wire g12285;
wire II31247;
wire g33009;
wire g8567;
wire g12857;
wire g34746;
wire g13209;
wire g19526;
wire g33697;
wire g27967;
wire g29969;
wire g19606;
wire g10151;
wire g18162;
wire II32834;
wire g18528;
wire II12746;
wire g23548;
wire g9535;
wire II14939;
wire g8751;
wire g25447;
wire g9498;
wire g15132;
wire g20372;
wire g13545;
wire II31791;
wire g29252;
wire g26094;
wire g32291;
wire g14037;
wire g25787;
wire g25154;
wire II14679;
wire g13115;
wire g33626;
wire g11356;
wire g16184;
wire g27242;
wire g29951;
wire g24130;
wire g19359;
wire g11173;
wire g19145;
wire g6856;
wire g17174;
wire g31170;
wire g24329;
wire II22800;
wire g14434;
wire g34209;
wire g15730;
wire g21366;
wire g17430;
wire II20895;
wire g10381;
wire g32031;
wire g26694;
wire g15049;
wire g30408;
wire g28650;
wire II14158;
wire II25244;
wire g24221;
wire g16098;
wire g26546;
wire g27382;
wire g6831;
wire II17780;
wire g22865;
wire g11429;
wire g16764;
wire g32368;
wire II13031;
wire g30274;
wire g32638;
wire g20173;
wire g25264;
wire g15162;
wire g34951;
wire g34261;
wire g11823;
wire g34841;
wire g28493;
wire g7027;
wire g10532;
wire g28188;
wire II18909;
wire g21759;
wire g33941;
wire II18822;
wire g12117;
wire g14003;
wire g16119;
wire gbuf106;
wire g22659;
wire g34596;
wire g32388;
wire g24204;
wire g30180;
wire g13325;
wire g32824;
wire g13868;
wire g29509;
wire g18769;
wire g21512;
wire g15139;
wire g9373;
wire g26337;
wire g21382;
wire g32900;
wire g34867;
wire g25928;
wire g32789;
wire g18434;
wire II27523;
wire g18485;
wire g30997;
wire g10677;
wire g13500;
wire g28308;
wire II14992;
wire g10756;
wire g22197;
wire g16960;
wire g15042;
wire g18944;
wire g22056;
wire II32195;
wire II18858;
wire g28202;
wire g18454;
wire II21210;
wire g7471;
wire g32450;
wire g18110;
wire g23918;
wire g32044;
wire g9472;
wire g24273;
wire g10057;
wire g17788;
wire II22717;
wire II22710;
wire g22523;
wire g27329;
wire g32784;
wire g32117;
wire g11797;
wire g21902;
wire g27704;
wire II21300;
wire g18553;
wire II13684;
wire g14758;
wire g28095;
wire II26051;
wire g34413;
wire g26314;
wire II24552;
wire g33688;
wire g34072;
wire II20460;
wire g17532;
wire II20816;
wire g12160;
wire g11959;
wire g32657;
wire II14576;
wire g30498;
wire g6873;
wire g18723;
wire g32322;
wire g25417;
wire g18783;
wire g34217;
wire g7620;
wire g12578;
wire g18378;
wire g32183;
wire g22095;
wire g27341;
wire g10946;
wire g29956;
wire g17481;
wire g30507;
wire II31126;
wire g18824;
wire g29949;
wire g21783;
wire g20532;
wire II20495;
wire g15902;
wire g18255;
wire g28481;
wire g15582;
wire II31081;
wire g32277;
wire g12195;
wire g16195;
wire II19851;
wire g26104;
wire g9434;
wire g26293;
wire g25901;
wire g28624;
wire g34434;
wire g33149;
wire g14790;
wire g21860;
wire g28219;
wire g24097;
wire g13020;
wire II23949;
wire g14567;
wire g18595;
wire g9575;
wire II14609;
wire g27994;
wire II32797;
wire g30347;
wire g9416;
wire g24915;
wire g11653;
wire g18338;
wire g32355;
wire g11740;
wire g33808;
wire g32985;
wire g31875;
wire g26235;
wire g25324;
wire g9291;
wire g33723;
wire g26782;
wire g25238;
wire g34527;
wire g34974;
wire g10120;
wire g32893;
wire g33822;
wire g30321;
wire g30444;
wire II12067;
wire II28185;
wire II15212;
wire g31816;
wire g23526;
wire g10139;
wire g27574;
wire g31486;
wire II24015;
wire g29716;
wire g25683;
wire g27300;
wire II31286;
wire g34400;
wire g29960;
wire g34066;
wire II12618;
wire g27666;
wire g16871;
wire g30605;
wire g34990;
wire g14188;
wire g26825;
wire g20239;
wire II11892;
wire g30431;
wire g19856;
wire II16455;
wire g8696;
wire g18592;
wire g17714;
wire g33690;
wire g21714;
wire g24971;
wire g9780;
wire g30084;
wire g19878;
wire II22177;
wire g10060;
wire g28749;
wire g34085;
wire g28812;
wire II24784;
wire g14599;
wire g6905;
wire g27153;
wire g12322;
wire g32567;
wire g20180;
wire g32471;
wire g18645;
wire II18568;
wire g24191;
wire g28658;
wire g20608;
wire g29180;
wire II22684;
wire g29328;
wire II13731;
wire g18178;
wire g11576;
wire g18393;
wire g20772;
wire g33736;
wire II14839;
wire g16129;
wire g31890;
wire g9552;
wire II14956;
wire II11746;
wire g10488;
wire g24787;
wire g13307;
wire g15574;
wire g14548;
wire g10683;
wire g34930;
wire II32820;
wire II29438;
wire g27320;
wire g22180;
wire g30417;
wire II14229;
wire g29635;
wire g14393;
wire II32525;
wire g21661;
wire g19402;
wire g7262;
wire g16966;
wire g24766;
wire g7693;
wire g17156;
wire g33608;
wire g30411;
wire II18421;
wire g12865;
wire g31221;
wire g17765;
wire g16719;
wire g17725;
wire g15054;
wire g8956;
wire g20390;
wire g33161;
wire g32765;
wire g29106;
wire g32614;
wire II26936;
wire g33125;
wire II18101;
wire II31041;
wire g28621;
wire g10086;
wire g21943;
wire II14602;
wire g15789;
wire g29540;
wire II21238;
wire g22317;
wire g31518;
wire g29172;
wire II22937;
wire g18140;
wire g17814;
wire g32305;
wire g12135;
wire g7597;
wire g28403;
wire g26387;
wire II18262;
wire II16489;
wire g18331;
wire g21726;
wire g32216;
wire II29303;
wire II16512;
wire g20056;
wire g12012;
wire g18800;
wire g33067;
wire g10873;
wire g21831;
wire g28048;
wire g9648;
wire g32167;
wire g23886;
wire g34108;
wire g33839;
wire g30024;
wire g9984;
wire g30489;
wire g12879;
wire g28538;
wire g27108;
wire g22868;
wire g7716;
wire g34365;
wire g19588;
wire g27415;
wire g19567;
wire g30113;
wire g33493;
wire g25960;
wire g23879;
wire g24308;
wire g33429;
wire g11950;
wire g20197;
wire g16816;
wire g25615;
wire II23917;
wire g32854;
wire g27305;
wire g28531;
wire II32364;
wire g18799;
wire g23488;
wire g27100;
wire g25113;
wire II24334;
wire g23942;
wire g23403;
wire g7533;
wire g34020;
wire g8515;
wire g34718;
wire g27367;
wire g6845;
wire II17585;
wire g8481;
wire g20575;
wire g11937;
wire g25594;
wire g18403;
wire g24393;
wire g25045;
wire g25892;
wire g16021;
wire g23006;
wire g33400;
wire g9620;
wire g28775;
wire II32228;
wire II33261;
wire g29672;
wire g24013;
wire g16278;
wire g21389;
wire g19792;
wire g34450;
wire g12905;
wire g30056;
wire g12856;
wire g24933;
wire g32036;
wire g25298;
wire g14336;
wire g21814;
wire g34912;
wire II18782;
wire g29811;
wire g25852;
wire g21969;
wire II24555;
wire g10569;
wire II22128;
wire g22058;
wire g18380;
wire g25172;
wire g32851;
wire g11862;
wire g33856;
wire II20499;
wire g24127;
wire g24354;
wire II32671;
wire g24765;
wire g13305;
wire g31668;
wire g31228;
wire g17410;
wire g16026;
wire g15112;
wire g32258;
wire g21770;
wire g23406;
wire II31157;
wire g28235;
wire g9834;
wire g25817;
wire g20531;
wire g24248;
wire g9621;
wire g16726;
wire g24433;
wire g8278;
wire g28628;
wire g34803;
wire II12013;
wire g21967;
wire II14222;
wire II20233;
wire g28112;
wire g29232;
wire g16925;
wire g27492;
wire g23809;
wire g24732;
wire g23047;
wire g14220;
wire g9338;
wire II14999;
wire g16740;
wire g28092;
wire g10695;
wire g7246;
wire g11192;
wire g26788;
wire g32779;
wire g30476;
wire g18366;
wire g25959;
wire g18615;
wire g18538;
wire g25048;
wire II15587;
wire g14337;
wire g17812;
wire g7440;
wire II30995;
wire g26603;
wire g30532;
wire g30458;
wire g7636;
wire g32180;
wire g21124;
wire g25662;
wire g7115;
wire g24911;
wire g8904;
wire II16847;
wire g34478;
wire g21852;
wire g10947;
wire g27301;
wire II27534;
wire g33428;
wire g23028;
wire g9901;
wire g33401;
wire gbuf10;
wire II14069;
wire II21978;
wire g18358;
wire g29856;
wire g31646;
wire g28436;
wire g9969;
wire g21559;
wire g32300;
wire II15542;
wire g9184;
wire g22178;
wire g23280;
wire g22063;
wire g9830;
wire g28138;
wire g18489;
wire g16186;
wire g32383;
wire g33290;
wire g16759;
wire g25873;
wire g13326;
wire g29868;
wire g34275;
wire g24059;
wire g30414;
wire g10877;
wire II15174;
wire g18339;
wire g10732;
wire g30038;
wire g9809;
wire g25605;
wire g29921;
wire g10872;
wire g11545;
wire g27283;
wire g26684;
wire II16040;
wire g15876;
wire g31188;
wire g34024;
wire g11250;
wire g24340;
wire g6818;
wire g20066;
wire g30445;
wire g10685;
wire g27685;
wire g15119;
wire II21285;
wire g26655;
wire g12874;
wire II26700;
wire g14384;
wire g32034;
wire g34260;
wire g32426;
wire g30328;
wire g9962;
wire g11980;
wire g32553;
wire g26721;
wire g32307;
wire g22514;
wire g11472;
wire g32544;
wire g33585;
wire g27800;
wire g20571;
wire g19631;
wire g30273;
wire g33851;
wire g15168;
wire g13866;
wire g31288;
wire g16844;
wire g22194;
wire g33242;
wire g33616;
wire g14544;
wire g27107;
wire II28908;
wire g14490;
wire g26091;
wire g12116;
wire g33800;
wire g18904;
wire g29145;
wire g29710;
wire g28380;
wire II32109;
wire g33714;
wire g32678;
wire g25126;
wire g30172;
wire g21511;
wire g24936;
wire g34960;
wire g34082;
wire g22756;
wire g24376;
wire g33484;
wire II31026;
wire gbuf89;
wire g32244;
wire g28318;
wire g23445;
wire g29963;
wire g21896;
wire g18786;
wire g22161;
wire g29034;
wire g21928;
wire g8219;
wire g31266;
wire II14705;
wire g27340;
wire g9246;
wire g25321;
wire g33037;
wire g14398;
wire g12018;
wire g24132;
wire g20642;
wire II15288;
wire g28625;
wire g19275;
wire g18257;
wire g17428;
wire g29683;
wire II22461;
wire g23362;
wire II20744;
wire g14642;
wire g33743;
wire g11117;
wire g32037;
wire II20584;
wire II32274;
wire g29060;
wire II16593;
wire g11829;
wire g34210;
wire g18196;
wire g8669;
wire g22903;
wire g18164;
wire g9451;
wire g28311;
wire g21944;
wire g14145;
wire g17502;
wire II18581;
wire g17753;
wire g27826;
wire g29195;
wire g29349;
wire II27368;
wire g14804;
wire g26656;
wire II26130;
wire g27205;
wire g18993;
wire g29652;
wire g27932;
wire g22652;
wire g18102;
wire g29938;
wire II26451;
wire g13996;
wire g31766;
wire g17488;
wire g22122;
wire g22031;
wire g23363;
wire g15716;
wire g28899;
wire II14271;
wire g20537;
wire g15058;
wire g11954;
wire g23522;
wire g11032;
wire g34633;
wire g23061;
wire g25116;
wire II15556;
wire II18839;
wire g22492;
wire g13462;
wire g24622;
wire g23909;
wire g26298;
wire g14405;
wire g33863;
wire g8461;
wire g18594;
wire g20917;
wire g15633;
wire g34041;
wire g26909;
wire II28838;
wire g23529;
wire g32398;
wire g20183;
wire II14186;
wire g31901;
wire g18191;
wire g30316;
wire II14351;
wire g24919;
wire g28535;
wire g21431;
wire g18462;
wire II14830;
wire II32518;
wire g23528;
wire II14518;
wire g26102;
wire g30558;
wire g12208;
wire g19544;
wire g32891;
wire g28020;
wire g11938;
wire g11953;
wire g9683;
wire II31523;
wire II14855;
wire g33523;
wire g32295;
wire II22761;
wire g10222;
wire g13383;
wire g27093;
wire g31316;
wire g10081;
wire g34073;
wire g31498;
wire g32187;
wire g8227;
wire g11006;
wire g23659;
wire II31642;
wire g12344;
wire g17767;
wire g17513;
wire g31940;
wire g20236;
wire g9374;
wire g24274;
wire II18151;
wire g20212;
wire g13484;
wire g34216;
wire g23577;
wire gbuf82;
wire II15042;
wire g6961;
wire g21058;
wire g24096;
wire II14854;
wire g34439;
wire g22593;
wire g21810;
wire g13505;
wire g13963;
wire g20627;
wire g28208;
wire g9295;
wire g17181;
wire g11163;
wire g15036;
wire g27244;
wire g15067;
wire g16963;
wire g29882;
wire g22860;
wire g32821;
wire g33990;
wire g28415;
wire g16855;
wire g18154;
wire g15882;
wire II31232;
wire g21178;
wire g33703;
wire II12861;
wire g13271;
wire g30916;
wire II24383;
wire g24298;
wire g34583;
wire g30926;
wire II17557;
wire g23756;
wire II14745;
wire g28207;
wire g32996;
wire g22449;
wire g16124;
wire g11697;
wire II32352;
wire g11491;
wire g30161;
wire g10152;
wire g25005;
wire g18112;
wire g33175;
wire g33931;
wire II32150;
wire g21741;
wire II14532;
wire g26837;
wire g7593;
wire g24661;
wire II20487;
wire g23913;
wire g25017;
wire g20588;
wire g10384;
wire g28682;
wire g33758;
wire g32869;
wire g21304;
wire g16164;
wire g19440;
wire g19503;
wire g20328;
wire g29250;
wire II26430;
wire g11820;
wire g17120;
wire g8891;
wire g24706;
wire g11931;
wire g34180;
wire II31161;
wire g33631;
wire g19501;
wire g25625;
wire g7018;
wire g29941;
wire g13210;
wire g28496;
wire g18556;
wire g31566;
wire g34945;
wire g13258;
wire g28566;
wire g12839;
wire g15086;
wire II16579;
wire g23724;
wire g19957;
wire g17747;
wire g24384;
wire g29805;
wire g7461;
wire g33005;
wire g25024;
wire g21296;
wire g33555;
wire g11224;
wire g29342;
wire g16325;
wire g28470;
wire g20051;
wire g27537;
wire g8565;
wire g29351;
wire g32901;
wire g34605;
wire g12136;
wire g10841;
wire g22867;
wire g33660;
wire g9989;
wire g34845;
wire g28453;
wire II22240;
wire g16093;
wire g12604;
wire g30110;
wire II21757;
wire g23259;
wire g24185;
wire g25733;
wire g26785;
wire g25196;
wire g9574;
wire g15571;
wire g20082;
wire g17225;
wire g20102;
wire g31781;
wire g19600;
wire g34204;
wire g13202;
wire g22520;
wire II30746;
wire g34616;
wire g27474;
wire g7474;
wire g25244;
wire g14754;
wire g10503;
wire g23856;
wire II31212;
wire g19362;
wire g33268;
wire g26993;
wire II12876;
wire g14203;
wire g21707;
wire g29554;
wire g29706;
wire II31843;
wire g17268;
wire g32960;
wire g24652;
wire g30251;
wire g23545;
wire g19776;
wire g18640;
wire g32152;
wire II17461;
wire g17815;
wire g9060;
wire g15136;
wire II14228;
wire g21364;
wire g29239;
wire g17588;
wire g24996;
wire g25070;
wire II22866;
wire g13507;
wire g34283;
wire g23824;
wire g20707;
wire g24802;
wire g32760;
wire g14596;
wire g21838;
wire g32635;
wire g15907;
wire g18138;
wire g25213;
wire g33905;
wire g29188;
wire g23762;
wire g32613;
wire g18572;
wire g10794;
wire g29664;
wire g27879;
wire g15098;
wire g33929;
wire g8854;
wire g23480;
wire g21395;
wire II28014;
wire g23613;
wire g29318;
wire g25268;
wire II31021;
wire g13003;
wire g32279;
wire g11869;
wire g32819;
wire g32812;
wire g34771;
wire g16581;
wire g21277;
wire g21766;
wire g19336;
wire g11114;
wire g23779;
wire g8037;
wire g16307;
wire g14044;
wire g16716;
wire g21981;
wire g7268;
wire g31830;
wire g19569;
wire g26395;
wire g30434;
wire g9158;
wire g29773;
wire g29567;
wire g23615;
wire g18593;
wire g25910;
wire g24404;
wire g25169;
wire g18131;
wire g28330;
wire g29166;
wire g18413;
wire g27708;
wire g16968;
wire g8540;
wire g31949;
wire g12909;
wire II17901;
wire g13937;
wire g28547;
wire g18775;
wire g18703;
wire g23990;
wire II28567;
wire g17640;
wire g25188;
wire g28257;
wire g7191;
wire g14219;
wire g17474;
wire g14581;
wire II17661;
wire g28664;
wire g9716;
wire g13983;
wire g20079;
wire g20675;
wire g34109;
wire g12812;
wire g14296;
wire g11046;
wire g24640;
wire II23951;
wire g25043;
wire g32757;
wire g29108;
wire g28328;
wire II13906;
wire II21766;
wire II15030;
wire g24978;
wire g23865;
wire g14032;
wire g34743;
wire II32909;
wire g16511;
wire g20569;
wire g14668;
wire g12449;
wire g35002;
wire g30272;
wire g10348;
wire g10177;
wire g28587;
wire g23877;
wire g31924;
wire g28260;
wire g26389;
wire gbuf108;
wire g20131;
wire g27117;
wire g12086;
wire g14256;
wire g23194;
wire g32485;
wire g18143;
wire g33257;
wire II31166;
wire g28683;
wire g21848;
wire gbuf72;
wire g24683;
wire g23424;
wire g29599;
wire g31987;
wire g23349;
wire II26503;
wire g24990;
wire g9595;
wire g12465;
wire II14816;
wire g20320;
wire g24216;
wire g13663;
wire g13795;
wire g32787;
wire g33058;
wire II31604;
wire g24231;
wire g33844;
wire g32259;
wire g23889;
wire g27659;
wire g13885;
wire g23646;
wire g34564;
wire g18879;
wire g19709;
wire g19954;
wire g8091;
wire g18400;
wire g11992;
wire g30731;
wire II28548;
wire g7972;
wire g23686;
wire g17190;
wire g26889;
wire II16821;
wire g19586;
wire g34345;
wire g34469;
wire g14639;
wire g9095;
wire II31550;
wire g16232;
wire g8418;
wire g20558;
wire g17328;
wire II11980;
wire g18809;
wire g13102;
wire g8883;
wire g28595;
wire g20553;
wire g18981;
wire g19784;
wire II23688;
wire g24167;
wire g18236;
wire g8362;
wire g10194;
wire g21349;
wire g12169;
wire g32951;
wire g16516;
wire g29269;
wire g34099;
wire g13945;
wire g7227;
wire g20006;
wire g29526;
wire g14908;
wire g30356;
wire g21984;
wire g17087;
wire g30076;
wire g18730;
wire g24759;
wire g11306;
wire g24953;
wire g28697;
wire g29898;
wire g17584;
wire II31466;
wire g32363;
wire g32541;
wire g34505;
wire g23385;
wire g21777;
wire g18487;
wire g31151;
wire g13109;
wire g24869;
wire g26963;
wire g11155;
wire g15105;
wire g34127;
wire g18521;
wire g27258;
wire g32217;
wire g7791;
wire g25290;
wire II18752;
wire g29588;
wire g15819;
wire II17668;
wire g11960;
wire g13954;
wire g32666;
wire g25337;
wire g22873;
wire g32265;
wire g18292;
wire g12910;
wire g33390;
wire g25751;
wire g10341;
wire g10624;
wire g27556;
wire g16237;
wire II32470;
wire g12080;
wire g17952;
wire II25680;
wire g33316;
wire g25034;
wire g24814;
wire g31933;
wire g13605;
wire g8681;
wire g34712;
wire g23217;
wire g11363;
wire g33526;
wire g18122;
wire II13499;
wire g31852;
wire g27092;
wire g28818;
wire g21956;
wire g34326;
wire g30366;
wire g20617;
wire g32371;
wire g14602;
wire g32782;
wire g13861;
wire g18129;
wire g23323;
wire g34071;
wire g27009;
wire g26629;
wire g27377;
wire g16639;
wire gbuf30;
wire g30103;
wire g9751;
wire g26312;
wire II17575;
wire g27347;
wire g20381;
wire g15848;
wire g13240;
wire g18891;
wire g30611;
wire g18548;
wire II25689;
wire g21662;
wire g9252;
wire g32724;
wire g26183;
wire g27212;
wire g27597;
wire g12920;
wire g27126;
wire g22942;
wire g16806;
wire g33507;
wire II28301;
wire g10581;
wire g30286;
wire g28850;
wire g25137;
wire II13067;
wire g32730;
wire g33692;
wire g22133;
wire g28722;
wire g32497;
wire II18713;
wire II24434;
wire g32234;
wire II18006;
wire g23307;
wire g33682;
wire g18119;
wire g34602;
wire g25835;
wire g26846;
wire g30147;
wire g32885;
wire II11877;
wire g30152;
wire g29293;
wire g7157;
wire g32598;
wire g14413;
wire g27487;
wire g20190;
wire II12764;
wire g22219;
wire g25181;
wire g14359;
wire II23357;
wire g30528;
wire g33028;
wire g21883;
wire g16280;
wire g22012;
wire g26946;
wire g22103;
wire g23796;
wire g26930;
wire g21733;
wire g23793;
wire g16773;
wire g31145;
wire g31849;
wire g32512;
wire II20369;
wire g30006;
wire g20671;
wire g29498;
wire g26917;
wire g15740;
wire g22214;
wire g28643;
wire g23261;
wire g25975;
wire g33989;
wire g21286;
wire g28578;
wire g21821;
wire g24225;
wire g18329;
wire g28755;
wire g10699;
wire g32153;
wire g25546;
wire g25952;
wire g18600;
wire g9598;
wire II22819;
wire g22209;
wire II14884;
wire g10999;
wire g21407;
wire g22006;
wire g24630;
wire g21884;
wire g23203;
wire II12263;
wire g27243;
wire g24887;
wire g26379;
wire g18757;
wire g8163;
wire g34953;
wire g28418;
wire g22001;
wire II13762;
wire g26230;
wire g34701;
wire g31826;
wire g25777;
wire g15224;
wire g31895;
wire g24794;
wire g31747;
wire g31970;
wire II33119;
wire g28087;
wire g33042;
wire g26130;
wire g25747;
wire g13267;
wire g7752;
wire g9742;
wire g14874;
wire g21561;
wire II29985;
wire g25081;
wire II22886;
wire g13314;
wire II22753;
wire g22540;
wire g33914;
wire g24465;
wire g32731;
wire g16047;
wire g25640;
wire g18322;
wire g6799;
wire g26892;
wire g14858;
wire g11431;
wire g32533;
wire g7487;
wire g33086;
wire g7544;
wire g23750;
wire g23607;
wire g16287;
wire g27977;
wire g29504;
wire g25482;
wire II27558;
wire g16052;
wire g10727;
wire g32703;
wire g33540;
wire g18277;
wire g28119;
wire g19756;
wire g33518;
wire g14755;
wire g23339;
wire g29364;
wire g32684;
wire g33812;
wire g18226;
wire g28451;
wire g22989;
wire g18663;
wire g8052;
wire g16877;
wire g29251;
wire g28703;
wire g15156;
wire g28352;
wire g13045;
wire g28744;
wire gbuf15;
wire g10287;
wire II17198;
wire g17092;
wire g34471;
wire g33559;
wire g30311;
wire g12225;
wire II18778;
wire g31961;
wire g19573;
wire g29043;
wire g34390;
wire g13761;
wire g32958;
wire g22759;
wire II28199;
wire g6754;
wire g19127;
wire g33365;
wire g34963;
wire g10229;
wire g34910;
wire II25511;
wire g24118;
wire g28153;
wire g33465;
wire g19676;
wire g24108;
wire g26817;
wire g27762;
wire g20700;
wire II31569;
wire g34882;
wire g19358;
wire g20594;
wire gbuf63;
wire g19684;
wire g30001;
wire g19666;
wire g29321;
wire g13059;
wire g34300;
wire II24710;
wire g32235;
wire II27546;
wire g26171;
wire g22721;
wire g24429;
wire g18700;
wire II17723;
wire g9092;
wire g30542;
wire g23843;
wire g28483;
wire g33583;
wire II33106;
wire II15942;
wire g11621;
wire g7836;
wire II15073;
wire II23339;
wire g22024;
wire g10181;
wire g16625;
wire g19672;
wire g30486;
wire g26544;
wire g13631;
wire g18318;
wire g12318;
wire g14420;
wire g34872;
wire g9298;
wire II16775;
wire g20534;
wire g34447;
wire g10308;
wire g29583;
wire g27057;
wire g9488;
wire g18416;
wire II24603;
wire g32877;
wire g27589;
wire gbuf5;
wire g20751;
wire II29207;
wire g6841;
wire g29618;
wire II17923;
wire II16535;
wire g26247;
wire II24385;
wire g17292;
wire g14918;
wire g11910;
wire g18498;
wire g7803;
wire g21925;
wire g30230;
wire g19267;
wire g15735;
wire g34301;
wire g24879;
wire g9776;
wire II31545;
wire g7400;
wire g14830;
wire g30459;
wire g22957;
wire g27260;
wire gbuf116;
wire g29754;
wire g20775;
wire g27013;
wire g27141;
wire II15365;
wire g33099;
wire g15580;
wire g27004;
wire g24544;
wire g30509;
wire g29067;
wire g23201;
wire g25300;
wire g9316;
wire II18078;
wire g28606;
wire g15371;
wire g29895;
wire g19557;
wire g18173;
wire g26574;
wire g13063;
wire II29278;
wire g14937;
wire g24602;
wire g9602;
wire g16654;
wire g33951;
wire g26254;
wire g8593;
wire g21426;
wire g34677;
wire II32803;
wire g9177;
wire g18495;
wire g17618;
wire g18698;
wire II31272;
wire g6838;
wire g9449;
wire g13628;
wire II22366;
wire g24775;
wire g12940;
wire g18949;
wire II14330;
wire g20506;
wire g10159;
wire g10350;
wire II29185;
wire II15667;
wire g32641;
wire g13177;
wire g23083;
wire g18422;
wire g9848;
wire g25673;
wire g13671;
wire II12823;
wire g25567;
wire g32611;
wire g15594;
wire g19439;
wire g12144;
wire II19348;
wire g24120;
wire g15832;
wire g31503;
wire g13927;
wire g22405;
wire g29875;
wire g11893;
wire II22852;
wire g31484;
wire g24982;
wire II31326;
wire g24790;
wire g27645;
wire g20163;
wire g19343;
wire g27221;
wire g25632;
wire g28371;
wire g23931;
wire g33564;
wire g29334;
wire g25690;
wire g33431;
wire g30396;
wire g19472;
wire g25207;
wire g23585;
wire g28642;
wire g24540;
wire g12038;
wire g12414;
wire g23491;
wire g33994;
wire II14428;
wire g34147;
wire g29531;
wire g32239;
wire g30378;
wire g29520;
wire g33696;
wire g32989;
wire g34520;
wire g10472;
wire g28443;
wire II17442;
wire g34092;
wire g29998;
wire g33281;
wire g13889;
wire g32832;
wire g33176;
wire g31252;
wire g29326;
wire g30213;
wire II16476;
wire g33750;
wire g7928;
wire g15995;
wire g8830;
wire g19604;
wire g12378;
wire g16072;
wire g24332;
wire g30421;
wire g7236;
wire g32916;
wire g32410;
wire g18533;
wire g34536;
wire g12577;
wire g23954;
wire g27827;
wire g9517;
wire g25598;
wire g33735;
wire g26275;
wire g32029;
wire g29355;
wire II31342;
wire g17364;
wire g24072;
wire g24719;
wire g22088;
wire g6849;
wire g23219;
wire g17138;
wire g34191;
wire g20041;
wire II21810;
wire g24495;
wire g17477;
wire g32665;
wire g16883;
wire g15706;
wire g11268;
wire g11963;
wire g18387;
wire g11039;
wire g23236;
wire g15591;
wire g27483;
wire g31271;
wire g32805;
wire g21068;
wire g25694;
wire g20271;
wire g29244;
wire II14610;
wire g18252;
wire g34978;
wire g29153;
wire II19796;
wire g12483;
wire g27565;
wire g23996;
wire II14749;
wire g32692;
wire II33288;
wire g18582;
wire g18198;
wire g23450;
wire g32345;
wire II11721;
wire g22199;
wire g9862;
wire g25104;
wire g30098;
wire g31854;
wire g27044;
wire g33092;
wire g24043;
wire g33727;
wire g25012;
wire g18568;
wire g27338;
wire g11875;
wire II18885;
wire g18672;
wire g9916;
wire II25845;
wire g32351;
wire g32882;
wire II31515;
wire g28654;
wire g27731;
wire g30300;
wire g18288;
wire II22922;
wire g8676;
wire g12886;
wire II13729;
wire g28342;
wire g15913;
wire g20193;
wire g24169;
wire g7535;
wire II32473;
wire g34032;
wire II31236;
wire g15914;
wire g32474;
wire II12580;
wire g25783;
wire g27182;
wire g28529;
wire II14593;
wire g26803;
wire g26755;
wire g12124;
wire g21798;
wire g30032;
wire g23474;
wire g14116;
wire II24781;
wire g31707;
wire g30226;
wire g8281;
wire g7960;
wire g34270;
wire II16111;
wire g28313;
wire g11018;
wire g24360;
wire g22901;
wire g6975;
wire g10160;
wire g31666;
wire g32281;
wire g15871;
wire g33235;
wire g10402;
wire g32506;
wire g25613;
wire g12120;
wire II33297;
wire g16802;
wire II12790;
wire g16856;
wire g29579;
wire g19513;
wire g12954;
wire g9364;
wire g9013;
wire g16191;
wire g17699;
wire g26834;
wire g30493;
wire g32430;
wire g7586;
wire g17706;
wire g21951;
wire II21258;
wire II30331;
wire g14343;
wire g13330;
wire g12043;
wire g17141;
wire II13805;
wire g32459;
wire g7777;
wire g33833;
wire g10570;
wire g25377;
wire g33494;
wire g20091;
wire g20167;
wire II31242;
wire gbuf144;
wire II15572;
wire g32941;
wire g26874;
wire g27521;
wire g12550;
wire g9036;
wire g34508;
wire g23987;
wire g32455;
wire g23589;
wire g25561;
wire g32629;
wire II26393;
wire g25725;
wire g28038;
wire g21918;
wire g29360;
wire g28843;
wire g6992;
wire g12235;
wire g23057;
wire g29926;
wire g25138;
wire g25531;
wire g32769;
wire g9971;
wire g26711;
wire g10058;
wire g8643;
wire g31473;
wire II16193;
wire g9547;
wire g21456;
wire II22298;
wire g18336;
wire g34130;
wire g34372;
wire g30505;
wire g19716;
wire g24438;
wire g18642;
wire g17679;
wire g13779;
wire g14686;
wire g27612;
wire g16030;
wire g9309;
wire g31800;
wire II26929;
wire g12889;
wire g17409;
wire g28054;
wire g17494;
wire g11686;
wire g23278;
wire g23558;
wire g19886;
wire g32562;
wire g30012;
wire g32912;
wire g28162;
wire g16181;
wire g21972;
wire II13872;
wire g23243;
wire g32858;
wire g28405;
wire g27929;
wire g33245;
wire g10232;
wire g34174;
wire II15600;
wire g20178;
wire g29080;
wire g15051;
wire g20065;
wire g31232;
wire g15170;
wire II16163;
wire g14139;
wire g24398;
wire g14536;
wire g26651;
wire g26736;
wire g11234;
wire g7616;
wire g31774;
wire g10709;
wire g14396;
wire g29848;
wire g25202;
wire g25411;
wire g24060;
wire gbuf126;
wire II22525;
wire II20609;
wire g13038;
wire g32770;
wire II18543;
wire g33604;
wire g19636;
wire g32020;
wire g6829;
wire g23487;
wire II30054;
wire g33594;
wire g32228;
wire g7163;
wire g26718;
wire g17692;
wire g17467;
wire g25884;
wire g31373;
wire g23500;
wire II29271;
wire g29177;
wire g23358;
wire II32309;
wire g25940;
wire g32949;
wire II32116;
wire g23552;
wire g32752;
wire g33804;
wire g18354;
wire g28927;
wire II15932;
wire g33578;
wire II14395;
wire g32314;
wire II33264;
wire g22299;
wire g21724;
wire II22762;
wire g23392;
wire g24557;
wire g28526;
wire g18201;
wire g23691;
wire g32849;
wire g34749;
wire g32828;
wire g33412;
wire g20036;
wire g16809;
wire g10760;
wire g23399;
wire g9806;
wire g27063;
wire g23457;
wire II23711;
wire g28718;
wire g26828;
wire g8133;
wire g28885;
wire g23538;
wire g29302;
wire g23569;
wire II31061;
wire II31672;
wire g29785;
wire g12629;
wire g33355;
wire g8806;
wire g11927;
wire g24239;
wire II15107;
wire g20764;
wire g34297;
wire g28291;
wire g26900;
wire II26508;
wire g33479;
wire II21838;
wire g18467;
wire g29078;
wire g9489;
wire g26612;
wire II26418;
wire g29886;
wire g23210;
wire II17143;
wire g33204;
wire g25720;
wire g29619;
wire g11326;
wire g20656;
wire g30130;
wire g28363;
wire g32584;
wire g30184;
wire g14968;
wire g11290;
wire g34316;
wire g23901;
wire II32960;
wire g25731;
wire g24716;
wire II25161;
wire g24550;
wire g29376;
wire II16328;
wire g9748;
wire g32991;
wire g34286;
wire g27429;
wire g32286;
wire g11414;
wire g13542;
wire g29857;
wire g23431;
wire g17672;
wire g32338;
wire II31800;
wire g23623;
wire g26634;
wire g18779;
wire g27774;
wire g25266;
wire g17792;
wire g10212;
wire g28147;
wire II33249;
wire g7110;
wire g22982;
wire g12143;
wire g13809;
wire g14914;
wire g29955;
wire g16482;
wire II22149;
wire g32209;
wire g16506;
wire g10115;
wire II18788;
wire II30756;
wire g7947;
wire g25872;
wire g30386;
wire g33094;
wire g8310;
wire g19363;
wire g34726;
wire g12367;
wire II32237;
wire g33329;
wire g24288;
wire g12294;
wire g10720;
wire II11835;
wire g28614;
wire g24872;
wire II12373;
wire g32602;
wire g9927;
wire g28303;
wire g27219;
wire g8623;
wire g34062;
wire g34674;
wire g19788;
wire g27710;
wire g23861;
wire g29835;
wire g34942;
wire g15101;
wire II15682;
wire g32114;
wire g19746;
wire g31750;
wire g14097;
wire g34139;
wire g15674;
wire g31928;
wire II31277;
wire II32678;
wire g7431;
wire g7315;
wire g16608;
wire II31051;
wire g7497;
wire II22353;
wire II29211;
wire II27513;
wire g34250;
wire g7275;
wire g34483;
wire II29221;
wire g27577;
wire g14075;
wire g9021;
wire g16769;
wire g7957;
wire g21465;
wire g30191;
wire g18451;
wire II18350;
wire g12526;
wire g27525;
wire g22051;
wire g31795;
wire g30984;
wire g23283;
wire g24005;
wire g30983;
wire g27996;
wire g22019;
wire g33976;
wire g11134;
wire g30609;
wire g33036;
wire g34748;
wire g20229;
wire g25905;
wire g7344;
wire g12830;
wire g19140;
wire g10967;
wire g24178;
wire II17892;
wire g12841;
wire g24156;
wire gbuf137;
wire g33623;
wire g19651;
wire g23800;
wire g19522;
wire g14320;
wire g16738;
wire g21803;
wire g34795;
wire II13637;
wire g19353;
wire g29255;
wire II11697;
wire II22785;
wire g31809;
wire g27673;
wire g7362;
wire g20110;
wire g26700;
wire g21066;
wire g22488;
wire g11346;
wire g23915;
wire g21703;
wire II14714;
wire g25539;
wire II16201;
wire g34446;
wire g28950;
wire g30264;
wire g25629;
wire g29945;
wire g26208;
wire g13024;
wire g20528;
wire g34591;
wire II18154;
wire g16731;
wire g27437;
wire g14307;
wire g10272;
wire g27613;
wire g31507;
wire II12568;
wire II22499;
wire g31003;
wire g24744;
wire g25495;
wire g20387;
wire II18177;
wire g20698;
wire g13716;
wire g21915;
wire g21333;
wire g12287;
wire g23725;
wire g29850;
wire g25576;
wire g18658;
wire g7397;
wire g10090;
wire g14519;
wire g20446;
wire g21737;
wire g24603;
wire g30157;
wire g30552;
wire g12342;
wire g29071;
wire g34244;
wire g13410;
wire g7648;
wire g33332;
wire g18375;
wire g17392;
wire g8282;
wire g30294;
wire II23601;
wire g13415;
wire g24255;
wire g14453;
wire II23120;
wire g17684;
wire II24448;
wire g12853;
wire g33133;
wire II27555;
wire g25453;
wire g34541;
wire g7139;
wire g27925;
wire g29573;
wire g24607;
wire g27964;
wire g18820;
wire g17654;
wire g15968;
wire g25879;
wire g25425;
wire II16762;
wire g33100;
wire g12890;
wire g21246;
wire g34460;
wire II25146;
wire g9259;
wire g16861;
wire g19399;
wire II19775;
wire g9800;
wire g9660;
wire g13077;
wire g14048;
wire g31944;
wire g18940;
wire g12188;
wire g30255;
wire g11878;
wire g19139;
wire g19801;
wire g32122;
wire g10827;
wire g28789;
wire g19063;
wire g13516;
wire g28441;
wire g25297;
wire g33377;
wire g20637;
wire g30534;
wire g12191;
wire g28076;
wire g29763;
wire g25407;
wire g18134;
wire g18283;
wire II29571;
wire g18829;
wire g34857;
wire g18712;
wire g12862;
wire g29742;
wire g27202;
wire II18446;
wire g7456;
wire g24979;
wire II13140;
wire g8356;
wire g33110;
wire g12046;
wire g17668;
wire g33968;
wire g12651;
wire g34813;
wire g34869;
wire g33902;
wire g33897;
wire g29712;
wire g33117;
wire II22576;
wire II14368;
wire g22079;
wire g33477;
wire g8296;
wire g23062;
wire g7522;
wire g10605;
wire g31866;
wire g22456;
wire g29512;
wire g19662;
wire g23484;
wire g30080;
wire g32979;
wire g33004;
wire g29109;
wire g34194;
wire g11126;
wire g27209;
wire g12794;
wire g32176;
wire g26880;
wire g27145;
wire g10363;
wire g18299;
wire g9669;
wire g33030;
wire g24485;
wire g25175;
wire g31995;
wire g18500;
wire g12511;
wire g27403;
wire g26156;
wire g31891;
wire g20151;
wire g34420;
wire g13514;
wire g15014;
wire g32583;
wire g31016;
wire II18531;
wire g13125;
wire II23324;
wire g21273;
wire g16637;
wire g30045;
wire g34864;
wire g23516;
wire g31019;
wire g10597;
wire g24579;
wire g9152;
wire g15712;
wire g26129;
wire g14528;
wire g8058;
wire g18181;
wire II12167;
wire g32674;
wire g18768;
wire g28532;
wire g26829;
wire g28100;
wire g9934;
wire g25502;
wire g12798;
wire g31821;
wire II23980;
wire g13959;
wire g23393;
wire g17720;
wire g15130;
wire g33081;
wire g10588;
wire g15841;
wire g19499;
wire g23254;
wire g22836;
wire g33717;
wire II16651;
wire g15825;
wire II18529;
wire g32713;
wire g11513;
wire g6984;
wire g12817;
wire g34778;
wire II20188;
wire g23711;
wire II24585;
wire g26122;
wire g27561;
wire g24482;
wire g33261;
wire g19764;
wire g15694;
wire g9264;
wire g11881;
wire g32465;
wire g34122;
wire g14701;
wire g14348;
wire g34766;
wire g33539;
wire g25055;
wire g28395;
wire g27546;
wire gbuf78;
wire g18566;
wire g18449;
wire g30463;
wire g27628;
wire g29983;
wire II13111;
wire II23342;
wire g12081;
wire g34764;
wire g30121;
wire g6957;
wire g27468;
wire g31513;
wire g28511;
wire g24991;
wire g28691;
wire g32112;
wire g14194;
wire II18297;
wire g30020;
wire g28269;
wire g34610;
wire g6926;
wire g19980;
wire g7097;
wire g23221;
wire g17775;
wire g24822;
wire g34621;
wire g15093;
wire g18543;
wire g25060;
wire g25669;
wire g8742;
wire g29612;
wire g29483;
wire g13031;
wire g12871;
wire g24670;
wire g33909;
wire g10375;
wire g16526;
wire g29012;
wire g22149;
wire g28516;
wire g23340;
wire g13708;
wire II22583;
wire g16311;
wire g11945;
wire g20841;
wire II17626;
wire g30350;
wire g17152;
wire g15145;
wire g21385;
wire g13855;
wire g24524;
wire g18737;
wire g13940;
wire g24283;
wire g28857;
wire g10369;
wire g33982;
wire g13676;
wire g24943;
wire g18602;
wire II22024;
wire g7625;
wire g33383;
wire g18232;
wire g32015;
wire g18637;
wire g34006;
wire g10887;
wire g29913;
wire II12242;
wire g26344;
wire g31298;
wire g15071;
wire g32521;
wire g33532;
wire g24570;
wire II30989;
wire g16521;
wire II16721;
wire g21933;
wire g28946;
wire g32972;
wire g30519;
wire g17414;
wire g30500;
wire g31525;
wire g27506;
wire g30063;
wire g21844;
wire g20150;
wire g18509;
wire g32276;
wire g32896;
wire g14247;
wire g9888;
wire g21188;
wire g34682;
wire g27579;
wire g21825;
wire g18241;
wire g8898;
wire g15816;
wire g24247;
wire g28172;
wire g34512;
wire g34353;
wire g34048;
wire g33447;
wire g32737;
wire g25965;
wire g31811;
wire II31312;
wire g25069;
wire g17689;
wire g15725;
wire g14041;
wire g15797;
wire g24503;
wire g23378;
wire g20681;
wire II12779;
wire g14514;
wire g14996;
wire g24420;
wire g15962;
wire g33450;
wire g33937;
wire g23814;
wire g18934;
wire g13086;
wire g34455;
wire g13132;
wire g16593;
wire g20207;
wire g27583;
wire g33422;
wire g25242;
wire g29227;
wire II18600;
wire g18433;
wire g7567;
wire g33790;
wire g34171;
wire II32699;
wire II14633;
wire g22547;
wire II11629;
wire g11202;
wire g31118;
wire g32939;
wire g33145;
wire g24241;
wire g27395;
wire g32088;
wire g20706;
wire g21685;
wire g12902;
wire g26859;
wire g26284;
wire g28864;
wire g25557;
wire g32096;
wire II27508;
wire g31885;
wire g30394;
wire g22038;
wire g23003;
wire g28116;
wire g13458;
wire g23894;
wire g30177;
wire g9538;
wire g29183;
wire g18688;
wire g16216;
wire g23572;
wire g26250;
wire g20994;
wire g32572;
wire g11709;
wire g20087;
wire g13040;
wire g28158;
wire g10262;
wire g10610;
wire g14575;
wire II27388;
wire g24987;
wire g7632;
wire g14210;
wire g13821;
wire g20782;
wire g21428;
wire g21721;
wire g29906;
wire g31753;
wire g18301;
wire g22927;
wire g11182;
wire g23021;
wire g8778;
wire g25225;
wire g14727;
wire g13493;
wire g34699;
wire g24583;
wire g25895;
wire II33167;
wire g15061;
wire g13898;
wire g32930;
wire g21182;
wire II15732;
wire g25985;
wire g11442;
wire II32690;
wire g24567;
wire g25931;
wire g34490;
wire g26325;
wire g22643;
wire g34695;
wire g17719;
wire g27970;
wire II21242;
wire g13249;
wire II31352;
wire II18625;
wire g10413;
wire II16502;
wire g17246;
wire g27375;
wire g28288;
wire g34305;
wire g33049;
wire II15609;
wire g18517;
wire g34136;
wire g17193;
wire II13443;
wire g18887;
wire II31776;
wire g21872;
wire g23497;
wire g15839;
wire II33210;
wire g12981;
wire g19697;
wire g14423;
wire g10038;
wire g30499;
wire g29261;
wire g19474;
wire g33048;
wire g16535;
wire g20578;
wire g27029;
wire g28056;
wire g27971;
wire g33890;
wire g18340;
wire g12820;
wire g12435;
wire II15079;
wire g9429;
wire g29222;
wire II24033;
wire g12204;
wire g22975;
wire g27832;
wire g10473;
wire g32791;
wire g10394;
wire II26649;
wire g14092;
wire g12022;
wire g24122;
wire II31482;
wire g33297;
wire II31077;
wire g9842;
wire g29190;
wire g34499;
wire II12214;
wire g23514;
wire g21352;
wire g25657;
wire g33123;
wire g33344;
wire g15650;
wire g34037;
wire g23324;
wire g32052;
wire g25255;
wire g32620;
wire II12451;
wire g19733;
wire g8343;
wire g29371;
wire g33569;
wire g19414;
wire g12938;
wire g12107;
wire g34404;
wire g20695;
wire g32358;
wire II14276;
wire g31783;
wire g26081;
wire g16220;
wire g23223;
wire g32699;
wire g32839;
wire II12289;
wire II23381;
wire g31283;
wire II16371;
wire g23172;
wire g15150;
wire II20846;
wire g21346;
wire g13475;
wire g20669;
wire g31139;
wire g9670;
wire g31916;
wire g32984;
wire g30233;
wire g18347;
wire g16674;
wire g15750;
wire g17525;
wire g27356;
wire g34920;
wire II13184;
wire g28633;
wire g24626;
wire g28820;
wire g19430;
wire g20871;
wire g18175;
wire g12896;
wire II15846;
wire g22683;
wire g15937;
wire II31817;
wire II13326;
wire g26925;
wire g34187;
wire g23103;
wire g9283;
wire g20160;
wire g22707;
wire g27989;
wire g9073;
wire g27277;
wire g22090;
wire g9212;
wire g11446;
wire g11425;
wire g23665;
wire g25708;
wire g21607;
wire g14004;
wire g22922;
wire g29632;
wire g18717;
wire g31293;
wire II26460;
wire g24024;
wire g29778;
wire II31112;
wire g32206;
wire g21905;
wire g25938;
wire g18370;
wire II18819;
wire g25446;
wire g24296;
wire g7051;
wire g27084;
wire g10206;
wire g24321;
wire II32639;
wire g20564;
wire g24085;
wire g25153;
wire g12686;
wire g16296;
wire g11769;
wire g25644;
wire g19208;
wire g22666;
wire II32187;
wire g26089;
wire II12605;
wire g24265;
wire g17527;
wire gbuf94;
wire g13914;
wire g31466;
wire g32539;
wire g12638;
wire g20171;
wire g22447;
wire g21758;
wire II32192;
wire g21762;
wire g7686;
wire gbuf133;
wire g28204;
wire g25553;
wire g12371;
wire g16762;
wire g14447;
wire g27457;
wire II15811;
wire g27248;
wire II25677;
wire g14978;
wire g24799;
wire g32394;
wire g9197;
wire g16125;
wire g28499;
wire g10533;
wire g8397;
wire g34671;
wire g21879;
wire g29199;
wire II18168;
wire g16610;
wire g16596;
wire g10110;
wire g21383;
wire II22289;
wire g32864;
wire g11143;
wire g25773;
wire g32746;
wire g20585;
wire g7596;
wire II23963;
wire g9456;
wire g33700;
wire II32756;
wire g11480;
wire g34267;
wire g10380;
wire g24092;
wire g23927;
wire g33707;
wire g11002;
wire II14668;
wire gbuf148;
wire g20106;
wire g9534;
wire II22028;
wire g14079;
wire g7751;
wire g24270;
wire g32825;
wire II31581;
wire g25621;
wire g22714;
wire g29644;
wire g34842;
wire g32382;
wire g31141;
wire g29793;
wire g25737;
wire g32138;
wire gbuf86;
wire g25020;
wire g18472;
wire g24229;
wire g29809;
wire g20216;
wire g19580;
wire g10108;
wire g19417;
wire g21689;
wire g25995;
wire II26381;
wire II16028;
wire II14257;
wire II12300;
wire g7918;
wire II16024;
wire g23939;
wire g8612;
wire g22526;
wire g24923;
wire g7543;
wire g34914;
wire g22539;
wire g8290;
wire g15021;
wire g13480;
wire g28457;
wire g30399;
wire g22071;
wire g16321;
wire g19467;
wire II14170;
wire g11291;
wire g34556;
wire g32954;
wire g14360;
wire g18547;
wire g22098;
wire g24961;
wire g16747;
wire g18599;
wire g25221;
wire g8655;
wire g27233;
wire g34206;
wire g7823;
wire g8390;
wire II13007;
wire g33816;
wire g16629;
wire II23336;
wire g31609;
wire g23658;
wire g22417;
wire g10890;
wire g20623;
wire g34077;
wire g34184;
wire II12203;
wire g31921;
wire g8774;
wire g9747;
wire g30825;
wire g12609;
wire II11785;
wire g29073;
wire g26024;
wire g26907;
wire g27159;
wire g13623;
wire g13216;
wire II24027;
wire g9415;
wire II20189;
wire g33404;
wire g21283;
wire g32221;
wire II12049;
wire g23821;
wire g7259;
wire g26549;
wire II18344;
wire g14127;
wire II20747;
wire gbuf47;
wire g12497;
wire g25571;
wire g22864;
wire g9444;
wire II31271;
wire II14902;
wire g32886;
wire g19455;
wire g34756;
wire g24853;
wire g15615;
wire g27602;
wire g34033;
wire g12181;
wire II24415;
wire g27387;
wire g21360;
wire g20657;
wire g29278;
wire g24788;
wire g32997;
wire g13223;
wire g28837;
wire II21860;
wire g10190;
wire g31222;
wire g26485;
wire g25077;
wire g17818;
wire g11148;
wire g31261;
wire g33406;
wire g17573;
wire g25570;
wire g17655;
wire g22081;
wire II14204;
wire II14653;
wire g32840;
wire g8626;
wire II25869;
wire g6802;
wire g18694;
wire g13116;
wire g32815;
wire g25103;
wire g33785;
wire g22173;
wire g29959;
wire II22685;
wire g34230;
wire g13255;
wire g19770;
wire II18259;
wire II18382;
wire g30989;
wire g30365;
wire g13277;
wire g20699;
wire g28715;
wire g10566;
wire g33972;
wire g28793;
wire g34849;
wire II15129;
wire g14888;
wire II18107;
wire g14207;
wire g18825;
wire II32970;
wire g29667;
wire g20187;
wire g25050;
wire g29235;
wire g27875;
wire g8236;
wire g14184;
wire g33000;
wire g29205;
wire g22046;
wire g30309;
wire g14750;
wire g33573;
wire g10632;
wire g12239;
wire II32455;
wire g29292;
wire g19435;
wire g7438;
wire II24048;
wire g9433;
wire g10613;
wire g23873;
wire II17420;
wire g26971;
wire g28490;
wire II14119;
wire g31494;
wire g17533;
wire g17872;
wire g17781;
wire g34284;
wire g20703;
wire g11754;
wire g8359;
wire g24355;
wire g20441;
wire g14838;
wire g26096;
wire g23127;
wire g32639;
wire II18662;
wire g33613;
wire g34524;
wire g22491;
wire g27982;
wire g27991;
wire g23525;
wire g16585;
wire g19263;
wire g31476;
wire g21901;
wire g12878;
wire g23539;
wire II29894;
wire g33665;
wire g11309;
wire g20055;
wire g30034;
wire II30728;
wire g33499;
wire g15703;
wire II12159;
wire g21459;
wire g27518;
wire g14984;
wire g11891;
wire II23306;
wire g25755;
wire g31869;
wire g24436;
wire g30554;
wire g34661;
wire g8439;
wire g25044;
wire g28955;
wire g30472;
wire II13968;
wire g28479;
wire g24728;
wire II25882;
wire g23899;
wire g11984;
wire g13772;
wire g29802;
wire g8195;
wire g10121;
wire g16814;
wire g18581;
wire II31600;
wire II11632;
wire g34368;
wire g21963;
wire g16669;
wire g9966;
wire g26269;
wire g24975;
wire g32254;
wire II12219;
wire g9864;
wire g23629;
wire g34010;
wire g32408;
wire g12492;
wire gbuf97;
wire g21856;
wire g17470;
wire g24655;
wire g6875;
wire g24309;
wire g34276;
wire g26294;
wire II14766;
wire g26812;
wire II31101;
wire g23409;
wire g23402;
wire g30389;
wire g30093;
wire g30221;
wire g18611;
wire g33480;
wire g24932;
wire g18806;
wire g17635;
wire g32402;
wire g20852;
wire g25307;
wire g29863;
wire g8466;
wire g23148;
wire g18108;
wire g32548;
wire g32694;
wire g24344;
wire g31859;
wire g19589;
wire g34224;
wire II15193;
wire g12767;
wire g19872;
wire g34681;
wire II17552;
wire g14813;
wire g28676;
wire g29975;
wire II20318;
wire g18405;
wire g23460;
wire II13759;
wire g26725;
wire g7232;
wire II22692;
wire g33278;
wire g27569;
wire g33273;
wire g30490;
wire g18707;
wire g27135;
wire g18363;
wire g34646;
wire g28583;
wire g30402;
wire g31376;
wire g33607;
wire g11563;
wire II33285;
wire g32304;
wire g14872;
wire g18789;
wire g24769;
wire g31184;
wire II31748;
wire g8812;
wire g18396;
wire g14981;
wire II28832;
wire g13028;
wire g21050;
wire II31973;
wire g28712;
wire g17723;
wire g28554;
wire g26967;
wire g23993;
wire g20511;
wire g26994;
wire g18534;
wire g12705;
wire g30506;
wire g24500;
wire g28629;
wire g13301;
wire g30412;
wire g7619;
wire g30466;
wire g14977;
wire g27344;
wire g18296;
wire g21345;
wire g30107;
wire g33068;
wire II26050;
wire g12040;
wire g29179;
wire g26857;
wire g28539;
wire g30380;
wire g30343;
wire g17146;
wire g29315;
wire II15264;
wire g19576;
wire g25609;
wire g29925;
wire g34028;
wire g26229;
wire II15190;
wire II20035;
wire g22066;
wire g26077;
wire g12941;
wire g10399;
wire g21940;
wire II27567;
wire g16614;
wire g22843;
wire g21715;
wire g23380;
wire g11957;
wire g7780;
wire g33910;
wire g26673;
wire g34279;
wire g27690;
wire g25097;
wire g29537;
wire g33710;
wire g27961;
wire g15831;
wire g26329;
wire g12593;
wire g21748;
wire g25866;
wire g31212;
wire g18384;
wire g27663;
wire g21413;
wire g28469;
wire g24949;
wire g8505;
wire g32047;
wire g14149;
wire g29141;
wire g24641;
wire g34928;
wire g21948;
wire g18192;
wire g32516;
wire g13566;
wire g25287;
wire g34401;
wire g30510;
wire g33732;
wire g17757;
wire g24184;
wire g20631;
wire g16204;
wire g17761;
wire g18428;
wire II14482;
wire g11527;
wire II15617;
wire g32630;
wire g32659;
wire II16357;
wire g16737;
wire g29196;
wire g27380;
wire g18782;
wire g13974;
wire g14854;
wire g24918;
wire g22330;
wire g22181;
wire II24008;
wire g32184;
wire g12155;
wire g7532;
wire g17615;
wire g25902;
wire g9413;
wire g14383;
wire g20533;
wire g31224;
wire g16967;
wire g9661;
wire g22223;
wire g12880;
wire g28216;
wire g11413;
wire g23543;
wire g23714;
wire g21729;
wire g20566;
wire g26234;
wire g17429;
wire g7394;
wire g26652;
wire g11973;
wire g34883;
wire II12577;
wire g21556;
wire g33597;
wire g32191;
wire g28622;
wire g26933;
wire g24400;
wire g27431;
wire g9995;
wire II16438;
wire g21053;
wire g25027;
wire g30390;
wire II13892;
wire g18125;
wire g28853;
wire g17783;
wire II31985;
wire g19919;
wire g26365;
wire g11934;
wire g14238;
wire g18588;
wire g27983;
wire g23532;
wire g14540;
wire g34257;
wire g12538;
wire g20668;
wire g32617;
wire g9542;
wire g13189;
wire g33075;
wire g12047;
wire g24049;
wire g8388;
wire g25121;
wire g33685;
wire gbuf101;
wire g24666;
wire g13530;
wire II31152;
wire g23448;
wire g34416;
wire II18888;
wire g25237;
wire g21979;
wire g21832;
wire g32558;
wire g34973;
wire g25618;
wire g32210;
wire g24710;
wire II17495;
wire g11958;
wire II15831;
wire g7502;
wire g29986;
wire g11949;
wire g8714;
wire g27097;
wire g33017;
wire g13765;
wire g11435;
wire g34408;
wire g24293;
wire g21340;
wire g31480;
wire g21953;
wire g18117;
wire g18325;
wire g28082;
wire g27411;
wire g11404;
wire II22931;
wire g14564;
wire g25665;
wire g22538;
wire g31312;
wire g34970;
wire g17625;
wire g12075;
wire II18086;
wire g20060;
wire g26340;
wire g28166;
wire g29280;
wire g13529;
wire g15755;
wire g8895;
wire g10520;
wire gbuf99;
wire g33063;
wire g15063;
wire g28244;
wire g33293;
wire g19354;
wire g22698;
wire g26941;
wire g23922;
wire g17716;
wire g25766;
wire g24263;
wire g21887;
wire g27089;
wire g11999;
wire g32689;
wire g26025;
wire g16308;
wire g27312;
wire g23309;
wire II22096;
wire g20070;
wire g18272;
wire g26681;
wire g21377;
wire g22985;
wire g23108;
wire g7374;
wire g26896;
wire g21293;
wire g17366;
wire g19931;
wire g28574;
wire g28334;
wire g24779;
wire g13923;
wire II14249;
wire g18633;
wire g15807;
wire g34394;
wire g20069;
wire g32680;
wire g18221;
wire g23749;
wire g29325;
wire II24439;
wire g25650;
wire g32157;
wire g6854;
wire g31806;
wire g22004;
wire g22669;
wire g14655;
wire g32145;
wire g18618;
wire g28748;
wire g30089;
wire g30565;
wire g25505;
wire g11380;
wire g7153;
wire g34142;
wire g19546;
wire g34088;
wire g26510;
wire g24590;
wire g24676;
wire g21904;
wire g15152;
wire g18667;
wire II17852;
wire g30315;
wire g23847;
wire g12405;
wire g11967;
wire II30124;
wire g6927;
wire g10359;
wire g22144;
wire g25144;
wire g12314;
wire g15756;
wire II18620;
wire II21042;
wire II29936;
wire g15116;
wire g19539;
wire g25743;
wire gbuf67;
wire II15041;
wire g6850;
wire g34634;
wire g24460;
wire g7150;
wire g32627;
wire g13742;
wire g27365;
wire g32501;
wire II31619;
wire g29759;
wire g12831;
wire gbuf11;
wire g24104;
wire g33461;
wire g32310;
wire g18753;
wire g14506;
wire g27215;
wire g7361;
wire g21817;
wire g20276;
wire g18491;
wire g19771;
wire g33054;
wire II17956;
wire g17742;
wire g9153;
wire g22342;
wire g29689;
wire g17384;
wire g24864;
wire g12148;
wire g29382;
wire g23046;
wire g29602;
wire g20622;
wire g21922;
wire g22935;
wire g12415;
wire g19428;
wire g29860;
wire g24425;
wire g27017;
wire g24638;
wire g25678;
wire g29994;
wire II14508;
wire g26259;
wire g32632;
wire II17118;
wire g32980;
wire g30137;
wire g29905;
wire g16259;
wire g22061;
wire g26895;
wire g19660;
wire g29587;
wire g14122;
wire g34713;
wire g33552;
wire g16211;
wire gbuf31;
wire g19914;
wire g16644;
wire g23153;
wire g14739;
wire g34486;
wire g12760;
wire II16747;
wire g20771;
wire g27742;
wire g31487;
wire g12093;
wire g18107;
wire g25915;
wire g20050;
wire g28636;
wire II30262;
wire g34135;
wire g9282;
wire g28279;
wire g12417;
wire g28536;
wire g27289;
wire g18746;
wire g24875;
wire g10261;
wire g27355;
wire g18526;
wire g19564;
wire g29548;
wire g29966;
wire g24688;
wire g18184;
wire g9083;
wire g14169;
wire g21422;
wire g18660;
wire g33016;
wire g24415;
wire g18208;
wire g32477;
wire g15108;
wire g31788;
wire g27677;
wire g18977;
wire g29329;
wire g10899;
wire g29840;
wire g19274;
wire II31127;
wire g25980;
wire g32906;
wire II32806;
wire g13873;
wire g11914;
wire g19500;
wire g20502;
wire g33560;
wire II22153;
wire II22124;
wire g10922;
wire gbuf112;
wire g7404;
wire g19683;
wire g23300;
wire g28669;
wire g15082;
wire II22944;
wire g13055;
wire g23421;
wire g33546;
wire g31066;
wire g9891;
wire g15614;
wire II21189;
wire g17507;
wire g29529;
wire g29535;
wire II17488;
wire g10014;
wire g22544;
wire g8476;
wire g34474;
wire g18471;
wire g17393;
wire II26799;
wire g29607;
wire g29871;
wire g26484;
wire g31007;
wire g19751;
wire g31822;
wire g30430;
wire g11397;
wire g23505;
wire g31880;
wire g13464;
wire g16580;
wire g13632;
wire g31986;
wire g20738;
wire g9591;
wire g19998;
wire g18576;
wire g11591;
wire g19688;
wire g20679;
wire g12863;
wire g24055;
wire II15727;
wire g24644;
wire g13600;
wire g32328;
wire g28962;
wire II18912;
wire g25002;
wire g29264;
wire II13206;
wire g16770;
wire g34636;
wire g30919;
wire g32783;
wire g8406;
wire g21789;
wire g34116;
wire g18874;
wire II25028;
wire g32413;
wire g34515;
wire II22302;
wire g23958;
wire g10289;
wire g12464;
wire II13401;
wire g33918;
wire g15744;
wire g24507;
wire g32889;
wire g18952;
wire g15784;
wire g22182;
wire g30539;
wire g20145;
wire g25184;
wire g13820;
wire g17411;
wire g11793;
wire g31912;
wire g34987;
wire II12783;
wire g33253;
wire g25179;
wire g12996;
wire II22131;
wire g24021;
wire g32873;
wire g31319;
wire g30929;
wire g31517;
wire II31281;
wire g27717;
wire II16120;
wire g18832;
wire g28265;
wire g9823;
wire g8092;
wire g30071;
wire g9762;
wire g23972;
wire g7898;
wire g22307;
wire g10884;
wire g20554;
wire g25108;
wire g21996;
wire g30197;
wire g18511;
wire g10556;
wire g10815;
wire g30935;
wire g24835;
wire g8958;
wire g13975;
wire g32374;
wire g14036;
wire g33722;
wire g16512;
wire g24212;
wire g23949;
wire g31479;
wire g21397;
wire g18733;
wire g14215;
wire g13958;
wire g9905;
wire g13729;
wire g14107;
wire g13120;
wire II19843;
wire g9805;
wire g34775;
wire II24616;
wire II28128;
wire g19767;
wire g34199;
wire g31020;
wire g23024;
wire g30455;
wire g18246;
wire g18805;
wire g33925;
wire g11019;
wire g18586;
wire g27113;
wire g21835;
wire g29837;
wire g11225;
wire II13317;
wire g29131;
wire g29899;
wire g21037;
wire II18810;
wire g28543;
wire g20324;
wire g25954;
wire g30461;
wire g7948;
wire gbuf151;
wire g8763;
wire g29892;
wire g11826;
wire g18559;
wire g19780;
wire g30064;
wire g22992;
wire g24457;
wire g27096;
wire g10372;
wire II13847;
wire g16236;
wire g6971;
wire g18620;
wire g22125;
wire g6868;
wire g26758;
wire g34560;
wire g32593;
wire g15881;
wire g17772;
wire g28121;
wire g8606;
wire g23031;
wire g16617;
wire g32106;
wire g18563;
wire g8441;
wire g19712;
wire g9654;
wire g9752;
wire II19762;
wire g22633;
wire g14362;
wire g25326;
wire g9557;
wire II17999;
wire II12887;
wire g34877;
wire g25831;
wire g10620;
wire g19693;
wire g17155;
wire g13006;
wire g26841;
wire g34730;
wire g7527;
wire g18237;
wire g20913;
wire g31937;
wire II27503;
wire g23483;
wire g18826;
wire g24967;
wire II25562;
wire g25971;
wire g31758;
wire g24200;
wire g30546;
wire g16640;
wire II19789;
wire g33543;
wire g24627;
wire g33872;
wire g7308;
wire g25340;
wire g32488;
wire g19960;
wire g30922;
wire g13824;
wire g21745;
wire g30143;
wire g14612;
wire II23950;
wire g25009;
wire g18132;
wire g24163;
wire II14517;
wire g34684;
wire g13730;
wire g18147;
wire II20951;
wire g17056;
wire g27549;
wire g19386;
wire g23345;
wire g22762;
wire g9853;
wire II12858;
wire g22496;
wire g14585;
wire g24313;
wire II15070;
wire g32642;
wire g8974;
wire g8989;
wire g14178;
wire g26105;
wire g31837;
wire g32177;
wire g24136;
wire g33635;
wire g22112;
wire g24209;
wire g20712;
wire g15096;
wire g27536;
wire g27390;
wire g32716;
wire g25686;
wire g9861;
wire g25385;
wire g34994;
wire II23585;
wire g33311;
wire g22847;
wire g20604;
wire g21895;
wire g32481;
wire g32728;
wire g13501;
wire g10602;
wire g32196;
wire g24284;
wire g28591;
wire g30118;
wire g21370;
wire g24818;
wire g14417;
wire g20373;
wire g27822;
wire g26870;
wire g21386;
wire II12097;
wire g18284;
wire g17224;
wire g30048;
wire g11940;
wire g27226;
wire g10801;
wire II12252;
wire g32261;
wire g11519;
wire g14316;
wire g27769;
wire g21652;
wire g25473;
wire g34094;
wire g20716;
wire g25869;
wire g8160;
wire g34501;
wire g30524;
wire g7993;
wire g9477;
wire g22016;
wire g32594;
wire g29297;
wire g9932;
wire g30734;
wire g24813;
wire g34438;
wire g34574;
wire g20039;
wire II15536;
wire g14179;
wire g19853;
wire g25839;
wire g22753;
wire g19453;
wire g25945;
wire g23138;
wire g34178;
wire g28057;
wire II13010;
wire g28610;
wire g31792;
wire g31905;
wire g34247;
wire g26204;
wire g33772;
wire g28050;
wire g6996;
wire g19791;
wire g29606;
wire g25263;
wire g19373;
wire g21179;
wire g14645;
wire g16486;
wire g12744;
wire g34967;
wire g28115;
wire g8216;
wire g12232;
wire g24142;
wire g22883;
wire g13712;
wire g23152;
wire g30060;
wire g24008;
wire g20540;
wire g16884;
wire g19372;
wire g32606;
wire g30134;
wire g23434;
wire g32844;
wire g29306;
wire g19527;
wire g10655;
wire g34521;
wire g18421;
wire II16779;
wire g23471;
wire g28942;
wire g21415;
wire g34688;
wire g33843;
wire g27452;
wire g26290;
wire g13834;
wire g12284;
wire g13124;
wire g17650;
wire g20581;
wire g15679;
wire g19578;
wire g33137;
wire g18818;
wire g28070;
wire g23828;
wire g26879;
wire g27231;
wire g33159;
wire II26094;
wire g32123;
wire II18411;
wire g8700;
wire II25327;
wire g33961;
wire g15089;
wire g25247;
wire g23131;
wire II12103;
wire g21791;
wire II26948;
wire g8334;
wire g29990;
wire g25674;
wire g25535;
wire II16168;
wire g24749;
wire g16958;
wire g20636;
wire g27651;
wire g24554;
wire g33680;
wire g13142;
wire II31147;
wire g12512;
wire g15008;
wire g15426;
wire g18801;
wire g12858;
wire II33176;
wire g7092;
wire II32173;
wire g17662;
wire g19656;
wire g23943;
wire g23415;
wire g24476;
wire g23786;
wire g7380;
wire g29372;
wire II32950;
wire g33441;
wire g24079;
wire g27050;
wire g28226;
wire g27461;
wire g8154;
wire g15161;
wire g8971;
wire g33033;
wire g25218;
wire g12402;
wire g31777;
wire g18211;
wire g30195;
wire g16272;
wire g28751;
wire g15748;
wire g34378;
wire g25514;
wire II18280;
wire g11640;
wire II25095;
wire g27573;
wire g7387;
wire g9827;
wire II20321;
wire g20665;
wire g7953;
wire g20201;
wire g29979;
wire g31469;
wire g28331;
wire g10040;
wire g24515;
wire g34868;
wire g30181;
wire II16498;
wire gbuf62;
wire g19779;
wire II32791;
wire g12356;
wire g8913;
wire g21828;
wire g24499;
wire g14741;
wire g22837;
wire II22444;
wire g31919;
wire g30202;
wire g20902;
wire g26850;
wire g15821;
wire g32118;
wire g20081;
wire g8492;
wire g16305;
wire II22275;
wire g18670;
wire g13745;
wire g10542;
wire g22722;
wire g34158;
wire g28148;
wire g10335;
wire g15861;
wire g23376;
wire g34659;
wire II14993;
wire g28201;
wire g32360;
wire g25723;
wire g28296;
wire g20783;
wire g21809;
wire g11110;
wire g23565;
wire g20501;
wire II12896;
wire g24001;
wire g25272;
wire g23748;
wire g18814;
wire g21225;
wire g25155;
wire g24205;
wire II14537;
wire g12522;
wire g28135;
wire g21867;
wire g28307;
wire g28043;
wire g28096;
wire II22873;
wire g18910;
wire g33979;
wire g32334;
wire g22055;
wire II14350;
wire g34013;
wire g18654;
wire g21337;
wire g33468;
wire g34464;
wire g21899;
wire II32461;
wire g21307;
wire g32809;
wire g14251;
wire g31276;
wire g30291;
wire g27543;
wire g30298;
wire g23396;
wire g34451;
wire g12431;
wire g14706;
wire g11804;
wire g22996;
wire g23419;
wire g24039;
wire g34153;
wire g28799;
wire g33638;
wire g19144;
wire g16448;
wire g14233;
wire g33425;
wire g17217;
wire g29950;
wire II21993;
wire g27591;
wire g13968;
wire g33130;
wire II25779;
wire g14793;
wire g34595;
wire II22892;
wire II14192;
wire g18540;
wire g18266;
wire g16279;
wire g21911;
wire g27968;
wire g24194;
wire g32649;
wire g32863;
wire g23016;
wire g12002;
wire g26241;
wire II31694;
wire g24535;
wire g27316;
wire g28045;
wire g15131;
wire g24251;
wire g11083;
wire g16245;
wire g28184;
wire g13091;
wire g11652;
wire g18379;
wire g33472;
wire II24694;
wire g33876;
wire g11043;
wire g10199;
wire g13411;
wire g29105;
wire II33037;
wire g25637;
wire g23290;
wire g29247;
wire g18350;
wire g33893;
wire g10497;
wire g14568;
wire II14735;
wire g33415;
wire g23495;
wire g30606;
wire g16870;
wire g20174;
wire g26751;
wire g19855;
wire II32305;
wire g27290;
wire g29173;
wire g31760;
wire g31122;
wire g10705;
wire g24721;
wire g26304;
wire g11122;
wire g16970;
wire g23774;
wire g24064;
wire g34998;
wire II22844;
wire g8016;
wire g18392;
wire g11035;
wire g21183;
wire g7582;
wire g19612;
wire g26938;
wire II27735;
wire g14392;
wire g16843;
wire g25654;
wire g14187;
wire g8691;
wire g12323;
wire II25598;
wire g32623;
wire g28346;
wire II14957;
wire g21738;
wire g21773;
wire g17613;
wire g31307;
wire g30425;
wire II18252;
wire g30996;
wire g20609;
wire g12374;
wire g10035;
wire g23478;
wire g29240;
wire g21752;
wire g9333;
wire g28448;
wire II33291;
wire g14735;
wire g34630;
wire g23878;
wire g27735;
wire g8864;
wire II27954;
wire g17135;
wire g34931;
wire g18724;
wire g21868;
wire g29812;
wire g29273;
wire II18148;
wire g7964;
wire g10511;
wire g32927;
wire g34787;
wire g18256;
wire g31878;
wire g22515;
wire g21062;
wire g8347;
wire g25148;
wire g32238;
wire g20600;
wire g29909;
wire II16479;
wire g22198;
wire g27186;
wire g17669;
wire g29330;
wire g18926;
wire g33126;
wire g8155;
wire gbuf57;
wire g26733;
wire g9162;
wire g18455;
wire g20208;
wire g7187;
wire g10323;
wire g17175;
wire g13944;
wire gbuf1;
wire g31303;
wire g24259;
wire g11235;
wire g9258;
wire II26705;
wire g34382;
wire g7851;
wire g21861;
wire g32354;
wire II28576;
wire g12806;
wire g33489;
wire g10403;
wire g25816;
wire g33239;
wire g34909;
wire II15168;
wire g16292;
wire g21206;
wire g26054;
wire g28824;
wire g22115;
wire g28183;
wire II15717;
wire g30497;
wire g8135;
wire g20380;
wire g19905;
wire g28248;
wire g14591;
wire g32656;
wire g13336;
wire g31129;
wire g34723;
wire II15223;
wire g17752;
wire g33104;
wire g25614;
wire g29930;
wire g28639;
wire g34376;
wire g33271;
wire g31274;
wire g9917;
wire g23836;
wire g28632;
wire g27331;
wire g13539;
wire g26779;
wire g24012;
wire II33075;
wire g33052;
wire g27416;
wire II14381;
wire g28776;
wire g33924;
wire g13437;
wire II31036;
wire g33983;
wire g29146;
wire g34717;
wire g19626;
wire g32247;
wire g7134;
wire g30164;
wire g26808;
wire g29782;
wire g28482;
wire II17104;
wire g28241;
wire g6814;
wire II17249;
wire II27579;
wire g26359;
wire II18536;
wire g18646;
wire g20590;
wire g29115;
wire g20181;
wire g20547;
wire g17726;
wire g11026;
wire g24394;
wire II31246;
wire g18813;
wire g7280;
wire g17675;
wire g32317;
wire g24825;
wire g33883;
wire g18261;
wire g7261;
wire g32945;
wire g25090;
wire g28410;
wire g32653;
wire g34531;
wire g20544;
wire g30057;
wire g33023;
wire g25593;
wire II32878;
wire g21782;
wire g13034;
wire g26714;
wire g33798;
wire g14547;
wire g30281;
wire g17713;
wire g10085;
wire g9978;
wire g10674;
wire g32661;
wire g24330;
wire II12336;
wire g12695;
wire II21006;
wire g29311;
wire II23119;
wire g22710;
wire g30069;
wire II11688;
wire g7660;
wire g19543;
wire g19401;
wire g28617;
wire g12211;
wire II18504;
wire g27293;
wire g9581;
wire g24703;
wire g27152;
wire II30641;
wire g15781;
wire g26271;
wire II14365;
wire g17498;
wire g24527;
wire g24266;
wire g32414;
wire g25565;
wire g9975;
wire g18163;
wire g34293;
wire g32566;
wire g17732;
wire g30207;
wire g16284;
wire g33838;
wire II15254;
wire g24363;
wire g12866;
wire g31815;
wire g28404;
wire g9490;
wire g18204;
wire g18444;
wire g22316;
wire g13782;
wire g16316;
wire g27385;
wire g27270;
wire g30346;
wire g26153;
wire g26388;
wire II24041;
wire g29636;
wire g23983;
wire g15788;
wire g24908;
wire g32168;
wire g18332;
wire g11815;
wire g25786;
wire II20647;
wire II29304;
wire g20739;
wire g32462;
wire g18793;
wire g7715;
wire g29797;
wire g23247;
wire g11205;
wire g22680;
wire g21429;
wire g25038;
wire g12887;
wire g26922;
wire g34004;
wire g23387;
wire g28154;
wire g9103;
wire II25846;
wire g32797;
wire g23007;
wire g32282;
wire g10614;
wire g28736;
wire g14771;
wire g9226;
wire II13183;
wire g25112;
wire g8871;
wire g29337;
wire II18891;
wire g16158;
wire g25935;
wire II14267;
wire g27139;
wire g23810;
wire g34113;
wire g24958;
wire g16577;
wire g30450;
wire g7004;
wire g27037;
wire II25613;
wire g15509;
wire g34494;
wire g33141;
wire g25804;
wire g23648;
wire g26218;
wire g22521;
wire g27026;
wire g27580;
wire g12906;
wire g13278;
wire g28959;
wire g21761;
wire g14821;
wire g32588;
wire g15055;
wire g22585;
wire g12780;
wire g11023;
wire g29367;
wire g14275;
wire g28884;
wire g10862;
wire g32499;
wire g23890;
wire g27370;
wire g26288;
wire g30405;
wire g34941;
wire g7922;
wire II12930;
wire II31459;
wire g28314;
wire g22648;
wire g26630;
wire g33490;
wire g11858;
wire g33956;
wire g34220;
wire g13707;
wire g31977;
wire g32934;
wire g32790;
wire g13871;
wire g21938;
wire g29046;
wire II31839;
wire g8743;
wire II26337;
wire g19619;
wire II21033;
wire g11674;
wire g16662;
wire g17595;
wire g18681;
wire II23390;
wire g16538;
wire g12026;
wire g29201;
wire g9070;
wire g10429;
wire g33603;
wire g13067;
wire II32441;
wire g7258;
wire g11395;
wire g25760;
wire g9959;
wire g32835;
wire g32967;
wire g32143;
wire II15002;
wire g27507;
wire II23918;
wire g9528;
wire g22043;
wire g8955;
wire g31889;
wire g24724;
wire g29592;
wire g23228;
wire g25697;
wire II14198;
wire g22094;
wire g34649;
wire g33148;
wire II31346;
wire g20384;
wire g18344;
wire g9899;
wire g32323;
wire g31657;
wire g17307;
wire g30016;
wire g29841;
wire II24524;
wire g32084;
wire g8182;
wire g10390;
wire g12891;
wire g27333;
wire g27030;
wire g30280;
wire g20560;
wire g11129;
wire II31486;
wire g26910;
wire g10830;
wire g24325;
wire g23510;
wire g19737;
wire g13911;
wire II33282;
wire g29630;
wire g9671;
wire g31257;
wire II33279;
wire g34691;
wire g24302;
wire g19368;
wire g33349;
wire g11608;
wire g14198;
wire g20267;
wire g19412;
wire g13050;
wire g12192;
wire g25963;
wire g26745;
wire g28987;
wire g17680;
wire g29748;
wire g24518;
wire g34799;
wire g13082;
wire g25522;
wire g33098;
wire g7788;
wire g9491;
wire g25991;
wire g34312;
wire g21734;
wire g29289;
wire g7738;
wire g26205;
wire g10608;
wire g33246;
wire g16623;
wire g32470;
wire g28562;
wire g19520;
wire g9985;
wire g22687;
wire g23333;
wire g34341;
wire g10073;
wire g19635;
wire g33689;
wire g27148;
wire g27286;
wire g29813;
wire g18179;
wire g18424;
wire II31564;
wire II31616;
wire g13016;
wire g20096;
wire g22400;
wire g30114;
wire g11849;
wire g32056;
wire g33565;
wire gbuf45;
wire g21247;
wire g13087;
wire g16677;
wire g29224;
wire g30085;
wire g31805;
wire II24675;
wire g9077;
wire II25909;
wire g9999;
wire g10418;
wire g21351;
wire g28648;
wire g32550;
wire II20461;
wire g14571;
wire II12935;
wire g31326;
wire g11987;
wire g23969;
wire g19949;
wire g15027;
wire II26682;
wire g20662;
wire g20597;
wire g29693;
wire g22662;
wire g32202;
wire g29626;
wire g23880;
wire g7340;
wire g31322;
wire g9247;
wire g14625;
wire II14885;
wire g10552;
wire g25719;
wire g26391;
wire II33179;
wire g12849;
wire g32741;
wire g23904;
wire g27160;
wire g27130;
wire g26519;
wire g17528;
wire g14556;
wire g13106;
wire g33522;
wire g28419;
wire g21358;
wire II13384;
wire g19537;
wire g27103;
wire gbuf38;
wire g18456;
wire g14008;
wire g23963;
wire g34442;
wire g21603;
wire g27886;
wire g29513;
wire g25906;
wire II12261;
wire g25704;
wire g8458;
wire g31992;
wire g28283;
wire II18408;
wire g31966;
wire g33821;
wire g32702;
wire g32988;
wire g24029;
wire g34352;
wire g14338;
wire g34049;
wire g15653;
wire g26955;
wire g15731;
wire g18605;
wire g34412;
wire g22075;
wire g13807;
wire gbuf40;
wire g7040;
wire g10916;
wire II18009;
wire g34856;
wire g33755;
wire II12270;
wire g33536;
wire g18482;
wire g20613;
wire g24409;
wire g12882;
wire II22539;
wire g13129;
wire g34735;
wire gbuf29;
wire g33648;
wire g34419;
wire g22218;
wire g33942;
wire g21256;
wire g9771;
wire g21659;
wire g13918;
wire II12666;
wire g29790;
wire g20680;
wire g25479;
wire g15738;
wire g33711;
wire g20874;
wire g16634;
wire g18311;
wire g29767;
wire g12170;
wire g28525;
wire g24575;
wire g15959;
wire g27649;
wire II23149;
wire g9731;
wire g28322;
wire gbuf22;
wire g18167;
wire g10360;
wire g23279;
wire g32554;
wire g18675;
wire g33373;
wire g28071;
wire g11889;
wire g12924;
wire g18476;
wire g34388;
wire II12903;
wire g28104;
wire g14062;
wire g30041;
wire II31117;
wire g18771;
wire g14496;
wire g18729;
wire g27502;
wire g8553;
wire g18945;
wire g31237;
wire II12842;
wire II31686;
wire II15053;
wire g17247;
wire II31858;
wire g30596;
wire g22151;
wire g14165;
wire g34760;
wire g23729;
wire g30372;
wire g22166;
wire g28376;
wire g32042;
wire g28786;
wire g34397;
wire g28725;
wire g21875;
wire g31169;
wire g19516;
wire g6978;
wire g14943;
wire g27668;
wire II25380;
wire g32587;
wire g26823;
wire g18504;
wire g12790;
wire g23919;
wire g30149;
wire g28062;
wire II19831;
wire g14442;
wire g13568;
wire g10389;
wire g31315;
wire g29487;
wire g28584;
wire g16177;
wire g28573;
wire II14187;
wire g7812;
wire g7827;
wire g25380;
wire g30248;
wire g11498;
wire g21712;
wire II25399;
wire g24648;
wire g19074;
wire g24335;
wire g19595;
wire g26604;
wire g22832;
wire g12950;
wire g27823;
wire g26883;
wire g23242;
wire g20027;
wire g27519;
wire g10047;
wire g33627;
wire g9050;
wire g24820;
wire g34626;
wire g6953;
wire g32721;
wire g25649;
wire g28353;
wire g34083;
wire g14344;
wire g13393;
wire g31540;
wire g23050;
wire g26884;
wire g34999;
wire g13699;
wire g29769;
wire g27533;
wire g32051;
wire II18337;
wire II15342;
wire g18622;
wire g19494;
wire g25713;
wire g27703;
wire g32774;
wire g34421;
wire II21115;
wire II31301;
wire g12822;
wire g19742;
wire g30363;
wire g24067;
wire g30354;
wire g7209;
wire g29475;
wire g31844;
wire g28515;
wire g11566;
wire g10185;
wire g24056;
wire g11426;
wire g25033;
wire g34227;
wire g24586;
wire g13680;
wire g13511;
wire g28253;
wire g30125;
wire g33387;
wire g25968;
wire g31247;
wire II22769;
wire g23216;
wire g28399;
wire II18398;
wire g25059;
wire g31123;
wire g28729;
wire g12977;
wire g15126;
wire g7074;
wire II12089;
wire g26862;
wire g27421;
wire g19427;
wire g16525;
wire g18443;
wire g11675;
wire g16645;
wire g26891;
wire g27633;
wire g12220;
wire g21308;
wire g33514;
wire g31209;
wire g34669;
wire II15003;
wire g30467;
wire g33849;
wire g7028;
wire g12351;
wire II12183;
wire g26125;
wire g13756;
wire g26348;
wire g26903;
wire g15792;
wire g26020;
wire g14408;
wire g19492;
wire II14510;
wire g32019;
wire g34057;
wire g12218;
wire g32461;
wire g19760;
wire g27253;
wire g28550;
wire g30266;
wire g32468;
wire g10119;
wire g11832;
wire II21744;
wire g16429;
wire g7196;
wire g23504;
wire g32492;
wire II18829;
wire II18051;
wire g23274;
wire g11276;
wire g34614;
wire g24471;
wire II15122;
wire g34666;
wire g33265;
wire g13295;
wire g21892;
wire II12767;
wire g24236;
wire II32467;
wire g30100;
wire g15729;
wire g10034;
wire g32369;
wire g26873;
wire g13044;
wire g9511;
wire g15141;
wire g22228;
wire g16475;
wire g19881;
wire g28860;
wire g7907;
wire g34745;
wire g11313;
wire g8457;
wire g16609;
wire g34103;
wire II25591;
wire g30454;
wire g30672;
wire g19396;
wire g21841;
wire g33454;
wire g28670;
wire II19772;
wire g27770;
wire g12166;
wire g14682;
wire g7498;
wire g13990;
wire g27542;
wire g15813;
wire g34894;
wire g15075;
wire g29290;
wire g24674;
wire II27742;
wire g7675;
wire II24597;
wire g25107;
wire g16223;
wire g22029;
wire g19652;
wire g13627;
wire g6819;
wire g29157;
wire g27499;
wire g13595;
wire g33262;
wire g25088;
wire g26543;
wire II13750;
wire g25524;
wire g23869;
wire II14866;
wire g9900;
wire g16075;
wire g33529;
wire g7892;
wire g25130;
wire g28686;
wire g33986;
wire g31948;
wire II11860;
wire g17317;
wire g7026;
wire g30206;
wire g18227;
wire g18601;
wire g29910;
wire g21968;
wire g21267;
wire g25672;
wire g33266;
wire g18240;
wire g20529;
wire g33382;
wire g20870;
wire g32712;
wire II12128;
wire g28268;
wire g19757;
wire gbuf105;
wire g12667;
wire g30077;
wire g27118;
wire g14971;
wire g21840;
wire g24450;
wire g18736;
wire g29268;
wire g15780;
wire II20355;
wire g20198;
wire g33487;
wire g26338;
wire g28009;
wire g24090;
wire II31469;
wire g9569;
wire g31872;
wire g31208;
wire gbuf93;
wire g20995;
wire g19486;
wire g29897;
wire gbuf117;
wire g17324;
wire g28634;
wire g23687;
wire g25525;
wire g24760;
wire g32540;
wire g28243;
wire g11238;
wire g27766;
wire g16226;
wire g21916;
wire g13806;
wire g15099;
wire g26400;
wire II31844;
wire g33227;
wire g30017;
wire g34586;
wire g10585;
wire g11467;
wire g16517;
wire II13392;
wire g11845;
wire g32959;
wire II12787;
wire g18111;
wire g15787;
wire g33556;
wire II19704;
wire II27552;
wire g18821;
wire g14598;
wire II17121;
wire II32617;
wire g15842;
wire g15798;
wire g28546;
wire g23251;
wire g24264;
wire g26990;
wire g31848;
wire g27974;
wire g29582;
wire g29107;
wire g28372;
wire g33512;
wire g18830;
wire g31311;
wire g27526;
wire g12870;
wire g32650;
wire g15811;
wire gbuf75;
wire g21189;
wire g10550;
wire g15106;
wire g24222;
wire g18093;
wire g21702;
wire g14669;
wire g34770;
wire II12355;
wire g22018;
wire g34055;
wire g8119;
wire g33021;
wire II21297;
wire g24791;
wire g32599;
wire g6958;
wire g14297;
wire g31867;
wire g27545;
wire g8170;
wire g28694;
wire g32990;
wire g29982;
wire g27383;
wire g12918;
wire g27654;
wire g23348;
wire g31249;
wire II30745;
wire g29834;
wire g10417;
wire g10349;
wire g18118;
wire II12877;
wire g28930;
wire II31796;
wire g24684;
wire g22148;
wire II12534;
wire g14358;
wire g21750;
wire g30513;
wire g30520;
wire g16690;
wire g9594;
wire g7064;
wire g18401;
wire g33331;
wire g13032;
wire g12065;
wire g17766;
wire g34603;
wire g34950;
wire g31375;
wire g13884;
wire g13294;
wire g16807;
wire II17131;
wire II22936;
wire g31989;
wire g13526;
wire g14569;
wire g18704;
wire II15205;
wire II29717;
wire g6837;
wire g21276;
wire g20134;
wire g20601;
wire g8075;
wire g31485;
wire g24338;
wire g14061;
wire g25923;
wire g33174;
wire g20078;
wire g25149;
wire g29495;
wire g6923;
wire g33502;
wire II31116;
wire g24776;
wire g15090;
wire g30583;
wire g25004;
wire g13248;
wire g27676;
wire g30730;
wire g33374;
wire g6994;
wire g32522;
wire g7450;
wire g34443;
wire g23306;
wire g27999;
wire g23088;
wire g21297;
wire g32181;
wire g26769;
wire g17619;
wire g32739;
wire g34737;
wire g21882;
wire g23453;
wire g31144;
wire II12199;
wire g7158;
wire g21417;
wire g8757;
wire g30062;
wire g30007;
wire g12196;
wire g14582;
wire g16238;
wire g21285;
wire g22833;
wire g26849;
wire g34792;
wire g28533;
wire g25648;
wire g18638;
wire g19857;
wire g18529;
wire II19012;
wire g33724;
wire g28471;
wire g24099;
wire g32655;
wire g23195;
wire g23795;
wire g25023;
wire g14412;
wire g11514;
wire g19488;
wire g34197;
wire g25180;
wire g18448;
wire g29352;
wire g6985;
wire g16077;
wire II21969;
wire g13076;
wire g7936;
wire g16194;
wire g20676;
wire g21057;
wire g7991;
wire g16636;
wire g26752;
wire II28458;
wire g10606;
wire g22013;
wire g7514;
wire g20054;
wire II29302;
wire g34098;
wire g29521;
wire g18585;
wire g32590;
wire g28086;
wire g17508;
wire g10828;
wire g20035;
wire g19387;
wire g8228;
wire g32952;
wire g32738;
wire g32926;
wire g11977;
wire g34711;
wire g28103;
wire II24396;
wire g30043;
wire g27094;
wire g20628;
wire g33065;
wire II14650;
wire g29907;
wire II12808;
wire g11357;
wire II28241;
wire II13498;
wire g18142;
wire g14206;
wire g30044;
wire g9485;
wire g25682;
wire g16123;
wire g8766;
wire g21957;
wire g34944;
wire gbuf46;
wire g28320;
wire g18306;
wire g28527;
wire g20327;
wire g25916;
wire g26628;
wire g33423;
wire g32484;
wire g11993;
wire II13802;
wire g29890;
wire g34141;
wire g30927;
wire g31804;
wire g26392;
wire g7219;
wire g22937;
wire g27162;
wire g31930;
wire g20129;
wire II29277;
wire g28743;
wire g30310;
wire g18742;
wire g34405;
wire g27366;
wire g23498;
wire g11401;
wire g28197;
wire g34812;
wire g30610;
wire II12288;
wire g20565;
wire g9072;
wire II11691;
wire g30025;
wire g33050;
wire g22030;
wire g24297;
wire g25953;
wire g18176;
wire g11469;
wire g23423;
wire g32538;
wire g22057;
wire g19677;
wire g28140;
wire g26926;
wire g22025;
wire g19673;
wire g21813;
wire g24107;
wire g18153;
wire g27765;
wire g8324;
wire g28484;
wire g27278;
wire II22400;
wire g21920;
wire g34487;
wire g19670;
wire g14820;
wire g22857;
wire g18608;
wire g9203;
wire g11833;
wire g30182;
wire II20985;
wire g28700;
wire g7222;
wire II13442;
wire g19534;
wire g22720;
wire g34411;
wire g19407;
wire g34472;
wire g24537;
wire g24082;
wire g22665;
wire g24100;
wire g25746;
wire g25089;
wire g32472;
wire g21560;
wire g27051;
wire g31810;
wire g7680;
wire g8479;
wire g33566;
wire g18484;
wire g24731;
wire g32207;
wire g25643;
wire II32440;
wire g30124;
wire g25341;
wire g31896;
wire II26972;
wire g29035;
wire g21927;
wire g29507;
wire g20161;
wire II18479;
wire II27941;
wire II15382;
wire g21331;
wire g11430;
wire g9935;
wire g30370;
wire II33149;
wire g22974;
wire g10925;
wire g22534;
wire g14627;
wire II27570;
wire g23769;
wire II14827;
wire g34736;
wire g23511;
wire g32357;
wire g14659;
wire g28118;
wire g27833;
wire g28563;
wire g21851;
wire g33913;
wire g34433;
wire g7379;
wire g10609;
wire g17327;
wire g30936;
wire g8741;
wire g18542;
wire g17432;
wire g16633;
wire g13476;
wire g23895;
wire g14191;
wire g24133;
wire g28047;
wire g10578;
wire g16876;
wire g18310;
wire g14791;
wire g27218;
wire g27058;
wire g29527;
wire g33330;
wire II18803;
wire g24861;
wire g18494;
wire g10831;
wire g11389;
wire g26598;
wire g33813;
wire g14211;
wire g15149;
wire II27385;
wire g14726;
wire g18664;
wire g20038;
wire g23104;
wire g29855;
wire g7328;
wire g30234;
wire g29702;
wire g8302;
wire g23930;
wire g34146;
wire g17648;
wire g32640;
wire g33591;
wire g15611;
wire g27374;
wire g34379;
wire g7424;
wire g18159;
wire g16097;
wire g19568;
wire g34645;
wire g17390;
wire g26103;
wire g12601;
wire g29731;
wire g24986;
wire g34091;
wire g29085;
wire g11962;
wire II14773;
wire g22167;
wire g8355;
wire g22718;
wire g18557;
wire II32161;
wire g30577;
wire g33430;
wire II26989;
wire g19438;
wire g23876;
wire II18487;
wire g14988;
wire g25874;
wire II12927;
wire g24541;
wire g10416;
wire g24647;
wire g28254;
wire g28657;
wire g34398;
wire g11892;
wire g33464;
wire II13124;
wire g22550;
wire g33012;
wire g12818;
wire g34750;
wire g32139;
wire g12903;
wire g34308;
wire g25691;
wire g32280;
wire g7828;
wire g24190;
wire II17675;
wire g22646;
wire g13852;
wire g18497;
wire g27229;
wire II18414;
wire g24123;
wire g32722;
wire g17610;
wire g15751;
wire g27445;
wire g25503;
wire g33695;
wire g29617;
wire II21831;
wire g29335;
wire g25467;
wire g14574;
wire g29603;
wire g32961;
wire g26824;
wire g27359;
wire g13066;
wire g16657;
wire g9480;
wire g29029;
wire g18697;
wire g13739;
wire g33298;
wire g33954;
wire g22632;
wire g18123;
wire g19477;
wire g19875;
wire g34309;
wire g31752;
wire g25656;
wire g19698;
wire g28719;
wire g26602;
wire g10474;
wire II22467;
wire g23813;
wire g32636;
wire g33936;
wire g34172;
wire II12076;
wire g18514;
wire g17505;
wire g31759;
wire g7162;
wire g30018;
wire g24545;
wire g20184;
wire g31008;
wire g31669;
wire g27882;
wire II18495;
wire g22850;
wire g26488;
wire g8470;
wire g32621;
wire g32892;
wire g32766;
wire g9460;
wire g12971;
wire g30290;
wire II23998;
wire g29532;
wire g18665;
wire g33437;
wire g33513;
wire g28827;
wire g31784;
wire g11773;
wire g24840;
wire g28553;
wire g26890;
wire g19885;
wire g31119;
wire g34528;
wire g34479;
wire g22298;
wire g26292;
wire g23649;
wire g16741;
wire g27557;
wire g18417;
wire g17297;
wire II16733;
wire g9797;
wire g33542;
wire II32800;
wire g26021;
wire g22037;
wire g26685;
wire g31884;
wire g27928;
wire g15068;
wire g34577;
wire II22114;
wire II24549;
wire g32250;
wire g28815;
wire g18643;
wire g15052;
wire g10851;
wire g24051;
wire g29867;
wire g11191;
wire g25105;
wire g13657;
wire g33291;
wire g14454;
wire g32853;
wire g9831;
wire g28924;
wire g11471;
wire II21977;
wire g23838;
wire g27509;
wire g30031;
wire g10684;
wire g28369;
wire g33364;
wire g32035;
wire II31610;
wire g29845;
wire g28605;
wire g32169;
wire g19506;
wire g27261;
wire g9636;
wire g25612;
wire g21059;
wire g24410;
wire g27686;
wire g6848;
wire g24350;
wire g24025;
wire g29874;
wire g20574;
wire g12672;
wire g28662;
wire g11546;
wire II31092;
wire g27282;
wire g33243;
wire g29718;
wire g32838;
wire g19572;
wire g31771;
wire g32427;
wire g30415;
wire g22170;
wire g18802;
wire g7650;
wire g24564;
wire g17693;
wire g9961;
wire g21992;
wire g25771;
wire g11111;
wire g26720;
wire g23184;
wire g12873;
wire g28833;
wire g19519;
wire II18191;
wire g12867;
wire g8507;
wire g28037;
wire g18355;
wire g9354;
wire g10318;
wire g25491;
wire g9245;
wire g10929;
wire g31976;
wire g22226;
wire g30111;
wire g20666;
wire g33923;
wire g34804;
wire g33832;
wire g13970;
wire g14956;
wire g13291;
wire II18165;
wire g30483;
wire g34589;
wire g22339;
wire g32241;
wire g28198;
wire g18530;
wire g26541;
wire g32751;
wire g11144;
wire g23405;
wire g25262;
wire g15111;
wire g33661;
wire II12240;
wire II31222;
wire g34081;
wire g21931;
wire g13459;
wire g32469;
wire g33807;
wire g23029;
wire g24494;
wire II24003;
wire g16199;
wire g20784;
wire g17418;
wire g12151;
wire g16304;
wire g24839;
wire g15171;
wire g24395;
wire II17970;
wire g9902;
wire g14395;
wire g17638;
wire g27450;
wire g15581;
wire g14113;
wire g29929;
wire g20854;
wire g7469;
wire g18104;
wire g17727;
wire g29649;
wire g19433;
wire g26099;
wire g33080;
wire g24929;
wire g13672;
wire g23060;
wire g18447;
wire g18103;
wire g26863;
wire g18507;
wire g8462;
wire g24785;
wire g11790;
wire g7251;
wire g24912;
wire II17406;
wire g33495;
wire g31472;
wire g26339;
wire g24206;
wire II12251;
wire II18882;
wire g30446;
wire g10311;
wire g30303;
wire g15721;
wire g31528;
wire g23521;
wire g34014;
wire g8863;
wire g24361;
wire g17427;
wire g10133;
wire g14803;
wire g27206;
wire g26804;
wire g21966;
wire g14407;
wire g7149;
wire g22121;
wire g13461;
wire II11701;
wire g27155;
wire g33681;
wire g28343;
wire g22087;
wire g15039;
wire g16854;
wire g23502;
wire g25115;
wire g20918;
wire II15289;
wire g30492;
wire g32883;
wire g7289;
wire g13137;
wire g8239;
wire g9629;
wire II14505;
wire g23486;
wire g25322;
wire g15719;
wire II31539;
wire g33041;
wire g27660;
wire g8164;
wire g25597;
wire II24704;
wire g13313;
wire g18822;
wire g29174;
wire g12110;
wire g12185;
wire g34042;
wire g22840;
wire g17363;
wire g24193;
wire g19545;
wire g23440;
wire g11251;
wire g15140;
wire g23527;
wire g27106;
wire II17374;
wire g32442;
wire g12377;
wire g28608;
wire II14185;
wire g10037;
wire II14702;
wire g32561;
wire g11952;
wire g27532;
wire g16628;
wire g7513;
wire g25782;
wire g12049;
wire g20535;
wire II17542;
wire g11154;
wire g23537;
wire II30861;
wire II13850;
wire g26780;
wire g19915;
wire II27529;
wire II20447;
wire II29270;
wire g32107;
wire g23296;
wire g21052;
wire g30437;
wire g6755;
wire g26827;
wire II26368;
wire g26092;
wire g30345;
wire g34757;
wire g21658;
wire II31151;
wire g17598;
wire g31761;
wire g30607;
wire g21406;
wire g17140;
wire g29150;
wire g26833;
wire g18333;
wire g27825;
wire g33734;
wire g32220;
wire g22076;
wire g15872;
wire g8105;
wire g20237;
wire g23444;
wire g29962;
wire g24795;
wire g18785;
wire g19601;
wire II16102;
wire g7595;
wire g26131;
wire g30257;
wire g34418;
wire g21510;
wire g25689;
wire g24707;
wire g15707;
wire g31187;
wire II14730;
wire g30395;
wire g26805;
wire g21462;
wire g9982;
wire g19715;
wire g8807;
wire g28626;
wire g18348;
wire g27669;
wire g34333;
wire g32359;
wire g17220;
wire II12061;
wire g8534;
wire g32344;
wire g12308;
wire g32761;
wire g9964;
wire g21877;
wire g26361;
wire g32685;
wire g30360;
wire g16219;
wire g10893;
wire g21945;
wire g10793;
wire g17600;
wire g16163;
wire g33789;
wire g18199;
wire g34606;
wire g18388;
wire II31241;
wire g14631;
wire II32953;
wire g17176;
wire II22865;
wire g33342;
wire g34594;
wire g27211;
wire g25883;
wire g27285;
wire g8663;
wire g7615;
wire g7592;
wire g26945;
wire g34263;
wire g10273;
wire g24715;
wire g17712;
wire g29258;
wire II30686;
wire g12598;
wire g33704;
wire g29233;
wire g20272;
wire g28236;
wire g29287;
wire g23322;
wire II32654;
wire g25575;
wire g10504;
wire g33639;
wire g31280;
wire g19860;
wire g7971;
wire g12341;
wire II22464;
wire g28388;
wire g28588;
wire g28495;
wire g26914;
wire II32464;
wire g25661;
wire g12967;
wire g18139;
wire g21305;
wire g8905;
wire g28596;
wire g8630;
wire g7148;
wire g34579;
wire g29640;
wire II11740;
wire g25626;
wire g29942;
wire II18609;
wire g23578;
wire g33127;
wire g21513;
wire g28302;
wire g26913;
wire II32158;
wire g20672;
wire g10383;
wire g34253;
wire g21839;
wire II18765;
wire g22670;
wire g28723;
wire g16743;
wire g18885;
wire g7913;
wire g27436;
wire g25976;
wire g13021;
wire g18372;
wire II32388;
wire g20909;
wire g29804;
wire g32115;
wire g29070;
wire g17609;
wire g24150;
wire g11939;
wire g10544;
wire g24171;
wire g16730;
wire g14377;
wire g14675;
wire g25993;
wire g6803;
wire g17651;
wire g25164;
wire g22201;
wire g14367;
wire g18464;
wire g11172;
wire II22901;
wire g33524;
wire g8399;
wire g7441;
wire g32188;
wire g30246;
wire g24275;
wire g20375;
wire g23282;
wire II17392;
wire g23940;
wire II31311;
wire g23616;
wire g29566;
wire II31027;
wire g10528;
wire g8925;
wire g13869;
wire g10197;
wire II31062;
wire g16765;
wire g32813;
wire g17123;
wire g21907;
wire g22624;
wire g26908;
wire g20000;
wire g23935;
wire II19719;
wire g33624;
wire g16622;
wire II14853;
wire g13483;
wire II20891;
wire g27132;
wire g19413;
wire g12628;
wire II18671;
wire g7733;
wire g25197;
wire g25452;
wire g33973;
wire g33579;
wire g13506;
wire g25061;
wire g23530;
wire g33427;
wire g10971;
wire g33402;
wire g17955;
wire g13281;
wire II27253;
wire g28478;
wire g6982;
wire g27554;
wire g12842;
wire g16751;
wire g34565;
wire II18245;
wire g21177;
wire g20591;
wire II22748;
wire II15214;
wire g19400;
wire g31917;
wire II13564;
wire g30999;
wire g21900;
wire g24044;
wire II31192;
wire g34205;
wire g14334;
wire g17487;
wire g27402;
wire g23916;
wire g28200;
wire g14072;
wire g25668;
wire II15862;
wire g12854;
wire g16750;
wire g22448;
wire g27348;
wire g16721;
wire g13778;
wire g19790;
wire II22846;
wire g34213;
wire II33267;
wire g31782;
wire g32473;
wire g21394;
wire g13508;
wire g12286;
wire g28191;
wire g29711;
wire II31593;
wire gbuf107;
wire g30592;
wire g31877;
wire g29310;
wire II19671;
wire g17589;
wire g22495;
wire g20653;
wire g10948;
wire g14974;
wire g17475;
wire g29954;
wire g21980;
wire g29207;
wire g32612;
wire II17747;
wire II31257;
wire II24625;
wire II18071;
wire g25296;
wire g33618;
wire g18597;
wire g27074;
wire g7655;
wire g34747;
wire g29707;
wire II17474;
wire g18573;
wire gbuf2;
wire g23076;
wire g30439;
wire g9835;
wire g18436;
wire g17929;
wire II15162;
wire g22050;
wire II23680;
wire g16717;
wire g32968;
wire g22116;
wire g27924;
wire g30560;
wire g28040;
wire g31831;
wire g26270;
wire g25757;
wire g11970;
wire g23614;
wire g31925;
wire g16584;
wire II32119;
wire II18589;
wire g9049;
wire g33352;
wire g17786;
wire g24972;
wire g14308;
wire g13004;
wire g30514;
wire g16931;
wire g27965;
wire g29662;
wire II23602;
wire g32271;
wire g24419;
wire g31289;
wire g27629;
wire g29590;
wire II23987;
wire II27514;
wire g33339;
wire g28454;
wire g13888;
wire g30256;
wire g32902;
wire g29479;
wire g30271;
wire g32420;
wire g23903;
wire II32594;
wire II22547;
wire II19484;
wire g18767;
wire g13211;
wire g12137;
wire g10537;
wire II18580;
wire g22042;
wire g18907;
wire g34343;
wire g16920;
wire g17512;
wire II25514;
wire g29077;
wire g34640;
wire g27576;
wire g27245;
wire II26419;
wire g27302;
wire g21710;
wire g20580;
wire g30185;
wire g16589;
wire g19481;
wire g9206;
wire g32574;
wire g29377;
wire g27409;
wire g20149;
wire II14932;
wire g10153;
wire g9599;
wire g7868;
wire g28109;
wire g13114;
wire g23801;
wire g34002;
wire g26356;
wire g24155;
wire g29359;
wire g10530;
wire g18762;
wire g30252;
wire g23546;
wire g29997;
wire g26212;
wire II33273;
wire II22031;
wire II25576;
wire g31017;
wire g31900;
wire II33300;
wire g34932;
wire g12982;
wire g28067;
wire g11885;
wire g31131;
wire g10582;
wire g26343;
wire g7975;
wire g34313;
wire II21291;
wire g26847;
wire g12930;
wire g22138;
wire g32377;
wire g20204;
wire g10376;
wire II19674;
wire g33520;
wire g32349;
wire g29516;
wire g13284;
wire g16242;
wire g7873;
wire II22872;
wire g20618;
wire g32496;
wire g21971;
wire II23360;
wire g26928;
wire g31502;
wire g18976;
wire g27505;
wire g13513;
wire g32675;
wire g33718;
wire g28444;
wire g8954;
wire g32536;
wire g15079;
wire II16135;
wire g25707;
wire g32010;
wire g31166;
wire g33451;
wire g28568;
wire g27220;
wire II14584;
wire g28325;
wire g20158;
wire g32669;
wire g22455;
wire g33446;
wire II31347;
wire g26888;
wire g29497;
wire II29284;
wire gbuf100;
wire g31941;
wire g33506;
wire II26296;
wire g8977;
wire g21976;
wire II11777;
wire g33393;
wire g30545;
wire g13948;
wire g14058;
wire g20191;
wire g15833;
wire g27698;
wire g33144;
wire g16213;
wire g33855;
wire g26931;
wire II22823;
wire g26918;
wire g27691;
wire g17013;
wire g10905;
wire g34861;
wire II12849;
wire II18813;
wire g15849;
wire g30447;
wire g34169;
wire II12279;
wire II20222;
wire g9386;
wire g22636;
wire g27550;
wire g13951;
wire g22457;
wire g14537;
wire g32097;
wire g20277;
wire g24015;
wire g34005;
wire g34359;
wire II23970;
wire g19069;
wire g31838;
wire g19694;
wire g31934;
wire II16521;
wire g22124;
wire g33003;
wire g30535;
wire g34327;
wire g34496;
wire g20912;
wire g33960;
wire g18249;
wire g17302;
wire g29741;
wire g21454;
wire g32268;
wire g7903;
wire g34966;
wire g27257;
wire g25456;
wire II26742;
wire g33040;
wire II18849;
wire g20159;
wire g9500;
wire g33637;
wire g32175;
wire g33531;
wire g33887;
wire g14601;
wire g22155;
wire g19800;
wire g24166;
wire g7096;
wire g33527;
wire g10364;
wire g32619;
wire g6987;
wire g23685;
wire g9061;
wire g26836;
wire g29482;
wire g20494;
wire g34852;
wire II14817;
wire g13762;
wire g12045;
wire g25925;
wire II15633;
wire g18522;
wire g13323;
wire g31013;
wire g12795;
wire II28566;
wire g32725;
wire g24653;
wire g11047;
wire II27713;
wire g27460;
wire g18711;
wire g33219;
wire g32014;
wire II33024;
wire g18982;
wire g27700;
wire g33683;
wire g34619;
wire II14690;
wire g31823;
wire II13020;
wire g24232;
wire g27114;
wire g14257;
wire II17636;
wire g31492;
wire g30028;
wire II31102;
wire g11214;
wire g27830;
wire g18217;
wire g10627;
wire g18508;
wire g12453;
wire g33379;
wire g18233;
wire g17413;
wire g29633;
wire g33901;
wire g25037;
wire g20434;
wire g28696;
wire g13667;
wire g34504;
wire g28297;
wire g14768;
wire g34468;
wire g14066;
wire g32511;
wire g25908;
wire g30518;
wire g29294;
wire g20587;
wire g15724;
wire g13796;
wire II31306;
wire g8899;
wire g17583;
wire g25399;
wire g28258;
wire g31294;
wire II14788;
wire g24246;
wire g29004;
wire g12490;
wire g16689;
wire g33089;
wire g7138;
wire g18732;
wire g21209;
wire II18233;
wire g10361;
wire g32275;
wire g25964;
wire II12776;
wire g19344;
wire g16772;
wire g11270;
wire g34354;
wire g11978;
wire g21987;
wire g14562;
wire II17228;
wire II26427;
wire g29279;
wire g33020;
wire II25356;
wire g10829;
wire gbuf73;
wire II29368;
wire II22822;
wire g33356;
wire g10761;
wire g13515;
wire g28880;
wire g31150;
wire II31491;
wire g26121;
wire g29613;
wire g21806;
wire g15122;
wire g28075;
wire g17213;
wire g14522;
wire g18725;
wire g31244;
wire g7897;
wire g18244;
wire g28663;
wire g34106;
wire g13660;
wire g29885;
wire g20213;
wire g32251;
wire g34783;
wire g33997;
wire g12015;
wire g25134;
wire g21716;
wire g16312;
wire g21674;
wire g34060;
wire g24578;
wire g34694;
wire g16706;
wire g12900;
wire g31653;
wire g30359;
wire g11715;
wire g13850;
wire g33517;
wire g13728;
wire g24262;
wire II13045;
wire g12147;
wire g16687;
wire g32872;
wire g27517;
wire g6815;
wire g21847;
wire g26119;
wire g25549;
wire II28390;
wire g24483;
wire II11866;
wire g9713;
wire g19422;
wire II31751;
wire g28949;
wire g12466;
wire g16527;
wire g13999;
wire g33258;
wire g28994;
wire II32693;
wire g13117;
wire II29236;
wire g26682;
wire g25769;
wire g29262;
wire g24568;
wire g8114;
wire g23884;
wire g25894;
wire II27314;
wire g22340;
wire g22684;
wire II21222;
wire g22100;
wire II31561;
wire g31962;
wire g11181;
wire g28053;
wire g34777;
wire g19471;
wire II13979;
wire g22642;
wire g26326;
wire g32149;
wire g34698;
wire g27490;
wire g25986;
wire g25930;
wire g23244;
wire g22325;
wire g16422;
wire g17705;
wire g23844;
wire g28287;
wire II31351;
wire g22928;
wire g14054;
wire g10182;
wire g29182;
wire II31586;
wire g30440;
wire gbuf125;
wire g24421;
wire g30175;
wire g16159;
wire g34709;
wire II14400;
wire g10724;
wire g15695;
wire g28373;
wire II33270;
wire g33315;
wire g34491;
wire g18886;
wire g32610;
wire g27821;
wire g10981;
wire g9906;
wire g13217;
wire II17380;
wire g18341;
wire g16202;
wire g29036;
wire g17091;
wire g24426;
wire g32527;
wire g32931;
wire II31814;
wire II22899;
wire g32831;
wire g13915;
wire II26785;
wire g28264;
wire g13320;
wire II14211;
wire g12039;
wire g18432;
wire g29629;
wire g32445;
wire g34456;
wire g16651;
wire g33343;
wire g8945;
wire g30216;
wire g22757;
wire g12079;
wire g21420;
wire g21425;
wire II21019;
wire g26749;
wire II13077;
wire g20168;
wire g23642;
wire g18692;
wire g34985;
wire g24664;
wire II32067;
wire g20705;
wire g26258;
wire g23229;
wire g10059;
wire g26952;
wire g28074;
wire g33072;
wire g28462;
wire g26960;
wire g10428;
wire g24240;
wire g31888;
wire g26257;
wire g25802;
wire II11816;
wire g27522;
wire II24054;
wire g11911;
wire II12910;
wire g17644;
wire g23004;
wire g16182;
wire g18680;
wire g18503;
wire g34678;
wire g28282;
wire g18685;
wire g23336;
wire g10050;
wire g27976;
wire g23222;
wire g26307;
wire II24679;
wire g12029;
wire g13062;
wire g27140;
wire g28310;
wire g26893;
wire g7633;
wire g32573;
wire g33116;
wire g19711;
wire g27955;
wire g15085;
wire g25163;
wire g24573;
wire II15300;
wire g31465;
wire g27354;
wire g14936;
wire g20086;
wire g15157;
wire g18170;
wire g8639;
wire II29297;
wire g24488;
wire II18734;
wire g33845;
wire g23966;
wire g34391;
wire g29044;
wire g28120;
wire g20643;
wire g33019;
wire g19649;
wire g25208;
wire g8539;
wire g27268;
wire g10281;
wire g11872;
wire II33140;
wire g12895;
wire g8984;
wire II11820;
wire g22899;
wire II12890;
wire g16673;
wire g12224;
wire g26082;
wire g28272;
wire g23690;
wire g13174;
wire g11445;
wire g33896;
wire g34038;
wire gbuf49;
wire g20509;
wire g24322;
wire II18530;
wire g32500;
wire g32804;
wire g24314;
wire g18065;
wire g10203;
wire g9213;
wire g16666;
wire II17401;
wire g14441;
wire g33306;
wire g34702;
wire g21163;
wire g19685;
wire g32364;
wire II32766;
wire g14005;
wire g27324;
wire g32200;
wire II19756;
wire g22384;
wire II17188;
wire g8396;
wire g25152;
wire II26406;
wire II13329;
wire g17524;
wire g12687;
wire g10430;
wire g23991;
wire g18631;
wire g33234;
wire II30735;
wire II14925;
wire g18756;
wire II23315;
wire g21776;
wire g20108;
wire g12021;
wire g34525;
wire II26356;
wire g13912;
wire g12246;
wire g21434;
wire g13083;
wire g14885;
wire g19462;
wire g14446;
wire g28420;
wire g27361;
wire g29794;
wire g11371;
wire g17526;
wire g28452;
wire g32771;
wire g28335;
wire g10393;
wire II12135;
wire g12100;
wire gbuf66;
wire g29320;
wire II29986;
wire g32327;
wire g18565;
wire g20525;
wire g9775;
wire g34219;
wire g9558;
wire g7998;
wire g26186;
wire g11691;
wire g32745;
wire g27016;
wire g24128;
wire g20092;
wire g30231;
wire II19863;
wire g32120;
wire g18223;
wire g10521;
wire g29259;
wire g22919;
wire g15808;
wire II32433;
wire g21730;
wire g21140;
wire g19732;
wire II25005;
wire g14807;
wire g27183;
wire II18131;
wire II23369;
wire II18674;
wire II14247;
wire g20778;
wire II16057;
wire g24589;
wire g34409;
wire g33561;
wire g24942;
wire II29314;
wire g24764;
wire g11127;
wire g10816;
wire g23171;
wire g22988;
wire g19415;
wire II24281;
wire g32715;
wire g16532;
wire II25541;
wire g25996;
wire g22589;
wire g24896;
wire g13013;
wire g29937;
wire g15634;
wire g31233;
wire g16190;
wire g18992;
wire II11750;
wire g9585;
wire II31072;
wire g26809;
wire g27730;
wire g17770;
wire g26300;
wire g25710;
wire II12403;
wire g27430;
wire g10408;
wire g24224;
wire g8677;
wire g26608;
wire g24287;
wire g22528;
wire g13329;
wire II13464;
wire g27294;
wire g18671;
wire g15915;
wire g34256;
wire g26176;
wire g15135;
wire g28677;
wire g12121;
wire g30099;
wire g29243;
wire g23778;
wire g32292;
wire g32395;
wire g24146;
wire g32505;
wire g13867;
wire g31756;
wire g26959;
wire g7534;
wire g25226;
wire g10233;
wire g28400;
wire g19409;
wire g9185;
wire g22191;
wire g11981;
wire g24068;
wire g12125;
wire g29346;
wire g20711;
wire g33091;
wire g33860;
wire g26571;
wire g16872;
wire II27784;
wire g28187;
wire g16803;
wire g9915;
wire g24770;
wire g24061;
wire g19869;
wire g14730;
wire g17149;
wire g7840;
wire g25125;
wire g33328;
wire g18650;
wire g29501;
wire g34900;
wire g30284;
wire g10377;
wire g32850;
wire g34190;
wire g22907;
wire g22876;
wire g23708;
wire g26816;
wire g11509;
wire g7296;
wire g34543;
wire g32915;
wire II30644;
wire g17738;
wire II27409;
wire g30367;
wire g17466;
wire g8381;
wire II18214;
wire g16611;
wire g28919;
wire g30477;
wire g12931;
wire g17226;
wire g34542;
wire g28362;
wire g24331;
wire g15864;
wire g18371;
wire g34507;
wire g11160;
wire II17808;
wire g9843;
wire g20248;
wire II27718;
wire g11994;
wire II17569;
wire g33108;
wire g23782;
wire g32411;
wire g12836;
wire g33676;
wire g24207;
wire g29480;
wire g6974;
wire g25556;
wire II19384;
wire g32547;
wire g28111;
wire g27482;
wire g28580;
wire g25752;
wire II18276;
wire g28309;
wire g8055;
wire II30761;
wire II16471;
wire g8280;
wire g9863;
wire g24372;
wire g11330;
wire g25096;
wire g14133;
wire g23550;
wire g20921;
wire g25288;
wire g14148;
wire g33411;
wire g31126;
wire g10295;
wire g32664;
wire g17469;
wire g27566;
wire g27386;
wire g31270;
wire g8756;
wire g13025;
wire g23857;
wire g18614;
wire g34934;
wire g21067;
wire II26459;
wire g21723;
wire g10028;
wire g10708;
wire g24052;
wire g29574;
wire g8316;
wire g22319;
wire g34021;
wire II32846;
wire g30420;
wire g27997;
wire g12622;
wire g21558;
wire g30104;
wire g24582;
wire g14231;
wire g21822;
wire g33272;
wire g28704;
wire g33932;
wire g9705;
wire g28044;
wire g21467;
wire g33586;
wire g32027;
wire II21002;
wire g26737;
wire g23551;
wire g11233;
wire g15059;
wire g34534;
wire g9285;
wire g13995;
wire g17671;
wire g17495;
wire II24600;
wire g32162;
wire g26856;
wire g17721;
wire g21897;
wire g33132;
wire g23277;
wire g26128;
wire g32670;
wire g19209;
wire II30055;
wire g12430;
wire g29675;
wire g24523;
wire g21871;
wire g14183;
wire g17718;
wire g33875;
wire II26670;
wire g8205;
wire g18399;
wire g26157;
wire g23872;
wire g29300;
wire g24341;
wire g31372;
wire g34535;
wire g26645;
wire g24754;
wire II32547;
wire g9972;
wire g7879;
wire g32021;
wire g30308;
wire g26719;
wire g29686;
wire II21288;
wire g29025;
wire g29097;
wire g14543;
wire g11010;
wire g24880;
wire g32911;
wire II29351;
wire g20447;
wire g10030;
wire II33255;
wire g23359;
wire II26667;
wire II32871;
wire g20570;
wire g20241;
wire g20548;
wire g14387;
wire g14431;
wire g30504;
wire g30072;
wire g34248;
wire g34104;
wire g9684;
wire g19902;
wire g32055;
wire II27391;
wire g24432;
wire g6810;
wire g34131;
wire g32227;
wire g34115;
wire g21123;
wire g33987;
wire g31579;
wire g11865;
wire g31819;
wire g32072;
wire II15043;
wire g26657;
wire g31253;
wire g13977;
wire g14898;
wire g18369;
wire g6993;
wire II28162;
wire g33829;
wire g14223;
wire g21878;
wire II26072;
wire II28174;
wire g25726;
wire g23985;
wire II12712;
wire g24405;
wire g24656;
wire g16507;
wire II14836;
wire g14641;
wire II20204;
wire II22327;
wire g23986;
wire g27548;
wire g24904;
wire g23953;
wire II31156;
wire g21455;
wire g11410;
wire g25233;
wire g15883;
wire g33483;
wire II32056;
wire g29142;
wire g22080;
wire g33139;
wire g25013;
wire II18452;
wire g34977;
wire g32995;
wire g11737;
wire g28163;
wire II22918;
wire II13995;
wire g23995;
wire g12370;
wire g10678;
wire g15877;
wire g20059;
wire g29361;
wire II12997;
wire g18796;
wire g33831;
wire g26635;
wire g29755;
wire g29609;
wire g28174;
wire g27614;
wire g16264;
wire g25400;
wire g11374;
wire g29317;
wire g11115;
wire g32337;
wire g7304;
wire g18209;
wire g26613;
wire g30285;
wire g10053;
wire g34675;
wire g33439;
wire II28579;
wire II24117;
wire g27033;
wire g17290;
wire g24170;
wire g34720;
wire g14028;
wire g33093;
wire g31524;
wire II14206;
wire g28223;
wire II31297;
wire g10510;
wire g24443;
wire g21932;
wire g32843;
wire g27962;
wire g13463;
wire g23860;
wire g17572;
wire II26676;
wire II12374;
wire g13908;
wire g30293;
wire g20085;
wire g16483;
wire g34517;
wire II32988;
wire II22921;
wire g8796;
wire g14021;
wire g24629;
wire II31202;
wire g25732;
wire g25513;
wire g32603;
wire g23010;
wire g33908;
wire g15094;
wire g33549;
wire g17284;
wire g17151;
wire g22999;
wire g34660;
wire g10721;
wire g18414;
wire g13499;
wire g28567;
wire g29281;
wire g25538;
wire g28340;
wire g23900;
wire g31279;
wire g18202;
wire g27759;
wire g32942;
wire g32199;
wire g23699;
wire g20767;
wire g6821;
wire g33474;
wire g8134;
wire g33880;
wire g24558;
wire g19787;
wire g22139;
wire g24016;
wire II31211;
wire g18186;
wire II12269;
wire g32829;
wire g12592;
wire g33025;
wire g23456;
wire g34245;
wire gbuf83;
wire g29303;
wire g26396;
wire II18694;
wire g24004;
wire g34123;
wire g24188;
wire II26523;
wire g9392;
wire g23411;
wire g10044;
wire g19370;
wire g25739;
wire II15333;
wire g12851;
wire g24604;
wire g30131;
wire II22264;
wire II31807;
wire g25530;
wire g16702;
wire g24551;
wire g23233;
wire g14844;
wire g29881;
wire g21332;
wire g29555;
wire g12008;
wire g24280;
wire g8951;
wire g28416;
wire g33678;
wire II23399;
wire g25139;
wire g16187;
wire g21414;
wire g14751;
wire II32458;
wire II22683;
wire g31506;
wire g25073;
wire g30263;
wire g8654;
wire g20710;
wire g13095;
wire II14171;
wire g10166;
wire II23345;
wire g10001;
wire g23771;
wire g18720;
wire g29974;
wire II14050;
wire II17460;
wire g27775;
wire g24960;
wire g28681;
wire g27413;
wire g30158;
wire g34076;
wire g29851;
wire g21769;
wire g18362;
wire g34725;
wire g12429;
wire II11793;
wire g33008;
wire II13565;
wire gbuf24;
wire g26295;
wire g11382;
wire g10617;
wire g29663;
wire g33055;
wire g33101;
wire g23726;
wire g25426;
wire g24704;
wire g24254;
wire g23655;
wire g18655;
wire g25480;
wire g25776;
wire g20388;
wire g26386;
wire g15127;
wire II16544;
wire g12347;
wire g23432;
wire g34296;
wire g7766;
wire II13152;
wire g10107;
wire g16306;
wire g12955;
wire g23531;
wire II32938;
wire g32384;
wire g11402;
wire g18810;
wire g16707;
wire g22177;
wire g32128;
wire g16929;
wire g28934;
wire g11763;
wire g17433;
wire g10112;
wire g24608;
wire g24743;
wire II12503;
wire g27878;
wire g25580;
wire g27458;
wire II27401;
wire g15965;
wire g33286;
wire g30336;
wire II15773;
wire g9807;
wire II31057;
wire g19747;
wire g30050;
wire g16324;
wire g15005;
wire g10338;
wire g15167;
wire II18066;
wire g29764;
wire g25408;
wire g31796;
wire II26693;
wire g32776;
wire g8059;
wire II32794;
wire II15144;
wire II31216;
wire g31497;
wire g24111;
wire g34870;
wire g7439;
wire II22712;
wire g34484;
wire g18262;
wire g11360;
wire g14379;
wire g18539;
wire g8255;
wire g8365;
wire g30011;
wire g19444;
wire g27330;
wire g23211;
wire g12525;
wire g19593;
wire g27596;
wire g31808;
wire g33570;
wire g28292;
wire g26690;
wire g32330;
wire g18894;
wire g13492;
wire g29511;
wire g15700;
wire g19352;
wire g8587;
wire g17182;
wire g14321;
wire g20103;
wire g33799;
wire g13901;
wire g25947;
wire g25099;
wire g6960;
wire II15295;
wire g18957;
wire g33035;
wire g26701;
wire g28732;
wire g13771;
wire g22590;
wire g10355;
wire g34582;
wire II14259;
wire g10029;
wire g28206;
wire g27337;
wire g7684;
wire g7475;
wire g31481;
wire g34280;
wire II32439;
wire g28357;
wire g14930;
wire g28488;
wire II13779;
wire g24137;
wire g18929;
wire g14871;
wire g31913;
wire g24201;
wire g28707;
wire g26935;
wire g34145;
wire II24067;
wire g24665;
wire g8273;
wire g34330;
wire g32983;
wire g28747;
wire g8912;
wire g22531;
wire g9056;
wire g13103;
wire g24466;
wire g30314;
wire g9829;
wire g15011;
wire g29692;
wire II14016;
wire g18157;
wire g34561;
wire g18634;
wire II31007;
wire g19533;
wire gbuf96;
wire g11381;
wire g22664;
wire g32068;
wire g19880;
wire g33361;
wire g33545;
wire g24303;
wire g11935;
wire g25748;
wire g25001;
wire g16813;
wire g31967;
wire g13528;
wire g9529;
wire g22936;
wire g32707;
wire g25160;
wire g16212;
wire g16283;
wire g27122;
wire II19927;
wire g33386;
wire II22622;
wire gbuf12;
wire II22046;
wire g22005;
wire g6825;
wire g29523;
wire g24408;
wire g12059;
wire g33955;
wire g28144;
wire g24103;
wire g7887;
wire g26923;
wire II14212;
wire g20077;
wire g13892;
wire g21127;
wire g18116;
wire g9391;
wire g19540;
wire II17938;
wire II18861;
wire g26672;
wire g29751;
wire g23334;
wire g34765;
wire g30614;
wire g34576;
wire g8889;
wire g10351;
wire g13017;
wire g34816;
wire g21954;
wire g9607;
wire g18326;
wire g33310;
wire II30192;
wire g19930;
wire g24591;
wire g8009;
wire g11405;
wire g23923;
wire g29879;
wire g22519;
wire g32104;
wire g20130;
wire g33580;
wire g27161;
wire g14613;
wire g18273;
wire g28157;
wire g21886;
wire g21735;
wire II25692;
wire g11490;
wire g12907;
wire g15115;
wire g23308;
wire g34588;
wire g22329;
wire g12311;
wire g19383;
wire g13555;
wire g34763;
wire g22647;
wire II15307;
wire g33917;
wire g16203;
wire g24687;
wire g18903;
wire g20007;
wire g26820;
wire g24966;
wire g24675;
wire g27854;
wire g25592;
wire g20598;
wire g29536;
wire g30115;
wire g18668;
wire g9590;
wire g18518;
wire II22557;
wire g14570;
wire g30373;
wire II18560;
wire g8808;
wire g24211;
wire II26638;
wire g10800;
wire g10921;
wire g10553;
wire g24115;
wire g25241;
wire g25870;
wire g25085;
wire g25981;
wire g33353;
wire g18185;
wire g15708;
wire g11966;
wire g25742;
wire g20577;
wire g32487;
wire g33460;
wire g28713;
wire g24729;
wire g9965;
wire g32142;
wire II30400;
wire g34367;
wire g20219;
wire g14959;
wire g9958;
wire g18278;
wire g29185;
wire g26253;
wire g33658;
wire g12074;
wire g23720;
wire g18470;
wire g28613;
wire g24548;
wire g33434;
wire II31031;
wire II12075;
wire g14027;
wire g28856;
wire g19786;
wire g29263;
wire II15577;
wire II16875;
wire g29608;
wire g13041;
wire g34475;
wire g25542;
wire g33621;
wire g29368;
wire g17741;
wire II12287;
wire g19890;
wire g23381;
wire g13299;
wire g28271;
wire g26954;
wire g34516;
wire g13300;
wire g18126;
wire g21924;
wire g27412;
wire g17501;
wire II22485;
wire g23388;
wire g15836;
wire II13182;
wire g8721;
wire g28214;
wire g29595;
wire II14301;
wire g20561;
wire II17446;
wire g18135;
wire II17671;
wire g16811;
wire g26287;
wire g13822;
wire II25612;
wire g8579;
wire g13010;
wire g28442;
wire g20028;
wire g23841;
wire II31162;
wire g21921;
wire g20268;
wire g29859;
wire g23682;
wire g32645;
wire g23427;
wire g12052;
wire g17239;
wire g24468;
wire g12152;
wire g9554;
wire g32509;
wire II15208;
wire g8442;
wire II12572;
wire g13675;
wire g34342;
wire g31488;
wire g29914;
wire g11373;
wire g11866;
wire g28892;
wire g30021;
wire g17614;
wire II15918;
wire g29274;
wire II20830;
wire g18490;
wire g25528;
wire g13312;
wire II24078;
wire g29154;
wire g34774;
wire g25047;
wire g32457;
wire g9564;
wire g33980;
wire g34873;
wire g18146;
wire II31096;
wire g33469;
wire g30081;
wire g26778;
wire g27933;
wire g33247;
wire g34667;
wire g25955;
wire g27264;
wire g26179;
wire g16233;
wire II22912;
wire II14550;
wire g32269;
wire II21992;
wire g12914;
wire g20058;
wire g28385;
wire g16964;
wire g12221;
wire g33335;
wire g33496;
wire g12997;
wire g32754;
wire g30002;
wire g19961;
wire g30240;
wire g18875;
wire g21697;
wire II12819;
wire II12538;
wire g23030;
wire g28107;
wire II18855;
wire g32595;
wire g27040;
wire g25217;
wire g11255;
wire g12381;
wire g34264;
wire II32186;
wire g18739;
wire g32648;
wire g8713;
wire g32303;
wire II31625;
wire g22107;
wire g28542;
wire g34807;
wire g15815;
wire g24843;
wire g30353;
wire II16575;
wire g18216;
wire g15812;
wire g6954;
wire g32955;
wire g8417;
wire g33381;
wire g17199;
wire g25348;
wire g19997;
wire g12864;
wire g27129;
wire g33368;
wire g22306;
wire II15814;
wire g28239;
wire g30277;
wire II17615;
wire g14664;
wire g13622;
wire g19062;
wire g27234;
wire g25877;
wire g30572;
wire g28602;
wire g23314;
wire g9478;
wire g16313;
wire g32686;
wire g34349;
wire g24925;
wire g18623;
wire II15036;
wire g31154;
wire II18872;
wire g10821;
wire g30186;
wire II25359;
wire g20323;
wire g17192;
wire g14663;
wire g29191;
wire g31985;
wire g9772;
wire g34573;
wire g34052;
wire g10288;
wire g17059;
wire g12477;
wire g27493;
wire g31246;
wire g29236;
wire g26377;
wire g21289;
wire g25109;
wire g14565;
wire g14416;
wire g34976;
wire II31859;
wire II12120;
wire g34988;
wire g25187;
wire g12939;
wire g33263;
wire g15743;
wire g24347;
wire g20194;
wire g18946;
wire g33084;
wire II17379;
wire g29788;
wire g29870;
wire gbuf7;
wire g26689;
wire g34878;
wire g13523;
wire g18953;
wire g15783;
wire g30517;
wire g8584;
wire g13156;
wire g13378;
wire g16866;
wire g22661;
wire g20977;
wire g34716;
wire g9822;
wire g27601;
wire g32735;
wire g28134;
wire g11149;
wire g18833;
wire g10928;
wire g8957;
wire g11929;
wire g30176;
wire g27650;
wire g34183;
wire g14761;
wire g16695;
wire g21988;
wire g22210;
wire g29491;
wire g13079;
wire g13322;
wire g6946;
wire g7891;
wire g26887;
wire g34567;
wire g23503;
wire g30129;
wire II18653;
wire g12014;
wire g25488;
wire g10033;
wire g7806;
wire g34613;
wire g9253;
wire g20869;
wire g33728;
wire g27045;
wire g24819;
wire g23084;
wire g29007;
wire g14170;
wire gbuf41;
wire g20717;
wire g8990;
wire II17125;
wire g25369;
wire g24957;
wire g20146;
wire II24060;
wire g8021;
wire g11037;
wire g23792;
wire II14797;
wire g13567;
wire g25886;
wire g14065;
wire g20605;
wire g27325;
wire g27541;
wire g32231;
wire g32834;
wire g14422;
wire g18763;
wire g14644;
wire g32480;
wire II14509;
wire g21282;
wire g9506;
wire g16300;
wire g34093;
wire g14848;
wire g11217;
wire g34639;
wire g17088;
wire g33047;
wire g18598;
wire g14586;
wire II16515;
wire g17771;
wire g15793;
wire g27098;
wire g34555;
wire g17399;
wire g16604;
wire II16345;
wire g19852;
wire g32195;
wire g21713;
wire g30225;
wire g23189;
wire g19594;
wire gbuf19;
wire g34796;
wire g7195;
wire g34322;
wire g23957;
wire g28690;
wire g32922;
wire g7526;
wire g7041;
wire g25008;
wire g22208;
wire g9381;
wire g18562;
wire g14363;
wire g28814;
wire g7932;
wire g17154;
wire g21403;
wire g27648;
wire g31541;
wire g27551;
wire g16618;
wire g21788;
wire II15677;
wire g22215;
wire II32613;
wire g33069;
wire gbuf54;
wire g11269;
wire g10802;
wire g34179;
wire g26625;
wire g29128;
wire II14935;
wire g14913;
wire g14497;
wire g29894;
wire g33686;
wire II22958;
wire g18297;
wire g34045;
wire g19968;
wire g28609;
wire g16239;
wire g25972;
wire g9754;
wire g20635;
wire g33370;
wire g29953;
wire g24416;
wire g30108;
wire g32681;
wire g11510;
wire g21808;
wire II22967;
wire g8389;
wire g19950;
wire g10589;
wire g9887;
wire g19147;
wire g23482;
wire g34940;
wire g28323;
wire g30040;
wire g15822;
wire II18385;
wire g31140;
wire g28726;
wire g33719;
wire g20283;
wire g18302;
wire g21272;
wire II12893;
wire g17287;
wire g33628;
wire g23573;
wire g21855;
wire g13583;
wire g27384;
wire g17816;
wire g31218;
wire g29985;
wire g14290;
wire g14432;
wire g28733;
wire g11384;
wire g29254;
wire g29569;
wire g15134;
wire g7046;
wire g34054;
wire g31223;
wire g20765;
wire g34207;
wire II33131;
wire g10002;
wire II22788;
wire II18571;
wire g20374;
wire g23017;
wire g27036;
wire g27240;
wire g9537;
wire g31269;
wire g7473;
wire g19719;
wire g29869;
wire g10156;
wire g20624;
wire g18546;
wire g34120;
wire g33943;
wire g9746;
wire II25242;
wire g26090;
wire g17709;
wire g8177;
wire g8748;
wire g32860;
wire g22159;
wire g32456;
wire g32706;
wire g10354;
wire g18604;
wire g21654;
wire g28458;
wire II28591;
wire g23266;
wire g22530;
wire g21514;
wire g13543;
wire g27572;
wire g9653;
wire g13596;
wire g15829;
wire g9014;
wire g16712;
wire g25498;
wire g21833;
wire g19565;
wire g34188;
wire g8833;
wire g11932;
wire g20089;
wire g22017;
wire II31869;
wire g31601;
wire g33584;
wire g15125;
wire g24498;
wire g17179;
wire g10111;
wire g24095;
wire g20330;
wire II14497;
wire g31929;
wire g25327;
wire g18551;
wire g31873;
wire II17094;
wire g24175;
wire g21329;
wire g22863;
wire g21380;
wire g32159;
wire II32234;
wire g24271;
wire g14609;
wire g8922;
wire g25849;
wire II13483;
wire g28819;
wire g13000;
wire g23944;
wire g28765;
wire g25192;
wire II14225;
wire g23350;
wire g24380;
wire g21011;
wire g18314;
wire g10775;
wire g20179;
wire g20080;
wire g28097;
wire g15699;
wire g24040;
wire g22054;
wire g34598;
wire g27594;
wire g23286;
wire g34271;
wire II29337;
wire g15803;
wire g25156;
wire g18253;
wire g24327;
wire g32089;
wire g32631;
wire g14679;
wire g34843;
wire g25396;
wire II32921;
wire g14773;
wire g24114;
wire g9852;
wire g13007;
wire g29719;
wire g13509;
wire g33701;
wire II18903;
wire g31284;
wire g32786;
wire g28306;
wire g21396;
wire g34162;
wire g14166;
wire g17471;
wire g12972;
wire g34287;
wire g34231;
wire g32285;
wire g32808;
wire g23285;
wire g27988;
wire g23617;
wire g24278;
wire g32424;
wire g22525;
wire g24659;
wire g34452;
wire g29880;
wire g9064;
wire g29331;
wire g14252;
wire g26793;
wire g25677;
wire g29993;
wire g19581;
wire g10612;
wire II21784;
wire II33246;
wire g20538;
wire g16595;
wire II16713;
wire g15590;
wire g27027;
wire g15673;
wire g32964;
wire II15663;
wire g24032;
wire g10856;
wire g19794;
wire g25093;
wire g29758;
wire g29891;
wire g13110;
wire II18265;
wire g30192;
wire g27020;
wire g15024;
wire g27969;
wire g26605;
wire II13276;
wire g16588;
wire g32124;
wire g20442;
wire g29657;
wire g22490;
wire g26261;
wire g21785;
wire II21100;
wire g22881;
wire g12859;
wire g14792;
wire g8818;
wire II12106;
wire g13856;
wire g34529;
wire g14905;
wire II26952;
wire g32816;
wire g17530;
wire g26548;
wire g28250;
wire g11610;
wire g32848;
wire g29775;
wire II11826;
wire II13715;
wire g9721;
wire g7541;
wire g29373;
wire g18577;
wire g25578;
wire g19468;
wire g28557;
wire g31908;
wire g23630;
wire g18619;
wire g26291;
wire II18063;
wire g27249;
wire g22135;
wire II20999;
wire g27225;
wire g23291;
wire g19450;
wire g26906;
wire g32847;
wire g34731;
wire II15263;
wire g24809;
wire g14333;
wire II15878;
wire g25141;
wire g8858;
wire g23087;
wire II22719;
wire g13394;
wire g23230;
wire g32130;
wire g9819;
wire g15859;
wire II25369;
wire g34068;
wire g29770;
wire g14278;
wire II14424;
wire g20905;
wire g17592;
wire g23653;
wire g7824;
wire g10541;
wire g14271;
wire II24414;
wire g31710;
wire gbuf39;
wire g13247;
wire g17579;
wire g12182;
wire g15739;
wire g7086;
wire II33134;
wire g26789;
wire g14024;
wire g34519;
wire g33405;
wire II12117;
wire g19528;
wire g33708;
wire g18468;
wire g33407;
wire g24143;
wire g29808;
wire II22542;
wire g24389;
wire g31260;
wire II15089;
wire g32400;
wire g34166;
wire g15056;
wire g23461;
wire g31183;
wire g30465;
wire g30413;
wire g32763;
wire g32403;
wire g11592;
wire g28046;
wire g30276;
wire g9816;
wire II21480;
wire II16698;
wire g23544;
wire g27959;
wire II22286;
wire g23360;
wire g32857;
wire g24789;
wire g32978;
wire g26724;
wire g14841;
wire g16023;
wire II13730;
wire g18395;
wire g29147;
wire g33606;
wire g26516;
wire g21143;
wire g25815;
wire II11903;
wire g32676;
wire II11908;
wire g29849;
wire g10022;
wire g29547;
wire g25711;
wire g33837;
wire g30418;
wire g24526;
wire g15109;
wire g10736;
wire g29381;
wire g19752;
wire g25785;
wire g26972;
wire g19553;
wire g19364;
wire g23721;
wire g33725;
wire g27682;
wire g30433;
wire g27102;
wire g32463;
wire g15165;
wire g31841;
wire g32971;
wire g13302;
wire g19772;
wire II29149;
wire g11997;
wire g23508;
wire g24865;
wire g25203;
wire g32165;
wire II30766;
wire g32616;
wire g21138;
wire g7063;
wire g18794;
wire gbuf113;
wire g15102;
wire g31785;
wire g10898;
wire II28588;
wire g13994;
wire g25026;
wire g24501;
wire g20510;
wire g21290;
wire g29170;
wire g19523;
wire g33595;
wire II17884;
wire g34215;
wire g28772;
wire g9180;
wire g18639;
wire II22792;
wire II17609;
wire g24508;
wire g13436;
wire g12114;
wire g7496;
wire g28986;
wire II23919;
wire II12204;
wire g24751;
wire g29586;
wire g12936;
wire g23420;
wire g16122;
wire g18351;
wire g27721;
wire g32826;
wire g15656;
wire g26160;
wire II32684;
wire g22060;
wire g24437;
wire g28347;
wire g23447;
wire II17590;
wire g25560;
wire g8450;
wire g16128;
wire g14391;
wire II18125;
wire g23777;
wire g22844;
wire g34680;
wire g19680;
wire II31221;
wire g30054;
wire g21962;
wire g20629;
wire g22072;
wire g30487;
wire g9099;
wire g7223;
wire g24931;
wire g26864;
wire g23401;
wire g28777;
wire g21816;
wire g24560;
wire g22189;
wire g30165;
wire g18150;
wire g16025;
wire g32409;
wire g33867;
wire gbuf104;
wire g28217;
wire g8561;
wire II23318;
wire g22311;
wire g29862;
wire g20230;
wire g25236;
wire g23581;
wire g22711;
wire g27451;
wire II12151;
wire g32565;
wire g27151;
wire g33904;
wire g11974;
wire II31874;
wire g10664;
wire g18781;
wire II23348;
wire g11280;
wire g24917;
wire g29197;
wire g32324;
wire g11153;
wire g24334;
wire g12019;
wire g32203;
wire g27203;
wire g24391;
wire g21862;
wire g26810;
wire II17496;
wire g26233;
wire g21555;
wire g8851;
wire g34415;
wire g17735;
wire g31813;
wire II19857;
wire g15904;
wire g14186;
wire g9662;
wire II22564;
wire g20982;
wire g25903;
wire II24438;
wire g32119;
wire g27727;
wire g18452;
wire g34070;
wire g34087;
wire II32758;
wire g28649;
wire II12761;
wire g15850;
wire g21949;
wire II16596;
wire g17780;
wire g29803;
wire g28114;
wire g32353;
wire g25617;
wire g29933;
wire g9614;
wire g27837;
wire g16885;
wire g33810;
wire g25381;
wire g30349;
wire g10671;
wire g12084;
wire g29688;
wire g30391;
wire g24364;
wire II24690;
wire g12189;
wire II31984;
wire II17355;
wire g19911;
wire II24700;
wire II31276;
wire II17744;
wire g28653;
wire II25743;
wire g6903;
wire g11735;
wire g30536;
wire g14831;
wire g21363;
wire g27343;
wire g27373;
wire g33270;
wire g9516;
wire g30562;
wire g29737;
wire g9968;
wire g31778;
wire g21344;
wire g11479;
wire g21466;
wire g32224;
wire g14587;
wire g22359;
wire g23303;
wire g18647;
wire g16222;
wire g26334;
wire g19854;
wire g25685;
wire g30335;
wire g9020;
wire g7649;
wire g33488;
wire g33294;
wire g18376;
wire g7109;
wire g24890;
wire g24939;
wire g11493;
wire II24576;
wire II33070;
wire g33784;
wire g24075;
wire g18109;
wire g34753;
wire g30496;
wire II31131;
wire g34018;
wire g24294;
wire g12646;
wire g33024;
wire g24718;
wire g31858;
wire g34402;
wire g28179;
wire g11036;
wire g17762;
wire g31892;
wire g20217;
wire II31042;
wire g32038;
wire II14734;
wire g13565;
wire II26439;
wire g8829;
wire g33590;
wire g34929;
wire g9334;
wire g27664;
wire g15064;
wire g25129;
wire g28475;
wire II31146;
wire g32046;
wire g15715;
wire g32907;
wire g32230;
wire g32551;
wire g7563;
wire g28867;
wire g25579;
wire g32515;
wire g29202;
wire g25449;
wire g27088;
wire g13706;
wire g23848;
wire II24674;
wire g29625;
wire g32935;
wire g17596;
wire g10142;
wire g11489;
wire g10421;
wire g21941;
wire g31286;
wire g27131;
wire g32580;
wire g11571;
wire g32517;
wire g9618;
wire II31659;
wire II22143;
wire g25836;
wire g34622;
wire g11941;
wire g11915;
wire g27351;
wire g27984;
wire g9779;
wire g33163;
wire II22470;
wire g7611;
wire g8181;
wire g29223;
wire g26766;
wire g11780;
wire g32148;
wire g16539;
wire g29637;
wire g9890;
wire g14313;
wire g24198;
wire g18682;
wire g34949;
wire II31810;
wire II24462;
wire g21728;
wire II24455;
wire g34648;
wire g31213;
wire g11607;
wire g30453;
wire II11726;
wire g26026;
wire g18345;
wire g23492;
wire g32822;
wire g23888;
wire g13058;
wire g18182;
wire II21226;
wire g32163;
wire II24278;
wire II30261;
wire g31789;
wire g31672;
wire g34003;
wire g15652;
wire g32218;
wire g28644;
wire g32729;
wire II22945;
wire g18776;
wire g19360;
wire g29842;
wire g10838;
wire g19266;
wire II30718;
wire g26483;
wire g30529;
wire g9104;
wire g28668;
wire II14516;
wire g34846;
wire g29798;
wire g14000;
wire g34226;
wire g7166;
wire g23008;
wire g8609;
wire g29902;
wire gbuf122;
wire g8594;
wire g27136;
wire g22129;
wire g22681;
wire g18133;
wire g7845;
wire II31727;
wire gbuf129;
wire g19644;
wire g24635;
wire g28286;
wire g25850;
wire II31770;
wire g26964;
wire g29747;
wire g12364;
wire g22853;
wire g13998;
wire II14923;
wire g31757;
wire g18626;
wire g32798;
wire g25111;
wire II32449;
wire II17314;
wire g29505;
wire g14093;
wire g34979;
wire g26226;
wire g24980;
wire g30212;
wire g6820;
wire g23354;
wire g8572;
wire g30138;
wire g20097;
wire II31071;
wire g30406;
wire g26842;
wire g33491;
wire g16349;
wire g20498;
wire g30171;
wire g26897;
wire II30123;
wire g24422;
wire g32946;
wire g29385;
wire g28958;
wire II17159;
wire II22755;
wire g33015;
wire g32660;
wire g11206;
wire g32749;
wire g25016;
wire g7994;
wire g25779;
wire g11988;
wire g21760;
wire g34655;
wire g15804;
wire II13382;
wire g29134;
wire g32449;
wire g34395;
wire g21421;
wire g25459;
wire g25653;
wire g18617;
wire g12249;
wire g25258;
wire g15669;
wire g32740;
wire II14570;
wire g14899;
wire g32156;
wire g15153;
wire g16291;
wire g12899;
wire g32732;
wire g28630;
wire II20462;
wire g24708;
wire g24299;
wire g12025;
wire II20954;
wire g22026;
wire II18633;
wire g25989;
wire g8346;
wire g9217;
wire g29324;
wire g29651;
wire g24028;
wire g13510;
wire g31327;
wire g32504;
wire g30918;
wire II25586;
wire g17846;
wire g22543;
wire II31820;
wire g28194;
wire g23575;
wire g20514;
wire g25703;
wire g25569;
wire g12035;
wire g26649;
wire g21359;
wire II17173;
wire g21348;
wire g22668;
wire g34432;
wire g28124;
wire II30740;
wire g24081;
wire g24994;
wire g27992;
wire g7980;
wire g19783;
wire II28851;
wire g9745;
wire g28247;
wire g26086;
wire II18135;
wire g33147;
wire g18457;
wire g23025;
wire g32624;
wire g27588;
wire g33820;
wire g14445;
wire g33814;
wire g19689;
wire g29650;
wire g16162;
wire II29233;
wire g31323;
wire g30566;
wire g29040;
wire g6928;
wire g30247;
wire II18681;
wire g25992;
wire g14681;
wire g29015;
wire g14515;
wire g33113;
wire II12218;
wire g34304;
wire g34495;
wire g20242;
wire g24585;
wire g34690;
wire g25962;
wire g8286;
wire g23858;
wire II22589;
wire g11398;
wire g13479;
wire g22537;
wire g22926;
wire g28637;
wire g12228;
wire g25056;
wire g27273;
wire g25700;
wire g31897;
wire g18752;
wire g34202;
wire g22069;
wire g24086;
wire g33892;
wire II22930;
wire g11123;
wire II29263;
wire g30095;
wire g11130;
wire g33587;
wire g24326;
wire II12468;
wire g8292;
wire g24258;
wire g18590;
wire II31474;
wire g32578;
wire g20505;
wire II15128;
wire g10812;
wire g19273;
wire II13862;
wire g26187;
wire II14790;
wire gbuf21;
wire g23864;
wire g17774;
wire g23816;
wire g32589;
wire g27434;
wire g26424;
wire II31046;
wire g29768;
wire g25765;
wire g30551;
wire g22093;
wire g11011;
wire g17520;
wire g31746;
wire g22984;
wire g26147;
wire g20774;
wire g28577;
wire g24290;
wire g17015;
wire II29981;
wire g33120;
wire g22688;
wire g18535;
wire g24269;
wire g29814;
wire g16842;
wire II13581;
wire g16643;
wire II24364;
wire g19521;
wire g22516;
wire g29989;
wire g24317;
wire g29967;
wire g13955;
wire g34800;
wire g14276;
wire II27238;
wire g19984;
wire g7888;
wire g18527;
wire g14720;
wire g20154;
wire g14177;
wire g21937;
wire g32264;
wire g18166;
wire g28592;
wire g24935;
wire g30549;
wire II15569;
wire II24331;
wire g32373;
wire g13933;
wire g31834;
wire g10883;
wire g33964;
wire g17763;
wire g25698;
wire g10601;
wire g21301;
wire g30067;
wire II27561;
wire g21975;
wire II22343;
wire II22180;
wire g11312;
wire II22972;
wire g30597;
wire g29486;
wire g28317;
wire II17650;
wire g11427;
wire g33640;
wire g34865;
wire g12461;
wire g15728;
wire g19865;
wire g19596;
wire g16178;
wire g24162;
wire g33314;
wire g8522;
wire g32050;
wire g18716;
wire g11497;
wire g33760;
wire g15752;
wire g22134;
wire g16246;
wire g23232;
wire g22487;
wire g26335;
wire g12357;
wire g33859;
wire g32296;
wire g32043;
wire g16299;
wire g31624;
wire g32679;
wire g18245;
wire g6867;
wire II26530;
wire g9229;
wire g32801;
wire g31945;
wire g7266;
wire g22450;
wire g28768;
wire g21802;
wire g31468;
wire g9880;
wire II13623;
wire g28133;
wire g24019;
wire g12119;
wire g28332;
wire g19393;
wire g10909;
wire g13289;
wire g33535;
wire g24667;
wire g6959;
wire g12042;
wire g21401;
wire g19556;
wire g16592;
wire g33455;
wire g34855;
wire g29889;
wire g33197;
wire g29519;
wire g31843;
wire g7858;
wire g33647;
wire g23258;
wire g12881;
wire g33712;
wire g25293;
wire g31994;
wire II33232;
wire g27376;
wire g12295;
wire g17010;
wire g27501;
wire g13919;
wire g13029;
wire gbuf32;
wire gbuf48;
wire g16476;
wire II29199;
wire g14707;
wire g23375;
wire g10623;
wire g9730;
wire g13823;
wire g18483;
wire g18088;
wire g11449;
wire gbuf28;
wire II23375;
wire II28925;
wire g22529;
wire g25926;
wire g33289;
wire g7343;
wire g10412;
wire g21757;
wire II22000;
wire II24759;
wire g34198;
wire gbuf87;
wire II15004;
wire g15138;
wire g21416;
wire g15344;
wire g21893;
wire g15097;
wire g7917;
wire g22150;
wire g28998;
wire g28699;
wire g14216;
wire g32018;
wire g31314;
wire g11846;
wire g16522;
wire g23058;
wire II23384;
wire g12471;
wire g16053;
wire II20116;
wire g10573;
wire g11252;
wire g18307;
wire g24504;
wire g33993;
wire g33449;
wire g33136;
wire g34058;
wire g26878;
wire II27749;
wire g24981;
wire g22227;
wire g32361;
wire gbuf154;
wire g29730;
wire g30671;
wire II29939;
wire g31857;
wire g27771;
wire g25729;
wire g17419;
wire g23868;
wire g21829;
wire g7369;
wire g24036;
wire g32899;
wire g10178;
wire g27364;
wire g33394;
wire g25173;
wire g34627;
wire g18721;
wire g20452;
wire g25523;
wire g16676;
wire g33440;
wire g28685;
wire g25761;
wire g32974;
wire gbuf140;
wire g22761;
wire g33850;
wire g13121;
wire g29298;
wire g23248;
wire g14347;
wire g14640;
wire g13035;
wire g21781;
wire II11716;
wire g28512;
wire gbuf59;
wire g34500;
wire g15074;
wire g24057;
wire g15678;
wire g12641;
wire g12821;
wire g28232;
wire g8405;
wire g19495;
wire g31639;
wire g21874;
wire g26347;
wire g29884;
wire g34448;
wire II33027;
wire g14921;
wire g31516;
wire g14546;
wire g10388;
wire g21670;
wire II21941;
wire g33254;
wire g15588;
wire g34119;
wire g30198;
wire g18749;
wire g28079;
wire g34982;
wire II29579;
wire II24508;
wire g18930;
wire g26852;
wire g6811;
wire g12976;
wire g17125;
wire g23678;
wire g8770;
wire g26182;
wire g18238;
wire g31069;
wire g28152;
wire g16599;
wire II14409;
wire g24757;
wire g31297;
wire g24773;
wire g19768;
wire g13907;
wire g12543;
wire g18512;
wire g34266;
wire g30144;
wire g24574;
wire g31520;
wire g23896;
wire g19577;
wire g11317;
wire g20040;
wire g34429;
wire g33359;
wire g15081;
wire g17312;
wire g8093;
wire g8300;
wire g25714;
wire g27796;
wire g34957;
wire g18222;
wire g29474;
wire g11888;
wire g6998;
wire g29570;
wire g21186;
wire g32249;
wire g21294;
wire g7517;
wire g26940;
wire II31106;
wire II18323;
wire g19493;
wire II31231;
wire II26095;
wire g30297;
wire g15088;
wire II29441;
wire g19482;
wire g23414;
wire g24491;
wire g23823;
wire g11283;
wire g17576;
wire g18815;
wire g12778;
wire g30244;
wire g25246;
wire g33928;
wire g25534;
wire g31241;
wire g17656;
wire g26671;
wire g11294;
wire g8792;
wire II31597;
wire g15103;
wire g10796;
wire g30101;
wire g17603;
wire g24671;
wire g11920;
wire g18442;
wire g24964;
wire g23477;
wire g25212;
wire g33884;
wire g31149;
wire g13133;
wire g27391;
wire g25079;
wire g14590;
wire g22995;
wire g23273;
wire g34984;
wire g29760;
wire g16959;
wire II15255;
wire g25631;
wire II15149;
wire g19653;
wire II12729;
wire g11753;
wire g23237;
wire g12755;
wire g18212;
wire g21279;
wire g29056;
wire g33574;
wire g22130;
wire g13929;
wire g29187;
wire g17926;
wire g14780;
wire g9280;
wire g13260;
wire II20753;
wire g26249;
wire g19657;
wire g29576;
wire II16741;
wire g28522;
wire g21990;
wire g14510;
wire II29913;
wire g24748;
wire g28227;
wire II13424;
wire g30289;
wire g29285;
wire g22172;
wire g18759;
wire g23132;
wire g22049;
wire II31361;
wire II22425;
wire g18410;
wire g9024;
wire II29313;
wire g29167;
wire g30591;
wire g27599;
wire g27238;
wire g8538;
wire g23239;
wire g26351;
wire g34285;
wire II15121;
wire g25076;
wire g18420;
wire g19200;
wire g29343;
wire g12219;
wire g7133;
wire g16430;
wire g29708;
wire g22097;
wire II14567;
wire g9250;
wire g17490;
wire g30135;
wire g23435;
wire g23695;
wire II14205;
wire II13606;
wire II31302;
wire II19786;
wire g23946;
wire g7870;
wire g25944;
wire g32311;
wire g19374;
wire g24660;
wire g23151;
wire g22884;
wire g18678;
wire g29307;
wire g10567;
wire II25219;
wire II17976;
wire g29275;
wire g10116;
wire g23319;
wire g32607;
wire g16782;
wire g21336;
wire g19466;
wire g28063;
wire g23014;
wire g32333;
wire g10654;
wire g17754;
wire g24555;
wire g10093;
wire II18434;
wire g27158;
wire II14727;
wire g26575;
wire g23938;
wire II12523;
wire g34522;
wire II29253;
wire g10590;
wire g13833;
wire g11303;
wire g9687;
wire II17148;
wire g17746;
wire g25574;
wire g22872;
wire g34729;
wire g22062;
wire II20488;
wire g25051;
wire g15566;
wire g8285;
wire g34463;
wire g24152;
wire II11825;
wire g11003;
wire g16320;
wire g25410;
wire g21742;
wire II11801;
wire g6808;
wire g30533;
wire g31493;
wire II17166;
wire II18089;
wire g28585;
wire g18918;
wire g29338;
wire g30339;
wire g28572;
wire II13057;
wire II32763;
wire g25420;
wire g18267;
wire gbuf80;
wire g34459;
wire II24237;
wire g25882;
wire g22113;
wire g34241;
wire g8085;
wire g17690;
wire g34703;
wire g21765;
wire II12884;
wire g7072;
wire g24892;
wire g23780;
wire g18651;
wire g22542;
wire g19743;
wire g33238;
wire g32577;
wire g16227;
wire g29068;
wire g33803;
wire g11044;
wire g14232;
wire g31922;
wire g19434;
wire g28672;
wire g18293;
wire g24071;
wire g33228;
wire g22991;
wire g26382;
wire g21912;
wire g12845;
wire g24534;
wire g12001;
wire g10198;
wire II26644;
wire g30600;
wire g28031;
wire g28752;
wire g18381;
wire g18205;
wire g23418;
wire g18463;
wire g24643;
wire g13239;
wire II12631;
wire g27313;
wire g29621;
wire II15299;
wire II13694;
wire g14069;
wire g8038;
wire II18104;
wire g25100;
wire II17456;
wire II15937;
wire g10336;
wire II12418;
wire II19802;
wire II14399;
wire II15080;
wire g25943;
wire II17964;
wire g30201;
wire II13705;
wire g16487;
wire II29977;
wire g25622;
wire g7952;
wire g9826;
wire g24000;
wire g24516;
wire g25273;
wire g29645;
wire g33060;
wire g21228;
wire g20200;
wire g27179;
wire g23566;
wire g23928;
wire g13414;
wire g14638;
wire g8914;
wire g28427;
wire g30237;
wire II29262;
wire g23820;
wire II31803;
wire g14361;
wire g27406;
wire II32956;
wire g20107;
wire g12945;
wire g31963;
wire g12951;
wire g24046;
wire II11734;
wire g29978;
wire g11323;
wire g20584;
wire g34480;
wire g25271;
wire g11118;
wire g24250;
wire g23747;
wire g20112;
wire g18772;
wire g16171;
wire g34387;
wire g25736;
wire g26399;
wire g32391;
wire g31238;
wire g14088;
wire II23962;
wire g29697;
wire g25724;
wire g34034;
wire g25604;
wire g29920;
wire g32071;
wire g34658;
wire g21866;
wire g12521;
wire g21606;
wire gbuf132;
wire g22898;
wire g33571;
wire g13594;
wire g13496;
wire g14696;
wire g21997;
wire g20500;
wire g33029;
wire II29444;
wire g13143;
wire g29476;
wire gbuf149;
wire g33323;
wire g34926;
wire g23719;
wire g16723;
wire g18479;
wire g11747;
wire g23260;
wire g25780;
wire g20545;
wire g24228;
wire g18693;
wire g28368;
wire g27734;
wire II20388;
wire g20073;
wire g12129;
wire g8650;
wire g7503;
wire g25120;
wire g20661;
wire g34938;
wire g22084;
wire g27187;
wire g18890;
wire II13751;
wire g34836;
wire gbuf58;
wire g13100;
wire g6772;
wire g28823;
wire g33601;
wire g31991;
wire g26653;
wire g32695;
wire g21252;
wire g30557;
wire g34786;
wire g25552;
wire g10966;
wire g7446;
wire g30381;
wire g23554;
wire g21061;
wire g21919;
wire g15860;
wire II15175;
wire g9733;
wire II15238;
wire g9693;
wire g16667;
wire g13943;
wire g18780;
wire g19690;
wire g31302;
wire g12805;
wire g31596;
wire g11912;
wire g23906;
wire g32532;
wire g32341;
wire g24713;
wire g19632;
wire g7659;
wire g30153;
wire g27486;
wire g11985;
wire II15788;
wire II33143;
wire g22653;
wire g13188;
wire g10409;
wire g10404;
wire g18149;
wire g28618;
wire g24836;
wire g16703;
wire g15704;
wire g17134;
wire g19906;
wire g10398;
wire g31227;
wire g31591;
wire g24369;
wire II31786;
wire II30468;
wire g9018;
wire g16896;
wire g33473;
wire II32601;
wire g31501;
wire g32190;
wire g13094;
wire g8136;
wire g25284;
wire g33744;
wire g13335;
wire g28182;
wire g8933;
wire g33074;
wire g26939;
wire g19443;
wire g20630;
wire g25222;
wire g24976;
wire g34043;
wire g33538;
wire g25636;
wire g32288;
wire II12411;
wire g11903;
wire g27738;
wire II14671;
wire II15148;
wire g9954;
wire g26051;
wire g26268;
wire g11164;
wire g34997;
wire g32919;
wire II31037;
wire g13655;
wire g27291;
wire g34631;
wire g30424;
wire g12009;
wire g13384;
wire g31779;
wire g22904;
wire g22190;
wire g9976;
wire II33276;
wire g23517;
wire II20223;
wire g31763;
wire g31306;
wire g17499;
wire g24065;
wire g26279;
wire g27699;
wire g15910;
wire g12749;
wire g22156;
wire II22665;
wire g29092;
wire g18197;
wire g25506;
wire g26759;
wire II31091;
wire g23298;
wire g33044;
wire g21772;
wire g9910;
wire g8506;
wire g22331;
wire g10130;
wire g24345;
wire g17137;
wire g24375;
wire g12944;
wire g21739;
wire g33414;
wire g34337;
wire g26715;
wire g33277;
wire g27426;
wire g10129;
wire g26830;
wire II29371;
wire II18301;
wire g17479;
wire g34424;
wire g13664;
wire g25230;
wire g15967;
wire g14382;
wire II31207;
wire g26511;
wire g21790;
wire g24924;
wire g24907;
wire g11560;
wire g28293;
wire g19050;
wire g24401;
wire g24900;
wire g29304;
wire g18819;
wire g8672;
wire g34538;
wire g23802;
wire II17857;
wire g32415;
wire g34292;
wire g11861;
wire g30222;
wire II16639;
wire g27722;
wire II12016;
wire g7542;
wire II28480;
wire g28210;
wire g7618;
wire g24319;
wire g12590;
wire II31974;
wire g34063;
wire g9543;
wire g34513;
wire g14227;
wire g34903;
wire g21690;
wire g33699;
wire g23982;
wire g14123;
wire g21794;
wire g30068;
wire g23139;
wire g13973;
wire II32976;
wire g34358;
wire g33817;
wire g30037;
wire g33846;
wire g27180;
wire g20924;
wire g31904;
wire g6997;
wire g29314;
wire g33879;
wire II23303;
wire g24758;
wire II20467;
wire g33617;
wire g25803;
wire II18224;
wire g26305;
wire g13986;
wire g31273;
wire g23837;
wire g20188;
wire g31194;
wire g30092;
wire g9657;
wire II30901;
wire II27533;
wire g17145;
wire g14136;
wire g32756;
wire g23026;
wire g34223;
wire g16758;
wire g28167;
wire g34277;
wire g26811;
wire g34724;
wire II23327;
wire g21747;
wire g26631;
wire g31851;
wire g22990;
wire g30473;
wire g29783;
wire g32248;
wire g18287;
wire g19575;
wire g9637;
wire g33105;
wire II31316;
wire g32865;
wire g29114;
wire II14713;
wire g31290;
wire g27336;
wire g12840;
wire g10704;
wire g31258;
wire g34373;
wire g21753;
wire g23111;
wire g30304;
wire g34025;
wire g24351;
wire g11025;
wire g33731;
wire g20541;
wire g32318;
wire II31226;
wire g28240;
wire g13191;
wire g30429;
wire g24183;
wire g13107;
wire g26280;
wire g34100;
wire g18807;
wire g33797;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g72 <= 0;
  else
    g72 <= g24166;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g73 <= 0;
  else
    g73 <= g24167;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g84 <= 0;
  else
    g84 <= g24168;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g90 <= 0;
  else
    g90 <= g24169;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g91 <= 0;
  else
    g91 <= g24170;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g92 <= 0;
  else
    g92 <= g24171;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g99 <= 0;
  else
    g99 <= g24172;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g100 <= 0;
  else
    g100 <= g24173;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g110 <= 0;
  else
    g110 <= g34848;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g112 <= 0;
  else
    g112 <= g34879;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g113 <= 0;
  else
    g113 <= g24174;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g114 <= 0;
  else
    g114 <= g24175;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g115 <= 0;
  else
    g115 <= g24176;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g116 <= 0;
  else
    g116 <= g24177;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g120 <= 0;
  else
    g120 <= g24178;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g124 <= 0;
  else
    g124 <= g24179;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g125 <= 0;
  else
    g125 <= g24180;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g126 <= 0;
  else
    g126 <= g24181;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g127 <= 0;
  else
    g127 <= g24182;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g134 <= 0;
  else
    g134 <= g24183;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g135 <= 0;
  else
    g135 <= g24184;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g44 <= 0;
  else
    g44 <= g24185;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g45 <= 0;
  else
    g45 <= g34990;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g46 <= 0;
  else
    g46 <= g34991;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g47 <= 0;
  else
    g47 <= g34992;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g48 <= 0;
  else
    g48 <= g34993;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g49 <= 0;
  else
    g49 <= g34994;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g50 <= 0;
  else
    g50 <= g34995;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g51 <= 0;
  else
    g51 <= g34996;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g52 <= 0;
  else
    g52 <= g34997;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g53 <= 0;
  else
    g53 <= g24161;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g54 <= 0;
  else
    g54 <= g24162;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g55 <= 0;
  else
    g55 <= g35002;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g56 <= 0;
  else
    g56 <= g24163;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g57 <= 0;
  else
    g57 <= g24164;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g58 <= 0;
  else
    g58 <= g30328;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g63 <= 0;
  else
    g63 <= g34847;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g71 <= 0;
  else
    g71 <= g34786;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g85 <= 0;
  else
    g85 <= g34717;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g93 <= 0;
  else
    g93 <= g34878;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g101 <= 0;
  else
    g101 <= g34787;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g111 <= 0;
  else
    g111 <= g34718;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g43 <= 0;
  else
    g43 <= g34789;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g64 <= 0;
  else
    g64 <= g24165;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g65 <= 0;
  else
    g65 <= g34785;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g70 <= 0;
  else
    g70 <= g18093;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4507 <= 0;
  else
    g4507 <= g30458;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4459 <= 0;
  else
    g4459 <= g34253;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4369 <= 0;
  else
    g4369 <= g26970;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4473 <= 0;
  else
    g4473 <= g34256;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4462 <= 0;
  else
    g4462 <= g34254;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4581 <= 0;
  else
    g4581 <= g26969;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4467 <= 0;
  else
    g4467 <= g34255;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4474 <= 0;
  else
    g4474 <= g10384;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4477 <= 0;
  else
    g4477 <= g26960;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4480 <= 0;
  else
    g4480 <= g31896;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4495 <= 0;
  else
    g4495 <= g33036;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4498 <= 0;
  else
    g4498 <= g33037;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4501 <= 0;
  else
    g4501 <= g33038;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4504 <= 0;
  else
    g4504 <= g33039;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4512 <= 0;
  else
    g4512 <= g33040;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4521 <= 0;
  else
    g4521 <= g26971;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4527 <= 0;
  else
    g4527 <= g28082;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4515 <= 0;
  else
    g4515 <= g26964;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4519 <= 0;
  else
    g4519 <= g33616;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4520 <= 0;
  else
    g4520 <= g6972;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4483 <= 0;
  else
    g4483 <= gbuf1;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4486 <= 0;
  else
    g4486 <= g26961;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4489 <= 0;
  else
    g4489 <= g26962;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4492 <= 0;
  else
    g4492 <= g26963;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4537 <= 0;
  else
    g4537 <= g34024;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4423 <= 0;
  else
    g4423 <= gbuf2;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4540 <= 0;
  else
    g4540 <= g31897;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4543 <= 0;
  else
    g4543 <= g33042;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4567 <= 0;
  else
    g4567 <= g33043;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4546 <= 0;
  else
    g4546 <= g33045;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4549 <= 0;
  else
    g4549 <= g33041;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4552 <= 0;
  else
    g4552 <= g33044;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4570 <= 0;
  else
    g4570 <= g33617;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4571 <= 0;
  else
    g4571 <= g6974;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4555 <= 0;
  else
    g4555 <= gbuf3;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4558 <= 0;
  else
    g4558 <= g26966;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4561 <= 0;
  else
    g4561 <= g26968;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4564 <= 0;
  else
    g4564 <= g26967;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4534 <= 0;
  else
    g4534 <= g34023;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4420 <= 0;
  else
    g4420 <= g26965;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4438 <= 0;
  else
    g4438 <= g26953;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4449 <= 0;
  else
    g4449 <= g26955;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4443 <= 0;
  else
    g4443 <= gbuf4;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4446 <= 0;
  else
    g4446 <= g26954;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4452 <= 0;
  else
    g4452 <= gbuf5;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4434 <= 0;
  else
    g4434 <= g26956;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4430 <= 0;
  else
    g4430 <= g26957;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4427 <= 0;
  else
    g4427 <= g26952;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4375 <= 0;
  else
    g4375 <= g26951;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4414 <= 0;
  else
    g4414 <= g26946;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4411 <= 0;
  else
    g4411 <= gbuf6;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4408 <= 0;
  else
    g4408 <= g26945;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4405 <= 0;
  else
    g4405 <= gbuf7;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4401 <= 0;
  else
    g4401 <= g26948;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4388 <= 0;
  else
    g4388 <= g26949;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4382 <= 0;
  else
    g4382 <= g26947;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4417 <= 0;
  else
    g4417 <= g31895;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4392 <= 0;
  else
    g4392 <= g26950;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4456 <= 0;
  else
    g4456 <= g25692;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4455 <= 0;
  else
    g4455 <= g26959;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1 <= 0;
  else
    g1 <= g26958;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4304 <= 0;
  else
    g4304 <= g24281;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4308 <= 0;
  else
    g4308 <= gbuf8;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2932 <= 0;
  else
    g2932 <= g24282;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4639 <= 0;
  else
    g4639 <= g34025;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4621 <= 0;
  else
    g4621 <= g34460;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4628 <= 0;
  else
    g4628 <= g34457;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4633 <= 0;
  else
    g4633 <= g34458;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4643 <= 0;
  else
    g4643 <= g34259;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4340 <= 0;
  else
    g4340 <= g34459;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4349 <= 0;
  else
    g4349 <= g34257;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4358 <= 0;
  else
    g4358 <= g34258;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g66 <= 0;
  else
    g66 <= g24334;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4531 <= 0;
  else
    g4531 <= g24335;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4311 <= 0;
  else
    g4311 <= g34449;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4322 <= 0;
  else
    g4322 <= g34450;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4332 <= 0;
  else
    g4332 <= g34455;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4584 <= 0;
  else
    g4584 <= g34451;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4593 <= 0;
  else
    g4593 <= g34452;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4601 <= 0;
  else
    g4601 <= g34453;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4608 <= 0;
  else
    g4608 <= g34454;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4616 <= 0;
  else
    g4616 <= g34456;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4366 <= 0;
  else
    g4366 <= g26944;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4372 <= 0;
  else
    g4372 <= g34882;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4836 <= 0;
  else
    g4836 <= g34265;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4864 <= 0;
  else
    g4864 <= g34034;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4871 <= 0;
  else
    g4871 <= g34035;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4878 <= 0;
  else
    g4878 <= g34036;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4843 <= 0;
  else
    g4843 <= g34466;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4849 <= 0;
  else
    g4849 <= g34465;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4854 <= 0;
  else
    g4854 <= g34467;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4859 <= 0;
  else
    g4859 <= g34468;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4917 <= 0;
  else
    g4917 <= g34638;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4922 <= 0;
  else
    g4922 <= g34639;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4907 <= 0;
  else
    g4907 <= g34640;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4912 <= 0;
  else
    g4912 <= g34641;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4927 <= 0;
  else
    g4927 <= g34642;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4931 <= 0;
  else
    g4931 <= g21904;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4932 <= 0;
  else
    g4932 <= g21905;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4572 <= 0;
  else
    g4572 <= g29279;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4578 <= 0;
  else
    g4578 <= g29278;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4999 <= 0;
  else
    g4999 <= g25694;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5002 <= 0;
  else
    g5002 <= gbuf9;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5005 <= 0;
  else
    g5005 <= gbuf10;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5008 <= 0;
  else
    g5008 <= gbuf11;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4983 <= 0;
  else
    g4983 <= g34041;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4991 <= 0;
  else
    g4991 <= g34038;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4966 <= 0;
  else
    g4966 <= g34039;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4975 <= 0;
  else
    g4975 <= g34037;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4899 <= 0;
  else
    g4899 <= g34040;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4894 <= 0;
  else
    g4894 <= g28087;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4888 <= 0;
  else
    g4888 <= g34266;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4939 <= 0;
  else
    g4939 <= g28088;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4933 <= 0;
  else
    g4933 <= g34267;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4950 <= 0;
  else
    g4950 <= g28089;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4944 <= 0;
  else
    g4944 <= g34268;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4961 <= 0;
  else
    g4961 <= g28090;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4955 <= 0;
  else
    g4955 <= g34269;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4646 <= 0;
  else
    g4646 <= g34260;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4674 <= 0;
  else
    g4674 <= g34026;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4681 <= 0;
  else
    g4681 <= g34027;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4688 <= 0;
  else
    g4688 <= g34028;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4653 <= 0;
  else
    g4653 <= g34462;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4659 <= 0;
  else
    g4659 <= g34461;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4664 <= 0;
  else
    g4664 <= g34463;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4669 <= 0;
  else
    g4669 <= g34464;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4727 <= 0;
  else
    g4727 <= g34633;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4732 <= 0;
  else
    g4732 <= g34634;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4717 <= 0;
  else
    g4717 <= g34635;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4722 <= 0;
  else
    g4722 <= g34636;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4737 <= 0;
  else
    g4737 <= g34637;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4741 <= 0;
  else
    g4741 <= g21902;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4742 <= 0;
  else
    g4742 <= g21903;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g59 <= 0;
  else
    g59 <= g29277;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4575 <= 0;
  else
    g4575 <= g29276;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4809 <= 0;
  else
    g4809 <= g25693;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4812 <= 0;
  else
    g4812 <= gbuf12;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4815 <= 0;
  else
    g4815 <= gbuf13;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4818 <= 0;
  else
    g4818 <= gbuf14;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4793 <= 0;
  else
    g4793 <= g34033;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4801 <= 0;
  else
    g4801 <= g34030;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4776 <= 0;
  else
    g4776 <= g34031;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4785 <= 0;
  else
    g4785 <= g34029;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4709 <= 0;
  else
    g4709 <= g34032;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4704 <= 0;
  else
    g4704 <= g28083;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4698 <= 0;
  else
    g4698 <= g34261;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4749 <= 0;
  else
    g4749 <= g28084;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4743 <= 0;
  else
    g4743 <= g34262;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4760 <= 0;
  else
    g4760 <= g28085;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4754 <= 0;
  else
    g4754 <= g34263;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4771 <= 0;
  else
    g4771 <= g28086;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4765 <= 0;
  else
    g4765 <= g34264;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5313 <= 0;
  else
    g5313 <= g24336;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5290 <= 0;
  else
    g5290 <= gbuf15;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5320 <= 0;
  else
    g5320 <= gbuf16;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5276 <= 0;
  else
    g5276 <= gbuf17;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5283 <= 0;
  else
    g5283 <= gbuf18;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5308 <= 0;
  else
    g5308 <= gbuf19;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5327 <= 0;
  else
    g5327 <= gbuf20;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5331 <= 0;
  else
    g5331 <= gbuf21;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5335 <= 0;
  else
    g5335 <= gbuf22;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5339 <= 0;
  else
    g5339 <= gbuf23;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5343 <= 0;
  else
    g5343 <= g24337;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5348 <= 0;
  else
    g5348 <= g24338;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5352 <= 0;
  else
    g5352 <= g24339;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5357 <= 0;
  else
    g5357 <= g33618;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5297 <= 0;
  else
    g5297 <= g33619;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5101 <= 0;
  else
    g5101 <= g25700;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5109 <= 0;
  else
    g5109 <= gbuf24;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5062 <= 0;
  else
    g5062 <= g25702;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5105 <= 0;
  else
    g5105 <= g25701;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5112 <= 0;
  else
    g5112 <= gbuf25;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5022 <= 0;
  else
    g5022 <= g25703;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5016 <= 0;
  else
    g5016 <= g31898;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5029 <= 0;
  else
    g5029 <= g31902;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5033 <= 0;
  else
    g5033 <= g31904;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5037 <= 0;
  else
    g5037 <= g31899;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5041 <= 0;
  else
    g5041 <= g31900;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5046 <= 0;
  else
    g5046 <= g31901;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5052 <= 0;
  else
    g5052 <= g31903;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5057 <= 0;
  else
    g5057 <= g33046;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5069 <= 0;
  else
    g5069 <= g28092;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5073 <= 0;
  else
    g5073 <= g28091;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5077 <= 0;
  else
    g5077 <= g25704;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5080 <= 0;
  else
    g5080 <= g25695;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5084 <= 0;
  else
    g5084 <= g25696;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5092 <= 0;
  else
    g5092 <= g25697;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5097 <= 0;
  else
    g5097 <= g25698;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g86 <= 0;
  else
    g86 <= g25699;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5164 <= 0;
  else
    g5164 <= g30459;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5170 <= 0;
  else
    g5170 <= g33047;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5176 <= 0;
  else
    g5176 <= g33048;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5180 <= 0;
  else
    g5180 <= g33049;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5188 <= 0;
  else
    g5188 <= g33050;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5196 <= 0;
  else
    g5196 <= g30460;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5224 <= 0;
  else
    g5224 <= g30464;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5240 <= 0;
  else
    g5240 <= g30468;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5256 <= 0;
  else
    g5256 <= g30472;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5204 <= 0;
  else
    g5204 <= g30476;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5200 <= 0;
  else
    g5200 <= g30461;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5228 <= 0;
  else
    g5228 <= g30465;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5244 <= 0;
  else
    g5244 <= g30469;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5260 <= 0;
  else
    g5260 <= g30473;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5212 <= 0;
  else
    g5212 <= g30477;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5208 <= 0;
  else
    g5208 <= g30462;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5232 <= 0;
  else
    g5232 <= g30466;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5248 <= 0;
  else
    g5248 <= g30470;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5264 <= 0;
  else
    g5264 <= g30474;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5220 <= 0;
  else
    g5220 <= g30478;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5216 <= 0;
  else
    g5216 <= g30463;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5236 <= 0;
  else
    g5236 <= g30467;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5252 <= 0;
  else
    g5252 <= g30471;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5268 <= 0;
  else
    g5268 <= g30475;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5272 <= 0;
  else
    g5272 <= g30479;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g128 <= 0;
  else
    g128 <= g28093;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5156 <= 0;
  else
    g5156 <= g29285;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5120 <= 0;
  else
    g5120 <= g25708;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5115 <= 0;
  else
    g5115 <= g29280;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5124 <= 0;
  else
    g5124 <= g29281;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5128 <= 0;
  else
    g5128 <= g25705;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5134 <= 0;
  else
    g5134 <= g29282;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5138 <= 0;
  else
    g5138 <= g29283;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5142 <= 0;
  else
    g5142 <= g29284;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5148 <= 0;
  else
    g5148 <= g25706;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5152 <= 0;
  else
    g5152 <= g25707;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5160 <= 0;
  else
    g5160 <= g34643;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5659 <= 0;
  else
    g5659 <= g24340;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5637 <= 0;
  else
    g5637 <= gbuf26;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5666 <= 0;
  else
    g5666 <= gbuf27;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5623 <= 0;
  else
    g5623 <= gbuf28;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5630 <= 0;
  else
    g5630 <= gbuf29;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5654 <= 0;
  else
    g5654 <= gbuf30;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5673 <= 0;
  else
    g5673 <= gbuf31;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5677 <= 0;
  else
    g5677 <= gbuf32;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5681 <= 0;
  else
    g5681 <= gbuf33;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5685 <= 0;
  else
    g5685 <= gbuf34;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5689 <= 0;
  else
    g5689 <= g24341;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5694 <= 0;
  else
    g5694 <= g24342;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5698 <= 0;
  else
    g5698 <= g24343;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5703 <= 0;
  else
    g5703 <= g33620;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5644 <= 0;
  else
    g5644 <= g33621;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5448 <= 0;
  else
    g5448 <= g25714;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5456 <= 0;
  else
    g5456 <= gbuf35;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5406 <= 0;
  else
    g5406 <= g25716;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5452 <= 0;
  else
    g5452 <= g25715;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5459 <= 0;
  else
    g5459 <= gbuf36;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5366 <= 0;
  else
    g5366 <= g25717;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5360 <= 0;
  else
    g5360 <= g31905;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5373 <= 0;
  else
    g5373 <= g31909;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5377 <= 0;
  else
    g5377 <= g31911;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5381 <= 0;
  else
    g5381 <= g31906;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5385 <= 0;
  else
    g5385 <= g31907;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5390 <= 0;
  else
    g5390 <= g31908;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5396 <= 0;
  else
    g5396 <= g31910;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5401 <= 0;
  else
    g5401 <= g33051;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5413 <= 0;
  else
    g5413 <= g28095;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5417 <= 0;
  else
    g5417 <= g28094;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5421 <= 0;
  else
    g5421 <= g25718;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5424 <= 0;
  else
    g5424 <= g25709;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5428 <= 0;
  else
    g5428 <= g25710;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5436 <= 0;
  else
    g5436 <= g25711;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5441 <= 0;
  else
    g5441 <= g25712;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5445 <= 0;
  else
    g5445 <= g25713;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5511 <= 0;
  else
    g5511 <= g30480;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5517 <= 0;
  else
    g5517 <= g33052;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5523 <= 0;
  else
    g5523 <= g33053;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5527 <= 0;
  else
    g5527 <= g33054;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5535 <= 0;
  else
    g5535 <= g33055;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5543 <= 0;
  else
    g5543 <= g30481;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5571 <= 0;
  else
    g5571 <= g30485;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5587 <= 0;
  else
    g5587 <= g30489;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5603 <= 0;
  else
    g5603 <= g30493;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5551 <= 0;
  else
    g5551 <= g30497;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5547 <= 0;
  else
    g5547 <= g30482;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5575 <= 0;
  else
    g5575 <= g30486;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5591 <= 0;
  else
    g5591 <= g30490;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5607 <= 0;
  else
    g5607 <= g30494;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5559 <= 0;
  else
    g5559 <= g30498;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5555 <= 0;
  else
    g5555 <= g30483;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5579 <= 0;
  else
    g5579 <= g30487;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5595 <= 0;
  else
    g5595 <= g30491;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5611 <= 0;
  else
    g5611 <= g30495;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5567 <= 0;
  else
    g5567 <= g30499;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5563 <= 0;
  else
    g5563 <= g30484;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5583 <= 0;
  else
    g5583 <= g30488;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5599 <= 0;
  else
    g5599 <= g30492;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5615 <= 0;
  else
    g5615 <= g30496;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5619 <= 0;
  else
    g5619 <= g30500;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4821 <= 0;
  else
    g4821 <= g28096;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5503 <= 0;
  else
    g5503 <= g29291;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5467 <= 0;
  else
    g5467 <= g25722;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5462 <= 0;
  else
    g5462 <= g29286;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5471 <= 0;
  else
    g5471 <= g29287;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5475 <= 0;
  else
    g5475 <= g25719;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5481 <= 0;
  else
    g5481 <= g29288;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5485 <= 0;
  else
    g5485 <= g29289;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5489 <= 0;
  else
    g5489 <= g29290;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5495 <= 0;
  else
    g5495 <= g25720;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5499 <= 0;
  else
    g5499 <= g25721;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5507 <= 0;
  else
    g5507 <= g34644;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6005 <= 0;
  else
    g6005 <= g24344;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5983 <= 0;
  else
    g5983 <= gbuf37;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6012 <= 0;
  else
    g6012 <= gbuf38;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5969 <= 0;
  else
    g5969 <= gbuf39;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5976 <= 0;
  else
    g5976 <= gbuf40;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6000 <= 0;
  else
    g6000 <= gbuf41;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6019 <= 0;
  else
    g6019 <= gbuf42;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6023 <= 0;
  else
    g6023 <= gbuf43;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6027 <= 0;
  else
    g6027 <= gbuf44;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6031 <= 0;
  else
    g6031 <= gbuf45;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6035 <= 0;
  else
    g6035 <= g24345;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6040 <= 0;
  else
    g6040 <= g24346;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6044 <= 0;
  else
    g6044 <= g24347;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6049 <= 0;
  else
    g6049 <= g33622;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5990 <= 0;
  else
    g5990 <= g33623;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5794 <= 0;
  else
    g5794 <= g25728;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5802 <= 0;
  else
    g5802 <= gbuf46;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5752 <= 0;
  else
    g5752 <= g25730;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5798 <= 0;
  else
    g5798 <= g25729;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5805 <= 0;
  else
    g5805 <= gbuf47;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5712 <= 0;
  else
    g5712 <= g25731;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5706 <= 0;
  else
    g5706 <= g31912;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5719 <= 0;
  else
    g5719 <= g31916;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5723 <= 0;
  else
    g5723 <= g31918;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5727 <= 0;
  else
    g5727 <= g31913;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5731 <= 0;
  else
    g5731 <= g31914;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5736 <= 0;
  else
    g5736 <= g31915;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5742 <= 0;
  else
    g5742 <= g31917;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5747 <= 0;
  else
    g5747 <= g33056;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5759 <= 0;
  else
    g5759 <= g28098;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5763 <= 0;
  else
    g5763 <= g28097;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5767 <= 0;
  else
    g5767 <= g25732;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5770 <= 0;
  else
    g5770 <= g25723;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5774 <= 0;
  else
    g5774 <= g25724;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5782 <= 0;
  else
    g5782 <= g25725;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5787 <= 0;
  else
    g5787 <= g25726;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5791 <= 0;
  else
    g5791 <= g25727;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5857 <= 0;
  else
    g5857 <= g30501;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5863 <= 0;
  else
    g5863 <= g33057;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5869 <= 0;
  else
    g5869 <= g33058;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5873 <= 0;
  else
    g5873 <= g33059;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5881 <= 0;
  else
    g5881 <= g33060;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5889 <= 0;
  else
    g5889 <= g30502;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5917 <= 0;
  else
    g5917 <= g30506;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5933 <= 0;
  else
    g5933 <= g30510;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5949 <= 0;
  else
    g5949 <= g30514;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5897 <= 0;
  else
    g5897 <= g30518;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5893 <= 0;
  else
    g5893 <= g30503;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5921 <= 0;
  else
    g5921 <= g30507;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5937 <= 0;
  else
    g5937 <= g30511;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5953 <= 0;
  else
    g5953 <= g30515;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5905 <= 0;
  else
    g5905 <= g30519;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5901 <= 0;
  else
    g5901 <= g30504;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5925 <= 0;
  else
    g5925 <= g30508;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5941 <= 0;
  else
    g5941 <= g30512;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5957 <= 0;
  else
    g5957 <= g30516;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5913 <= 0;
  else
    g5913 <= g30520;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5909 <= 0;
  else
    g5909 <= g30505;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5929 <= 0;
  else
    g5929 <= g30509;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5945 <= 0;
  else
    g5945 <= g30513;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5961 <= 0;
  else
    g5961 <= g30517;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5965 <= 0;
  else
    g5965 <= g30521;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4831 <= 0;
  else
    g4831 <= g28099;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5849 <= 0;
  else
    g5849 <= g29297;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5813 <= 0;
  else
    g5813 <= g25736;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5808 <= 0;
  else
    g5808 <= g29292;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5817 <= 0;
  else
    g5817 <= g29293;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5821 <= 0;
  else
    g5821 <= g25733;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5827 <= 0;
  else
    g5827 <= g29294;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5831 <= 0;
  else
    g5831 <= g29295;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5835 <= 0;
  else
    g5835 <= g29296;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5841 <= 0;
  else
    g5841 <= g25734;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5845 <= 0;
  else
    g5845 <= g25735;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5853 <= 0;
  else
    g5853 <= g34645;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6351 <= 0;
  else
    g6351 <= g24348;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6329 <= 0;
  else
    g6329 <= gbuf48;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6358 <= 0;
  else
    g6358 <= gbuf49;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6315 <= 0;
  else
    g6315 <= gbuf50;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6322 <= 0;
  else
    g6322 <= gbuf51;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6346 <= 0;
  else
    g6346 <= gbuf52;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6365 <= 0;
  else
    g6365 <= gbuf53;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6369 <= 0;
  else
    g6369 <= gbuf54;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6373 <= 0;
  else
    g6373 <= gbuf55;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6377 <= 0;
  else
    g6377 <= gbuf56;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6381 <= 0;
  else
    g6381 <= g24349;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6386 <= 0;
  else
    g6386 <= g24350;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6390 <= 0;
  else
    g6390 <= g24351;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6395 <= 0;
  else
    g6395 <= g33624;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6336 <= 0;
  else
    g6336 <= g33625;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6140 <= 0;
  else
    g6140 <= g25742;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6148 <= 0;
  else
    g6148 <= gbuf57;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6098 <= 0;
  else
    g6098 <= g25744;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6144 <= 0;
  else
    g6144 <= g25743;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6151 <= 0;
  else
    g6151 <= gbuf58;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6058 <= 0;
  else
    g6058 <= g25745;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6052 <= 0;
  else
    g6052 <= g31919;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6065 <= 0;
  else
    g6065 <= g31923;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6069 <= 0;
  else
    g6069 <= g31925;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6073 <= 0;
  else
    g6073 <= g31920;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6077 <= 0;
  else
    g6077 <= g31921;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6082 <= 0;
  else
    g6082 <= g31922;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6088 <= 0;
  else
    g6088 <= g31924;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6093 <= 0;
  else
    g6093 <= g33061;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6105 <= 0;
  else
    g6105 <= g28101;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6109 <= 0;
  else
    g6109 <= g28100;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6113 <= 0;
  else
    g6113 <= g25746;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6116 <= 0;
  else
    g6116 <= g25737;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6120 <= 0;
  else
    g6120 <= g25738;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6128 <= 0;
  else
    g6128 <= g25739;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6133 <= 0;
  else
    g6133 <= g25740;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6137 <= 0;
  else
    g6137 <= g25741;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6203 <= 0;
  else
    g6203 <= g30522;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6209 <= 0;
  else
    g6209 <= g33062;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6215 <= 0;
  else
    g6215 <= g33063;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6219 <= 0;
  else
    g6219 <= g33064;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6227 <= 0;
  else
    g6227 <= g33065;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6235 <= 0;
  else
    g6235 <= g30523;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6263 <= 0;
  else
    g6263 <= g30527;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6279 <= 0;
  else
    g6279 <= g30531;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6295 <= 0;
  else
    g6295 <= g30535;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6243 <= 0;
  else
    g6243 <= g30539;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6239 <= 0;
  else
    g6239 <= g30524;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6267 <= 0;
  else
    g6267 <= g30528;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6283 <= 0;
  else
    g6283 <= g30532;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6299 <= 0;
  else
    g6299 <= g30536;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6251 <= 0;
  else
    g6251 <= g30540;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6247 <= 0;
  else
    g6247 <= g30525;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6271 <= 0;
  else
    g6271 <= g30529;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6287 <= 0;
  else
    g6287 <= g30533;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6303 <= 0;
  else
    g6303 <= g30537;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6259 <= 0;
  else
    g6259 <= g30541;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6255 <= 0;
  else
    g6255 <= g30526;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6275 <= 0;
  else
    g6275 <= g30530;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6291 <= 0;
  else
    g6291 <= g30534;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6307 <= 0;
  else
    g6307 <= g30538;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6311 <= 0;
  else
    g6311 <= g30542;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4826 <= 0;
  else
    g4826 <= g28102;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6195 <= 0;
  else
    g6195 <= g29303;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6159 <= 0;
  else
    g6159 <= g25750;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6154 <= 0;
  else
    g6154 <= g29298;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6163 <= 0;
  else
    g6163 <= g29299;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6167 <= 0;
  else
    g6167 <= g25747;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6173 <= 0;
  else
    g6173 <= g29300;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6177 <= 0;
  else
    g6177 <= g29301;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6181 <= 0;
  else
    g6181 <= g29302;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6187 <= 0;
  else
    g6187 <= g25748;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6191 <= 0;
  else
    g6191 <= g25749;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6199 <= 0;
  else
    g6199 <= g34646;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6697 <= 0;
  else
    g6697 <= g24352;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6675 <= 0;
  else
    g6675 <= gbuf59;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6704 <= 0;
  else
    g6704 <= gbuf60;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6661 <= 0;
  else
    g6661 <= gbuf61;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6668 <= 0;
  else
    g6668 <= gbuf62;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6692 <= 0;
  else
    g6692 <= gbuf63;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6711 <= 0;
  else
    g6711 <= gbuf64;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6715 <= 0;
  else
    g6715 <= gbuf65;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6719 <= 0;
  else
    g6719 <= gbuf66;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6723 <= 0;
  else
    g6723 <= gbuf67;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6727 <= 0;
  else
    g6727 <= g24353;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6732 <= 0;
  else
    g6732 <= g24354;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6736 <= 0;
  else
    g6736 <= g24355;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6741 <= 0;
  else
    g6741 <= g33626;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6682 <= 0;
  else
    g6682 <= g33627;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6486 <= 0;
  else
    g6486 <= g25756;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6494 <= 0;
  else
    g6494 <= gbuf68;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6444 <= 0;
  else
    g6444 <= g25758;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6490 <= 0;
  else
    g6490 <= g25757;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6497 <= 0;
  else
    g6497 <= gbuf69;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6404 <= 0;
  else
    g6404 <= g25759;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6398 <= 0;
  else
    g6398 <= g31926;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6411 <= 0;
  else
    g6411 <= g31930;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6415 <= 0;
  else
    g6415 <= g31932;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6419 <= 0;
  else
    g6419 <= g31927;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6423 <= 0;
  else
    g6423 <= g31928;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6428 <= 0;
  else
    g6428 <= g31929;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6434 <= 0;
  else
    g6434 <= g31931;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6439 <= 0;
  else
    g6439 <= g33066;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6451 <= 0;
  else
    g6451 <= g28104;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6455 <= 0;
  else
    g6455 <= g28103;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6459 <= 0;
  else
    g6459 <= g25760;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6462 <= 0;
  else
    g6462 <= g25751;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6466 <= 0;
  else
    g6466 <= g25752;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6474 <= 0;
  else
    g6474 <= g25753;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6479 <= 0;
  else
    g6479 <= g25754;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6483 <= 0;
  else
    g6483 <= g25755;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6549 <= 0;
  else
    g6549 <= g30543;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6555 <= 0;
  else
    g6555 <= g33067;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6561 <= 0;
  else
    g6561 <= g33068;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6565 <= 0;
  else
    g6565 <= g33069;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6573 <= 0;
  else
    g6573 <= g33070;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6581 <= 0;
  else
    g6581 <= g30544;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6609 <= 0;
  else
    g6609 <= g30548;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6625 <= 0;
  else
    g6625 <= g30552;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6641 <= 0;
  else
    g6641 <= g30556;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6589 <= 0;
  else
    g6589 <= g30560;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6585 <= 0;
  else
    g6585 <= g30545;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6613 <= 0;
  else
    g6613 <= g30549;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6629 <= 0;
  else
    g6629 <= g30553;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6645 <= 0;
  else
    g6645 <= g30557;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6597 <= 0;
  else
    g6597 <= g30561;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6593 <= 0;
  else
    g6593 <= g30546;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6617 <= 0;
  else
    g6617 <= g30550;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6633 <= 0;
  else
    g6633 <= g30554;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6649 <= 0;
  else
    g6649 <= g30558;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6605 <= 0;
  else
    g6605 <= g30562;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6601 <= 0;
  else
    g6601 <= g30547;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6621 <= 0;
  else
    g6621 <= g30551;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6637 <= 0;
  else
    g6637 <= g30555;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6653 <= 0;
  else
    g6653 <= g30559;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6657 <= 0;
  else
    g6657 <= g30563;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5011 <= 0;
  else
    g5011 <= g28105;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6541 <= 0;
  else
    g6541 <= g29309;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6505 <= 0;
  else
    g6505 <= g25764;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6500 <= 0;
  else
    g6500 <= g29304;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6509 <= 0;
  else
    g6509 <= g29305;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6513 <= 0;
  else
    g6513 <= g25761;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6519 <= 0;
  else
    g6519 <= g29306;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6523 <= 0;
  else
    g6523 <= g29307;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6527 <= 0;
  else
    g6527 <= g29308;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6533 <= 0;
  else
    g6533 <= g25762;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6537 <= 0;
  else
    g6537 <= g25763;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6545 <= 0;
  else
    g6545 <= g34647;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3303 <= 0;
  else
    g3303 <= g24267;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3281 <= 0;
  else
    g3281 <= gbuf70;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3310 <= 0;
  else
    g3310 <= gbuf71;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3267 <= 0;
  else
    g3267 <= gbuf72;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3274 <= 0;
  else
    g3274 <= gbuf73;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3298 <= 0;
  else
    g3298 <= gbuf74;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3317 <= 0;
  else
    g3317 <= gbuf75;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3321 <= 0;
  else
    g3321 <= gbuf76;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3325 <= 0;
  else
    g3325 <= gbuf77;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3329 <= 0;
  else
    g3329 <= gbuf78;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3338 <= 0;
  else
    g3338 <= g24268;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3343 <= 0;
  else
    g3343 <= g24269;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3347 <= 0;
  else
    g3347 <= g24270;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3352 <= 0;
  else
    g3352 <= g33609;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3288 <= 0;
  else
    g3288 <= g33610;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3092 <= 0;
  else
    g3092 <= g25648;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3100 <= 0;
  else
    g3100 <= gbuf79;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3050 <= 0;
  else
    g3050 <= g25650;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3096 <= 0;
  else
    g3096 <= g25649;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3103 <= 0;
  else
    g3103 <= gbuf80;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3010 <= 0;
  else
    g3010 <= g25651;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3004 <= 0;
  else
    g3004 <= g31873;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3017 <= 0;
  else
    g3017 <= g31877;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3021 <= 0;
  else
    g3021 <= g31879;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3025 <= 0;
  else
    g3025 <= g31874;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3029 <= 0;
  else
    g3029 <= g31875;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3034 <= 0;
  else
    g3034 <= g31876;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3040 <= 0;
  else
    g3040 <= g31878;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3045 <= 0;
  else
    g3045 <= g33020;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3057 <= 0;
  else
    g3057 <= g28062;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3061 <= 0;
  else
    g3061 <= g28061;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3065 <= 0;
  else
    g3065 <= g25652;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3068 <= 0;
  else
    g3068 <= g25643;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3072 <= 0;
  else
    g3072 <= g25644;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3080 <= 0;
  else
    g3080 <= g25645;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3085 <= 0;
  else
    g3085 <= g25646;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3089 <= 0;
  else
    g3089 <= g25647;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3155 <= 0;
  else
    g3155 <= g30393;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3161 <= 0;
  else
    g3161 <= g33021;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3167 <= 0;
  else
    g3167 <= g33022;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3171 <= 0;
  else
    g3171 <= g33023;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3179 <= 0;
  else
    g3179 <= g33024;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3187 <= 0;
  else
    g3187 <= g30394;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3215 <= 0;
  else
    g3215 <= g30398;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3231 <= 0;
  else
    g3231 <= g30402;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3247 <= 0;
  else
    g3247 <= g30406;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3195 <= 0;
  else
    g3195 <= g30410;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3191 <= 0;
  else
    g3191 <= g30395;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3219 <= 0;
  else
    g3219 <= g30399;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3235 <= 0;
  else
    g3235 <= g30403;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3251 <= 0;
  else
    g3251 <= g30407;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3203 <= 0;
  else
    g3203 <= g30411;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3199 <= 0;
  else
    g3199 <= g30396;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3223 <= 0;
  else
    g3223 <= g30400;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3239 <= 0;
  else
    g3239 <= g30404;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3255 <= 0;
  else
    g3255 <= g30408;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3211 <= 0;
  else
    g3211 <= g30412;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3207 <= 0;
  else
    g3207 <= g30397;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3227 <= 0;
  else
    g3227 <= g30401;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3243 <= 0;
  else
    g3243 <= g30405;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3259 <= 0;
  else
    g3259 <= g30409;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3263 <= 0;
  else
    g3263 <= g30413;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3333 <= 0;
  else
    g3333 <= g28063;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3147 <= 0;
  else
    g3147 <= g29262;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3111 <= 0;
  else
    g3111 <= g25656;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3106 <= 0;
  else
    g3106 <= g29257;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3115 <= 0;
  else
    g3115 <= g29258;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3119 <= 0;
  else
    g3119 <= g25653;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3125 <= 0;
  else
    g3125 <= g29259;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3129 <= 0;
  else
    g3129 <= g29260;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3133 <= 0;
  else
    g3133 <= g29261;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3139 <= 0;
  else
    g3139 <= g25654;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3143 <= 0;
  else
    g3143 <= g25655;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3151 <= 0;
  else
    g3151 <= g34625;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3654 <= 0;
  else
    g3654 <= g24271;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3632 <= 0;
  else
    g3632 <= gbuf81;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3661 <= 0;
  else
    g3661 <= gbuf82;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3618 <= 0;
  else
    g3618 <= gbuf83;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3625 <= 0;
  else
    g3625 <= gbuf84;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3649 <= 0;
  else
    g3649 <= gbuf85;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3668 <= 0;
  else
    g3668 <= gbuf86;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3672 <= 0;
  else
    g3672 <= gbuf87;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3676 <= 0;
  else
    g3676 <= gbuf88;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3680 <= 0;
  else
    g3680 <= gbuf89;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3689 <= 0;
  else
    g3689 <= g24272;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3694 <= 0;
  else
    g3694 <= g24273;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3698 <= 0;
  else
    g3698 <= g24274;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3703 <= 0;
  else
    g3703 <= g33611;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3639 <= 0;
  else
    g3639 <= g33612;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3443 <= 0;
  else
    g3443 <= g25662;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3451 <= 0;
  else
    g3451 <= gbuf90;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3401 <= 0;
  else
    g3401 <= g25664;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3447 <= 0;
  else
    g3447 <= g25663;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3454 <= 0;
  else
    g3454 <= gbuf91;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3361 <= 0;
  else
    g3361 <= g25665;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3355 <= 0;
  else
    g3355 <= g31880;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3368 <= 0;
  else
    g3368 <= g31884;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3372 <= 0;
  else
    g3372 <= g31886;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3376 <= 0;
  else
    g3376 <= g31881;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3380 <= 0;
  else
    g3380 <= g31882;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3385 <= 0;
  else
    g3385 <= g31883;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3391 <= 0;
  else
    g3391 <= g31885;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3396 <= 0;
  else
    g3396 <= g33025;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3408 <= 0;
  else
    g3408 <= g28065;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3412 <= 0;
  else
    g3412 <= g28064;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3416 <= 0;
  else
    g3416 <= g25666;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3419 <= 0;
  else
    g3419 <= g25657;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3423 <= 0;
  else
    g3423 <= g25658;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3431 <= 0;
  else
    g3431 <= g25659;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3436 <= 0;
  else
    g3436 <= g25660;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3440 <= 0;
  else
    g3440 <= g25661;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3506 <= 0;
  else
    g3506 <= g30414;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3512 <= 0;
  else
    g3512 <= g33026;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3518 <= 0;
  else
    g3518 <= g33027;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3522 <= 0;
  else
    g3522 <= g33028;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3530 <= 0;
  else
    g3530 <= g33029;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3538 <= 0;
  else
    g3538 <= g30415;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3566 <= 0;
  else
    g3566 <= g30419;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3582 <= 0;
  else
    g3582 <= g30423;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3598 <= 0;
  else
    g3598 <= g30427;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3546 <= 0;
  else
    g3546 <= g30431;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3542 <= 0;
  else
    g3542 <= g30416;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3570 <= 0;
  else
    g3570 <= g30420;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3586 <= 0;
  else
    g3586 <= g30424;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3602 <= 0;
  else
    g3602 <= g30428;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3554 <= 0;
  else
    g3554 <= g30432;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3550 <= 0;
  else
    g3550 <= g30417;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3574 <= 0;
  else
    g3574 <= g30421;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3590 <= 0;
  else
    g3590 <= g30425;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3606 <= 0;
  else
    g3606 <= g30429;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3562 <= 0;
  else
    g3562 <= g30433;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3558 <= 0;
  else
    g3558 <= g30418;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3578 <= 0;
  else
    g3578 <= g30422;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3594 <= 0;
  else
    g3594 <= g30426;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3610 <= 0;
  else
    g3610 <= g30430;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3614 <= 0;
  else
    g3614 <= g30434;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3684 <= 0;
  else
    g3684 <= g28066;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3498 <= 0;
  else
    g3498 <= g29268;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3462 <= 0;
  else
    g3462 <= g25670;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3457 <= 0;
  else
    g3457 <= g29263;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3466 <= 0;
  else
    g3466 <= g29264;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3470 <= 0;
  else
    g3470 <= g25667;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3476 <= 0;
  else
    g3476 <= g29265;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3480 <= 0;
  else
    g3480 <= g29266;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3484 <= 0;
  else
    g3484 <= g29267;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3490 <= 0;
  else
    g3490 <= g25668;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3494 <= 0;
  else
    g3494 <= g25669;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3502 <= 0;
  else
    g3502 <= g34626;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4005 <= 0;
  else
    g4005 <= g24275;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3983 <= 0;
  else
    g3983 <= gbuf92;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4012 <= 0;
  else
    g4012 <= gbuf93;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3969 <= 0;
  else
    g3969 <= gbuf94;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3976 <= 0;
  else
    g3976 <= gbuf95;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4000 <= 0;
  else
    g4000 <= gbuf96;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4019 <= 0;
  else
    g4019 <= gbuf97;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4023 <= 0;
  else
    g4023 <= gbuf98;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4027 <= 0;
  else
    g4027 <= gbuf99;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4031 <= 0;
  else
    g4031 <= gbuf100;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4040 <= 0;
  else
    g4040 <= g24276;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4045 <= 0;
  else
    g4045 <= g24277;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4049 <= 0;
  else
    g4049 <= g24278;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4054 <= 0;
  else
    g4054 <= g33613;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3990 <= 0;
  else
    g3990 <= g33614;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3794 <= 0;
  else
    g3794 <= g25676;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3802 <= 0;
  else
    g3802 <= gbuf101;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3752 <= 0;
  else
    g3752 <= g25678;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3798 <= 0;
  else
    g3798 <= g25677;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3805 <= 0;
  else
    g3805 <= gbuf102;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3712 <= 0;
  else
    g3712 <= g25679;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3706 <= 0;
  else
    g3706 <= g31887;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3719 <= 0;
  else
    g3719 <= g31891;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3723 <= 0;
  else
    g3723 <= g31893;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3727 <= 0;
  else
    g3727 <= g31888;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3731 <= 0;
  else
    g3731 <= g31889;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3736 <= 0;
  else
    g3736 <= g31890;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3742 <= 0;
  else
    g3742 <= g31892;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3747 <= 0;
  else
    g3747 <= g33030;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3759 <= 0;
  else
    g3759 <= g28068;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3763 <= 0;
  else
    g3763 <= g28067;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3767 <= 0;
  else
    g3767 <= g25680;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3770 <= 0;
  else
    g3770 <= g25671;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3774 <= 0;
  else
    g3774 <= g25672;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3782 <= 0;
  else
    g3782 <= g25673;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3787 <= 0;
  else
    g3787 <= g25674;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3791 <= 0;
  else
    g3791 <= g25675;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3857 <= 0;
  else
    g3857 <= g30435;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3863 <= 0;
  else
    g3863 <= g33031;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3869 <= 0;
  else
    g3869 <= g33032;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3873 <= 0;
  else
    g3873 <= g33033;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3881 <= 0;
  else
    g3881 <= g33034;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3889 <= 0;
  else
    g3889 <= g30436;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3917 <= 0;
  else
    g3917 <= g30440;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3933 <= 0;
  else
    g3933 <= g30444;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3949 <= 0;
  else
    g3949 <= g30448;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3897 <= 0;
  else
    g3897 <= g30452;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3893 <= 0;
  else
    g3893 <= g30437;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3921 <= 0;
  else
    g3921 <= g30441;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3937 <= 0;
  else
    g3937 <= g30445;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3953 <= 0;
  else
    g3953 <= g30449;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3905 <= 0;
  else
    g3905 <= g30453;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3901 <= 0;
  else
    g3901 <= g30438;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3925 <= 0;
  else
    g3925 <= g30442;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3941 <= 0;
  else
    g3941 <= g30446;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3957 <= 0;
  else
    g3957 <= g30450;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3913 <= 0;
  else
    g3913 <= g30454;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3909 <= 0;
  else
    g3909 <= g30439;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3929 <= 0;
  else
    g3929 <= g30443;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3945 <= 0;
  else
    g3945 <= g30447;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3961 <= 0;
  else
    g3961 <= g30451;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3965 <= 0;
  else
    g3965 <= g30455;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4035 <= 0;
  else
    g4035 <= g28069;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3849 <= 0;
  else
    g3849 <= g29274;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3813 <= 0;
  else
    g3813 <= g25684;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3808 <= 0;
  else
    g3808 <= g29269;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3817 <= 0;
  else
    g3817 <= g29270;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3821 <= 0;
  else
    g3821 <= g25681;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3827 <= 0;
  else
    g3827 <= g29271;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3831 <= 0;
  else
    g3831 <= g29272;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3835 <= 0;
  else
    g3835 <= g29273;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3841 <= 0;
  else
    g3841 <= g25682;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3845 <= 0;
  else
    g3845 <= g25683;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3853 <= 0;
  else
    g3853 <= g34627;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4165 <= 0;
  else
    g4165 <= g28079;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4169 <= 0;
  else
    g4169 <= g28080;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4125 <= 0;
  else
    g4125 <= g28081;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4072 <= 0;
  else
    g4072 <= g25691;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4064 <= 0;
  else
    g4064 <= g25685;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4057 <= 0;
  else
    g4057 <= g25686;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4141 <= 0;
  else
    g4141 <= g25687;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4082 <= 0;
  else
    g4082 <= g26938;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4076 <= 0;
  else
    g4076 <= g28070;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4087 <= 0;
  else
    g4087 <= g29275;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4093 <= 0;
  else
    g4093 <= g30456;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4098 <= 0;
  else
    g4098 <= g31894;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4108 <= 0;
  else
    g4108 <= g33035;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4104 <= 0;
  else
    g4104 <= g33615;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4145 <= 0;
  else
    g4145 <= g26939;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4112 <= 0;
  else
    g4112 <= g28071;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4116 <= 0;
  else
    g4116 <= g28072;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4119 <= 0;
  else
    g4119 <= g28073;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4122 <= 0;
  else
    g4122 <= g28074;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4153 <= 0;
  else
    g4153 <= g30457;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4164 <= 0;
  else
    g4164 <= g26940;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4129 <= 0;
  else
    g4129 <= g28075;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4132 <= 0;
  else
    g4132 <= g28076;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4135 <= 0;
  else
    g4135 <= g28077;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4138 <= 0;
  else
    g4138 <= g28078;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4172 <= 0;
  else
    g4172 <= g34733;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4176 <= 0;
  else
    g4176 <= g34734;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4146 <= 0;
  else
    g4146 <= g34628;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4157 <= 0;
  else
    g4157 <= g34629;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4258 <= 0;
  else
    g4258 <= g21893;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4264 <= 0;
  else
    g4264 <= g21894;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4269 <= 0;
  else
    g4269 <= g21895;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4273 <= 0;
  else
    g4273 <= g24280;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4239 <= 0;
  else
    g4239 <= g21892;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4294 <= 0;
  else
    g4294 <= g21900;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4297 <= 0;
  else
    g4297 <= gbuf103;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4300 <= 0;
  else
    g4300 <= g34735;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4253 <= 0;
  else
    g4253 <= g34630;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4249 <= 0;
  else
    g4249 <= g34631;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4245 <= 0;
  else
    g4245 <= g34632;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4277 <= 0;
  else
    g4277 <= g21896;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4281 <= 0;
  else
    g4281 <= gbuf104;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4284 <= 0;
  else
    g4284 <= g21897;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4287 <= 0;
  else
    g4287 <= g21898;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4291 <= 0;
  else
    g4291 <= gbuf105;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2946 <= 0;
  else
    g2946 <= g21899;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4191 <= 0;
  else
    g4191 <= g21901;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4188 <= 0;
  else
    g4188 <= gbuf106;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4194 <= 0;
  else
    g4194 <= gbuf107;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4197 <= 0;
  else
    g4197 <= gbuf108;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4200 <= 0;
  else
    g4200 <= gbuf109;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4204 <= 0;
  else
    g4204 <= gbuf110;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4207 <= 0;
  else
    g4207 <= gbuf111;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4210 <= 0;
  else
    g4210 <= gbuf112;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4180 <= 0;
  else
    g4180 <= gbuf113;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4185 <= 0;
  else
    g4185 <= g21891;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4213 <= 0;
  else
    g4213 <= gbuf114;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4216 <= 0;
  else
    g4216 <= gbuf115;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4219 <= 0;
  else
    g4219 <= gbuf116;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4222 <= 0;
  else
    g4222 <= gbuf117;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4226 <= 0;
  else
    g4226 <= gbuf118;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4229 <= 0;
  else
    g4229 <= gbuf119;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4232 <= 0;
  else
    g4232 <= gbuf120;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4235 <= 0;
  else
    g4235 <= gbuf121;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4242 <= 0;
  else
    g4242 <= g24279;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g305 <= 0;
  else
    g305 <= g26880;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g311 <= 0;
  else
    g311 <= g26881;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g336 <= 0;
  else
    g336 <= g26886;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g324 <= 0;
  else
    g324 <= g26887;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g316 <= 0;
  else
    g316 <= g26883;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g319 <= 0;
  else
    g319 <= g26882;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g329 <= 0;
  else
    g329 <= g26885;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g333 <= 0;
  else
    g333 <= g26884;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g344 <= 0;
  else
    g344 <= g26890;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g347 <= 0;
  else
    g347 <= gbuf122;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g351 <= 0;
  else
    g351 <= g26891;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g355 <= 0;
  else
    g355 <= g26892;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g74 <= 0;
  else
    g74 <= g26893;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g106 <= 0;
  else
    g106 <= g26889;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g341 <= 0;
  else
    g341 <= g26888;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g637 <= 0;
  else
    g637 <= g24212;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g640 <= 0;
  else
    g640 <= gbuf123;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g559 <= 0;
  else
    g559 <= gbuf124;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g562 <= 0;
  else
    g562 <= g25613;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g568 <= 0;
  else
    g568 <= g26895;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g572 <= 0;
  else
    g572 <= g28045;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g586 <= 0;
  else
    g586 <= g29224;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g577 <= 0;
  else
    g577 <= g30334;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g582 <= 0;
  else
    g582 <= g31866;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g590 <= 0;
  else
    g590 <= g32978;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g595 <= 0;
  else
    g595 <= g33538;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g599 <= 0;
  else
    g599 <= g33964;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g604 <= 0;
  else
    g604 <= g34251;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g608 <= 0;
  else
    g608 <= g34438;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g613 <= 0;
  else
    g613 <= g34599;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g617 <= 0;
  else
    g617 <= g34724;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g622 <= 0;
  else
    g622 <= g34790;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g626 <= 0;
  else
    g626 <= g34849;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g632 <= 0;
  else
    g632 <= g34880;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g859 <= 0;
  else
    g859 <= g26900;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g869 <= 0;
  else
    g869 <= gbuf125;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g875 <= 0;
  else
    g875 <= gbuf126;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g878 <= 0;
  else
    g878 <= gbuf127;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g881 <= 0;
  else
    g881 <= gbuf128;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g884 <= 0;
  else
    g884 <= gbuf129;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g887 <= 0;
  else
    g887 <= gbuf130;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g872 <= 0;
  else
    g872 <= gbuf131;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g225 <= 0;
  else
    g225 <= g26901;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g255 <= 0;
  else
    g255 <= g26902;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g232 <= 0;
  else
    g232 <= g26903;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g262 <= 0;
  else
    g262 <= g26904;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g239 <= 0;
  else
    g239 <= g26905;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g269 <= 0;
  else
    g269 <= g26906;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g246 <= 0;
  else
    g246 <= g26907;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g446 <= 0;
  else
    g446 <= g26908;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g890 <= 0;
  else
    g890 <= g34440;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g862 <= 0;
  else
    g862 <= g26909;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g896 <= 0;
  else
    g896 <= g26910;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g901 <= 0;
  else
    g901 <= g25620;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g391 <= 0;
  else
    g391 <= g26911;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g365 <= 0;
  else
    g365 <= g25595;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g358 <= 0;
  else
    g358 <= gbuf132;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g370 <= 0;
  else
    g370 <= g25597;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g376 <= 0;
  else
    g376 <= g25596;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g385 <= 0;
  else
    g385 <= g25598;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g203 <= 0;
  else
    g203 <= g25599;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g854 <= 0;
  else
    g854 <= g32980;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g847 <= 0;
  else
    g847 <= g24216;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g703 <= 0;
  else
    g703 <= g24214;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g837 <= 0;
  else
    g837 <= g24215;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g843 <= 0;
  else
    g843 <= g25619;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g812 <= 0;
  else
    g812 <= g26898;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g817 <= 0;
  else
    g817 <= g25617;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g832 <= 0;
  else
    g832 <= g25618;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g822 <= 0;
  else
    g822 <= g26899;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g827 <= 0;
  else
    g827 <= g28055;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g723 <= 0;
  else
    g723 <= g29229;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g645 <= 0;
  else
    g645 <= g28046;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g681 <= 0;
  else
    g681 <= g28047;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g699 <= 0;
  else
    g699 <= g28053;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g650 <= 0;
  else
    g650 <= g28049;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g655 <= 0;
  else
    g655 <= g28050;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g718 <= 0;
  else
    g718 <= g28051;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g661 <= 0;
  else
    g661 <= g28052;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g728 <= 0;
  else
    g728 <= g28054;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g79 <= 0;
  else
    g79 <= g26896;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g691 <= 0;
  else
    g691 <= g28048;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g686 <= 0;
  else
    g686 <= g25614;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g667 <= 0;
  else
    g667 <= g25615;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g671 <= 0;
  else
    g671 <= g29225;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g676 <= 0;
  else
    g676 <= g29226;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g714 <= 0;
  else
    g714 <= g29227;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g499 <= 0;
  else
    g499 <= g25609;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g504 <= 0;
  else
    g504 <= g25610;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g513 <= 0;
  else
    g513 <= g25611;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g518 <= 0;
  else
    g518 <= g25612;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g528 <= 0;
  else
    g528 <= g26894;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g482 <= 0;
  else
    g482 <= g28044;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g490 <= 0;
  else
    g490 <= g29223;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g417 <= 0;
  else
    g417 <= g24209;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g411 <= 0;
  else
    g411 <= g29222;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g424 <= 0;
  else
    g424 <= g24202;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g475 <= 0;
  else
    g475 <= g24208;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g441 <= 0;
  else
    g441 <= g24207;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g437 <= 0;
  else
    g437 <= g24206;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g433 <= 0;
  else
    g433 <= g24205;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g429 <= 0;
  else
    g429 <= g24204;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g401 <= 0;
  else
    g401 <= g24203;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g392 <= 0;
  else
    g392 <= g24200;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g405 <= 0;
  else
    g405 <= g24201;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g182 <= 0;
  else
    g182 <= g25602;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g174 <= 0;
  else
    g174 <= g25601;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g168 <= 0;
  else
    g168 <= g25600;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g460 <= 0;
  else
    g460 <= g25605;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g452 <= 0;
  else
    g452 <= g25604;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g457 <= 0;
  else
    g457 <= g25603;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g471 <= 0;
  else
    g471 <= g25608;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g464 <= 0;
  else
    g464 <= g25607;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g468 <= 0;
  else
    g468 <= g25606;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g479 <= 0;
  else
    g479 <= g24210;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g102 <= 0;
  else
    g102 <= g33962;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g496 <= 0;
  else
    g496 <= g33963;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g732 <= 0;
  else
    g732 <= g25616;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g753 <= 0;
  else
    g753 <= g26897;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g799 <= 0;
  else
    g799 <= g24213;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g802 <= 0;
  else
    g802 <= gbuf133;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g736 <= 0;
  else
    g736 <= gbuf134;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g739 <= 0;
  else
    g739 <= g29228;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g744 <= 0;
  else
    g744 <= g30335;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g749 <= 0;
  else
    g749 <= g31867;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g758 <= 0;
  else
    g758 <= g32979;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g763 <= 0;
  else
    g763 <= g33539;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g767 <= 0;
  else
    g767 <= g33965;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g772 <= 0;
  else
    g772 <= g34252;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g776 <= 0;
  else
    g776 <= g34439;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g781 <= 0;
  else
    g781 <= g34600;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g785 <= 0;
  else
    g785 <= g34725;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g790 <= 0;
  else
    g790 <= g34791;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g794 <= 0;
  else
    g794 <= g34850;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g807 <= 0;
  else
    g807 <= g34881;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g554 <= 0;
  else
    g554 <= g34911;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g538 <= 0;
  else
    g538 <= g34719;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g546 <= 0;
  else
    g546 <= g34722;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g542 <= 0;
  else
    g542 <= g24211;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g534 <= 0;
  else
    g534 <= g34723;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g550 <= 0;
  else
    g550 <= g34720;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g136 <= 0;
  else
    g136 <= g34598;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g199 <= 0;
  else
    g199 <= g34721;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g278 <= 0;
  else
    g278 <= g25594;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g283 <= 0;
  else
    g283 <= g28043;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g287 <= 0;
  else
    g287 <= g31865;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g291 <= 0;
  else
    g291 <= g32977;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g294 <= 0;
  else
    g294 <= g33535;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g298 <= 0;
  else
    g298 <= g33961;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g142 <= 0;
  else
    g142 <= g34250;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g146 <= 0;
  else
    g146 <= g30333;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g164 <= 0;
  else
    g164 <= g31864;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g150 <= 0;
  else
    g150 <= g32976;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g153 <= 0;
  else
    g153 <= g33534;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g157 <= 0;
  else
    g157 <= g33960;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g160 <= 0;
  else
    g160 <= g34249;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g301 <= 0;
  else
    g301 <= g33536;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g222 <= 0;
  else
    g222 <= g33537;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g194 <= 0;
  else
    g194 <= g25592;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g191 <= 0;
  else
    g191 <= gbuf135;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g209 <= 0;
  else
    g209 <= g25593;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g215 <= 0;
  else
    g215 <= g25591;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g218 <= 0;
  else
    g218 <= gbuf136;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1249 <= 0;
  else
    g1249 <= g24247;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1266 <= 0;
  else
    g1266 <= g25630;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1280 <= 0;
  else
    g1280 <= g26919;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1252 <= 0;
  else
    g1252 <= g28058;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1256 <= 0;
  else
    g1256 <= g29235;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1259 <= 0;
  else
    g1259 <= g30342;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1263 <= 0;
  else
    g1263 <= g31870;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1270 <= 0;
  else
    g1270 <= g32984;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1274 <= 0;
  else
    g1274 <= g33542;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1277 <= 0;
  else
    g1277 <= g32985;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1418 <= 0;
  else
    g1418 <= g24254;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1422 <= 0;
  else
    g1422 <= gbuf137;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1426 <= 0;
  else
    g1426 <= gbuf138;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1430 <= 0;
  else
    g1430 <= gbuf139;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1548 <= 0;
  else
    g1548 <= g24260;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1564 <= 0;
  else
    g1564 <= g24262;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1559 <= 0;
  else
    g1559 <= g25638;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1554 <= 0;
  else
    g1554 <= g25637;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1570 <= 0;
  else
    g1570 <= g24258;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1585 <= 0;
  else
    g1585 <= gbuf140;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1589 <= 0;
  else
    g1589 <= g24261;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1576 <= 0;
  else
    g1576 <= g24255;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1579 <= 0;
  else
    g1579 <= gbuf141;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1339 <= 0;
  else
    g1339 <= g24259;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1500 <= 0;
  else
    g1500 <= g24256;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1582 <= 0;
  else
    g1582 <= gbuf142;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1333 <= 0;
  else
    g1333 <= gbuf143;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1399 <= 0;
  else
    g1399 <= g24257;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1459 <= 0;
  else
    g1459 <= gbuf144;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1322 <= 0;
  else
    g1322 <= gbuf145;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1514 <= 0;
  else
    g1514 <= g30344;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1526 <= 0;
  else
    g1526 <= g30345;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1521 <= 0;
  else
    g1521 <= g24252;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1306 <= 0;
  else
    g1306 <= g25636;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1532 <= 0;
  else
    g1532 <= g24253;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1536 <= 0;
  else
    g1536 <= g26925;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1542 <= 0;
  else
    g1542 <= g30346;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1413 <= 0;
  else
    g1413 <= g30347;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1395 <= 0;
  else
    g1395 <= g25634;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1404 <= 0;
  else
    g1404 <= g26921;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1319 <= 0;
  else
    g1319 <= g24248;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1312 <= 0;
  else
    g1312 <= g25631;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1351 <= 0;
  else
    g1351 <= g25632;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1345 <= 0;
  else
    g1345 <= g28059;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1361 <= 0;
  else
    g1361 <= g30343;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1367 <= 0;
  else
    g1367 <= g31871;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1373 <= 0;
  else
    g1373 <= g32986;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1379 <= 0;
  else
    g1379 <= g33543;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1384 <= 0;
  else
    g1384 <= g25633;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1389 <= 0;
  else
    g1389 <= g26920;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1489 <= 0;
  else
    g1489 <= g24249;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1495 <= 0;
  else
    g1495 <= g24250;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1442 <= 0;
  else
    g1442 <= g24251;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1437 <= 0;
  else
    g1437 <= g29236;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1478 <= 0;
  else
    g1478 <= g26924;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1454 <= 0;
  else
    g1454 <= g29239;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1448 <= 0;
  else
    g1448 <= g26922;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1467 <= 0;
  else
    g1467 <= g29237;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1472 <= 0;
  else
    g1472 <= g26923;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1484 <= 0;
  else
    g1484 <= g29238;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1300 <= 0;
  else
    g1300 <= g25635;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1291 <= 0;
  else
    g1291 <= g34602;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1296 <= 0;
  else
    g1296 <= g34729;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1283 <= 0;
  else
    g1283 <= g34730;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1287 <= 0;
  else
    g1287 <= g34731;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1311 <= 0;
  else
    g1311 <= g21724;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g929 <= 0;
  else
    g929 <= g21725;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g904 <= 0;
  else
    g904 <= g24231;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g921 <= 0;
  else
    g921 <= g25621;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g936 <= 0;
  else
    g936 <= g26912;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g907 <= 0;
  else
    g907 <= g28056;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g911 <= 0;
  else
    g911 <= g29230;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g914 <= 0;
  else
    g914 <= g30336;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g918 <= 0;
  else
    g918 <= g31868;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g925 <= 0;
  else
    g925 <= g32981;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g930 <= 0;
  else
    g930 <= g33540;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g933 <= 0;
  else
    g933 <= g32982;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1075 <= 0;
  else
    g1075 <= g24238;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1079 <= 0;
  else
    g1079 <= gbuf146;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1083 <= 0;
  else
    g1083 <= gbuf147;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1087 <= 0;
  else
    g1087 <= gbuf148;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1205 <= 0;
  else
    g1205 <= g24244;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1221 <= 0;
  else
    g1221 <= g24246;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1216 <= 0;
  else
    g1216 <= g25629;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1211 <= 0;
  else
    g1211 <= g25628;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1227 <= 0;
  else
    g1227 <= g24242;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1242 <= 0;
  else
    g1242 <= gbuf149;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1246 <= 0;
  else
    g1246 <= g24245;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1233 <= 0;
  else
    g1233 <= g24239;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1236 <= 0;
  else
    g1236 <= gbuf150;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g996 <= 0;
  else
    g996 <= g24243;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1157 <= 0;
  else
    g1157 <= g24240;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1239 <= 0;
  else
    g1239 <= gbuf151;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g990 <= 0;
  else
    g990 <= gbuf152;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1056 <= 0;
  else
    g1056 <= g24241;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1116 <= 0;
  else
    g1116 <= gbuf153;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g979 <= 0;
  else
    g979 <= gbuf154;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1171 <= 0;
  else
    g1171 <= g30338;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1183 <= 0;
  else
    g1183 <= g30339;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1178 <= 0;
  else
    g1178 <= g24236;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g962 <= 0;
  else
    g962 <= g25627;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1189 <= 0;
  else
    g1189 <= g24237;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1193 <= 0;
  else
    g1193 <= g26918;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1199 <= 0;
  else
    g1199 <= g30340;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1070 <= 0;
  else
    g1070 <= g30341;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1052 <= 0;
  else
    g1052 <= g25625;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1061 <= 0;
  else
    g1061 <= g26914;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g976 <= 0;
  else
    g976 <= g24232;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g969 <= 0;
  else
    g969 <= g25622;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1008 <= 0;
  else
    g1008 <= g25623;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1002 <= 0;
  else
    g1002 <= g28057;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1018 <= 0;
  else
    g1018 <= g30337;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1024 <= 0;
  else
    g1024 <= g31869;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1030 <= 0;
  else
    g1030 <= g32983;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1036 <= 0;
  else
    g1036 <= g33541;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1041 <= 0;
  else
    g1041 <= g25624;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1046 <= 0;
  else
    g1046 <= g26913;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1146 <= 0;
  else
    g1146 <= g24233;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1152 <= 0;
  else
    g1152 <= g24234;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1099 <= 0;
  else
    g1099 <= g24235;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1094 <= 0;
  else
    g1094 <= g29231;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1135 <= 0;
  else
    g1135 <= g26917;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1111 <= 0;
  else
    g1111 <= g29234;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1105 <= 0;
  else
    g1105 <= g26915;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1124 <= 0;
  else
    g1124 <= g29232;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1129 <= 0;
  else
    g1129 <= g26916;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1141 <= 0;
  else
    g1141 <= g29233;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g956 <= 0;
  else
    g956 <= g25626;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g947 <= 0;
  else
    g947 <= g34601;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g952 <= 0;
  else
    g952 <= g34726;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g939 <= 0;
  else
    g939 <= g34727;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g943 <= 0;
  else
    g943 <= g34728;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g967 <= 0;
  else
    g967 <= g21722;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g968 <= 0;
  else
    g968 <= g21723;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1592 <= 0;
  else
    g1592 <= g33544;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1644 <= 0;
  else
    g1644 <= g33551;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1636 <= 0;
  else
    g1636 <= g33545;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1668 <= 0;
  else
    g1668 <= g33546;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1682 <= 0;
  else
    g1682 <= g33971;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1687 <= 0;
  else
    g1687 <= g33547;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1604 <= 0;
  else
    g1604 <= g33972;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1600 <= 0;
  else
    g1600 <= g33966;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1608 <= 0;
  else
    g1608 <= g33967;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1620 <= 0;
  else
    g1620 <= g33970;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1616 <= 0;
  else
    g1616 <= g33969;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1612 <= 0;
  else
    g1612 <= g33968;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1632 <= 0;
  else
    g1632 <= g30348;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1624 <= 0;
  else
    g1624 <= g32987;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1648 <= 0;
  else
    g1648 <= g32988;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1664 <= 0;
  else
    g1664 <= g32990;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1657 <= 0;
  else
    g1657 <= g32989;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1677 <= 0;
  else
    g1677 <= g29240;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1691 <= 0;
  else
    g1691 <= g29241;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1696 <= 0;
  else
    g1696 <= g30349;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1700 <= 0;
  else
    g1700 <= g30350;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1706 <= 0;
  else
    g1706 <= g33548;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1710 <= 0;
  else
    g1710 <= g33549;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1714 <= 0;
  else
    g1714 <= g33550;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1720 <= 0;
  else
    g1720 <= g30351;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1724 <= 0;
  else
    g1724 <= g30352;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1728 <= 0;
  else
    g1728 <= g33552;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1779 <= 0;
  else
    g1779 <= g33559;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1772 <= 0;
  else
    g1772 <= g33553;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1802 <= 0;
  else
    g1802 <= g33554;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1816 <= 0;
  else
    g1816 <= g33978;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1821 <= 0;
  else
    g1821 <= g33555;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1740 <= 0;
  else
    g1740 <= g33979;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1736 <= 0;
  else
    g1736 <= g33973;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1744 <= 0;
  else
    g1744 <= g33974;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1756 <= 0;
  else
    g1756 <= g33977;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1752 <= 0;
  else
    g1752 <= g33976;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1748 <= 0;
  else
    g1748 <= g33975;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1768 <= 0;
  else
    g1768 <= g30353;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1760 <= 0;
  else
    g1760 <= g32991;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1783 <= 0;
  else
    g1783 <= g32992;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1798 <= 0;
  else
    g1798 <= g32994;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1792 <= 0;
  else
    g1792 <= g32993;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1811 <= 0;
  else
    g1811 <= g29242;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1825 <= 0;
  else
    g1825 <= g29243;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1830 <= 0;
  else
    g1830 <= g30354;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1834 <= 0;
  else
    g1834 <= g30355;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1840 <= 0;
  else
    g1840 <= g33556;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1844 <= 0;
  else
    g1844 <= g33557;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1848 <= 0;
  else
    g1848 <= g33558;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1854 <= 0;
  else
    g1854 <= g30356;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1858 <= 0;
  else
    g1858 <= g30357;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1862 <= 0;
  else
    g1862 <= g33560;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1913 <= 0;
  else
    g1913 <= g33567;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1906 <= 0;
  else
    g1906 <= g33561;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1936 <= 0;
  else
    g1936 <= g33562;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1950 <= 0;
  else
    g1950 <= g33985;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1955 <= 0;
  else
    g1955 <= g33563;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1874 <= 0;
  else
    g1874 <= g33986;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1870 <= 0;
  else
    g1870 <= g33980;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1878 <= 0;
  else
    g1878 <= g33981;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1890 <= 0;
  else
    g1890 <= g33984;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1886 <= 0;
  else
    g1886 <= g33983;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1882 <= 0;
  else
    g1882 <= g33982;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1902 <= 0;
  else
    g1902 <= g30358;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1894 <= 0;
  else
    g1894 <= g32995;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1917 <= 0;
  else
    g1917 <= g32996;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1932 <= 0;
  else
    g1932 <= g32998;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1926 <= 0;
  else
    g1926 <= g32997;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1945 <= 0;
  else
    g1945 <= g29244;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1959 <= 0;
  else
    g1959 <= g29245;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1964 <= 0;
  else
    g1964 <= g30359;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1968 <= 0;
  else
    g1968 <= g30360;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1974 <= 0;
  else
    g1974 <= g33564;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1978 <= 0;
  else
    g1978 <= g33565;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1982 <= 0;
  else
    g1982 <= g33566;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1988 <= 0;
  else
    g1988 <= g30361;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1992 <= 0;
  else
    g1992 <= g30362;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1996 <= 0;
  else
    g1996 <= g33568;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2047 <= 0;
  else
    g2047 <= g33575;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2040 <= 0;
  else
    g2040 <= g33569;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2070 <= 0;
  else
    g2070 <= g33570;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2084 <= 0;
  else
    g2084 <= g33992;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2089 <= 0;
  else
    g2089 <= g33571;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2008 <= 0;
  else
    g2008 <= g33993;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2004 <= 0;
  else
    g2004 <= g33987;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2012 <= 0;
  else
    g2012 <= g33988;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2024 <= 0;
  else
    g2024 <= g33991;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2020 <= 0;
  else
    g2020 <= g33990;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2016 <= 0;
  else
    g2016 <= g33989;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2036 <= 0;
  else
    g2036 <= g30363;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2028 <= 0;
  else
    g2028 <= g32999;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2051 <= 0;
  else
    g2051 <= g33000;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2066 <= 0;
  else
    g2066 <= g33002;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2060 <= 0;
  else
    g2060 <= g33001;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2079 <= 0;
  else
    g2079 <= g29246;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2093 <= 0;
  else
    g2093 <= g29247;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2098 <= 0;
  else
    g2098 <= g30364;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2102 <= 0;
  else
    g2102 <= g30365;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2108 <= 0;
  else
    g2108 <= g33572;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2112 <= 0;
  else
    g2112 <= g33573;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2116 <= 0;
  else
    g2116 <= g33574;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2122 <= 0;
  else
    g2122 <= g30366;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2126 <= 0;
  else
    g2126 <= g30367;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2130 <= 0;
  else
    g2130 <= g34603;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2138 <= 0;
  else
    g2138 <= g34604;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2145 <= 0;
  else
    g2145 <= g34605;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2151 <= 0;
  else
    g2151 <= g18421;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2152 <= 0;
  else
    g2152 <= g18422;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2153 <= 0;
  else
    g2153 <= g33576;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2204 <= 0;
  else
    g2204 <= g33583;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2197 <= 0;
  else
    g2197 <= g33577;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2227 <= 0;
  else
    g2227 <= g33578;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2241 <= 0;
  else
    g2241 <= g33999;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2246 <= 0;
  else
    g2246 <= g33579;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2165 <= 0;
  else
    g2165 <= g34000;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2161 <= 0;
  else
    g2161 <= g33994;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2169 <= 0;
  else
    g2169 <= g33995;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2181 <= 0;
  else
    g2181 <= g33998;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2177 <= 0;
  else
    g2177 <= g33997;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2173 <= 0;
  else
    g2173 <= g33996;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2193 <= 0;
  else
    g2193 <= g30368;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2185 <= 0;
  else
    g2185 <= g33003;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2208 <= 0;
  else
    g2208 <= g33004;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2223 <= 0;
  else
    g2223 <= g33006;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2217 <= 0;
  else
    g2217 <= g33005;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2236 <= 0;
  else
    g2236 <= g29248;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2250 <= 0;
  else
    g2250 <= g29249;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2255 <= 0;
  else
    g2255 <= g30369;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2259 <= 0;
  else
    g2259 <= g30370;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2265 <= 0;
  else
    g2265 <= g33580;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2269 <= 0;
  else
    g2269 <= g33581;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2273 <= 0;
  else
    g2273 <= g33582;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2279 <= 0;
  else
    g2279 <= g30371;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2283 <= 0;
  else
    g2283 <= g30372;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2287 <= 0;
  else
    g2287 <= g33584;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2338 <= 0;
  else
    g2338 <= g33591;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2331 <= 0;
  else
    g2331 <= g33585;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2361 <= 0;
  else
    g2361 <= g33586;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2375 <= 0;
  else
    g2375 <= g34006;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2380 <= 0;
  else
    g2380 <= g33587;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2299 <= 0;
  else
    g2299 <= g34007;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2295 <= 0;
  else
    g2295 <= g34001;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2303 <= 0;
  else
    g2303 <= g34002;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2315 <= 0;
  else
    g2315 <= g34005;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2311 <= 0;
  else
    g2311 <= g34004;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2307 <= 0;
  else
    g2307 <= g34003;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2327 <= 0;
  else
    g2327 <= g30373;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2319 <= 0;
  else
    g2319 <= g33007;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2342 <= 0;
  else
    g2342 <= g33008;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2357 <= 0;
  else
    g2357 <= g33010;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2351 <= 0;
  else
    g2351 <= g33009;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2370 <= 0;
  else
    g2370 <= g29250;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2384 <= 0;
  else
    g2384 <= g29251;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2389 <= 0;
  else
    g2389 <= g30374;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2393 <= 0;
  else
    g2393 <= g30375;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2399 <= 0;
  else
    g2399 <= g33588;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2403 <= 0;
  else
    g2403 <= g33589;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2407 <= 0;
  else
    g2407 <= g33590;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2413 <= 0;
  else
    g2413 <= g30376;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2417 <= 0;
  else
    g2417 <= g30377;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2421 <= 0;
  else
    g2421 <= g33592;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2472 <= 0;
  else
    g2472 <= g33599;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2465 <= 0;
  else
    g2465 <= g33593;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2495 <= 0;
  else
    g2495 <= g33594;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2509 <= 0;
  else
    g2509 <= g34013;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2514 <= 0;
  else
    g2514 <= g33595;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2433 <= 0;
  else
    g2433 <= g34014;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2429 <= 0;
  else
    g2429 <= g34008;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2437 <= 0;
  else
    g2437 <= g34009;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2449 <= 0;
  else
    g2449 <= g34012;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2445 <= 0;
  else
    g2445 <= g34011;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2441 <= 0;
  else
    g2441 <= g34010;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2461 <= 0;
  else
    g2461 <= g30378;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2453 <= 0;
  else
    g2453 <= g33011;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2476 <= 0;
  else
    g2476 <= g33012;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2491 <= 0;
  else
    g2491 <= g33014;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2485 <= 0;
  else
    g2485 <= g33013;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2504 <= 0;
  else
    g2504 <= g29252;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2518 <= 0;
  else
    g2518 <= g29253;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2523 <= 0;
  else
    g2523 <= g30379;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2527 <= 0;
  else
    g2527 <= g30380;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2533 <= 0;
  else
    g2533 <= g33596;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2537 <= 0;
  else
    g2537 <= g33597;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2541 <= 0;
  else
    g2541 <= g33598;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2547 <= 0;
  else
    g2547 <= g30381;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2551 <= 0;
  else
    g2551 <= g30382;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2555 <= 0;
  else
    g2555 <= g33600;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2606 <= 0;
  else
    g2606 <= g33607;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2599 <= 0;
  else
    g2599 <= g33601;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2629 <= 0;
  else
    g2629 <= g33602;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2643 <= 0;
  else
    g2643 <= g34020;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2648 <= 0;
  else
    g2648 <= g33603;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2567 <= 0;
  else
    g2567 <= g34021;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2563 <= 0;
  else
    g2563 <= g34015;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2571 <= 0;
  else
    g2571 <= g34016;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2583 <= 0;
  else
    g2583 <= g34019;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2579 <= 0;
  else
    g2579 <= g34018;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2575 <= 0;
  else
    g2575 <= g34017;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2595 <= 0;
  else
    g2595 <= g30383;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2587 <= 0;
  else
    g2587 <= g33015;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2610 <= 0;
  else
    g2610 <= g33016;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2625 <= 0;
  else
    g2625 <= g33018;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2619 <= 0;
  else
    g2619 <= g33017;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2638 <= 0;
  else
    g2638 <= g29254;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2652 <= 0;
  else
    g2652 <= g29255;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2657 <= 0;
  else
    g2657 <= g30384;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2661 <= 0;
  else
    g2661 <= g30385;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2667 <= 0;
  else
    g2667 <= g33604;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2671 <= 0;
  else
    g2671 <= g33605;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2675 <= 0;
  else
    g2675 <= g33606;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2681 <= 0;
  else
    g2681 <= g30386;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2685 <= 0;
  else
    g2685 <= g30387;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2689 <= 0;
  else
    g2689 <= g34606;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2697 <= 0;
  else
    g2697 <= g34607;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2704 <= 0;
  else
    g2704 <= g34608;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2710 <= 0;
  else
    g2710 <= g18527;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2711 <= 0;
  else
    g2711 <= g18528;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2837 <= 0;
  else
    g2837 <= g26935;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2841 <= 0;
  else
    g2841 <= g26936;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2712 <= 0;
  else
    g2712 <= g26937;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2715 <= 0;
  else
    g2715 <= g24263;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2719 <= 0;
  else
    g2719 <= g25639;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2724 <= 0;
  else
    g2724 <= g26926;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2729 <= 0;
  else
    g2729 <= g28060;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2735 <= 0;
  else
    g2735 <= g29256;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2741 <= 0;
  else
    g2741 <= g30388;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2748 <= 0;
  else
    g2748 <= g31872;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2756 <= 0;
  else
    g2756 <= g33019;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2759 <= 0;
  else
    g2759 <= g33608;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2763 <= 0;
  else
    g2763 <= g34022;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2767 <= 0;
  else
    g2767 <= g26927;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2779 <= 0;
  else
    g2779 <= g26928;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2791 <= 0;
  else
    g2791 <= g26929;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2795 <= 0;
  else
    g2795 <= g26930;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2787 <= 0;
  else
    g2787 <= g34444;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2783 <= 0;
  else
    g2783 <= g34442;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2775 <= 0;
  else
    g2775 <= g34443;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2771 <= 0;
  else
    g2771 <= g34441;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2831 <= 0;
  else
    g2831 <= g30391;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g121 <= 0;
  else
    g121 <= g30389;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2799 <= 0;
  else
    g2799 <= g26931;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2811 <= 0;
  else
    g2811 <= g26932;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2823 <= 0;
  else
    g2823 <= g26933;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2827 <= 0;
  else
    g2827 <= g26934;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2819 <= 0;
  else
    g2819 <= g34448;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2815 <= 0;
  else
    g2815 <= g34446;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2807 <= 0;
  else
    g2807 <= g34447;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2803 <= 0;
  else
    g2803 <= g34445;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2834 <= 0;
  else
    g2834 <= g30392;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g117 <= 0;
  else
    g117 <= g30390;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2999 <= 0;
  else
    g2999 <= g34805;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2994 <= 0;
  else
    g2994 <= g34732;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2988 <= 0;
  else
    g2988 <= g34624;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2868 <= 0;
  else
    g2868 <= g34616;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2873 <= 0;
  else
    g2873 <= g34615;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2890 <= 0;
  else
    g2890 <= g34799;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2844 <= 0;
  else
    g2844 <= g34609;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2852 <= 0;
  else
    g2852 <= g34610;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2860 <= 0;
  else
    g2860 <= g34611;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2894 <= 0;
  else
    g2894 <= g34612;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g37 <= 0;
  else
    g37 <= g34613;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g94 <= 0;
  else
    g94 <= g34614;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2848 <= 0;
  else
    g2848 <= g34792;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2856 <= 0;
  else
    g2856 <= g34793;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2864 <= 0;
  else
    g2864 <= g34794;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2898 <= 0;
  else
    g2898 <= g34795;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2882 <= 0;
  else
    g2882 <= g34796;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2878 <= 0;
  else
    g2878 <= g34797;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2886 <= 0;
  else
    g2886 <= g34798;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2980 <= 0;
  else
    g2980 <= g34800;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2984 <= 0;
  else
    g2984 <= g34980;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2907 <= 0;
  else
    g2907 <= g34617;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2912 <= 0;
  else
    g2912 <= g34618;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2922 <= 0;
  else
    g2922 <= g34619;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2936 <= 0;
  else
    g2936 <= g34620;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2950 <= 0;
  else
    g2950 <= g34621;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2960 <= 0;
  else
    g2960 <= g34622;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2970 <= 0;
  else
    g2970 <= g34623;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2902 <= 0;
  else
    g2902 <= g34801;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2917 <= 0;
  else
    g2917 <= g34802;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2927 <= 0;
  else
    g2927 <= g34803;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2941 <= 0;
  else
    g2941 <= g34806;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2955 <= 0;
  else
    g2955 <= g34807;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2965 <= 0;
  else
    g2965 <= g34808;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2975 <= 0;
  else
    g2975 <= g34804;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3003 <= 0;
  else
    g3003 <= g21726;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5 <= 0;
  else
    g5 <= g12833;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6 <= 0;
  else
    g6 <= g34589;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g7 <= 0;
  else
    g7 <= g34590;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g8 <= 0;
  else
    g8 <= g34591;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g9 <= 0;
  else
    g9 <= g34592;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g16 <= 0;
  else
    g16 <= g34593;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g19 <= 0;
  else
    g19 <= g34594;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g28 <= 0;
  else
    g28 <= g34595;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g31 <= 0;
  else
    g31 <= g34596;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g34 <= 0;
  else
    g34 <= g34877;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g12 <= 0;
  else
    g12 <= g30326;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g22 <= 0;
  else
    g22 <= g29209;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g25 <= 0;
  else
    g25 <= g15048;
assign g18281 = (g1373&g16136);
assign II28897 = ((~g30155));
assign g20592 = ((~g15277));
assign II26071 = ((~g26026))|((~II26070));
assign g24124 = ((~g21209));
assign g31542 = (g19050&g29814);
assign g31799 = ((~g29385));
assign II13463 = ((~g2380))|((~II13462));
assign g30503 = (g30243)|(g22024);
assign g22225 = (g21332)|(g17654);
assign g24850 = ((~II24022));
assign g32057 = ((~g31003))|((~g13297));
assign g10306 = ((~II13726));
assign g17674 = ((~II18647));
assign g13491 = (g6999&g12160);
assign g28911 = ((~g27907))|((~g7456))|((~g2465));
assign g14745 = ((~g12423));
assign II15363 = ((~g10182))|((~g2675));
assign II15147 = ((~g9864))|((~g5659));
assign g30086 = (g28536&g20704);
assign g24362 = ((~g21370))|((~g22136));
assign g21718 = (g370&g21037);
assign g8508 = ((~g3827));
assign II14712 = ((~g9671))|((~g5128));
assign g30484 = (g30154)|(g21980);
assign g32453 = ((~II29981));
assign g33602 = (g33425)|(g18511);
assign g29928 = ((~g28871));
assign g20549 = ((~g15277));
assign g34089 = (g22957&g9104&g33744);
assign g9977 = ((~g2667));
assign g27059 = ((~g7577)&(~g25895));
assign g20649 = ((~g18065));
assign g21930 = (g5180&g18997);
assign g9700 = ((~g2361)&(~g2287));
assign g17417 = ((~g14804));
assign g32491 = ((~g31566));
assign II32535 = ((~g34296));
assign g30384 = (g30101)|(g18517);
assign g24396 = ((~g22885));
assign g31471 = (g29754&g23399);
assign g32767 = ((~g30735));
assign g21693 = ((~II21254));
assign g19524 = ((~g15695));
assign g34351 = ((~g34174));
assign g34132 = ((~g33831));
assign II18509 = ((~g5623));
assign g24600 = (g22591&g19652);
assign g16508 = ((~II17704));
assign g22712 = ((~g18957))|((~g2864));
assign g13626 = ((~g11273));
assign g22527 = ((~g19546));
assign g28160 = (g26309&g27463);
assign II12994 = ((~g6748));
assign g27547 = (g26549&g17759);
assign g24903 = (g128&g23889);
assign g21458 = ((~g15758));
assign g16530 = ((~g14454));
assign g26632 = ((~g25473));
assign g7252 = ((~g1592));
assign g22719 = ((~II22024));
assign II20203 = ((~g16246))|((~g11147));
assign g32879 = ((~g31327));
assign g34370 = (g34067&g10554);
assign g32226 = (g31145)|(g29645);
assign II21802 = ((~g21308));
assign g8938 = ((~g4899));
assign g32852 = ((~g30614));
assign g23609 = ((~g21611));
assign g18644 = (g15098&g17125);
assign g24985 = ((~g23586));
assign g25907 = (g24799&g22519);
assign II13240 = ((~g5794));
assign g34643 = (g34554)|(g18752);
assign g15647 = ((~g11924)&(~g14248));
assign g14394 = ((~g12116)&(~g9414));
assign g28840 = ((~g27858))|((~g7380))|((~g2287));
assign II20542 = ((~g16508));
assign g33470 = (g32528&II31046&II31047);
assign II12041 = ((~g2741));
assign g7521 = ((~g5630));
assign g29308 = (g28612)|(g18815);
assign g33097 = ((~g31950)&(~g4628));
assign II18307 = ((~g12977));
assign g32274 = (g31256&g20447);
assign g17296 = ((~II18280));
assign g29740 = (g2648&g29154);
assign g12855 = ((~g10430)&(~g6854));
assign g32910 = ((~g31327)&(~II30468)&(~II30469));
assign g33592 = (g33412)|(g18475);
assign g21780 = (g3391&g20391);
assign g31239 = ((~g29916));
assign g15348 = ((~II17111));
assign g31883 = (g31132)|(g21777);
assign g12193 = ((~g2342)&(~g8316));
assign g25200 = ((~g5742))|((~g23642));
assign g22036 = (g5937&g19147);
assign II16526 = ((~g10430));
assign g32438 = ((~g30991));
assign g19765 = ((~g16897));
assign II21047 = ((~g17429));
assign g17694 = ((~g12435)&(~g12955));
assign g22220 = ((~II21802));
assign g12300 = ((~II15144));
assign g29295 = (g28663)|(g18780);
assign g28186 = (g27209)|(g27185)|(g27161)|(g27146);
assign gbuf3 = (g4571);
assign g23276 = (g19681)|(g16161);
assign g28773 = (g27535)|(g16803);
assign g28619 = (g27358)|(g16517);
assign g8106 = ((~g3133));
assign g10230 = ((~II13694));
assign g29301 = (g28686)|(g18797);
assign g19449 = (g15567)|(g12939);
assign g32943 = ((~g31710));
assign g11232 = ((~g4966)&(~g7898)&(~g9064));
assign g6847 = ((~g2283));
assign g33669 = ((~g33378))|((~g862));
assign g31772 = (g30035)|(g28654);
assign g10882 = ((~g7601));
assign g27481 = (g26400&g14630);
assign g19638 = ((~g17324));
assign g29873 = ((~g6875)&(~g28458));
assign g22625 = (g18910)|(g18933);
assign g25317 = ((~g9766)&(~g23782));
assign g20573 = ((~g17384));
assign g15809 = (g3917&g14154);
assign g23984 = ((~g19210));
assign g15053 = ((~g12836)&(~g13350));
assign II32225 = ((~g34121));
assign II12070 = ((~g785));
assign g18334 = (g1696&g17873);
assign g6827 = ((~g1277));
assign g29846 = ((~g28391));
assign g34706 = (g34496&g10570);
assign g14764 = ((~g7738))|((~g12798));
assign g8130 = ((~g4515));
assign II13509 = ((~g2089))|((~g2093));
assign g20240 = ((~g17847));
assign g23183 = (g19545)|(g15911);
assign g24196 = (g333&g22722);
assign g32772 = ((~g31327));
assign g24906 = ((~g8743))|((~g23088));
assign g29336 = (g4704&g28363);
assign g25544 = ((~g22594));
assign g30376 = (g30112)|(g18471);
assign g8123 = ((~g3808));
assign g25630 = (g24532)|(g18263);
assign g12868 = ((~g10377));
assign g33874 = ((~II31724));
assign g34249 = (g34110)|(g21702);
assign g30608 = (g13604)|(g29736);
assign g32803 = ((~g31376));
assign g16066 = ((~g10929)&(~g13307));
assign g11907 = ((~g7170)&(~g7184));
assign g8032 = ((~II12355));
assign g18465 = (g2384&g15224);
assign g23297 = (g19692)|(g16178);
assign g25564 = ((~g22312));
assign g17652 = ((~g15033));
assign g11584 = ((~g8229)&(~g8172));
assign g23313 = ((~g21070));
assign g13413 = ((~g11737));
assign g32663 = ((~g30673));
assign g32510 = ((~g31194));
assign II26880 = ((~g27527));
assign g19432 = ((~g15885));
assign g32343 = (g31473&g20710);
assign II23321 = ((~g21693));
assign g34544 = ((~II32613));
assign g21876 = (g4119&g19801);
assign g33694 = (g32402)|(g33429);
assign g18250 = (g6821&g16897);
assign II17919 = ((~g14609));
assign g30219 = (g28698&g23887);
assign g31762 = (g30011)|(g30030);
assign g30423 = (g29887)|(g21807);
assign g32131 = (g24495)|(g30926);
assign II11682 = ((~g2756));
assign g21657 = ((~g17657));
assign g25639 = (g25122)|(g18530);
assign g28052 = (g27710)|(g18167);
assign g34193 = (g33809)|(g33814);
assign g19903 = ((~g13707))|((~g16319))|((~g8227));
assign g14489 = ((~g12126))|((~g5084));
assign g29575 = (g2066&g28604);
assign g34833 = ((~II33047));
assign g12921 = ((~g12228));
assign g33675 = (g33164&g10727&g22332);
assign g17821 = ((~II18829));
assign g32914 = ((~g31672));
assign g31278 = (g29716&g23302);
assign g34334 = (g34090&g19865);
assign g32312 = (g31302&g20591);
assign g27523 = (g26549&g17718);
assign g11900 = ((~II14708));
assign g29151 = ((~g27858));
assign g17136 = ((~g14348));
assign g10217 = ((~g2102));
assign g23051 = ((~g7960)&(~g19427));
assign g34112 = (g22957&g9104&g33778);
assign g32557 = ((~g31376));
assign II29218 = ((~g30304));
assign g25232 = ((~g22228));
assign g10117 = ((~g2509));
assign g8804 = ((~g4035));
assign g33088 = ((~g31997)&(~g7224));
assign g20273 = ((~g17128));
assign g22142 = (g7957&g19140);
assign g29246 = (g28710)|(g18406);
assign g28361 = (g27153)|(g15839);
assign g34272 = ((~g34229));
assign g23994 = ((~g19277));
assign II14332 = ((~g9966))|((~II14330));
assign g27479 = ((~g9056)&(~g26616));
assign g32830 = ((~g31327));
assign g15148 = ((~g13716)&(~g12893));
assign g28059 = (g27042)|(g18276);
assign g33729 = ((~II31586));
assign g7297 = ((~g6069));
assign II11753 = ((~g4492));
assign II17207 = ((~g13835));
assign g11811 = ((~g9724));
assign g32211 = (g31124)|(g29603);
assign II16460 = ((~g10430));
assign g18994 = (g16303)|(g13632);
assign g23337 = ((~g20924));
assign g32987 = (g32311)|(g18323);
assign g16701 = (g5547&g14845);
assign g30469 = (g30153)|(g21940);
assign g24796 = (g7097&g23714);
assign g33233 = (g32094&g23005);
assign g24189 = (g324&g22722);
assign g7132 = ((~g4558));
assign g30333 = (g29834)|(g21699);
assign g32933 = ((~g31376));
assign g26277 = (g2547&g25400);
assign g32895 = ((~g30673));
assign g18389 = (g1974&g15171);
assign g27138 = (g26055&g16607);
assign g30302 = ((~g28924));
assign g9360 = ((~g3372));
assign g34406 = (g34184)|(g25123);
assign g17790 = ((~g6311))|((~g14575))|((~g6322))|((~g10003));
assign g30150 = ((~g28846)&(~g7424));
assign g10400 = ((~g7002));
assign g26301 = (g2145&g25244);
assign g24946 = (g22360)|(g22409)|(g8130);
assign g22638 = ((~g18957))|((~g2886));
assign g27184 = (g26628&g13756);
assign g18349 = (g1768&g17955);
assign g8678 = ((~g376))|((~g358));
assign g18391 = (g1982&g15171);
assign g9011 = ((~g1422));
assign g12804 = ((~g9927));
assign g20496 = ((~g17929));
assign g8137 = ((~g411));
assign g10405 = ((~g7064));
assign g22855 = ((~g20391));
assign II14893 = ((~g9819));
assign g28151 = (g8426&g27295);
assign g12179 = (g9745&g10027);
assign II22845 = ((~g12113))|((~II22844));
assign g24565 = (g22309)|(g19275);
assign g29362 = (g27379&g28307);
assign g7537 = ((~g311));
assign g28344 = (g27136)|(g15820);
assign g32283 = (g31259&g20506);
assign g16661 = ((~g14454));
assign g10099 = ((~g6682));
assign g9582 = ((~g703));
assign g22086 = (g6299&g19210);
assign g24149 = ((~g19338));
assign g30491 = (g30178)|(g21987);
assign g13656 = (g278&g11144);
assign g15720 = ((~g5917))|((~g14497))|((~g6019))|((~g9935));
assign g26606 = (g1018&g24510);
assign g33888 = ((~g33346));
assign g24069 = ((~g19968));
assign g31301 = (g30170&g27907);
assign g33109 = ((~g31997)&(~g4584));
assign g17637 = ((~g12933));
assign II29720 = ((~g30931));
assign g9914 = ((~g2533));
assign g33090 = ((~g31997)&(~g4593));
assign g13047 = (g8534&g11042);
assign g15867 = ((~g14714))|((~g9417))|((~g9340));
assign g34880 = (g34867)|(g18153);
assign g24427 = (g4961&g22919);
assign g32356 = (g2704&g31710);
assign g16179 = (g6187&g14321);
assign g25740 = (g25164)|(g22055);
assign g12126 = ((~g9989)&(~g5069));
assign g11169 = ((~II14229))|((~II14230));
assign g12041 = ((~II14905));
assign g33128 = ((~g4653)&(~g32057));
assign g13138 = ((~II15765));
assign g25781 = ((~g24510));
assign g29948 = ((~g28853));
assign g12122 = ((~g9705));
assign II26004 = ((~g26818));
assign g20614 = ((~g15426));
assign g16795 = ((~II18009));
assign II22900 = ((~g12193))|((~II22899));
assign g6900 = ((~g3440));
assign g22117 = (g6597&g19277);
assign g30228 = (g28715&g23903);
assign g18803 = (g15161&g15480);
assign g18531 = (g2719&g15277);
assign g33881 = (g33292&g20586);
assign g11344 = ((~g9015));
assign g30245 = (g28733&g23935);
assign g24300 = (g15123&g22228);
assign g23917 = (g1472&g19428);
assign g17954 = ((~g832)&(~g14279));
assign g27575 = (g26147)|(g24731);
assign g28753 = ((~II27235));
assign g26357 = (g22547&g25525);
assign g16767 = ((~II17989));
assign g34728 = (g34661)|(g18214);
assign g17740 = ((~g5945))|((~g14497))|((~g6012))|((~g12351));
assign g27693 = ((~g25216))|((~g26752));
assign g30998 = ((~g29719));
assign g33935 = ((~II31817));
assign g26667 = ((~g23642)&(~g25175));
assign g34252 = (g34146)|(g18180);
assign g25106 = (g17391&g23506);
assign g29485 = (g28535)|(g27594);
assign g16766 = (g6649&g12915);
assign g34152 = ((~II32109));
assign II26440 = ((~g14271))|((~II26438));
assign g9825 = ((~II13391))|((~II13392));
assign g13477 = ((~II15954));
assign g27401 = ((~II26094))|((~II26095));
assign g27635 = (g23032&g26281&g26424&g24996);
assign g14376 = ((~g12126));
assign g8373 = ((~g2485));
assign g18263 = (g1249&g16000);
assign g12217 = ((~II15070));
assign g34242 = ((~II32225));
assign g32609 = ((~g30735));
assign g11045 = (g5787&g9883);
assign g16800 = (g13436)|(g11027);
assign g24003 = ((~g21514));
assign II13054 = ((~g6744));
assign g18954 = ((~g17427));
assign g25032 = ((~g23639));
assign g25946 = (g24496&g19537);
assign g24088 = ((~g21209));
assign g30265 = ((~g7051)&(~g29036));
assign g25131 = ((~g23699));
assign g15911 = (g3111&g13530);
assign g14443 = ((~II16596));
assign II15702 = ((~g12217));
assign II12314 = ((~g1500));
assign g18286 = (g1404&g16164);
assign g29996 = ((~g28962));
assign g34566 = (g34376&g17489);
assign g33625 = (g33373)|(g18809);
assign g31803 = ((~g29385));
assign g33974 = (g33846)|(g18345);
assign g21248 = ((~g15224));
assign g10373 = ((~g6917));
assign g11924 = ((~g7187)&(~g7209));
assign g24045 = ((~g21193));
assign g18917 = ((~g16077));
assign g26161 = (g2518&g25139);
assign g30550 = (g30226)|(g22121);
assign II29447 = ((~g30729));
assign II23971 = ((~g490))|((~II23969));
assign g23215 = ((~g20785));
assign g23563 = ((~g20682));
assign g9200 = ((~g1548));
assign g14785 = ((~g12629));
assign g29973 = (g28981&g9206);
assign g10762 = ((~g8470));
assign g30568 = ((~g29339));
assign g8915 = ((~II12884));
assign g24359 = ((~g22550));
assign g16752 = ((~II17976));
assign g29257 = (g28228)|(g18600);
assign g12233 = ((~g10338));
assign II18143 = ((~g13350));
assign g18268 = (g1280&g16000);
assign g30344 = (g29630)|(g18298);
assign II18285 = ((~g13638));
assign g34001 = (g33844)|(g18450);
assign II20167 = ((~g990))|((~II20165));
assign II16679 = ((~g12039));
assign g27133 = (g25788)|(g24392);
assign g30010 = (g29035&g9274);
assign g26145 = (g11962&g25131);
assign g17809 = (g7873&g13125);
assign II28594 = ((~g29379));
assign g17608 = ((~g5953))|((~g12067))|((~g5969))|((~g14701));
assign g15966 = (g3462&g13555);
assign g33287 = (g32146)|(g29586);
assign g31797 = ((~g29385));
assign g33778 = ((~II31625));
assign g16886 = ((~II18078));
assign g18427 = (g2181&g18008);
assign g30526 = (g30181)|(g22072);
assign g32441 = ((~II29969));
assign II26960 = (g24995&g26424&g22698);
assign g26614 = ((~g25426));
assign II13374 = ((~g6490));
assign II31256 = (g31021&g31841&g32824&g32825);
assign g27508 = (g26549&g17684);
assign g30296 = ((~g28889));
assign g18884 = ((~g15938));
assign g24034 = ((~g19968));
assign II11992 = ((~g763));
assign g17778 = ((~II18778));
assign g30403 = (g29750)|(g21762);
assign g26206 = (g2523&g25495);
assign g18791 = (g6044&g15634);
assign g13098 = ((~g5933))|((~g12129))|((~g6023))|((~g9935));
assign g20133 = ((~g17668))|((~g17634))|((~g17597))|((~g14569));
assign g30288 = ((~g7087)&(~g29073));
assign g10616 = (g7998&g174);
assign g32085 = (g27253&g31021);
assign g25788 = (g8010&g24579);
assign g12340 = ((~g4888))|((~g8984));
assign g10543 = (g8238&g437);
assign g25977 = (g25236&g20875);
assign g7495 = ((~g4375));
assign g29175 = ((~g6227)&(~g26977));
assign g27317 = ((~g24793))|((~g26255));
assign g29943 = (g2165&g28765);
assign g25627 = (g24503)|(g18247);
assign g18656 = (g15120&g17128);
assign g12505 = ((~g9444)&(~g9381));
assign g24257 = (g22938)|(g18310);
assign g34311 = ((~g34097));
assign g28211 = (g27029)|(g27034);
assign g20526 = ((~g15171));
assign g23489 = ((~g21468));
assign g10165 = ((~g5698));
assign II25606 = ((~g25465));
assign g17793 = (g6772&g11592&g6789&II18803);
assign g26872 = ((~g25411)&(~g25371));
assign g16708 = ((~II17916));
assign g32742 = ((~g31021));
assign g33131 = ((~g4659)&(~g32057));
assign g26826 = (g24907&g15747);
assign g14309 = (g10320)|(g11048);
assign II13889 = ((~g7598));
assign g7049 = ((~g5853));
assign g19861 = ((~g17096));
assign g34462 = (g34334)|(g18685);
assign II27492 = ((~g27511));
assign g33056 = (g32327)|(g22004);
assign g25261 = (g23348)|(g20193);
assign g18811 = (g6500&g15483);
assign g25994 = ((~g24575));
assign g27298 = (g26573&g23026);
assign g30159 = ((~g28799)&(~g14589));
assign g33322 = (g32202&g20450);
assign g8844 = ((~II12826));
assign g34593 = ((~II32687));
assign g34980 = (g34969)|(g18587);
assign g17157 = ((~g13350));
assign g13022 = ((~g11894));
assign g33823 = ((~g8774)&(~g33306)&(~g11083));
assign g34221 = ((~II32192));
assign g18373 = (g1890&g15171);
assign g29288 = (g28630)|(g18762);
assign g18653 = (g4176&g16249);
assign II19759 = ((~g17767));
assign g33102 = (g32399&g18978);
assign gbuf130 = (g884);
assign g16733 = (g5893&g14889);
assign g31861 = ((~II29441));
assign II29973 = ((~g31213));
assign g29641 = (g28520&g14237);
assign g17248 = ((~II18262));
assign g6977 = ((~II11753));
assign II15088 = ((~g9832))|((~II15087));
assign g25165 = (g14062&g23570);
assign g27590 = (g26179)|(g24764);
assign g31839 = ((~g29385));
assign g21939 = (g5224&g18997);
assign II18373 = ((~g13011));
assign g16484 = (g5244&g14755);
assign II15052 = ((~g9759))|((~II15051));
assign II15782 = ((~g10430));
assign g26902 = (g26378)|(g24219);
assign g32498 = ((~g31566));
assign g29478 = (g28111)|(g22160);
assign II14427 = ((~g8595))|((~g4005));
assign II12278 = ((~g1467))|((~II12277));
assign g24237 = (g22515)|(g18242);
assign g25596 = (g24865)|(g21718);
assign g11324 = ((~g7542));
assign g10140 = ((~g19));
assign II15213 = ((~g10035))|((~II15212));
assign g14616 = ((~II16733));
assign g6804 = ((~g490));
assign gbuf35 = (g5448);
assign g34769 = ((~II32953));
assign g31658 = ((~II29242));
assign g7908 = ((~g4157));
assign g28220 = (g23495)|(II26741)|(II26742);
assign g23781 = ((~II22937))|((~II22938));
assign g32483 = ((~g30673));
assign II23587 = ((~g4332))|((~II23585));
assign g33492 = (g32686&II31156&II31157);
assign g19782 = ((~II20188))|((~II20189));
assign g33868 = (g33278&g20542);
assign g24846 = (g3361&g23555&II24018);
assign g21913 = (g5069&g21468);
assign II32840 = ((~g34480));
assign g27310 = (g26574&g23059);
assign g28612 = (g27524&g20539);
assign g24673 = (g22659&g19748);
assign II19487 = ((~g15125));
assign II27927 = ((~g28803));
assign g23863 = ((~g19210));
assign g23476 = ((~g21468));
assign g18188 = (g807&g17328);
assign g28918 = ((~g27832));
assign g23289 = ((~g20924));
assign g19686 = ((~g17062));
assign II32815 = ((~g34470));
assign g15562 = ((~g14943));
assign g13251 = ((~II15814));
assign g28761 = (g21434&g26424&g25299&g27416);
assign II16855 = ((~g10473));
assign II31056 = (g30735&g31805&g32536&g32537);
assign II22894 = ((~g21228))|((~II22892));
assign g10043 = ((~g1632));
assign g28524 = (g6821&g27084);
assign g10653 = ((~g10204))|((~g10042));
assign g28903 = ((~g27800))|((~g2197))|((~g7280));
assign g23941 = ((~g19074));
assign II17140 = ((~g13835));
assign g28977 = ((~g27937))|((~g2629))|((~g2555));
assign g18402 = (g2047&g15373);
assign g28108 = (g7975&g27237);
assign II15334 = ((~g10152))|((~II15333));
assign g27252 = (g26733&g26703);
assign g19720 = ((~II20130));
assign g8026 = ((~g3857));
assign g25833 = (g8228&g24626);
assign g33796 = (g33117&g25267);
assign g23234 = ((~g20375));
assign g34314 = (g25831)|(g34061);
assign g17597 = ((~g3191))|((~g13700))|((~g3303))|((~g8481));
assign II14455 = ((~g10197));
assign g25924 = (g24976&g16846);
assign g9305 = ((~g5381));
assign g24725 = (g19587&g23012);
assign g20385 = ((~g18008));
assign g17491 = ((~g12983));
assign g17578 = ((~g5212))|((~g14399))|((~g5283))|((~g12497));
assign g34124 = ((~g33819));
assign g27772 = ((~g7297)&(~g25839));
assign g23433 = ((~g21562));
assign g22980 = ((~II22153));
assign II27429 = (g25562&g26424&g22698);
assign II16613 = ((~g10430));
assign g25517 = ((~g22228));
assign II18120 = ((~g13350));
assign g29181 = ((~g6573)&(~g26994));
assign g17177 = (g6657&g14984);
assign g33809 = (g33432&g30184);
assign g24973 = ((~g21272))|((~g23462));
assign g32575 = ((~g31170));
assign g29093 = ((~g27858));
assign g31926 = (g31765)|(g22090);
assign g8131 = ((~g4776)&(~g4801)&(~g4793));
assign g18439 = (g2250&g18008);
assign g15118 = (g4253&g14454);
assign g17844 = ((~II18832));
assign g16646 = ((~g13437)&(~g11020)&(~g11372));
assign g8426 = ((~g3045));
assign g19710 = ((~g17059));
assign g15747 = ((~g13307));
assign g29267 = (g28257)|(g18622);
assign g25533 = ((~g22550));
assign g19371 = ((~II19857));
assign g33619 = (g33359)|(g18758);
assign g30200 = (g28665&g23862);
assign g24411 = (g4584&g22161);
assign g34672 = ((~II32800));
assign g34288 = (g26846)|(g34217);
assign g23352 = ((~g20924));
assign g13909 = ((~g11396))|((~g8847))|((~g11674))|((~g8803));
assign g13498 = ((~g12577))|((~g12522))|((~g12462))|((~g12416));
assign g26610 = (g14198&g24405);
assign g18777 = (g5808&g18065);
assign g31850 = ((~g29385));
assign II13723 = ((~g3167));
assign II33152 = ((~g34900));
assign g21609 = ((~g18008));
assign g21755 = (g3203&g20785);
assign g22045 = (g6069&g21611);
assign g29591 = (g28552&g11346);
assign g13540 = (g10822)|(g10827);
assign g20004 = ((~g17249));
assign g26572 = (g7443&g24439);
assign g32600 = ((~g31542));
assign II32074 = ((~g33670));
assign g23410 = ((~g21562));
assign g8434 = ((~g3080))|((~g3072));
assign g18719 = (g4894&g16795);
assign g9048 = ((~II12963));
assign g18939 = ((~g16077));
assign g34295 = (g34057&g19370);
assign g23252 = ((~II22353));
assign g21993 = (g5603&g19074);
assign g23436 = (g676&g20375);
assign g14993 = ((~g12695))|((~g12453));
assign g14516 = ((~g12227)&(~g9704));
assign g25067 = (g4722&g22885);
assign gbuf121 = (g4232);
assign II16629 = ((~g11987));
assign g34497 = (g34275&g33072);
assign g15843 = ((~g7922))|((~g7503))|((~g13264));
assign g27692 = (g26392&g20697);
assign g18726 = (g4927&g16077);
assign g21306 = ((~g15582));
assign g25057 = (g23275&g20511);
assign g24014 = (g7933&g19063);
assign g28693 = ((~g27837));
assign g20265 = ((~g17821));
assign II17750 = ((~g14383));
assign g33553 = (g33403)|(g18350);
assign II31500 = ((~g33176));
assign g34793 = (g34744)|(g18570);
assign g14094 = ((~g8770)&(~g11083));
assign II23118 = ((~g20076))|((~g417));
assign g20516 = ((~II20609));
assign g19397 = ((~g16449));
assign g21746 = (g3045&g20330);
assign g16670 = (g5953&g14999);
assign II32096 = ((~g33641));
assign g32182 = (g31753&g27937);
assign g14173 = ((~g12076));
assign g29005 = ((~g5164)&(~g7704)&(~g27999));
assign gbuf23 = (g5335);
assign g32336 = (g31596&g11842);
assign g22869 = ((~g20875));
assign g25715 = (g25071)|(g21966);
assign g28255 = (g8515&g27983);
assign g30521 = (g29331)|(g22042);
assign g33511 = (g32823&II31251&II31252);
assign g22147 = ((~g18997));
assign g12847 = ((~g6838)&(~g10430));
assign g7869 = ((~II12252))|((~II12253));
assign g10102 = ((~g6727));
assign g22179 = ((~g19210));
assign II23378 = ((~g23426));
assign g16524 = ((~g13822))|((~g13798));
assign gbuf76 = (g3317);
assign II30537 = ((~g32027));
assign g19421 = ((~g16326));
assign g34738 = (g34660&g33442);
assign g10175 = ((~g28));
assign II12141 = ((~g599));
assign g18541 = (g2767&g15277);
assign g15121 = ((~g12874)&(~g13605));
assign g31374 = (g29748&g23390);
assign g18203 = (g911&g15938);
assign g30026 = (g28476&g25064);
assign g25667 = (g24682)|(g18619);
assign g30123 = ((~g28768)&(~g7328));
assign g34069 = (g8774&g33797);
assign g30593 = ((~g29970));
assign g32013 = (g8673&g30614);
assign g31527 = (g7553&g29343);
assign g8531 = ((~g3288));
assign g27653 = (g26549&g15562);
assign g26154 = (g1830&g25426);
assign g22862 = (g1570&g19673);
assign g32651 = ((~g31376));
assign g27675 = ((~II26309));
assign g19490 = ((~g16489));
assign g32054 = (g10890&g30735);
assign g16688 = ((~g14045));
assign g15810 = (g3937&g14055);
assign g21751 = (g3167&g20785);
assign g31248 = (g25970)|(g29522);
assign g14192 = ((~g11385));
assign g7095 = ((~g6545));
assign g26124 = (g1811&g25116);
assign g16839 = (g13473)|(g11035);
assign g34922 = ((~II33158));
assign g11884 = ((~g8125));
assign g17687 = ((~g15042));
assign II15340 = ((~g10154))|((~g2541));
assign g27086 = (g25836&g22495);
assign g25967 = (g9373&g24986);
assign g14014 = ((~g3199))|((~g11217))|((~g3298))|((~g11519));
assign g13972 = (g11232)|(g11203);
assign g34850 = (g34841)|(g18185);
assign II22419 = ((~g19638));
assign g6995 = ((~g4944));
assign g29638 = (g2583&g29025);
assign g30382 = (g30137)|(g18498);
assign g27570 = (g26126)|(g24722);
assign II31307 = (g32898&g32899&g32900&g32901);
assign g10918 = ((~g1532)&(~g7751)&(~g7778));
assign g11989 = ((~II14839));
assign g29911 = ((~g28780));
assign g13432 = ((~g4793))|((~g10831));
assign g34971 = (g34869)|(g34962);
assign II18634 = ((~g2504))|((~II18633));
assign g9040 = ((~g499));
assign g22660 = ((~g19140));
assign g29515 = (g28888&g22342);
assign g10204 = ((~g2685));
assign g21268 = ((~g15680));
assign g11834 = ((~g8938)&(~g8822));
assign g21970 = (g5401&g21514);
assign g17416 = ((~g14956));
assign g33385 = ((~g32038));
assign g32523 = ((~g30825));
assign g8620 = ((~g3065));
assign g18735 = (g4983&g16826);
assign g21812 = (g3586&g20924);
assign g34444 = (g34389)|(g18546);
assign II22965 = ((~g12288))|((~g21228));
assign g32750 = ((~g30937));
assign g16225 = ((~g13544))|((~g13528))|((~g13043));
assign g33267 = (g32115)|(g29535);
assign II13391 = ((~g1821))|((~II13390));
assign g21823 = (g3731&g20453);
assign g11237 = ((~II14305));
assign g30061 = (g1036&g28188);
assign g24009 = (g19671&g10971);
assign g11248 = ((~g7953)&(~g4991)&(~g4983));
assign g21977 = (g5535&g19074);
assign g33984 = (g33881)|(g18374);
assign g30205 = (g28671&g23869);
assign g12978 = ((~II15593));
assign g7926 = ((~g3423));
assign g28518 = (g27281)|(g26158);
assign g15723 = ((~g10775))|((~g13104));
assign II12773 = ((~g4204));
assign g31207 = (g30252&g20739);
assign g8069 = ((~II12373))|((~II12374));
assign g27907 = (g17424)|(g26770);
assign II20130 = ((~g15748));
assign g13853 = (g4549&g10620);
assign g14782 = ((~g12755))|((~g10491));
assign g15799 = ((~g13110));
assign g18228 = (g1061&g16129);
assign g23459 = ((~g21611));
assign g24160 = ((~II23324));
assign g25758 = (g25151)|(g22105);
assign g34514 = (g34286&g19480);
assign g14521 = ((~g12170))|((~g5428));
assign g20199 = ((~g16815))|((~g13968))|((~g16749))|((~g13907));
assign g29661 = (g1687&g29015);
assign g33051 = (g32316)|(g21958);
assign g14738 = ((~II16821));
assign g33357 = (g32247&g20775);
assign g15073 = ((~g12844)&(~g13416));
assign g8187 = ((~g1657));
assign g16930 = (g239&g13132);
assign II12770 = ((~g4200));
assign g28242 = (g27769&g23626);
assign g20053 = ((~g17328));
assign g28938 = ((~g27796))|((~g8205));
assign g27119 = (g25877&g22542);
assign g21846 = (g3897&g21070);
assign g33500 = (g32744&II31196&II31197);
assign II26195 = ((~g26260));
assign g14573 = ((~g9506))|((~g12249));
assign g30670 = (g11330&g29359);
assign g14933 = ((~g12700))|((~g12571));
assign g27435 = (g26549&g17585);
assign g14680 = (g12024&g12053);
assign g10902 = (g7858&g1129);
assign g20639 = ((~g15224));
assign g11033 = ((~g8500));
assign g20209 = ((~g17821));
assign g26753 = (g16024&g24452);
assign g33138 = ((~g32287)&(~g31514));
assign g33066 = (g32341)|(g22096);
assign g16479 = ((~g14719)&(~g12490));
assign g13075 = ((~II15705));
assign g32252 = (g31183)|(g31206);
assign g25706 = (g25030)|(g18748);
assign g33424 = ((~g32415));
assign II12841 = ((~g4222))|((~II12840));
assign g23009 = (g20196&g14219);
assign g12796 = ((~g4467))|((~g6961));
assign g23854 = (g4093&g19506);
assign g10365 = ((~g6867));
assign g28102 = (g27995)|(g22089);
assign g25526 = (g23720&g21400);
assign g31623 = ((~g29669));
assign g31505 = (g30195&g24379);
assign g32208 = (g31120)|(g29584);
assign g30042 = (g29142&g12601);
assign g18714 = (g4864&g15915);
assign II33182 = ((~g34910));
assign g34851 = ((~II33075));
assign II22316 = ((~g19361));
assign II11865 = ((~g4434))|((~II11864));
assign II31701 = ((~g33164));
assign g16193 = (g6533&g14348);
assign g13518 = ((~g3719)&(~g11903));
assign g12884 = ((~g10392));
assign g32348 = (g2145&g31672);
assign g17122 = ((~g14348));
assign g6986 = ((~g4743));
assign II15105 = ((~g9780))|((~g5313));
assign g25451 = ((~g22228));
assign g28466 = (g27960&g17637);
assign g16681 = ((~II17884))|((~II17885));
assign II27738 = ((~g28140));
assign II32947 = ((~g34659));
assign g33002 = (g32304)|(g18419);
assign g26835 = ((~II25555));
assign II12583 = (g1157)|(g1239)|(g990);
assign g22154 = ((~g19074));
assign g34789 = ((~II32997));
assign g18303 = (g1536&g16489);
assign g26957 = (g26517)|(g24295);
assign II33034 = ((~g34769));
assign g9214 = ((~g617));
assign g26330 = ((~g8631)&(~g24825));
assign g33827 = ((~II31672));
assign g10607 = ((~g10233));
assign II29961 = ((~g30984));
assign g33992 = (g33900)|(g18408);
assign g30229 = (g28716&g23904);
assign g34986 = ((~II33258));
assign g24998 = (g17412&g23408);
assign g29761 = (g28310&g23228);
assign g24078 = ((~g20857));
assign g32925 = ((~g31327));
assign g28997 = ((~g27903))|((~g8324));
assign g17404 = ((~II18337));
assign g26882 = (g26650)|(g24188);
assign g15124 = (g13605)|(g4581);
assign g32711 = ((~g31070));
assign g9630 = ((~g6527));
assign g12337 = ((~g9340));
assign g25110 = (g10427&g23509);
assign g26821 = (g24821&g13103);
assign g18183 = (g781&g17328);
assign g28381 = ((~g27074))|((~g13621));
assign g21673 = ((~II21234));
assign g21335 = ((~II21067));
assign g24172 = ((~II23360));
assign II31142 = (g32661&g32662&g32663&g32664);
assign g25022 = ((~g714)&(~g23324));
assign g30598 = (g18898&g29862);
assign II15474 = ((~g10364));
assign II19707 = ((~g17590));
assign g21275 = ((~g15426));
assign II31002 = (g32459&g32460&g32461&g32462);
assign g12645 = ((~g4467)&(~g6961));
assign g6941 = ((~g3990));
assign g20720 = ((~g17847)&(~g9299));
assign g19613 = (g1437&g16713);
assign g24714 = (g6173&g23699);
assign II30741 = (g32085)|(g32030)|(g32224)|(g32013);
assign g14882 = ((~g12558))|((~g12453));
assign g33715 = (g33135&g19416);
assign g29510 = (g28856&g22342);
assign g32932 = ((~g31327));
assign g32260 = (g31250&g20385);
assign g13280 = ((~II15846));
assign g32581 = ((~g31070));
assign g9766 = ((~g2748));
assign II15533 = ((~g11867));
assign g24337 = (g23540)|(g18754);
assign g15091 = ((~g13177)&(~g12863));
assign g21298 = (g7697&g15825);
assign g16579 = ((~g13267));
assign g25019 = ((~g20055))|((~g23172));
assign g32174 = (g31708&g27837);
assign g27236 = (g24620)|(g25974);
assign g25922 = (g24959&g20065);
assign g10586 = ((~g7380))|((~g7418));
assign II27232 = ((~g27993));
assign g25239 = ((~g23972));
assign g19597 = ((~g1199))|((~g15995));
assign g34196 = (g33682&g24485);
assign II26531 = (g24099&g24100&g24101&g24102);
assign g12197 = ((~g7296))|((~g5290));
assign g10475 = ((~g8844));
assign g23052 = ((~g8334)&(~g19916));
assign g20157 = ((~g16886));
assign g31868 = (g30600)|(g18204);
assign g31832 = ((~g29385));
assign g25655 = (g24645)|(g18607);
assign g9257 = ((~g5115));
assign g33375 = ((~g32377));
assign g24180 = ((~II23384));
assign g16635 = (g5607&g14959);
assign g26390 = (g4423&g25554);
assign g33341 = (g32223&g20640);
assign g19932 = ((~g3376)&(~g16296));
assign II21930 = ((~g21297));
assign g24726 = (g15965&g23015);
assign g23452 = ((~g21468));
assign g26920 = (g25865)|(g18283);
assign g31121 = ((~g4776)&(~g29540));
assign g32116 = (g31658&g29929);
assign gbuf55 = (g6369);
assign g32622 = ((~g31376));
assign g18607 = (g3139&g16987);
assign g24098 = ((~g19984));
assign g32229 = (g31148)|(g29652);
assign g13805 = (g11489&g11394&g11356&II16129);
assign g27697 = (g25785&g23649);
assign II21849 = ((~g19620));
assign g33501 = (g32751&II31201&II31202);
assign g31014 = (g29367)|(g28160);
assign g22834 = (g102&g19630);
assign g34947 = ((~g34938));
assign g14597 = ((~II16713));
assign g12819 = ((~g9848))|((~g6961));
assign g26487 = (g15702&g24359);
assign g13621 = ((~g10573));
assign g25600 = (g24650)|(g18111);
assign g10935 = ((~g1459))|((~g7352));
assign g22923 = ((~II22124));
assign g9442 = ((~g5424))|((~g5428));
assign g33877 = (g33287&g20563);
assign g33121 = (g8748&g32212);
assign g27315 = (g12022&g26709);
assign g17529 = ((~g15039));
assign g29226 = (g28455)|(g18159);
assign g10019 = ((~g6479));
assign g14002 = ((~g8681)&(~g11083));
assign g24536 = (g19516&g22635);
assign g30937 = (g22626&g29814);
assign g24022 = ((~g20982));
assign g22973 = ((~g20330));
assign g8341 = ((~g3119));
assign g21354 = ((~g11468))|((~g17157));
assign g27032 = (g7704&g5180&g5188&g26200);
assign g17188 = ((~II18224));
assign g10515 = ((~g10337))|((~g5022));
assign g10427 = ((~g10053));
assign g23746 = ((~g20902));
assign g10649 = ((~g1183)&(~g8407));
assign g11669 = ((~g3863)&(~g8026));
assign g24154 = ((~II23306));
assign II33155 = ((~g34897));
assign g21330 = ((~g11401))|((~g17157));
assign g26686 = ((~g23678)&(~g25189));
assign g25642 = ((~II24787));
assign g12947 = ((~g7184))|((~g10561));
assign II22711 = ((~g11915))|((~II22710));
assign II21776 = ((~g21308));
assign g7201 = ((~II11865))|((~II11866));
assign g29192 = (g27163&g10290);
assign II12344 = ((~g3106))|((~g3111));
assign g24588 = (g5142&g23590);
assign g29508 = (g28152)|(g27041);
assign g19206 = (g460&g16206);
assign g20663 = ((~g15373));
assign II15167 = ((~g9904))|((~II15166));
assign g31128 = (g12187&g30016);
assign g26948 = (g26399)|(g24286);
assign g26022 = (g25271&g20751);
assign g28316 = (g27113)|(g15804);
assign g10396 = ((~g6997));
assign g17431 = ((~II18376));
assign II24474 = ((~g22546));
assign II31337 = (g32942&g32943&g32944&g32945);
assign g12024 = ((~g8381))|((~g8418));
assign g33240 = (g32052)|(g32068);
assign g30371 = (g30099)|(g18445);
assign g29888 = (g28418&g23352);
assign g34457 = (g34394)|(g18670);
assign g29220 = ((~II27576));
assign g23512 = ((~g20248));
assign g33899 = (g32132&g33335);
assign g13896 = ((~g3227))|((~g11194))|((~g3281))|((~g11350));
assign g28249 = (g27152&g19677);
assign g11316 = ((~g8967));
assign II24705 = (g24064&g24065&g24066&g24067);
assign g8005 = ((~g3025));
assign II14647 = ((~g7717));
assign g15873 = (g3550&g14072);
assign g24572 = (g5462&g23393);
assign g32537 = ((~g30825));
assign g22685 = (g11891&g20192);
assign g26323 = (g10262&g25273);
assign g27369 = (g25894&g25324);
assign g26083 = ((~g24809));
assign g29494 = (g9073&g28479);
assign g29018 = ((~g9586))|((~g27742));
assign II12189 = ((~g5869));
assign g16986 = (g246&g13142);
assign g17755 = ((~g5619))|((~g14522))|((~g5630))|((~g9864));
assign g19736 = (g12136&g17136);
assign g13297 = ((~g10831));
assign g8354 = ((~g4815));
assign g34768 = ((~II32950));
assign g24083 = ((~g19984));
assign II31477 = ((~g33391));
assign g27279 = ((~g26330));
assign g14189 = ((~II16391));
assign g29639 = (g28510&g11618);
assign II12735 = ((~g4572));
assign g27251 = (g26721&g26694);
assign g13469 = ((~g4983))|((~g10862));
assign g34488 = (g34417&g18988);
assign g18741 = (g15143&g17384);
assign g32793 = ((~g31021));
assign g33966 = (g33837)|(g18318);
assign g15935 = (g13029)|(g10665);
assign g31931 = (g31494)|(g22095);
assign g14744 = ((~g12578));
assign g18177 = (g749&g17328);
assign g31295 = (g26090)|(g29598);
assign II26687 = ((~g27880));
assign g25151 = (g17719&g23549);
assign g26927 = (g26711)|(g18539);
assign g28631 = (g27372)|(g16534);
assign g29049 = ((~g9640))|((~g27779));
assign g13939 = ((~g4899)&(~g8822)&(~g11173));
assign g33231 = (g32032)|(g32036);
assign g8690 = (g2941&g2936);
assign II31267 = (g32840&g32841&g32842&g32843);
assign g28141 = (g10831&g11797&g11261&g27163);
assign g19542 = ((~g16349));
assign g30242 = (g28730&g23927);
assign II31724 = ((~g33076));
assign g21859 = (g3941&g21070);
assign g28421 = ((~g27074))|((~g13715));
assign g31230 = (g30285&g20751);
assign g17682 = (g9742&g14637);
assign g25770 = ((~g25417)&(~g25377));
assign g24037 = ((~g21127));
assign II31187 = (g32726&g32727&g32728&g32729);
assign II22380 = ((~g21156));
assign g9672 = ((~g5390));
assign g31320 = (g26125)|(g29632);
assign g21356 = ((~g15780))|((~g15752))|((~g15743))|((~g13118));
assign g27544 = (g26087)|(g24671);
assign g28439 = (g27273&g10233);
assign g23245 = ((~g20785));
assign gbuf124 = (g640);
assign g13969 = (g11448)|(g8913);
assign g16672 = (g6295&g15008);
assign g22858 = ((~g20751));
assign g13738 = (g8880&g10572);
assign g8238 = ((~II12469))|((~II12470));
assign g25448 = (g11202&g22680);
assign g29556 = ((~g28349))|((~g13486));
assign g34481 = (g34404&g18916);
assign g24267 = (g23439)|(g18611);
assign g14740 = ((~g5913))|((~g12129))|((~g6031))|((~g12614));
assign II17114 = ((~g14358));
assign II21922 = ((~g21335));
assign g32637 = ((~g30735));
assign g19369 = ((~g15995));
assign g22092 = (g6419&g18833);
assign g18409 = (g2084&g15373);
assign g34011 = (g33884)|(g18479);
assign g27408 = (g26519&g17523);
assign g19351 = ((~g17367));
assign II25907 = ((~g26256))|((~g24782));
assign g13638 = ((~II16057));
assign II29269 = ((~g29486))|((~g12050));
assign gbuf92 = (g4005);
assign g30239 = (g28728&g23923);
assign g33140 = ((~g7693)&(~g32072));
assign g18710 = (g15135&g17302);
assign II27543 = ((~g28187));
assign g32982 = (g31948)|(g18208);
assign g20779 = ((~g15509));
assign g28078 = (g27140)|(g21880);
assign g10675 = (g3436&g8500);
assign g31751 = (g29975)|(g29990);
assign g28359 = (g27151)|(g15838);
assign g19874 = ((~g13665))|((~g16299))|((~g8163));
assign II33173 = ((~g34887));
assign II12463 = ((~g4812));
assign g16533 = ((~II17733));
assign II11737 = ((~g4467));
assign g32744 = ((~g31327));
assign g29628 = (g27924&g28648);
assign g19535 = (g15651)|(g13020);
assign g23964 = ((~g19147));
assign II18865 = ((~g14314));
assign g9100 = ((~g3752)&(~g3712));
assign g20733 = ((~g14406))|((~g17290))|((~g9509));
assign II13078 = ((~g5462))|((~II13077));
assign g18160 = (g645&g17433);
assign g12078 = ((~g8187))|((~g8093));
assign g29791 = (g28233)|(g22859);
assign g7161 = ((~II11843));
assign g19699 = ((~II20116));
assign II12545 = ((~g191))|((~II12544));
assign II33041 = ((~g34772));
assign II22571 = ((~g20097));
assign g13134 = ((~g11134))|((~g8470));
assign II14896 = ((~g9820));
assign g17647 = ((~g5905))|((~g14497))|((~g5976))|((~g12614));
assign g22885 = ((~g9104))|((~g20154));
assign g27582 = ((~g10857))|((~g26131))|((~g26105));
assign g33806 = ((~II31650));
assign g9496 = ((~g3303));
assign g18773 = (g5694&g15615);
assign g21205 = ((~g15656));
assign g22588 = (g79&g20078);
assign g31814 = ((~g29385));
assign g24243 = (g22992)|(g18254);
assign g18515 = (g2643&g15509);
assign g30019 = ((~g29060));
assign g7002 = ((~g5160));
assign II24051 = (g3380&g3385&g8492);
assign g28552 = ((~g10295)&(~g27602));
assign g31975 = (g31761&g22177);
assign g14861 = ((~g12744))|((~g10341));
assign g29283 = (g28627)|(g18746);
assign g9369 = ((~g5084));
assign g25837 = ((~g25064));
assign g11707 = ((~g8718))|((~g4864));
assign g12108 = ((~II14964));
assign II20165 = ((~g16246))|((~g990));
assign II17324 = ((~g14119));
assign g11762 = ((~g7964));
assign g33115 = (g32397)|(g32401);
assign g23812 = ((~g18997));
assign g28069 = (g27564)|(g21865);
assign g11207 = ((~g3639)&(~g6905));
assign g18898 = ((~g15566));
assign II28540 = ((~g28954));
assign g27271 = (g24547)|(g26053);
assign g19560 = (g15832&g1157&g10893);
assign g22120 = (g6585&g19277);
assign g14234 = ((~g9177))|((~g11881));
assign II30971 = ((~g32015));
assign g11336 = ((~g7620));
assign g19476 = ((~g16326));
assign g18008 = ((~II18868));
assign g23499 = ((~g20785));
assign g34811 = (g14165&g34766);
assign g34436 = ((~II32479));
assign g31254 = (g25981)|(g29534);
assign g34762 = (g34687)|(g34524);
assign g33788 = (g33122)|(g32041);
assign g32370 = (g29882)|(g31312);
assign g29908 = ((~g6918)&(~g28471));
assign g32795 = ((~g31327));
assign g21819 = (g3614&g20924);
assign g24897 = (g3401&g23223&II24064);
assign II21074 = ((~g17766));
assign g24310 = (g4495&g22228);
assign g30030 = (g29198&g12347);
assign g17568 = ((~II18486))|((~II18487));
assign gbuf43 = (g6019);
assign g28598 = ((~g27717));
assign g19518 = ((~g16239));
assign g21946 = (g5252&g18997);
assign g8526 = ((~g1526));
assign g18506 = (g2571&g15509);
assign g34173 = (g33679&g24368);
assign g14817 = ((~g12711))|((~g12622));
assign g25983 = (g2476&g25009);
assign g13065 = ((~g10476));
assign g20436 = ((~II20569));
assign g20175 = ((~II20433));
assign g19277 = ((~II19813));
assign II12415 = ((~g48));
assign g24199 = (g355&g22722);
assign g34307 = ((~g34087));
assign g34693 = (g34513)|(g34310);
assign g16096 = ((~g13530));
assign g32008 = (g31781&g22223);
assign g24581 = (g5124&g23590);
assign g31993 = (g31774&g22214);
assign g34381 = (g34166&g20594);
assign II28434 = ((~g28114));
assign g8301 = ((~g1399));
assign g25699 = (g25125)|(g21918);
assign g27228 = (g26055&g16773);
assign g10415 = ((~g7109));
assign g32219 = (g31131)|(g29620);
assign II17436 = ((~g13416));
assign g32049 = (g10902&g30735);
assign g25010 = (g23267)|(g2932);
assign g7174 = ((~g6052));
assign g10420 = ((~g9239));
assign g26958 = (g26395)|(g24297);
assign g11216 = ((~g7998)&(~g8037));
assign g25086 = (g13941&g23488);
assign g29749 = (g28295&g23214);
assign g7423 = ((~g2433));
assign II14924 = ((~g9558))|((~II14923));
assign g12904 = ((~g10410));
assign g29270 = (g28258)|(g18635);
assign g10036 = ((~g1816));
assign g21180 = ((~g18008));
assign g16658 = ((~g14157));
assign g27973 = ((~g7187)&(~g25839));
assign g31671 = ((~II29262))|((~II29263));
assign g22929 = ((~g19773)&(~g12970));
assign g13033 = ((~g11917));
assign g28656 = ((~g27742));
assign g22645 = (g18982)|(g15633);
assign g34628 = (g34493)|(g18653);
assign g13835 = ((~II16150));
assign g33842 = (g33255&g20322);
assign g33164 = (g32203)|(II30727)|(II30728);
assign g28513 = (g27276)|(g26123);
assign II15647 = ((~g12109));
assign g12540 = ((~g2587)&(~g8381));
assign g32837 = ((~g31327));
assign g28281 = (g7362&g1936&g27440);
assign g34697 = ((~g34545));
assign g10147 = ((~g728));
assign g34399 = (g34178)|(g25067);
assign g22875 = ((~g20516))|((~g2980));
assign g10378 = ((~g6926));
assign II11743 = ((~g4564));
assign II15130 = ((~g2527))|((~II15128));
assign II27777 = ((~g29043));
assign g18788 = (g6031&g15634);
assign II16555 = ((~g10430));
assign g11537 = ((~g8229)&(~g3873));
assign g32425 = (g31668&g21604);
assign II13511 = ((~g2093))|((~II13509));
assign g30392 = (g30091)|(g18558);
assign g14082 = ((~g11697))|((~g11537));
assign II26367 = ((~g26400))|((~II26366));
assign g13008 = ((~g11855));
assign g24378 = (g3106&g22718);
assign g29736 = (g28522&g10233);
assign g31125 = (g29502&g22973);
assign g22754 = ((~g20114))|((~g19376));
assign g32108 = (g31631&g29913);
assign g18649 = (g4049&g17271);
assign g34363 = (g34148&g20389);
assign II21234 = ((~g16540));
assign g22848 = (g19449&g19649);
assign II22801 = ((~g21434))|((~II22799));
assign II13335 = ((~g1687))|((~II13334));
assign g9274 = ((~g5857));
assign g24386 = ((~g22594));
assign g18193 = (g837&g17821);
assign g18790 = (g6040&g15634);
assign g28678 = ((~g27800));
assign g16601 = ((~II17783));
assign g20920 = ((~g15426));
assign g27820 = (g7670&g25932);
assign g28349 = ((~g27074))|((~g24770))|((~g27187))|((~g19644));
assign g12932 = ((~II15550));
assign g12111 = ((~g847))|((~g9166));
assign g20185 = ((~g16772))|((~g13928))|((~g16723))|((~g13882));
assign g34758 = (g34683&g19657);
assign g33011 = (g32338)|(g18481);
assign g30058 = (g29180&g12950);
assign g24208 = (g23404)|(g18121);
assign g15711 = (g460&g13437);
assign g34993 = ((~II33279));
assign g26815 = (g4108&g24528);
assign g28600 = (g27339)|(g16427);
assign g28581 = (g27329)|(g26276);
assign II12437 = ((~g4999));
assign g10027 = ((~g6523));
assign g23443 = ((~g21468));
assign g29965 = ((~g28903));
assign g21433 = ((~g17792))|((~g14830))|((~g17765))|((~g14750));
assign II33218 = ((~g34955));
assign g26869 = ((~g24842));
assign II23372 = ((~g23361));
assign g15757 = (g3207&g14066);
assign g34808 = (g34765)|(g18599);
assign g29143 = (g27650)|(g17146);
assign g23301 = ((~g21037));
assign g30361 = (g30109)|(g18391);
assign g25289 = ((~g22228));
assign g14924 = ((~g12558))|((~g12505));
assign g9963 = ((~g7));
assign g33275 = (g32127)|(g29564);
assign g22650 = ((~g7888))|((~g19581));
assign g8944 = ((~g370));
assign g24782 = (g23857)|(g23872);
assign II32516 = ((~g34424))|((~g34422));
assign g14147 = ((~II16357));
assign g24841 = (g21420)|(g23998);
assign g22908 = ((~g9104))|((~g20175));
assign g26951 = (g26390)|(g24289);
assign g29872 = (g28401&g23333);
assign g25316 = ((~g22763));
assign II11620 = ((~g1));
assign g20901 = ((~II20867));
assign g14895 = ((~g7766))|((~g12571));
assign II12987 = ((~g12));
assign g24223 = (g239&g22594);
assign g17486 = ((~II18411));
assign g20508 = ((~g15277));
assign g20644 = ((~g14342))|((~g17220))|((~g9372));
assign II18740 = (g13156&g11450&g11498);
assign g20232 = ((~g16931));
assign g18259 = (g15068&g16000);
assign g34962 = (g34945&g23020);
assign g27958 = (g25950&g22449);
assign g27414 = (g255&g26827);
assign g18991 = ((~g16136));
assign g32924 = ((~g30937));
assign II11635 = ((~g9));
assign g26609 = ((~g146)&(~g24732));
assign g16198 = ((~g9247)&(~g13574));
assign g21012 = (g16304&g4688);
assign g14125 = ((~II16345));
assign g26976 = ((~g5016)&(~g25791));
assign g11956 = (g2070&g7411);
assign g34687 = (g14181&g34543);
assign g34714 = ((~II32874));
assign g14794 = ((~g12492))|((~g12772));
assign g19408 = ((~g16066));
assign II21486 = ((~g18727));
assign g13460 = ((~II15942));
assign II20819 = ((~g17088));
assign g7528 = ((~g930));
assign g25147 = (g20202&g23542);
assign g24999 = ((~g23626));
assign g25123 = (g4732&g22885);
assign g23182 = ((~g21389));
assign g32396 = (g4698&g30983);
assign g24475 = (g3831&g23139);
assign g13486 = ((~g10862))|((~g4983))|((~g4966));
assign g26019 = (g5507&g25032);
assign g12708 = ((~g9518)&(~g9462));
assign g29347 = (g29176&g22201);
assign g17663 = ((~g10205)&(~g12983));
assign g25124 = (g4917&g22908);
assign g7985 = ((~g3506));
assign g25215 = ((~II24384))|((~II24385));
assign g12186 = (g1178&g7519);
assign g33599 = (g33087)|(g18500);
assign g27540 = (g26576&g17746);
assign g24778 = ((~g23286));
assign g27288 = (g26515&g23013);
assign g33575 = (g33086)|(g18420);
assign g20234 = ((~g17140)&(~g14207));
assign g29563 = (g1616&g28853);
assign g22841 = ((~g20391));
assign g34526 = (g34300&g19569);
assign g17785 = (g13341&g10762);
assign g25388 = ((~g22763));
assign g30235 = (g28723&g23915);
assign g17531 = ((~II18476));
assign g8171 = ((~g3817));
assign g29685 = (g2084&g28711);
assign g33861 = (g33271&g20502);
assign g23129 = (g19500)|(g15863);
assign g25688 = (g24812)|(g21887);
assign g34417 = (g27678)|(g34196);
assign g21362 = ((~g17873));
assign g31767 = (g30031)|(g30043);
assign g11631 = ((~g8595));
assign g17148 = ((~g827)&(~g14279));
assign g15718 = ((~g13858)&(~g11330));
assign g9311 = ((~g5523));
assign g34635 = (g34485)|(g18692);
assign g14386 = ((~II16544));
assign g24431 = ((~g22722));
assign g28923 = ((~g27775))|((~g8195));
assign g22192 = ((~g19801));
assign II31016 = (g30825&g31798&g32478&g32479);
assign g24053 = ((~g21256));
assign g24406 = (g13623&g22860);
assign II32222 = ((~g34118));
assign g26232 = (g2193&g25396);
assign g20780 = ((~g15509));
assign g10319 = ((~II13740));
assign g8647 = ((~g3416));
assign g31818 = ((~g29385));
assign g27455 = (g26488&g17603);
assign II12112 = ((~g794));
assign g9536 = (g1351)|(g1312);
assign g27207 = (g26055&g16692);
assign g7549 = ((~g1018))|((~g1030));
assign g9818 = ((~g6490));
assign g33988 = (g33861)|(g18397);
assign g34105 = (g33778&g9104&g18957);
assign g11200 = ((~g8592))|((~g3798));
assign g31186 = (g2375&g30088);
assign g25555 = ((~g22550));
assign g21903 = ((~II21480));
assign g28661 = (g27406)|(g16611);
assign II32752 = ((~g34510));
assign II17405 = ((~g13378))|((~II17404));
assign g7442 = ((~g896))|((~g890));
assign g21405 = (g13377&g15811);
assign g14222 = (g8655&g11826);
assign g16024 = ((~g14216)&(~g11890));
assign II21199 = ((~g17501));
assign g28192 = (g8891&g27415);
assign g33828 = (g33090&g24411);
assign g23952 = ((~g19277));
assign g17769 = (g1146&g13188);
assign g23408 = ((~g21468));
assign g32125 = (g30918)|(g29376);
assign II16181 = ((~g3672));
assign g21998 = (g5712&g21562);
assign g17810 = (g1495&g13246);
assign g13026 = ((~g11018));
assign g25664 = (g24681)|(g21789);
assign g10754 = ((~g7936))|((~g7913))|((~g8411));
assign g9839 = ((~g2724));
assign g28073 = (g27097)|(g21875);
assign g11736 = ((~g8165));
assign g33830 = (g33382&g20166);
assign II22111 = ((~g19919));
assign g29316 = (g28528&g6875&g3288);
assign g24930 = (g4826&g23948);
assign II32881 = ((~g34688));
assign g7634 = ((~II12123));
assign g27661 = (g26576&g15568);
assign g29866 = (g1906&g29116);
assign g24913 = (g4821&g23908);
assign g15114 = (g4239&g14454);
assign g30478 = (g30248)|(g21949);
assign g24367 = ((~g22550));
assign g21850 = (g3893&g21070);
assign g19795 = ((~g13600))|((~g16275));
assign g25681 = (g24710)|(g18636);
assign g28816 = (g27547)|(g16843);
assign g30073 = (g1379&g28194);
assign g18356 = (g1802&g17955);
assign g17606 = ((~g14999));
assign g30326 = ((~II28579));
assign g32466 = ((~g31070));
assign g32777 = ((~g31710));
assign II20562 = ((~g16525));
assign g18368 = (g1728&g17955);
assign g26165 = (g11980&g25153);
assign II11896 = ((~g4446));
assign g28237 = (g9492&g27597);
assign g14182 = (g11741)|(g11721)|(g753);
assign g24763 = (g17569&g22457);
assign g31515 = ((~g4983)&(~g29556));
assign g23351 = ((~g20924));
assign g10741 = ((~g8411));
assign g32759 = ((~g31376));
assign g7178 = ((~g4392));
assign g28477 = (g27966&g17676);
assign g17586 = ((~g14638))|((~g14601));
assign g24730 = (g6177&g23699);
assign g17643 = (g9681&g14599);
assign g34805 = (g34748)|(g18594);
assign g34262 = (g34075)|(g18697);
assign g27303 = (g11996&g26681);
assign g16022 = (g13048)|(g10707);
assign g9832 = ((~g2399));
assign g32762 = ((~g31672));
assign g33463 = (g32477&II31011&II31012);
assign g21965 = (g15149&g21514);
assign g34039 = (g33743)|(g18736);
assign g33766 = ((~II31619));
assign g11029 = (g5782&g9103);
assign g31268 = (g29552)|(g28266);
assign g18613 = (g3338&g17200);
assign II15705 = ((~g12218));
assign II29182 = ((~g30012));
assign g17717 = ((~g14937));
assign g10154 = ((~g2547));
assign g32032 = (g31373&g16515);
assign g32546 = ((~g31170));
assign II24579 = (g5731&g5736&g9875);
assign g26120 = (g9809&g25293);
assign g32671 = ((~g31528));
assign g30105 = ((~II28336));
assign g9903 = ((~g681));
assign g21709 = (g283&g20283);
assign g27266 = (g26789&g26770);
assign g21468 = ((~II21181));
assign g34022 = (g33873)|(g18538);
assign g17722 = ((~II18709));
assign II26100 = ((~g26365));
assign II30980 = ((~g32132));
assign g24921 = (g23721&g20739);
assign II31282 = (g32863&g32864&g32865&g32866);
assign II12758 = ((~g4093));
assign g25227 = ((~g22763));
assign g23170 = ((~g20046));
assign g8086 = ((~g168)&(~g174)&(~g182));
assign g27937 = (g14506)|(g26793);
assign g18398 = (g2020&g15373);
assign g24522 = ((~g22689));
assign g27281 = (g9830&g26615);
assign g22077 = (g6263&g19210);
assign g32309 = (g5160&g31528);
assign g27683 = (g25770&g23567);
assign g8011 = ((~g3167));
assign g28110 = (g27974&g18886);
assign g28680 = (g27427)|(g16633);
assign g31770 = (g30034)|(g30047);
assign g25589 = (g21690)|(g24159);
assign g30460 = (g30207)|(g21931);
assign g16660 = ((~g3953))|((~g11225))|((~g3969))|((~g13933));
assign g14950 = ((~g7812))|((~g12632));
assign II27576 = ((~g28173));
assign g26158 = (g2255&g25432);
assign g9174 = ((~g1205));
assign g26855 = (g2960&g24535);
assign g21870 = (g4093&g19801);
assign g33482 = (g32614&II31106&II31107);
assign g11796 = ((~g7985));
assign g27105 = (g26026&g16511);
assign g18909 = (g16226&g13570);
assign g20853 = ((~g15595));
assign g26127 = (g2236&g25119);
assign g21665 = ((~II21226));
assign g12112 = ((~g8139))|((~g1624));
assign g26860 = ((~II25594));
assign g24342 = (g23691)|(g18772);
assign g7244 = ((~g4408));
assign g34663 = (g32028)|(g34500);
assign g9186 = ((~II13010));
assign g11190 = ((~g8539))|((~g3447));
assign g18745 = (g5128&g17847);
assign g13303 = ((~II15869));
assign g18493 = (g2514&g15426);
assign g11998 = ((~g8324))|((~g8373));
assign g11933 = ((~g837))|((~g9334))|((~g7197));
assign g11470 = ((~g7625));
assign g20715 = ((~g15277));
assign g25194 = ((~g22763));
assign g29118 = ((~g27886))|((~g9755));
assign g27345 = ((~g9360)&(~g26636));
assign II20650 = ((~g17010));
assign g9223 = ((~g1216));
assign g14018 = ((~g10323))|((~g11483));
assign g12785 = ((~g9472)&(~g6549));
assign g34259 = (g34066)|(g18679);
assign g10737 = ((~g6961))|((~g9848));
assign g29771 = (g28322&g23242);
assign g18187 = (g794&g17328);
assign g25603 = (g24698)|(g18114);
assign g19437 = ((~g16349));
assign g33610 = (g33242)|(g18616);
assign g27980 = (g26105)|(g26131);
assign g21387 = ((~II21115));
assign g25738 = (g25059)|(g22053);
assign g29565 = (g1932&g28590);
assign g21717 = (g15051&g21037);
assign g24187 = (g305&g22722);
assign g33900 = (g33316&g20913);
assign g21894 = (g20112)|(g15107);
assign g32489 = ((~g30614));
assign g30563 = (g29347)|(g22134);
assign g32814 = ((~g31021));
assign II12205 = ((~g1135))|((~II12203));
assign g13887 = (g5204&g12402);
assign g24119 = ((~g19935));
assign g8720 = ((~g358)&(~g365));
assign g25062 = ((~g21403))|((~g23363));
assign g34599 = (g34542)|(g18149);
assign g27535 = (g26519&g17737);
assign g24182 = ((~II23390));
assign g32842 = ((~g31710));
assign g28687 = (g27434)|(g16638);
assign g30525 = (g30266)|(g22071);
assign g34916 = ((~II33140));
assign g31491 = ((~g8938)&(~g29725));
assign g17737 = ((~g14810));
assign II12046 = ((~g613));
assign g21222 = ((~g17430));
assign g14205 = ((~g12381));
assign g8400 = ((~g4836));
assign g11194 = ((~g3288)&(~g6875));
assign II15915 = ((~g10430));
assign g25072 = ((~g23630));
assign g21411 = ((~g15426));
assign g32401 = (g31116&g13432);
assign g33677 = (g33443&g31937);
assign g32302 = (g31279&g23485);
assign II18555 = ((~g5630));
assign II17111 = ((~g13809));
assign g34281 = (g34043&g19276);
assign g30119 = ((~g28761)&(~g7315));
assign g18458 = (g2357&g15224);
assign g28498 = ((~g8172)&(~g27635));
assign g13346 = ((~g4854))|((~g11012));
assign g14752 = ((~g12540)&(~g10040));
assign g12852 = ((~g6847)&(~g10430));
assign g29776 = (g28225)|(g22846);
assign g28537 = (g6832&g27089);
assign g20768 = ((~g17955));
assign g10106 = ((~g16));
assign II14480 = ((~g10074))|((~g655));
assign g31210 = (g2509&g30100);
assign g10857 = ((~g8712));
assign g28259 = ((~g10504))|((~g26987))|((~g26973));
assign g33907 = (g23088&g33219&g9104);
assign g28607 = (g27342)|(g26303);
assign g29734 = (g28201)|(g15872);
assign g11411 = ((~g9713))|((~g3625));
assign g24804 = ((~g19916))|((~g23105));
assign g34008 = (g33849)|(g18476);
assign g12051 = ((~g9595));
assign g20433 = ((~g17929));
assign g16875 = ((~g3223))|((~g13765))|((~g3317))|((~g11519));
assign g17150 = (g8579&g12995);
assign g29756 = (g22717)|(g28223);
assign II26581 = ((~g26942));
assign g20919 = ((~g15224));
assign II22864 = ((~g12146))|((~g21228));
assign g32780 = ((~g31327)&(~II30330)&(~II30331));
assign g34518 = (g34292&g19503);
assign g13273 = ((~g1459))|((~g10699));
assign g29666 = (g28980&g22498);
assign g8967 = ((~g4264))|((~g4258));
assign g7512 = ((~g5283));
assign g27024 = (g26826)|(g17692);
assign g8631 = ((~g283));
assign g29601 = (g1890&g28955);
assign g24147 = ((~g19402));
assign II23986 = ((~g22182))|((~II23985));
assign g24444 = (g10890)|(g22400);
assign g14335 = ((~g12045)&(~g9283));
assign g20539 = ((~g15483));
assign g17128 = ((~II18180));
assign g14776 = ((~g12780))|((~g12622));
assign g28212 = (g27030)|(g27035);
assign g25832 = (g8219&g24625);
assign g21983 = (g5555&g19074);
assign g11971 = ((~g8249))|((~g8302));
assign g29164 = ((~g9444)&(~g28010));
assign g10501 = (g1233&g9007);
assign g22143 = (g19568&g10971);
assign g18596 = (g2941&g16349);
assign g24807 = ((~II23979))|((~II23980));
assign g32633 = ((~g31154));
assign g34331 = (g27121)|(g34072);
assign g17571 = ((~g8579))|((~g14367));
assign g20084 = (g11591&g16609);
assign g25819 = (g25323)|(g23836);
assign g18827 = ((~g16000));
assign g30253 = (g28746&g23943);
assign II29582 = ((~g30591));
assign g26783 = (g25037&g21048);
assign g34237 = (g32715)|(g33955);
assign g24233 = (g22590)|(g18236);
assign g8795 = ((~II12793));
assign II31878 = ((~g33696));
assign g18897 = ((~g15509));
assign g14317 = ((~g5033))|((~g11862));
assign g33403 = (g32352&g21396);
assign g31847 = ((~g29385));
assign g23610 = ((~g18833));
assign g20586 = ((~g15171));
assign g14011 = ((~g10295))|((~g11473));
assign g13976 = ((~g11130));
assign g7841 = ((~g904));
assign g34826 = (g34742)|(g34685);
assign g31001 = (g29360)|(g28151);
assign g23011 = ((~g20330));
assign g18570 = (g2848&g16349);
assign g19912 = ((~g17328));
assign g16583 = ((~g14069));
assign g18415 = (g2108&g15373);
assign II13851 = ((~g862))|((~II13850));
assign g11855 = ((~II14671));
assign g34233 = (g32455)|(g33951);
assign g6870 = ((~g3089));
assign g15578 = ((~g7216)&(~g14279));
assign g14673 = ((~II16770));
assign g11979 = ((~g9861))|((~g5452));
assign g29353 = ((~II27713));
assign g27504 = (g26519&g17680);
assign g14694 = ((~II16795));
assign g9920 = ((~g4322));
assign g10897 = ((~g7601));
assign g18558 = (g2803&g15277);
assign g23524 = ((~g21562));
assign g10061 = ((~II13581));
assign g7285 = ((~g4643));
assign g16612 = (g5603&g14927);
assign g34581 = (g22864&g34312);
assign II17276 = ((~g13605));
assign gbuf84 = (g3618);
assign II32782 = ((~g34571));
assign g11048 = ((~II14158));
assign g26814 = ((~g25221));
assign g28569 = (g27453&g20433);
assign g28982 = (g27163&g12687&g20682&II27349);
assign g33026 = (g32307)|(g21795);
assign g33426 = ((~g32017));
assign g14104 = ((~g11514))|((~g8864));
assign g23507 = ((~g21562));
assign g19592 = ((~II20035));
assign g15701 = (g3821&g13584);
assign g23012 = ((~g20330));
assign g30512 = (g30191)|(g22033);
assign g24276 = (g23083)|(g18646);
assign g33970 = (g33868)|(g18322);
assign g28199 = (g27479&g16684);
assign g22110 = (g15167&g19277);
assign II12608 = ((~g1582));
assign g14378 = ((~g11979))|((~g9731));
assign g7916 = ((~II12300));
assign g32700 = ((~g31579));
assign g25158 = ((~g22228));
assign g34410 = (g34204&g21427);
assign g16275 = ((~g9291))|((~g13480));
assign g22546 = ((~II21918));
assign g25098 = ((~g22369));
assign II13718 = ((~g890));
assign g13290 = (g3897&g11534);
assign g20379 = ((~g17821));
assign g27595 = (g26733&g26703);
assign g30004 = (g28521&g25837);
assign g10356 = ((~g6819));
assign g21836 = (g3805&g20453);
assign g33705 = ((~II31550));
assign g14503 = ((~g12256));
assign II31296 = (g30937&g31848&g32882&g32883);
assign g25775 = (g2922&g24568);
assign g31482 = ((~g8883)&(~g29697));
assign g18578 = (g2873&g16349);
assign g25753 = (g25165)|(g22100);
assign g9450 = ((~g5817));
assign g15065 = ((~g13394)&(~g12840));
assign II18667 = ((~g6661));
assign g11366 = (g5016&g10338);
assign II29139 = ((~g29382));
assign g30051 = (g28513&g20604);
assign g27246 = (g26690&g26673);
assign g11030 = ((~g8292));
assign g18797 = (g6173&g15348);
assign g15880 = (g3211&g13980);
assign g23389 = (g9072&g19757);
assign g8997 = ((~g577));
assign g34212 = (g33761&g22689);
assign g10970 = (g854&g9582);
assign II23671 = ((~g23202));
assign g18136 = (g550&g17249);
assign II20937 = ((~g16967));
assign g20210 = ((~g16897));
assign g24620 = ((~g22902))|((~g22874));
assign II18248 = ((~g12938));
assign II14258 = ((~g8154))|((~II14257));
assign g27039 = (g7738&g5527&g5535&g26223);
assign g34050 = (g33772&g22942);
assign g26055 = ((~II25115));
assign II33197 = ((~g34930));
assign II31022 = (g32487&g32488&g32489&g32490);
assign g23770 = (g20188)|(g16868);
assign g34075 = (g33692&g19517);
assign II17491 = ((~g13416));
assign g7661 = ((~g1211)&(~g1216)&(~g1221)&(~g1205));
assign g22591 = (g18893)|(g18909);
assign II18762 = (g13156&g6767&g11498);
assign II17475 = ((~g13336))|((~II17474));
assign g29807 = (g28359&g23272);
assign g14563 = ((~II16676));
assign g11543 = ((~g9714))|((~g3969));
assign II15765 = ((~g10823));
assign II12402 = ((~g3808))|((~II12401));
assign g30915 = (g29886&g24778);
assign g9194 = ((~g827));
assign g32579 = ((~g30735));
assign g12983 = ((~II15600));
assign g29234 = (g28415)|(g18239);
assign g32688 = ((~g30735));
assign g31871 = (g30596)|(g18279);
assign g10896 = (g1205&g8654);
assign II18114 = ((~g14509));
assign II21483 = ((~g18726));
assign g16804 = (g5905&g14813);
assign g33064 = (g31993)|(g22067);
assign g10386 = ((~g6982));
assign g31489 = (g2204&g30305);
assign g32709 = ((~g30735));
assign g14029 = ((~g11283));
assign g12346 = ((~g9931)&(~g9933));
assign g26097 = (g5821&g25092);
assign II32757 = ((~g34469))|((~II32756));
assign g25510 = (g6444&g22300&II24619);
assign g21343 = ((~g16428));
assign g21056 = ((~g15426));
assign g28935 = ((~g27800))|((~g2227))|((~g7328));
assign g16309 = ((~II17639));
assign g22176 = ((~g18997));
assign g32293 = (g2827&g30593);
assign g18906 = (g13568&g16264);
assign g20625 = ((~g15348));
assign g15874 = (g3893&g14079);
assign II17741 = (g14988&g11450&g11498);
assign g17511 = (g14396)|(g14365)|(g11976)|(II18452);
assign g30337 = (g29334)|(g18220);
assign g29130 = ((~g27907));
assign g24305 = (g4477&g22228);
assign g22065 = (g6203&g19210);
assign g31281 = (g30106&g27742);
assign g32178 = (g31747&g27886);
assign g10000 = ((~g6151));
assign g10960 = ((~g9007));
assign g28099 = (g27992)|(g22043);
assign II22830 = (g21429)|(g21338)|(g21307);
assign g11383 = ((~g9061));
assign g28230 = (g27669)|(g14261);
assign g14732 = ((~g12662))|((~g12515));
assign g18290 = (g1467&g16449);
assign g14674 = ((~g5941))|((~g12067))|((~g6023))|((~g12614));
assign g13947 = ((~g8948)&(~g11083));
assign g31942 = ((~g8977)&(~g30583));
assign g30604 = (g18911&g29878);
assign g19617 = ((~g16349));
assign g10776 = ((~II14033));
assign II18588 = ((~g2370))|((~II18587));
assign g24112 = ((~g19935));
assign g7598 = ((~II12075))|((~II12076));
assign g23570 = ((~g18833));
assign g16846 = (g14034&g12591&g11185);
assign g33007 = (g32331)|(g18455);
assign g11171 = ((~g8088)&(~g9226)&(~g9200)&(~g9091));
assign g11403 = ((~g7595));
assign g30448 = (g29809)|(g21857);
assign g7591 = ((~g6668));
assign g33818 = (g33236&g20113);
assign g16176 = (g14596&g11779);
assign g23656 = ((~II22800))|((~II22801));
assign g16472 = ((~g14098));
assign g12752 = ((~g9576)&(~g9529));
assign g21288 = ((~g14616))|((~g17492));
assign g33528 = (g32946&II31336&II31337);
assign g16076 = (g13081)|(g10736);
assign g30279 = (g28637)|(g27668);
assign g34168 = (g33787)|(g19784);
assign g16323 = ((~II17653));
assign g14600 = ((~g9564))|((~g12311));
assign g25183 = ((~g22763));
assign g14538 = ((~g11973)&(~g9828));
assign g7809 = ((~g4864));
assign g18748 = (g5142&g17847);
assign g19489 = ((~g16449));
assign g14031 = ((~II16289));
assign g19674 = (g2819&g15867);
assign II33067 = ((~g34812));
assign g25956 = ((~g1413)&(~g24609));
assign g22010 = (g5787&g21562);
assign g12998 = ((~g11829));
assign g21805 = (g3550&g20924);
assign g34328 = ((~g34096));
assign g15506 = ((~II17131));
assign g30008 = (g29191&g12297);
assign II33050 = ((~g34777));
assign II12848 = ((~g4281))|((~g4277));
assign g24812 = (g19662&g22192);
assign g25036 = ((~g23733));
assign g16261 = (g7898)|(g13469);
assign g34782 = (g34711&g33888);
assign g10626 = (g4057&g7927);
assign g24179 = ((~II23381));
assign g24669 = (g22653&g19742);
assign g34550 = ((~g626))|((~g34359))|((~g12323));
assign g22123 = (g6609&g19277);
assign g14364 = ((~g12083)&(~g9415));
assign g14708 = (g74&g12369);
assign g32267 = (g31208)|(g31218);
assign g19384 = (g667&g16310);
assign g24165 = ((~II23339));
assign g31935 = ((~g30583)&(~g4349));
assign g25007 = ((~g22457));
assign g8765 = ((~g3333));
assign g16619 = (g6629&g14947);
assign g21705 = (g209&g20283);
assign g27687 = ((~g25200))|((~g26714));
assign II17416 = ((~g13806));
assign g13324 = (g854&g11326);
assign g26264 = (g24688&g8812&g8778&g10627);
assign II31176 = (g31579&g31827&g32708&g32709);
assign g18975 = ((~g15938));
assign g27256 = (g25937&g19698);
assign g19695 = ((~g17015));
assign g32591 = ((~g30614));
assign g27558 = (g26576&g17776);
assign II32827 = ((~g34477));
assign g8542 = ((~II12644));
assign g26078 = (g5128&g25055);
assign g18761 = (g5471&g17929);
assign g9753 = ((~g1890));
assign g34719 = (g34701)|(g18133);
assign g32618 = ((~g31154));
assign g22635 = ((~g19801));
assign II18879 = ((~g13267));
assign g9690 = ((~g732));
assign g34600 = (g34538)|(g18182);
assign g20495 = ((~g17926));
assign g20551 = ((~g17302));
assign g30249 = ((~g5297)&(~g28982));
assign g29045 = ((~g27779));
assign g6988 = ((~g4765));
assign g30262 = ((~g5644)&(~g29008));
assign g20619 = ((~g14317))|((~g17217));
assign g18523 = (g2675&g15509);
assign g34618 = (g34527)|(g18580);
assign g33684 = (g33139&g13565);
assign g34392 = ((~g34202));
assign g33248 = (g32131&g19996);
assign g26848 = (g2950&g24526);
assign g12419 = ((~g9402)&(~g9326));
assign g12255 = ((~g9958))|((~g6140));
assign g10808 = ((~g8509)&(~g7611));
assign g25671 = (g24637)|(g21828);
assign g10079 = ((~g1950));
assign II11879 = ((~g4430))|((~II11877));
assign g30544 = (g30257)|(g22115);
assign g31147 = (g12286&g30054);
assign g11916 = (g2227&g7328);
assign g32668 = ((~g31070));
assign g34056 = ((~II31984))|((~II31985));
assign II22871 = ((~g12150))|((~g21228));
assign g29496 = (g28567)|(g27615);
assign g30166 = (g28621&g23792);
assign g14415 = ((~g12147)&(~g9590));
assign g22131 = (g6641&g19277);
assign g13564 = (g4480&g12820);
assign g23196 = ((~g20785));
assign g25135 = ((~g22457));
assign g24356 = ((~g22594));
assign g30269 = (g28778&g23970);
assign g32514 = ((~g30735));
assign g33505 = (g32779&II31221&II31222);
assign g28720 = (g27486)|(g16704);
assign g9269 = ((~g5517));
assign g21881 = (g4064&g19801);
assign II26584 = ((~g26943));
assign g24451 = (g3476&g23112);
assign g8666 = ((~g3703));
assign gbuf50 = (g6358);
assign II22729 = ((~g21308));
assign g12970 = ((~g10555)&(~g10510)&(~g10488));
assign II12654 = ((~g1585));
assign g26929 = (g26635)|(g18543);
assign g21656 = ((~g17700));
assign II14800 = ((~g10107));
assign g33436 = ((~II30962));
assign g26854 = (g2868&g24534);
assign g32198 = (g4253&g31327);
assign g34996 = ((~II33288));
assign g7939 = ((~g1280));
assign g20602 = (g10803&g15580);
assign g32920 = ((~g30825));
assign II22989 = ((~g21175));
assign g20673 = ((~g15277));
assign g26932 = (g26684)|(g18549);
assign g10136 = ((~g6113));
assign gbuf118 = (g4222);
assign g25000 = ((~g23630));
assign g18320 = (g1616&g17873);
assign g22105 = (g6494&g18833);
assign g13737 = (g4501&g10571);
assign g12925 = (g8928)|(g10511);
assign g26213 = (g25357&g11724&g7586&g7558);
assign g33318 = (g31969)|(g32434);
assign II22824 = ((~g21434))|((~II22822));
assign II13403 = ((~g2250))|((~II13401));
assign g22002 = (g5706&g21562);
assign g25366 = (g7733&g22406);
assign g21768 = (g3243&g20785);
assign II14789 = ((~g9891))|((~II14788));
assign g8102 = ((~g3072));
assign g33334 = (g32219&g20613);
assign g20034 = (g15902)|(g13299);
assign g9741 = ((~II13317));
assign g12306 = ((~g7394))|((~g5666));
assign II23354 = ((~g23277));
assign g34476 = (g34399&g18891);
assign g31167 = (g10080&g30076);
assign g29282 = (g28617)|(g18745);
assign g26919 = (g25951)|(g18267);
assign g30733 = (g13807)|(g29773);
assign g27214 = (g26026&g13901);
assign II12345 = ((~g3106))|((~II12344));
assign g25581 = (g19338&g24150);
assign g15033 = ((~g12806))|((~g7142));
assign II31066 = (g31070&g31807&g32550&g32551);
assign g33392 = (g32344&g21362);
assign g21889 = (g4169&g19801);
assign g28896 = ((~g27837))|((~g1936))|((~g1862));
assign g16736 = (g6303&g15036);
assign g16513 = (g8345&g13708);
assign g14665 = ((~g12604))|((~g12798));
assign g8364 = ((~g1585));
assign g12915 = ((~g12806))|((~g12632));
assign g15786 = (g13940&g11233);
assign g19964 = ((~g17200));
assign g28716 = (g27481)|(g13887);
assign g27516 = ((~g9180)&(~g26657));
assign g19070 = ((~g16957)&(~g11720));
assign g31243 = ((~g29933));
assign g25249 = ((~g22228));
assign g27363 = (g10231&g26812);
assign g32543 = ((~g31376));
assign g18243 = (g1189&g16431);
assign g9821 = ((~g115));
assign g7418 = ((~g2361));
assign g9883 = ((~g5782))|((~g5774));
assign g24951 = ((~g199))|((~g23088));
assign g12491 = ((~g7285))|((~g4462))|((~g6961));
assign g34107 = (g33710)|(g33121);
assign II31171 = (g31528&g31826&g32701&g32702);
assign g28695 = (g27580&g20666);
assign g25349 = ((~g22432))|((~g12051));
assign g28545 = (g27301)|(g26230);
assign g25856 = (g25518)|(g25510)|(g25488)|(g25462);
assign g13574 = ((~II16024));
assign g34572 = (g34387&g33326);
assign g24681 = (g16653&g22988);
assign g10123 = ((~g4294)&(~g4297));
assign g20011 = ((~g3731))|((~g16476));
assign g26514 = (g7400&g25564);
assign g16725 = ((~g13963));
assign g18141 = (g568&g17533);
assign g27099 = (g14094&g26352);
assign g13989 = ((~g8697)&(~g11309));
assign g24218 = (g872&g22594);
assign g28954 = ((~g27830));
assign II18117 = ((~g13302));
assign g32644 = ((~g30735));
assign g13661 = ((~g528)&(~g11185));
assign g16694 = ((~g3905))|((~g13772))|((~g3976))|((~g11631));
assign II19238 = ((~g15079));
assign g27115 = (g26026&g16526);
assign g24091 = ((~g20720));
assign g20322 = ((~g17873));
assign g25374 = (g5366&g23789&II24527);
assign g16810 = (g13461)|(g11032);
assign g14542 = ((~g3582))|((~g11238))|((~g3672))|((~g8542));
assign g16208 = (g3965&g14085);
assign g24920 = ((~II24089));
assign g10039 = ((~g2273));
assign g31310 = (g30157&g27886);
assign g19338 = ((~g16031)&(~g1306));
assign g27090 = (g25997&g16423);
assign g7601 = ((~g1322)&(~g1333));
assign gbuf74 = (g3274);
assign II13390 = ((~g1821))|((~g1825));
assign g28500 = ((~g590))|((~g27629))|((~g12323));
assign g9714 = ((~g4012));
assign II30962 = ((~g32021));
assign g18406 = (g2060&g15373);
assign II21294 = ((~g18274));
assign g30358 = (g30108)|(g18381);
assign g26100 = (g1677&g25097);
assign g12463 = ((~g7513))|((~g6322));
assign g15847 = (g3191&g14005);
assign g20556 = ((~g15483));
assign g23347 = ((~II22444));
assign g28267 = (g7328&g2227&g27421);
assign g26944 = (g26130)|(g18658);
assign g34140 = (g33931&g23802);
assign g20522 = (g691)|(g16893);
assign g33259 = (g32109)|(g29521);
assign g24219 = (g225&g22594);
assign II17606 = (g14988&g11450&g6756);
assign II29228 = ((~g30314));
assign g31654 = (g29325&g13062);
assign g24654 = (g11735&g22922);
assign g34554 = (g34347&g20495);
assign g30223 = (g28702&g23895);
assign II32391 = ((~g34153));
assign g34965 = (g34949&g23084);
assign g33438 = ((~g31950)&(~g4621));
assign g28131 = ((~g27051))|((~g25838));
assign g32726 = ((~g31672));
assign g13287 = (g1221&g11472);
assign g18239 = (g1135&g16326);
assign g16518 = (g5571&g14956);
assign II17679 = ((~g13416));
assign g13851 = ((~g8224))|((~g11360));
assign g30087 = ((~g29121));
assign g18983 = ((~g16077));
assign g34347 = (g25986)|(g34102);
assign g24984 = (g22929&g12818);
assign g25814 = (g24760&g13323);
assign g12476 = ((~g7498))|((~g6704));
assign II21792 = ((~g21308));
assign g8097 = ((~g3029));
assign g18218 = (g1008&g16100);
assign g20998 = ((~g18065)&(~g9450));
assign g23022 = ((~g20283));
assign g14767 = ((~g10130)&(~g12204));
assign g7779 = ((~g1413));
assign g28068 = (g27310)|(g21838);
assign II14563 = ((~g802));
assign g16926 = (g14061)|(g11804)|(g11780);
assign g19682 = ((~g17015));
assign g19778 = ((~g16268)&(~g1061));
assign g18661 = ((~II19487));
assign g12016 = ((~g1648))|((~g8093));
assign II14290 = ((~g8282))|((~II14289));
assign g18234 = (g1129&g16326);
assign g30140 = (g28600&g23749);
assign g11559 = ((~II14509))|((~II14510));
assign g19769 = ((~g16987));
assign g11213 = ((~g4776)&(~g7892)&(~g9030));
assign g16771 = ((~g14018));
assign g26866 = (g20204)|(g20242)|(g24363);
assign g34467 = (g34341)|(g18717);
assign g23197 = (g19571)|(g15966);
assign g17582 = ((~g14768));
assign g16812 = ((~g13555));
assign g28298 = ((~g10533))|((~g26131))|((~g26990));
assign g14614 = (g11975&g11997);
assign g28508 = ((~II26989));
assign g7802 = ((~g324));
assign g30074 = ((~g29046));
assign g11842 = ((~II14660));
assign g19487 = (g499&g16680);
assign g28301 = (g27224&g19750);
assign g18731 = (g15140&g16861);
assign II15194 = ((~g9935))|((~II15193));
assign g21453 = (g16713&g13625);
assign g24093 = ((~g20998));
assign g13797 = ((~g8102))|((~g11273));
assign g28597 = (g27515&g20508);
assign g17085 = ((~g14238));
assign g18316 = (g1564&g16931);
assign II24064 = (g3385&g3391&g8492);
assign g21986 = (g5575&g19074);
assign g26970 = (g26308)|(g24332);
assign g30029 = (g29164&g12936);
assign g22309 = (g1478&g19751);
assign g16893 = ((~g10685))|((~g13252))|((~g703));
assign g19345 = ((~g17591));
assign g24678 = ((~g22994))|((~g23010));
assign II22561 = ((~g20841));
assign g8241 = ((~g1792));
assign g8575 = ((~g291));
assign g24546 = (g22447&g19523);
assign g27007 = ((~g5706)&(~g25821));
assign g17616 = ((~g14309));
assign g8478 = ((~g3103));
assign g19555 = (g15672)|(g13030);
assign g18092 = ((~II18882));
assign II15987 = ((~g12381));
assign gbuf119 = (g4226);
assign g25550 = ((~g22763));
assign g15373 = ((~II17118));
assign g18115 = (g460&g17015);
assign g15852 = (g13820&g13223);
assign g23383 = (g19756)|(g16222);
assign g24139 = (g17619&g21653);
assign g25275 = ((~g22342))|((~g11991));
assign II15650 = ((~g12110));
assign g32658 = ((~g31579));
assign g8443 = ((~g3736));
assign g18152 = (g613&g17533);
assign g25282 = ((~g22763));
assign g9559 = ((~g6077));
assign g12662 = ((~g5863)&(~g9274));
assign g17058 = ((~II18148));
assign g8595 = ((~II12666));
assign g26308 = (g6961&g25289);
assign g30174 = (g28628&g23812);
assign g20169 = (g16184)|(g13460);
assign g18171 = (g728&g17433);
assign g30480 = (g29321)|(g21972);
assign g27389 = (g26519&g17503);
assign II14663 = ((~g9747));
assign g11702 = ((~g6928));
assign g26256 = ((~g23873)&(~g25479));
assign g25820 = ((~g25051));
assign g30232 = (g28719&g23912);
assign g21281 = ((~g16286));
assign II15243 = ((~g6351))|((~II15241));
assign g32887 = ((~g30614));
assign g15785 = (g3558&g14107);
assign g34679 = (g14093&g34539);
assign g27269 = (g25943&g19734);
assign g20911 = ((~g15171));
assign g23684 = ((~II22819));
assign g29291 = (g28660)|(g18767);
assign g29528 = (g2429&g28874);
assign g18418 = (g2122&g15373);
assign g30342 = (g29330)|(g18261);
assign gbuf33 = (g5677);
assign g14055 = ((~g11697))|((~g11763));
assign g13061 = ((~g10981));
assign g20136 = ((~II20399));
assign g32222 = (g31141)|(g29636);
assign g32446 = ((~g31596));
assign g21175 = ((~II20951));
assign g34644 = (g34555)|(g18769);
assign g19661 = (g5489&g16969);
assign g15084 = (g2710&g12983);
assign g12099 = (g9619&g9888);
assign g34879 = ((~II33109));
assign g18270 = (g1291&g16031);
assign g27881 = ((~II26430));
assign II13149 = ((~g6745));
assign II17494 = ((~g13378))|((~g1448));
assign g16642 = (g6633&g14981);
assign g33541 = (g33101)|(g18223);
assign II21036 = ((~g17221));
assign g27018 = ((~II25750));
assign g11721 = ((~g10074));
assign g23883 = ((~g2779)&(~g21067));
assign g34149 = (g33760)|(g19674);
assign g25209 = ((~g22763));
assign g6809 = ((~g341));
assign g24642 = (g8290&g22898);
assign II32089 = ((~g33665));
assign g24777 = (g11345&g23066);
assign g15830 = ((~g13432));
assign g20777 = ((~g15224));
assign gbuf17 = (g5320);
assign g8784 = ((~II12764));
assign g23761 = ((~II22893))|((~II22894));
assign g12833 = ((~II15448));
assign g23429 = ((~g20453));
assign g32232 = (g31241&g20266);
assign g10725 = ((~g7846));
assign g13118 = ((~g5897))|((~g12067))|((~g6031))|((~g9935));
assign g30168 = (g28623&g23794);
assign g33305 = (g31935&g17811);
assign g25692 = ((~II24839));
assign g30364 = (g30086)|(g18411);
assign g29538 = (g2563&g28914);
assign g8803 = ((~g128))|((~g4646));
assign g34897 = (g34861)|(g21682);
assign g29072 = ((~g9402)&(~g26977));
assign II14967 = ((~g9964));
assign g22407 = ((~g19455));
assign g27046 = ((~g7544)&(~g25888));
assign g29924 = (g13031&g29190);
assign g25608 = (g24643)|(g18120);
assign g10583 = ((~g7475))|((~g862));
assign g23875 = ((~g18997));
assign g16282 = ((~g4933))|((~g13939))|((~g12088));
assign II32482 = ((~g34304));
assign g29597 = ((~g28444));
assign g26800 = (g24922)|(g24929);
assign g18496 = (g2537&g15426);
assign g25432 = ((~g12374))|((~g22384));
assign g19602 = ((~g16349));
assign g29522 = (g28923&g22369);
assign g34755 = ((~II32929));
assign g25599 = (g24914)|(g21721);
assign g19470 = ((~g16000));
assign g8249 = ((~g1917));
assign g30576 = (g18898&g29800);
assign g17320 = ((~II18297));
assign g11890 = (g7499&g9155);
assign g20610 = ((~g18008));
assign II12083 = ((~g568));
assign g34340 = (g34100&g19950);
assign g29206 = (g24124&II27528&II27529);
assign g8712 = ((~II12712));
assign g34143 = (g33934&g23828);
assign g17301 = ((~g14454));
assign g24315 = (g4521&g22228);
assign g27015 = ((~g26869));
assign g27154 = (g26055&g16630);
assign g12440 = ((~g9985));
assign g18385 = (g1959&g15171);
assign g32528 = ((~g31554));
assign g23992 = ((~g19210));
assign g8477 = ((~g3061));
assign g16652 = ((~g13892));
assign g20658 = (g1389&g15800);
assign II21934 = ((~g21273));
assign g8046 = ((~g528));
assign g12412 = ((~g10044))|((~g5297))|((~g5348));
assign g24698 = (g22664&g19761);
assign g34503 = (g34278&g19437);
assign g12146 = ((~g1783)&(~g8241));
assign g28640 = (g27384)|(g16590);
assign g29581 = (g28462&g11796);
assign g20567 = ((~g15426));
assign II14326 = ((~g8607));
assign g10183 = ((~g2595));
assign g11370 = (g8807)|(g550);
assign g29266 = (g28330)|(g18621);
assign g27360 = (g26488&g17417);
assign g15158 = ((~g13782)&(~g12901));
assign g22987 = ((~g20391));
assign g13014 = ((~g11872));
assign g23602 = ((~g9672)&(~g20979));
assign g14654 = (g7178&g10476);
assign g17710 = ((~g14764));
assign g19678 = ((~g16752));
assign g12729 = ((~g1657)&(~g8139));
assign g12101 = ((~g6336)&(~g7074));
assign g16868 = (g5813&g14297);
assign g26943 = ((~II25695));
assign g7395 = ((~g6005));
assign g25950 = ((~g1070)&(~g24591));
assign II33079 = ((~g34809));
assign g22008 = (g5774&g21562);
assign g11692 = ((~g8021)&(~g7985));
assign g20063 = (g15978)|(g13313);
assign g30930 = (g29915&g23342);
assign g22715 = ((~g20114))|((~g2999));
assign g31893 = (g31490)|(g21837);
assign g10715 = ((~g8526)&(~g8466));
assign g31749 = (g29974)|(g29988);
assign g25143 = (g4922&g22908);
assign g23715 = ((~g20764));
assign g21731 = (g3029&g20330);
assign g12245 = ((~g7344))|((~g5637));
assign g31828 = ((~g29385));
assign g17590 = ((~II18523));
assign g13763 = ((~g10971));
assign g18279 = (g1361&g16136);
assign g25439 = ((~g22498))|((~g12122));
assign g13377 = ((~g7873)&(~g10762));
assign II31848 = (g33479)|(g33480)|(g33481)|(g33482);
assign g34218 = (g33744&g22670);
assign g33581 = (g33333)|(g18443);
assign II27528 = (g20998&g24118&g24119&g24120);
assign g18708 = (g4818&g16782);
assign g7750 = ((~g1070));
assign g17758 = ((~g14861));
assign g23768 = ((~g18997));
assign g16289 = ((~g13223));
assign g34030 = (g33727)|(g18704);
assign g13876 = ((~g11432));
assign g23920 = (g4135&g19549);
assign g8165 = ((~g3530));
assign g18327 = (g1636&g17873);
assign g13525 = (g10019&g11911);
assign g14876 = ((~g12492))|((~g12443));
assign g13980 = ((~g10295))|((~g11435));
assign g22033 = (g5925&g19147);
assign g28555 = (g27429&g20373);
assign g18580 = (g2907&g16349);
assign g32189 = (g30824&g25369);
assign g28336 = ((~g27064))|((~g24756))|((~g27163))|((~g19644));
assign g17642 = ((~g14691));
assign g10072 = ((~g9));
assign g11995 = ((~g9645)&(~g7410));
assign g25990 = (g9461&g25017);
assign g10498 = ((~g7161));
assign g28705 = (g27460)|(g16672);
assign g6789 = ((~II11635));
assign g26683 = ((~g25514));
assign g31132 = (g29504&g22987);
assign g29502 = (g28139)|(g25871);
assign g33350 = (g32235&g20702);
assign II27495 = ((~g27961));
assign g14810 = ((~g12700))|((~g10312));
assign g12632 = ((~g9631)&(~g6565));
assign g24463 = ((~g23578));
assign g23264 = ((~g21037));
assign g10619 = (g3080&g7907);
assign II18360 = ((~g1426));
assign II24685 = (g24036&g24037&g24038&g24039);
assign g31475 = (g29756&g23406);
assign g32682 = ((~g30825));
assign g12292 = ((~g4698))|((~g8933));
assign g25768 = (g2912&g24560);
assign g11965 = ((~II14797));
assign II14169 = ((~g8389))|((~g3119));
assign g22022 = (g5873&g19147);
assign g12223 = ((~g2051)&(~g8365));
assign g17365 = (g7650&g13036);
assign g32962 = ((~g30735));
assign g26364 = ((~II25327));
assign g11714 = ((~g8107));
assign g28746 = (g27520)|(g16762);
assign g15938 = ((~II17401));
assign g22165 = (g15594&g18903);
assign II31332 = (g32935&g32936&g32937&g32938);
assign g32376 = (g2689&g31710);
assign g33916 = ((~II31776));
assign g34650 = ((~II32757))|((~II32758));
assign g18224 = (g1036&g16100);
assign g18524 = (g2681&g15509);
assign g33363 = (g32262&g20918);
assign g25157 = ((~g22498));
assign g20128 = ((~g17533));
assign g15480 = ((~II17125));
assign g23422 = ((~g21611));
assign g28080 = ((~II26581));
assign g28701 = (g27455)|(g16669);
assign g24959 = ((~g8858)&(~g23324));
assign g28273 = (g27927&g23729);
assign g27323 = (g26268&g23086);
assign g8719 = ((~II12719));
assign g26961 = (g26280)|(g24306);
assign g32956 = ((~g30825));
assign g32535 = ((~g31554));
assign g22070 = (g6243&g19210);
assign g33071 = (g31591&g32404);
assign g16749 = ((~g3957))|((~g13772))|((~g4027))|((~g11631));
assign g19571 = (g3498&g16812);
assign g24106 = ((~g19984));
assign g23956 = ((~g18957)&(~g18918)&(~g20136)&(~g20114));
assign g25978 = (g9391&g25001);
assign g21775 = (g3372&g20391);
assign g20100 = ((~II20369));
assign g29604 = (g2315&g28966);
assign II20870 = ((~g16216));
assign II31261 = (g30937&g31842&g32831&g32832);
assign II18709 = ((~g6668));
assign g25745 = (g25150)|(g22060);
assign g14713 = ((~g12483)&(~g9974));
assign g7785 = ((~g4621));
assign g28081 = ((~II26584));
assign g18755 = (g5343&g15595);
assign g27235 = (g25910&g19579);
assign g18158 = (g667&g17433);
assign g31950 = ((~g7285))|((~g30573));
assign g18120 = (g457&g17015);
assign g18475 = (g12853&g15426);
assign g34449 = (g34279)|(g18662);
assign II17925 = ((~g1478))|((~II17923));
assign g32690 = ((~g31070));
assign g22472 = (g7753&g9285&g21289);
assign g9155 = ((~II12997));
assign g22939 = (g9708&g21062);
assign g7685 = (g4382&g4375);
assign g12054 = ((~g7690));
assign g12952 = ((~II15572));
assign g18876 = ((~g15373));
assign g23377 = ((~g21070));
assign g28036 = ((~g26365));
assign g21826 = (g3742&g20453);
assign g32158 = (g31658&g30022);
assign g25140 = ((~g22228));
assign g25092 = ((~g23666));
assign g23417 = ((~g20391));
assign II31868 = (g33515)|(g33516)|(g33517)|(g33518);
assign g14714 = ((~g11405));
assign g15851 = (g3953&g14157);
assign gbuf65 = (g6711);
assign g14202 = (g869&g10632);
assign g28305 = (g27103)|(g15793);
assign g27571 = (g26127)|(g24723);
assign g18552 = (g2815&g15277);
assign g11409 = ((~g9842))|((~g3298));
assign g33922 = (g33448&g7202);
assign g8350 = ((~g4646));
assign g20785 = ((~II20846));
assign g8659 = ((~g2815));
assign g20389 = ((~g15277));
assign g24176 = ((~II23372));
assign II23163 = (g20982)|(g21127)|(g21193)|(g21256);
assign II22718 = ((~g11916))|((~II22717));
assign g30204 = (g28670&g23868);
assign g21605 = (g13005&g15695);
assign g7470 = ((~g5623));
assign g10939 = ((~g7352))|((~g1459));
assign g13473 = (g9797&g11841);
assign g18213 = (g952&g15979);
assign II20781 = ((~g17155));
assign g6888 = ((~II11701));
assign g18480 = (g2437&g15426);
assign II12541 = ((~g194));
assign g14425 = ((~g5644)&(~g12656));
assign II31853 = (g33488)|(g33489)|(g33490)|(g33491);
assign g27615 = (g26789&g26770);
assign g23698 = ((~g21611));
assign g30120 = (g28576&g21051);
assign g24328 = (g4567&g22228);
assign g11928 = ((~II14742));
assign g12459 = ((~g7437))|((~g5623));
assign g34875 = (g34836&g20073);
assign g23112 = ((~g21024))|((~g10733));
assign g28203 = ((~g12546))|((~g27985))|((~g27977));
assign g29008 = (g27163&g12730&g20739&II27364);
assign g27467 = (g269&g26832);
assign g13665 = ((~g11306));
assign g20904 = ((~g17433));
assign g29784 = (g28331&g23247);
assign g31272 = (g30117&g27742);
assign g30109 = (g28562&g20912);
assign g34657 = (g33114)|(g34497);
assign g19146 = ((~g15574));
assign g27593 = ((~g24972))|((~g24950))|((~g24906))|((~g26861));
assign g25274 = ((~g22763));
assign g15568 = ((~g14984));
assign g13495 = ((~g1008))|((~g11786))|((~g7972));
assign g12524 = ((~g7074))|((~g7087))|((~g10212));
assign g20638 = ((~g15224));
assign gbuf26 = (g5659);
assign g29660 = ((~g28448))|((~g9582));
assign g21339 = ((~g15725))|((~g13084))|((~g15713))|((~g13050));
assign g34157 = (g33794&g20159);
assign g19730 = ((~g17062));
assign g16956 = ((~g3925))|((~g13824))|((~g4019))|((~g11631));
assign II18579 = ((~g1945))|((~g14678));
assign g14253 = ((~g10032)&(~g12259)&(~g9217));
assign g23214 = ((~g20785));
assign g13139 = ((~g6589))|((~g12137))|((~g6723))|((~g10061));
assign g10519 = ((~g9326));
assign g32564 = ((~g31376));
assign g31864 = (g31271)|(g21703);
assign g18950 = (g11193&g16123);
assign g34466 = (g34337)|(g18716);
assign g29313 = (g28284)|(g27270);
assign II12483 = ((~g3096));
assign II31252 = (g32819&g32820&g32821&g32822);
assign g29952 = (g23576&g28939);
assign g31509 = ((~g599))|((~g29933))|((~g12323));
assign g28734 = (g27508)|(g16736);
assign g18469 = (g2399&g15224);
assign g34015 = (g33858)|(g18502);
assign g15567 = (g392&g13312);
assign g24623 = ((~g23076));
assign g13175 = ((~g10909));
assign g15133 = ((~g12883)&(~g13638));
assign g25485 = (g6098&g22220&II24600);
assign g19749 = (g732&g16646);
assign g16183 = ((~g9223)&(~g13545));
assign II24363 = ((~g23687))|((~g14320));
assign g25423 = ((~II24558));
assign g29571 = (g28452&g11762);
assign g27295 = ((~g24776))|((~g26208));
assign g15742 = ((~g5575))|((~g12093))|((~g5637))|((~g14669));
assign g15727 = (g13383)|(g13345)|(g13333)|(g11010);
assign g30982 = (g8895&g29933);
assign g14185 = (g8686&g11744);
assign g28571 = (g27458&g20435);
assign g18282 = (g1379&g16136);
assign g27392 = (g26576&g17507);
assign g14291 = ((~g9839)&(~g12155));
assign g23272 = ((~g20924));
assign g13011 = ((~II15623));
assign g27028 = (g26342&g1157);
assign II14991 = ((~g9685))|((~g6527));
assign g33419 = ((~g31978)&(~g7627));
assign g27439 = (g232&g26831);
assign g18880 = ((~g15656));
assign II25243 = ((~g490))|((~II25242));
assign g18652 = (g4172&g16249);
assign II13454 = ((~g1959))|((~II13452));
assign II32651 = ((~g34375));
assign g30407 = (g29794)|(g21766);
assign g23485 = ((~g20785));
assign g29550 = (g28990&g22457);
assign g30283 = (g28851&g23993);
assign g30187 = (g28643&g23840);
assign g10003 = ((~II13539));
assign g24926 = ((~g20172))|((~g20163))|((~g23357))|((~g13995));
assign g34830 = ((~II33044));
assign g14120 = ((~g11780))|((~g4907));
assign g26693 = ((~g25300));
assign g32861 = ((~g31376));
assign II12096 = ((~g1339))|((~g1322));
assign g19654 = ((~g16931));
assign g8859 = ((~g772));
assign g22994 = ((~g20436));
assign g17153 = (g6311&g14943);
assign g24286 = (g4405&g22550);
assign g24062 = ((~g19968));
assign g31219 = (g30265&g20875);
assign g33944 = ((~II31829));
assign g12937 = ((~g12419));
assign g11385 = ((~g8021)&(~g7985));
assign g27314 = (g12436&g26702);
assign g28970 = (g17405&g25196&g26424&g27445);
assign g31794 = ((~II29368));
assign g33458 = ((~II30992));
assign g14433 = ((~g12035))|((~g9890));
assign g23105 = ((~g8097))|((~g19887));
assign g29148 = (g27651)|(g26606);
assign g24609 = ((~g22850))|((~g22650));
assign g25265 = ((~II24455));
assign g15048 = ((~II16969));
assign g8737 = ((~II12729))|((~II12730));
assign g15077 = (g2138&g12955);
assign g9300 = ((~g5180));
assign g24253 = (g22525)|(g18300);
assign II12172 = ((~g2715));
assign g33389 = (g32272)|(g29964);
assign g18648 = (g4045&g17271);
assign II25351 = ((~g24466));
assign g23970 = ((~g19277));
assign g25577 = (g24143)|(g24144);
assign g31250 = (g25972)|(g29526);
assign g17715 = ((~II18700));
assign g31817 = ((~g29385));
assign g26840 = ((~II25562));
assign g19375 = ((~II19863));
assign g32846 = ((~g31376));
assign II22793 = ((~g11956))|((~II22792));
assign g10274 = ((~g976));
assign g28065 = (g27299)|(g21792);
assign g25730 = (g25107)|(g22013);
assign g27927 = ((~g9621)&(~g25856));
assign g24144 = (g17727&g21660);
assign g24173 = ((~II23363));
assign g24365 = ((~g22594));
assign g24842 = (g7804)|(g22669);
assign g32785 = ((~g31710));
assign g22896 = ((~g21012));
assign g33841 = (g33254&g20268);
assign g18206 = (g918&g15938);
assign g7540 = ((~II12026));
assign g10657 = (g8451&g4064);
assign g30442 = (g29797)|(g21851);
assign g34323 = ((~g34105));
assign g6973 = ((~II11743));
assign g30132 = ((~g28789)&(~g7362));
assign II32204 = ((~g33670))|((~II32202));
assign g26209 = ((~g23124)&(~g24779));
assign g34453 = (g34410)|(g18666);
assign g13554 = ((~g11336))|((~g7582))|((~g1351));
assign g32525 = ((~g31170));
assign II11809 = ((~g6741));
assign g24559 = (g22993&g19567);
assign g34299 = ((~g34080));
assign g18435 = (g2173&g18008);
assign g17221 = ((~II18245));
assign g7184 = ((~g5706))|((~g5752));
assign g8583 = (g2917&g2912);
assign g24041 = ((~g19968));
assign g28098 = (g27683)|(g22016);
assign g24388 = ((~g22885));
assign g12289 = ((~g9978))|((~g9766))|((~g9708));
assign g24605 = ((~g23139));
assign g24497 = ((~g23533)&(~g23553));
assign g28137 = ((~II26638));
assign g25216 = ((~g6088))|((~g23678));
assign g19529 = ((~g16349));
assign II17302 = ((~g14044));
assign g26731 = ((~g25470));
assign g32807 = ((~g31021));
assign g29253 = (g28697)|(g18490);
assign g18264 = (g1263&g16000);
assign II21058 = ((~g17747));
assign g31907 = (g31492)|(g21954);
assign g12252 = ((~g9995)&(~g10185));
assign g29305 = (g28602)|(g18811);
assign II16117 = ((~g10430));
assign g22041 = (g5957&g19147);
assign g18361 = (g1821&g17955);
assign g19451 = ((~g15938));
assign g14965 = ((~g12609))|((~g12571));
assign g26877 = (g21658)|(g25577);
assign g28171 = (g27016&g19385);
assign g11320 = ((~g4633))|((~g4621))|((~g7202));
assign g23871 = ((~g2811)&(~g21348));
assign g16488 = ((~g13697)&(~g13656));
assign g33410 = (g32360&g21409);
assign g24552 = (g22487&g19538);
assign g17593 = ((~II18537))|((~II18538));
assign g29082 = ((~g27837))|((~g9694));
assign g14130 = ((~g11621))|((~g8906));
assign II17008 = ((~g12857));
assign g33326 = ((~g32318));
assign II13452 = ((~g1955))|((~g1959));
assign g32284 = (g31260&g20507);
assign g9698 = ((~g2181));
assign II21013 = ((~g15806));
assign g29260 = (g28315)|(g18604);
assign g20269 = ((~g15844));
assign g33304 = (g32427&g31971);
assign g27527 = ((~II26195));
assign g25721 = (g25057)|(g18766);
assign g14038 = ((~g11514))|((~g11435));
assign g23788 = ((~g18997));
assign g33096 = ((~g31997)&(~g4608));
assign g15672 = (g433&g13458);
assign g23284 = ((~g20785));
assign II31052 = (g32531&g32532&g32533&g32534);
assign II32675 = ((~g34427));
assign II26664 = ((~g27708));
assign g9407 = ((~g6549));
assign II32982 = ((~g34749));
assign g26576 = ((~II25399));
assign II28062 = ((~g29194));
assign II12056 = ((~g2748));
assign g26260 = ((~g24759));
assign g20732 = ((~g15595));
assign g28990 = ((~g27882))|((~g8310));
assign g10799 = ((~g347)&(~g7541));
assign g23413 = ((~g21012));
assign II32812 = ((~g34588));
assign g20195 = ((~g16931));
assign g25611 = (g24931)|(g18128);
assign II13110 = ((~g5808))|((~II13109));
assign II30399 = (g29385)|(g31376)|(g30735)|(g30825);
assign g14781 = ((~g6259))|((~g12173))|((~g6377))|((~g12672));
assign g34114 = (g33920&g23742);
assign g18679 = (g4633&g15758);
assign g23978 = ((~g572))|((~g21389))|((~g12323));
assign g25949 = (g24701&g19559);
assign g18441 = (g2246&g18008);
assign g29992 = (g29012&g10490);
assign g20766 = ((~g17433));
assign g25676 = (g24668)|(g21833);
assign g26178 = (g2389&g25473);
assign g23238 = ((~g20924));
assign II13597 = ((~g4417));
assign g24747 = (g17510&g22417);
assign g22851 = (g496&g19654);
assign II15623 = ((~g12040));
assign g20172 = ((~g16876))|((~g8131));
assign II18370 = ((~g14873));
assign g12975 = ((~g12752));
assign g28224 = (g27163&g22763&g27064);
assign g32476 = ((~g30673));
assign g23945 = ((~g21611));
assign g28907 = ((~g27858))|((~g2361))|((~g2287));
assign g30193 = (g28650&g23848);
assign g29709 = (g2116&g29121);
assign II16676 = ((~g10588));
assign g23567 = ((~g21562));
assign g12369 = ((~g9049))|((~g637));
assign g12861 = ((~g10367));
assign g12428 = ((~g7472))|((~g6358));
assign g32290 = (g31267&g20525);
assign g28652 = (g27282&g10288);
assign g26832 = ((~g24850));
assign g10980 = ((~g9051));
assign g19793 = ((~g16292)&(~g1404));
assign g24478 = (g11003)|(g22450);
assign g20088 = ((~g17533));
assign II29245 = ((~g29491));
assign g16763 = (g6239&g14937);
assign g10169 = ((~g6395));
assign g23135 = ((~g16476)&(~g19981));
assign g8416 = ((~II12580));
assign g31876 = (g31125)|(g21731);
assign II12850 = ((~g4277))|((~II12848));
assign g33967 = (g33842)|(g18319);
assign g28966 = ((~g27858))|((~g2361))|((~g7380));
assign g8451 = ((~g4057));
assign g18744 = (g5124&g17847);
assign g20857 = ((~g17929)&(~g9380));
assign g13190 = ((~g10939));
assign g16209 = ((~g13478)&(~g4749));
assign g34065 = (g33813&g23148);
assign g22200 = ((~g19277));
assign II30760 = (g31778)|(g32295)|(g32046)|(g32050);
assign g6904 = ((~g3494));
assign g30322 = ((~g28431));
assign g16720 = ((~g14234));
assign g34137 = (g33928&g23802);
assign g30022 = ((~g29001));
assign g9284 = ((~g2161));
assign g21797 = (g3518&g20924);
assign g15631 = (g168&g13437);
assign g19658 = ((~g16987));
assign g30488 = (g30197)|(g21984);
assign g12589 = ((~g7591))|((~g6692));
assign g26702 = ((~g25309));
assign II20864 = ((~g16960));
assign II16417 = ((~g875));
assign g30238 = (g28727&g23922);
assign g27779 = (g17317)|(g26694);
assign g25537 = ((~g22763))|((~g2873));
assign g30055 = ((~g29157));
assign II26710 = ((~g27511));
assign II14761 = ((~g7753));
assign II12793 = ((~g4578));
assign g26712 = (g24508&g24463);
assign II14531 = ((~g8840))|((~II14530));
assign g15017 = (g10776)|(g8703);
assign g31775 = (g30048)|(g30059);
assign g10658 = ((~II13979));
assign g23989 = (g20581)|(g17179);
assign gbuf150 = (g1233);
assign II13990 = ((~g7636));
assign II14970 = ((~g9965));
assign g19753 = ((~g16987));
assign g20542 = ((~g17873));
assign g22300 = ((~II21815));
assign g32947 = ((~g31376));
assign g10397 = ((~g7018));
assign g17734 = ((~g5272))|((~g14490))|((~g5283))|((~g9780));
assign g31153 = (g12336&g30068);
assign g7239 = ((~g5033));
assign g34533 = (g34318&g19731);
assign g10219 = ((~g2697));
assign II16969 = ((~g13943));
assign g18674 = (g4340&g15758);
assign g30428 = (g29807)|(g21812);
assign g33836 = (g33096&g27020);
assign g22983 = ((~g979)&(~g16268)&(~g19853));
assign II14619 = ((~g4185));
assign g8514 = ((~g4258));
assign g32245 = (g31167)|(g29684);
assign g34530 = ((~II32591));
assign g24561 = (II23755)|(II23756);
assign g28778 = (g27540)|(g16808);
assign g24392 = (g3115&g23067);
assign g27454 = (g26488&g17602);
assign II25190 = ((~g25423));
assign II18310 = ((~g12978));
assign g19681 = (g5835&g17014);
assign g33596 = (g33341)|(g18494);
assign g13832 = (g8880&g10612);
assign g23654 = ((~g20248));
assign II13037 = ((~g4304));
assign g32332 = (g31325&g23558);
assign II23099 = ((~g20682));
assign g33835 = (g4340&g33413);
assign g27427 = (g26400&g17575);
assign g25082 = ((~g22342));
assign II17885 = ((~g1135))|((~II17883));
assign g29900 = ((~g3639)&(~g28471));
assign g25128 = (g17418&g23525);
assign g12843 = ((~g10359));
assign g25727 = (g25163)|(g22010);
assign g33106 = (g32408&g18990);
assign g14549 = ((~g9992)&(~g12705));
assign g17677 = ((~g14882));
assign II18417 = (g14444)|(g14414)|(g14392);
assign g23473 = ((~g20785));
assign g10096 = ((~g5767));
assign g32315 = (g31306&g23517);
assign g10676 = (g8506&g3774);
assign g9321 = ((~g5863));
assign g32604 = ((~g31154));
assign g29624 = (g28491&g8070);
assign g20650 = ((~g15348));
assign gbuf114 = (g4185);
assign g27705 = ((~g25237))|((~g26782));
assign g33878 = (g33288&g20565);
assign g26679 = ((~g25385));
assign g27562 = (g26102)|(g24703);
assign g8284 = ((~g5002));
assign g25591 = (g24642)|(g21705);
assign g18394 = (g1862&g15171);
assign g32103 = (g31609&g29905);
assign g22360 = ((~II21849));
assign g32464 = ((~g30735));
assign g9973 = ((~g2112));
assign g21784 = (g3423&g20391);
assign g26517 = (g15708&g24367);
assign g32278 = (g2811&g30572);
assign g28480 = ((~g8059)&(~g27602));
assign g15164 = ((~g13835)&(~g12906));
assign g32070 = (g10967&g30825);
assign g32977 = (g32169)|(g21710);
assign g6816 = ((~g933));
assign g28615 = ((~g27817));
assign g22310 = (g19662&g20235);
assign g18519 = (g2648&g15509);
assign II17639 = ((~g13350));
assign g10087 = ((~II13597));
assign g32856 = ((~g31021));
assign g28164 = (g8651&g27528);
assign g32024 = ((~II29582));
assign g22998 = ((~g20391));
assign g18323 = (g1632&g17873);
assign g28041 = (g24145)|(g26878);
assign g34810 = ((~II33020));
assign g25909 = (g8745&g24875);
assign g32970 = ((~g30825));
assign g33811 = (g33439&g17573);
assign g13093 = ((~g10649))|((~g7661))|((~g979))|((~g1061));
assign II15800 = ((~g11607));
assign g34291 = (g34055&g19366);
assign g24993 = ((~g22384));
assign g14927 = ((~g12695))|((~g10281));
assign g26345 = (g13051&g25505);
assign g7118 = ((~g832));
assign II29285 = ((~g29489))|((~II29284));
assign II22640 = ((~g21256));
assign g30154 = (g28611&g23769);
assign II31076 = (g30614&g31809&g32564&g32565);
assign g32855 = ((~g30825));
assign g14892 = ((~g12700))|((~g12515));
assign g14142 = ((~g11715))|((~g8958));
assign g27181 = (g26026&g16655);
assign g7411 = ((~g2040));
assign g25712 = (g25126)|(g21963);
assign g24705 = (g2890)|(g23267);
assign g30209 = (g28682&g23876);
assign g31824 = ((~g29385));
assign g25942 = (g24422)|(g22298);
assign g29117 = ((~g27886));
assign g24525 = ((~g22670));
assign II22488 = ((~g18984));
assign g17724 = (g11547&g11592&g11640&II18713);
assign g9613 = ((~g5062));
assign II20957 = ((~g16228));
assign g6832 = ((~II11665));
assign g16704 = (g5957&g15018);
assign g23018 = ((~g19801));
assign II20569 = ((~g16486));
assign g32166 = (g31007&g23029);
assign g19552 = ((~g16856));
assign g32495 = ((~g31070));
assign g19718 = ((~g17015));
assign g28406 = ((~g27064))|((~g13675));
assign II27449 = ((~g27737));
assign g28055 = (g27560)|(g18190);
assign g7519 = ((~g1157));
assign g27567 = (g26121)|(g24714);
assign g26306 = (g13087&g25286);
assign g18352 = (g1798&g17955);
assign g25228 = ((~g23828));
assign g9397 = ((~g6088));
assign II14733 = ((~g9732))|((~g5475));
assign g17465 = ((~g12955));
assign g25119 = ((~g22384));
assign g25635 = (g24504)|(g18293);
assign II17733 = ((~g14844));
assign g32418 = (g31126&g16239);
assign g24533 = ((~g22876));
assign g33871 = (g33281&g20546);
assign II31287 = (g32870&g32871&g32872&g32873);
assign g24192 = (g311&g22722);
assign g14588 = (g11957&g11974);
assign g19605 = (g15707)|(g13063);
assign g27485 = (g26519&g17644);
assign g24891 = ((~g23231));
assign g29249 = (g28658)|(g18438);
assign g9681 = ((~g5798));
assign II33189 = ((~g34929));
assign g10401 = ((~g7041));
assign g17464 = (g14334)|(g14313)|(g11935)|(II18385);
assign g20576 = ((~g18065));
assign g18377 = (g1894&g15171);
assign g28117 = (g8075&g27245);
assign g10540 = ((~g9392));
assign g15144 = ((~g13716)&(~g12890));
assign g30334 = (g29837)|(g18143);
assign g7846 = ((~g4843))|((~g4878));
assign g26819 = (g106&g24490);
assign g14254 = ((~g11968))|((~g11933))|((~g11951));
assign g17133 = (g10683&g13222);
assign g11028 = (g9730&g5428);
assign II14833 = ((~g10142));
assign g17670 = ((~g3893))|((~g13772))|((~g4005))|((~g8595));
assign g28870 = ((~g27796))|((~g14588));
assign g18683 = (g4674&g15885);
assign g6846 = ((~g2152));
assign g24281 = (g23397)|(g18656);
assign g23292 = (g19879&g16726);
assign g24074 = ((~g21193));
assign g23394 = ((~II22499));
assign g28367 = ((~II26880));
assign g9828 = ((~g2024));
assign II31111 = (g31070&g31815&g32615&g32616);
assign g32677 = ((~g30673));
assign g10080 = ((~g1982));
assign g33237 = (g32394&g25198);
assign g34785 = ((~II32985));
assign II14611 = ((~g8678))|((~II14609));
assign g10564 = ((~g9462));
assign II15929 = ((~g10430));
assign g27737 = ((~g26718));
assign g27150 = (g25804)|(g24400);
assign g28877 = ((~g27937))|((~g7490))|((~g7431));
assign g33417 = (g32371&g21424);
assign g25231 = ((~g22228));
assign II14818 = ((~g6513))|((~II14816));
assign g34374 = (g26294)|(g34139);
assign g29327 = (g29070&g22156);
assign g11496 = (g4382&g7495);
assign g19761 = ((~g17015));
assign II28336 = ((~g29147));
assign g29242 = (g28674)|(g18354);
assign g13942 = (g5897&g12512);
assign g21181 = ((~g15426));
assign g9911 = ((~g2384));
assign II15824 = ((~g1116));
assign g32121 = (g31616&g29942);
assign g34151 = ((~II32106));
assign g34144 = ((~II32093));
assign g7581 = ((~g1379));
assign II32648 = ((~g34371));
assign g19952 = ((~g15915));
assign g15057 = ((~g6810)&(~g13350));
assign g29332 = (g29107&g22170);
assign g23553 = (g19413&g11875);
assign g19907 = ((~g16210)&(~g13676));
assign II20205 = ((~g11147))|((~II20203));
assign g30427 = (g29796)|(g21811);
assign g7443 = ((~g914));
assign g30096 = (g28546&g20770);
assign g34933 = ((~g34916));
assign g29577 = (g2441&g28946);
assign g27083 = (g25819&g22456);
assign II33146 = ((~g34903));
assign II31873 = (g33524)|(g33525)|(g33526)|(g33527);
assign g28294 = ((~g27295));
assign g32940 = ((~g31376));
assign g33977 = (g33876)|(g18348);
assign g18254 = (g1236&g16897);
assign g16841 = (g5913&g14858);
assign g31309 = (g30132&g27837);
assign g18699 = (g4760&g16816);
assign II32855 = ((~g34540));
assign g10078 = ((~g1854));
assign g21793 = (g3412&g20391);
assign g28348 = (g27139)|(g15823);
assign g33903 = (g33447&g19146);
assign g12321 = ((~g9637));
assign g22517 = ((~g19720)&(~g1345));
assign g26765 = ((~g25309));
assign g11107 = ((~g9095)&(~g9177));
assign g18453 = (g2315&g15224);
assign g23999 = ((~g21468));
assign g23776 = ((~g21177));
assign g20247 = ((~g17015));
assign g8267 = ((~g2342));
assign g31305 = (g29741&g23354);
assign g25616 = (g25096)|(g18172);
assign g7631 = ((~g74));
assign g8297 = ((~g142));
assign g18337 = (g1706&g17873);
assign II13065 = ((~g4308))|((~g4304));
assign g21863 = (g3957&g21070);
assign g21653 = ((~g17663));
assign g19748 = ((~g17015));
assign g12083 = ((~g2217))|((~g8205));
assign g27733 = ((~g9305)&(~g25805));
assign g19559 = ((~g16129));
assign g31840 = ((~g29385));
assign g21452 = (g16119&g13624);
assign g15863 = (g13762&g13223);
assign g11741 = ((~g10033));
assign g32352 = (g29852)|(g31282);
assign g13334 = ((~g11048));
assign g9586 = ((~g1668)&(~g1592));
assign g23265 = (g20069&g20132);
assign g21720 = (g376&g21037);
assign g30537 = (g30246)|(g22083);
assign g9015 = ((~g3050)&(~g3010));
assign g18997 = ((~II19756));
assign g33327 = (g32208&g20561);
assign II13749 = ((~g4608))|((~g4584));
assign g30479 = (g29320)|(g21950);
assign g8697 = ((~g3694));
assign g8150 = ((~g2185));
assign g29370 = ((~g28585)&(~g28599));
assign g25382 = ((~g12333))|((~g22342));
assign g7886 = ((~g1442));
assign g17708 = ((~g5216))|((~g14490))|((~g5313))|((~g12497));
assign g29687 = (g2407&g29097);
assign g18346 = (g1752&g17955);
assign g32437 = ((~II29965));
assign g34921 = ((~II33155));
assign II17876 = ((~g13070));
assign g26079 = (g6199&g25060);
assign g23534 = ((~II22665));
assign g7293 = ((~g4452));
assign g14879 = ((~g12646))|((~g10266));
assign g13913 = ((~g8859)&(~g11083));
assign II33030 = ((~g34768));
assign g23382 = ((~g20682));
assign g28181 = ((~II26700));
assign II31528 = ((~g33219));
assign II26479 = ((~g25771));
assign g33567 = (g33081)|(g18394);
assign g29552 = (g2223&g28579);
assign g13018 = ((~II15636));
assign g26087 = (g5475&g25072);
assign g25031 = (g20675&g23432);
assign g14262 = ((~g10838));
assign g34064 = (g33919)|(g33922);
assign g30341 = (g29380)|(g18246);
assign II32665 = ((~g34386));
assign g19637 = (g5142&g16958);
assign g10392 = ((~g6989));
assign g30156 = ((~g28789)&(~g14587));
assign II30983 = ((~g32433));
assign g11443 = ((~g9916))|((~g3649));
assign II18476 = ((~g14031));
assign g18889 = ((~g15509));
assign g13625 = ((~g10971));
assign g20094 = (g8872&g16631);
assign g26423 = (g19488&g24356);
assign II32479 = ((~g34302));
assign g24158 = ((~II23318));
assign g6826 = ((~g218));
assign g19731 = ((~g17093));
assign II18627 = ((~g14712))|((~II18625));
assign g20599 = ((~g18065));
assign g28467 = (g26993&g12295);
assign g17779 = ((~g6637))|((~g14556))|((~g6704))|((~g12471));
assign g7690 = ((~g4669))|((~g4659))|((~g4653));
assign g7697 = ((~g4087));
assign g34386 = (g10800&g34060);
assign g26743 = ((~g25476));
assign g30495 = (g30222)|(g21991);
assign II12991 = ((~g6752));
assign g9856 = ((~g5343));
assign g29014 = ((~g27742));
assign g34623 = (g34525)|(g18585);
assign g11203 = ((~g4966)&(~g4991)&(~g9064));
assign g23335 = ((~g20391));
assign g28228 = (g27126&g19636);
assign g25749 = (g25094)|(g18800);
assign g8635 = ((~g2783));
assign g23582 = ((~II22729));
assign g21736 = (g3065&g20330);
assign g33609 = (g33239)|(g18615);
assign g8234 = (g4515&g4521);
assign g24584 = ((~g22852))|((~g22836))|((~g22715));
assign II33109 = ((~g34851));
assign g21779 = (g3385&g20391);
assign g24027 = ((~g20014));
assign g7050 = ((~g5845));
assign g22689 = (g18918&g9104);
assign g10032 = ((~g562));
assign g33124 = (g8945&g32296);
assign g27679 = ((~g25186))|((~g26685));
assign g21463 = ((~g15588));
assign g11183 = ((~g8135));
assign g14630 = ((~g12402));
assign g14940 = ((~g12744))|((~g12581));
assign g34700 = (g34535&g20129);
assign g31990 = (g31772&g18945);
assign g8180 = ((~g262));
assign g25717 = (g25106)|(g21968);
assign II18906 = ((~g16963));
assign g25132 = (g10497&g23528);
assign g11244 = (g8346&g8566);
assign g32748 = ((~g31710));
assign g32204 = (g4245&g31327);
assign g30579 = (g30173)|(g14571);
assign g23716 = (g9194)|(g20905);
assign g21353 = ((~g11467))|((~g17157));
assign g14064 = ((~g9214)&(~g12259));
assign g31914 = (g31499)|(g22000);
assign g33761 = ((~II31616));
assign g27500 = (g26400&g17672);
assign g19365 = ((~g16249));
assign g14902 = ((~g7791))|((~g12581));
assign g14444 = ((~g11936)&(~g9692));
assign g16632 = ((~g14454));
assign g17523 = ((~g14732));
assign g33646 = (g33389&g18876);
assign g9055 = (g2606)|(g2625);
assign g28981 = ((~g9234)&(~g27999));
assign g21010 = ((~g15634));
assign g15160 = ((~g12903)&(~g13809));
assign g23754 = (g14816&g21189);
assign g21049 = ((~g17433));
assign g30268 = (g28777&g23969);
assign g24631 = ((~g20516)&(~g20436)&(~g20219)&(~g22957));
assign g7909 = ((~g936));
assign g26080 = (g19393)|(g24502);
assign g34664 = ((~II32782));
assign g28178 = (g27019&g19397);
assign g31708 = ((~II29278))|((~II29279));
assign II29013 = ((~g29705));
assign g19479 = ((~g16449));
assign g24323 = (g4546&g22228);
assign g32615 = ((~g31376));
assign g23042 = ((~g16581)&(~g19462)&(~g10685));
assign g24125 = ((~g19890));
assign II21477 = ((~g18695));
assign g29923 = ((~g28874));
assign g25607 = (g24773)|(g18118);
assign g7121 = ((~II11820));
assign g33687 = (g33132&g4878);
assign g17569 = (g14416)|(g14394)|(g11995)|(II18492);
assign II16538 = ((~g10417));
assign g33346 = ((~g32132));
assign g31968 = (g31757&g22168);
assign g32792 = ((~g31710));
assign g32164 = (g30733&g25171);
assign g32918 = ((~g31327));
assign g24407 = ((~g22594));
assign II28582 = ((~g30116));
assign g23742 = (g19128&g9104);
assign g28425 = ((~g27493)&(~g26351));
assign g28215 = (g9264&g27565);
assign gbuf95 = (g3969);
assign g25702 = (g25068)|(g21921);
assign g13104 = ((~g1404))|((~g10794));
assign g20562 = ((~g17955));
assign g9555 = ((~II13206));
assign g31324 = (g30171&g27937);
assign g27372 = (g26488&g17476);
assign gbuf136 = (g215);
assign g28358 = (g27149)|(g15837);
assign g22053 = (g6116&g21611);
assign g18610 = (g15088&g17059);
assign g24261 = (g22862)|(g18314);
assign g33456 = ((~II30986));
assign g27990 = ((~g26770));
assign g34350 = (g26048)|(g34106);
assign g29795 = (g28344&g23257);
assign g34580 = (g29539&g34311);
assign g16675 = ((~II17873));
assign g19410 = ((~g16449));
assign g19530 = ((~g15829))|((~g10841));
assign g13084 = ((~g5587))|((~g12093))|((~g5677))|((~g9864));
assign g26286 = (g2126&g25389);
assign g19061 = ((~II19762));
assign g32799 = ((~g31710));
assign g28285 = (g9657&g27717);
assign g33119 = (g32420)|(g32428);
assign g30083 = (g28533&g20698);
assign g11415 = ((~g8080)&(~g8026));
assign II18367 = ((~g13010));
assign g25709 = (g25014)|(g21960);
assign g30452 = (g29891)|(g21861);
assign g10710 = ((~II14006));
assign g17096 = ((~II18168));
assign II27518 = (g20720&g24104&g24105&g24106);
assign g12885 = ((~g10382));
assign g27012 = ((~g6398)&(~g25856));
assign g29171 = ((~g27937));
assign II29002 = ((~g29675));
assign g12908 = ((~g10414));
assign g12028 = ((~II14884))|((~II14885));
assign II32696 = ((~g34434));
assign g18988 = ((~g15979));
assign g15814 = (g3574&g13920);
assign g19394 = ((~g16326));
assign II14046 = ((~g9900));
assign g27147 = (g25802)|(g24399);
assign g24018 = ((~II23162)&(~II23163));
assign gbuf128 = (g878);
assign g28900 = ((~g27886))|((~g7451))|((~g2040));
assign g29081 = ((~g27837));
assign g8873 = ((~II12849))|((~II12850));
assign g32965 = ((~g31710));
assign g28312 = (g27828&g26608);
assign g18715 = (g4871&g15915);
assign II23684 = ((~g23230));
assign g11372 = (g490)|(g482)|(g8038);
assign g23249 = ((~g21070));
assign g34492 = (g34272&g33430);
assign g13298 = ((~II15862));
assign g10290 = (g4358&g4349);
assign g14001 = ((~g739)&(~g11083));
assign II12826 = ((~g4349));
assign g30052 = ((~g29018));
assign g11279 = ((~g8504))|((~g3443));
assign g28727 = (g27500)|(g16729);
assign II32062 = ((~g33653));
assign g18382 = (g1936&g15171);
assign g13042 = (g433&g11048);
assign II14499 = ((~g8737))|((~II14497));
assign g33895 = ((~II31751));
assign II21787 = ((~g19422));
assign II29204 = ((~g29505));
assign g9617 = ((~II13240));
assign g9402 = ((~g6209));
assign g32570 = ((~g31554));
assign g24989 = ((~g21345))|((~g23363));
assign g29915 = ((~g6941)&(~g28484));
assign g33864 = (g33274&g20524);
assign g13311 = ((~II15878));
assign g17014 = ((~g14297));
assign g11867 = ((~II14679));
assign g31667 = ((~g30142));
assign g14277 = ((~II16455));
assign g24011 = (g7939&g19524);
assign g29594 = (g28529&g14192);
assign g14212 = ((~g5373)&(~g10537));
assign II15308 = ((~g2407))|((~II15306));
assign II29296 = ((~g29495))|((~II29295));
assign g33112 = ((~g31240)&(~g32194));
assign g29369 = (g28209&g22341);
assign g18230 = (g1111&g16326);
assign g13069 = ((~g5889))|((~g12067))|((~g6000))|((~g9935));
assign g34862 = (g16540&g34830);
assign g27586 = ((~g24924))|((~g24916))|((~g24905))|((~g26863));
assign g32833 = ((~g30825));
assign g25015 = ((~g23662));
assign g14342 = ((~g12163));
assign g23849 = ((~g19277));
assign g10207 = ((~g6315))|((~g6358))|((~g6329))|((~g6351));
assign g16290 = ((~g13260));
assign g30374 = (g30078)|(g18465);
assign g8345 = ((~g3794));
assign g8745 = ((~g744));
assign g10554 = ((~g8974));
assign g18766 = (g5495&g17929);
assign g29216 = ((~II27564));
assign g34707 = (g34544&g20579);
assign g24304 = (g12875&g22228);
assign g34338 = (g34099&g19905);
assign g30729 = ((~II28883));
assign g12222 = ((~g8310))|((~g2028));
assign g28280 = (g23761&g27724);
assign II13473 = ((~g4157));
assign g25240 = ((~g23650));
assign g19128 = ((~II19778));
assign g24881 = (g3050&g23211&II24048);
assign II33161 = ((~g34894));
assign g30387 = (g30151)|(g18524);
assign g16605 = ((~g13955));
assign g30179 = (g28634&g23819);
assign g7927 = ((~g4064));
assign g33657 = (g30991&g33443);
assign g33244 = (g32190&g23152);
assign II13548 = ((~g94));
assign II18492 = (g14538)|(g14513)|(g14446);
assign II15195 = ((~g6005))|((~II15193));
assign g32325 = (g31316&g23538);
assign g12020 = ((~g2028))|((~g8365));
assign g27328 = (g12482&g26736);
assign g16536 = (g5917&g14996);
assign g26274 = (g2130&g25210);
assign g26252 = (g2283&g25309);
assign II12719 = ((~g365));
assign g19785 = ((~g16987));
assign g25647 = (g24725)|(g21740);
assign g13264 = ((~g11869))|((~g11336))|((~g11849));
assign g28455 = (g27289&g20103);
assign g32141 = (g31639&g29963);
assign g26327 = (g8462)|(g24591);
assign g34428 = ((~II32455));
assign g33958 = (g33532)|(II31873)|(II31874);
assign g27342 = (g12592&g26792);
assign g25695 = (g24998)|(g21914);
assign g33360 = (g32253&g20869);
assign g21427 = ((~g17367));
assign g9390 = ((~g5808));
assign II32994 = ((~g34739));
assign g29970 = ((~II28199));
assign g31997 = ((~g22306))|((~g30580));
assign g22096 = (g6434&g18833);
assign g18342 = (g1592&g17873);
assign g32693 = ((~g31579));
assign II32997 = ((~g34760));
assign g13993 = ((~g3961))|((~g11255))|((~g3969))|((~g11419));
assign g25541 = ((~g22763));
assign II18304 = ((~g14790));
assign II24582 = (g9809&g9397&g6093);
assign g32672 = ((~g31579));
assign g33367 = (g32271&g21053);
assign g18629 = (g3680&g17226);
assign II16610 = ((~g10981));
assign g25762 = (g25095)|(g18816);
assign g14228 = ((~g5719)&(~g10561));
assign g24357 = ((~g22325));
assign g12824 = ((~g5881)&(~g9451));
assign g31245 = (g25964)|(g29516);
assign g26968 = (g26307)|(g24321);
assign II14644 = ((~g7717));
assign g28517 = (g27280)|(g26154);
assign II18320 = ((~g13605));
assign g26244 = (g24688&g8812&g10658&g8757);
assign g34371 = (g7450&g34044);
assign g33504 = (g32772&II31216&II31217);
assign g34981 = ((~g34973));
assign g29129 = ((~g27858));
assign g18979 = ((~g16136));
assign g7087 = ((~g6336));
assign g11012 = ((~g7693)&(~g7846));
assign g26346 = ((~g8522)&(~g24825));
assign g24033 = ((~g19919));
assign g33620 = (g33360)|(g18774);
assign II15593 = ((~g11989));
assign g14511 = (g10685)|(g546);
assign g24893 = ((~II24060));
assign g34975 = (g34871)|(g34964);
assign g34721 = (g34696)|(g18135);
assign g31523 = (g7528&g29333);
assign g28601 = (g27506&g20514);
assign II33214 = ((~g34954));
assign g16528 = ((~g14154));
assign g13597 = (g9247)|(g11149);
assign g28730 = (g27503)|(g13912);
assign g34046 = (g33906)|(g33908);
assign g20450 = ((~g15277));
assign g8740 = ((~II12735));
assign g24234 = (g22622)|(g18237);
assign g34059 = ((~g33658));
assign g32520 = ((~g31554)&(~II30054)&(~II30055));
assign g10822 = (g4264&g8514);
assign g12478 = ((~II15299))|((~II15300));
assign g23893 = ((~g19074));
assign II22619 = ((~g21193));
assign g20978 = ((~g15595));
assign II19235 = ((~g15078));
assign g20697 = ((~g17433));
assign g32736 = ((~g30937));
assign II16770 = ((~g6023));
assign g10367 = ((~g6870));
assign g24756 = ((~g22763));
assign g24700 = (g645&g23512);
assign g24950 = ((~g19442))|((~g23154));
assign g33516 = (g32860&II31276&II31277);
assign g15823 = (g3945&g14116);
assign g8057 = ((~g3068));
assign II24365 = ((~g14320))|((~II24363));
assign g13727 = ((~g174))|((~g203))|((~g168))|((~g12812));
assign g24489 = ((~II23694));
assign g14098 = ((~g11566))|((~g8864));
assign II13044 = ((~g5115))|((~II13043));
assign g18816 = (g6527&g15483);
assign g18624 = (g3490&g17062);
assign g11677 = ((~g7689));
assign g22641 = (g18974)|(g15631);
assign II17834 = ((~g14977));
assign g28739 = (g21434&g26424&g25274&g27395);
assign g32367 = (g29880)|(g31309);
assign g26393 = (g19467&g25558);
assign g26770 = (g24471)|(g10732);
assign g20682 = (g16238&g4646);
assign g7349 = ((~g1270));
assign g23059 = ((~g20453));
assign g25046 = ((~g23729));
assign g17634 = ((~g3219))|((~g11217))|((~g3281))|((~g13877));
assign g21678 = ((~g16540));
assign g26777 = ((~g25439));
assign II24445 = ((~g22923));
assign g26936 = ((~II25680));
assign g27121 = (g136&g26326);
assign g33934 = ((~II31814));
assign II20399 = ((~g16205));
assign g16243 = (g6483&g14275);
assign g14520 = ((~g9369))|((~g12163));
assign II11864 = ((~g4434))|((~g4401));
assign g33250 = ((~g32186));
assign g23835 = ((~g2791)&(~g21303));
assign g25041 = (g23261&g20494);
assign II25221 = ((~g24718))|((~II25219));
assign g27696 = (g25800&g23647);
assign g27265 = (g26785&g26759);
assign g20648 = ((~g15615));
assign g29110 = (g27187&g12687&g20751&II27429);
assign g32458 = ((~g30825));
assign g16777 = ((~II18003));
assign g18430 = (g2204&g18008);
assign g15655 = ((~g13202));
assign g16684 = ((~g14223));
assign II24505 = (g9607&g9229&g5057);
assign g32017 = ((~g31504)&(~g23475));
assign g14643 = (g11998&g12023);
assign g27559 = (g26576&g17777);
assign g21974 = (g5517&g19074);
assign II16660 = ((~g10981));
assign II14764 = ((~g9808))|((~g5821));
assign g16423 = ((~g14066));
assign II32185 = ((~g33665))|((~g33661));
assign g32569 = ((~g30673));
assign g20057 = ((~g16349));
assign g13857 = ((~II16163));
assign g16965 = (g269&g13140);
assign g24650 = (g22641&g19718);
assign g17683 = ((~g15027));
assign g28299 = (g9716&g27670);
assign gbuf79 = (g3092);
assign g12460 = ((~g10093))|((~g5644))|((~g5694));
assign g30127 = (g28494)|(g16805);
assign g23165 = (g13954&g19964);
assign g25937 = (g24406)|(g22216);
assign g11428 = ((~g7615));
assign g17198 = ((~g9282)&(~g14279));
assign g21843 = (g3869&g21070);
assign g30352 = (g30094)|(g18340);
assign g33260 = (g32110)|(g29524);
assign g12198 = ((~g9797)&(~g9800));
assign g34954 = ((~II33210));
assign g25101 = ((~g22384));
assign g32387 = (g31489)|(g29952);
assign g34510 = ((~g34418));
assign II18845 = ((~g6711));
assign g28251 = (g27826&g23662);
assign g27670 = ((~g25172))|((~g26666));
assign g12656 = ((~g7028));
assign g34612 = (g34514)|(g18566);
assign g33380 = (g32234)|(g29926);
assign g23356 = ((~g21070));
assign g25529 = ((~g22763));
assign gbuf145 = (g1459);
assign g20093 = (g15372&g14584);
assign g24245 = (g22849)|(g18256);
assign g33143 = ((~g32293)&(~g31518));
assign g31887 = (g31292)|(g21820);
assign g19335 = ((~g15717))|((~g1056));
assign g18727 = (g4931&g16077);
assign g15736 = ((~g6295))|((~g14575))|((~g6373))|((~g10003));
assign g9992 = ((~g5990));
assign gbuf51 = (g6315);
assign g30215 = (g28690&g23881);
assign g9691 = ((~g1706));
assign II13539 = ((~g6381));
assign g34751 = (g34674&g19543);
assign g21807 = (g3566&g20924);
assign g19541 = ((~g16136));
assign g28064 = (g27298)|(g21781);
assign g34860 = (g16540&g34823);
assign g32871 = ((~g30937));
assign g24577 = (g2856)|(g22531);
assign g10362 = ((~g6850));
assign g27128 = (g25997&g16583);
assign g18686 = (g4659&g15885);
assign g27829 = ((~g7345)&(~g25856));
assign g15159 = ((~g13809)&(~g12902));
assign g32937 = ((~g31021));
assign g34440 = (g34364)|(g24226);
assign g9749 = ((~g1691));
assign g16867 = (g13493)|(g11045);
assign g14999 = ((~g12739))|((~g12824));
assign II14899 = ((~g10198));
assign g34733 = (g34678)|(g18651);
assign g20025 = ((~g17271));
assign g17309 = ((~g9305)&(~g14344));
assign g22108 = (g6439&g18833);
assign g13798 = ((~g11280))|((~g3423));
assign g34111 = (g33733&g22936);
assign g19951 = ((~g16219)&(~g13709));
assign II18716 = (g13156&g11450&g6756);
assign g13697 = (g11166&g8608);
assign gbuf8 = (g4304);
assign II29965 = ((~g31189));
assign g27647 = ((~g3004)&(~g26616));
assign g28324 = (g9875&g27687);
assign g15120 = ((~g12873)&(~g13605));
assign II31107 = (g32610&g32611&g32612&g32613);
assign g16760 = (g5559&g14764);
assign g34943 = ((~II33197));
assign g24772 = (g16287&g23061);
assign g18313 = (g1430&g16931);
assign g28106 = ((~g7812)&(~g26994));
assign g25988 = (g9510&g25016);
assign g34597 = ((~II32699));
assign II32051 = ((~g33631));
assign g29518 = (g28906&g22384);
assign g32172 = (g2767&g31608);
assign g18169 = (g676&g17433);
assign g12898 = ((~g10405));
assign g31296 = (g30119&g27779);
assign g34935 = ((~II33189));
assign g33288 = (g32147)|(g29587);
assign g32921 = ((~g31672));
assign g28156 = ((~II26667));
assign g22216 = (g13660&g20000);
assign g33371 = (g32280&g21155);
assign g21402 = ((~g17757))|((~g14740))|((~g17716))|((~g14674));
assign g33534 = (g33186)|(g21700);
assign II31782 = ((~g33219));
assign gbuf27 = (g5637);
assign II13510 = ((~g2089))|((~II13509));
assign g6955 = ((~II11726));
assign g21936 = (g5200&g18997);
assign g10379 = ((~g6953));
assign II12372 = ((~g3457))|((~g3462));
assign g30541 = (g30281)|(g22087);
assign g30082 = (g29181&g12752);
assign g29765 = ((~II28014));
assign g25409 = ((~g22228));
assign g33376 = (g32294&g21268);
assign g32508 = ((~g30825));
assign g29489 = (g28550)|(g27601);
assign g17400 = ((~II18333));
assign gbuf20 = (g5308);
assign g32040 = (g14122&g31243);
assign g23967 = ((~g19210));
assign g9576 = ((~g6565));
assign II26578 = ((~g26941));
assign g30047 = (g29109&g9407);
assign II21029 = ((~g15816));
assign g33420 = (g32373&g21454);
assign g16700 = (g5208&g14838);
assign g18947 = ((~g16136));
assign g13409 = ((~II15918));
assign g22153 = ((~g18997));
assign g11293 = ((~g7527));
assign g20153 = ((~g16782));
assign gbuf42 = (g6000);
assign II12382 = ((~g47));
assign g27484 = (g25988)|(g24628);
assign g33885 = (g33296&g20609);
assign g27035 = (g26348&g1500);
assign g13252 = (g11561&g11511&g11469&g699);
assign g13544 = ((~g7972))|((~g10521))|((~g7549))|((~g1008));
assign g22830 = ((~g20283));
assign g15794 = (g3239&g14008);
assign II31006 = (g31376&g31796&g32464&g32465);
assign g33046 = (g32308)|(g21912);
assign g33858 = (g33268&g20448);
assign g24722 = (g17618&g22417);
assign g34858 = (g16540&g34816);
assign g14160 = ((~g11626))|((~g8958));
assign g34310 = (g14003&g34162);
assign g32585 = ((~g31542)&(~II30123)&(~II30124));
assign g18603 = (g3119&g16987);
assign g33083 = ((~g7805))|((~g32118));
assign g7301 = ((~g925));
assign II15051 = ((~g9759))|((~g2259));
assign g22682 = ((~g19379));
assign g18722 = (g4917&g16077);
assign g29744 = ((~g28431));
assign g34797 = (g34747)|(g18574);
assign g33702 = ((~II31545));
assign g14167 = ((~II16371));
assign g28560 = (g27311)|(g26249);
assign g21865 = (g3965&g21070);
assign g18545 = (g2783&g15277);
assign g29057 = ((~g27800))|((~g9649));
assign g33443 = ((~II30971));
assign g20770 = ((~g17955));
assign II12963 = ((~g640));
assign II12530 = ((~g4815));
assign g34182 = (g33691&g24384);
assign II18538 = ((~g14642))|((~II18536));
assign g30594 = (g18898&g29846);
assign II27364 = (g25541&g26424&g22698);
assign g23850 = ((~g12185))|((~g19462));
assign g26886 = (g26651)|(g24192);
assign g22158 = (g13698&g19609);
assign g28374 = (g27181)|(g15850);
assign II32935 = ((~g34657));
assign g32150 = (g31624&g29995);
assign g11178 = (g6682&g7097&g6668&g10061);
assign g29168 = (g27658)|(g26613);
assign g15856 = (g9056&g14223);
assign g12846 = ((~g6837)&(~g10430));
assign g19566 = ((~g16136));
assign g30481 = (g30221)|(g21977);
assign g29616 = (g1974&g29085);
assign g31070 = (g29814&g25985);
assign g22104 = (g6444&g18833);
assign g11302 = ((~g9496))|((~g3281));
assign g22083 = (g6287&g19210);
assign g21156 = ((~g17247));
assign g16431 = ((~II17675));
assign g14272 = ((~g6411)&(~g10598));
assign g21271 = ((~II21002));
assign g20005 = ((~g17433));
assign g25071 = (g12804&g23478);
assign g22048 = (g6052&g21611);
assign g27349 = ((~g26352));
assign g33282 = (g32143)|(g29577);
assign g26352 = ((~g744))|((~g24875))|((~g11679));
assign g6756 = ((~II11623));
assign g18096 = ((~II18894));
assign g32719 = ((~g31672));
assign g23947 = ((~g19210));
assign g33802 = (g33097&g14545);
assign g15732 = (g13411)|(g13384)|(g13349)|(g11016);
assign g30436 = (g29860)|(g21845);
assign g14163 = ((~g8997)&(~g12259));
assign II25366 = ((~g24477));
assign II27564 = ((~g28166));
assign II11878 = ((~g4388))|((~II11877));
assign g29032 = ((~g9300)&(~g27999));
assign g14209 = ((~g11415));
assign g29186 = ((~g27051))|((~g4507));
assign g31148 = (g2661&g30055);
assign g29968 = (g2433&g28843);
assign g32811 = ((~g30735));
assign g29276 = (g28616)|(g18709);
assign g10568 = ((~g7328))|((~g7374));
assign g25095 = (g23319&g20556);
assign g21399 = ((~g15224));
assign g29861 = (g28390&g23313);
assign g20164 = ((~g16826));
assign g25750 = (g25543)|(g18802);
assign g27600 = (g26755&g26725);
assign g34773 = ((~II32963));
assign II12026 = ((~g344));
assign g21302 = (g956&g15731);
assign g11511 = ((~II14481))|((~II14482));
assign g18365 = (g1848&g17955);
assign II15262 = ((~g10081))|((~g2273));
assign g17242 = ((~g14454));
assign g18696 = (g4741&g16053);
assign g12259 = (g9480&g640);
assign g25573 = (II24704&II24705);
assign II27730 = ((~g28752));
assign g26905 = (g26397)|(g24222);
assign g17745 = ((~g14978));
assign g25198 = ((~g22228));
assign g31285 = (g30134&g27800);
assign g15800 = (g10821)|(g13242);
assign g23547 = ((~g21611));
assign g23932 = ((~g7051))|((~g20875));
assign g33299 = ((~g608))|((~g32296))|((~g12323));
assign II25786 = ((~g26424));
assign g23611 = ((~g18833));
assign g14279 = ((~g12111))|((~g9246));
assign g34568 = (g34379&g17512);
assign g11418 = ((~II14424));
assign g7392 = ((~g4438));
assign g34160 = ((~II32119));
assign II12611 = (g1500)|(g1582)|(g1333);
assign g28559 = ((~g27700));
assign g21743 = (g3100&g20330);
assign g12779 = ((~g9444));
assign g21854 = (g3921&g21070);
assign II19917 = ((~g18088));
assign g18987 = (g182&g16162);
assign g8791 = ((~II12787));
assign g21890 = (g4125&g19801);
assign g17817 = (g11547&g6782&g11640&II18819);
assign g7643 = ((~g4322));
assign g13144 = ((~II15773));
assign g26267 = ((~g8033)&(~g24732));
assign g16260 = ((~g4888))|((~g13910))|((~g12088));
assign g33927 = (g33094&g21412);
assign g20371 = ((~g16956))|((~g14088))|((~g16694))|((~g16660));
assign g27930 = ((~II26451));
assign g29028 = ((~g27933))|((~g8381));
assign g21193 = ((~g15348)&(~g12135));
assign g28521 = ((~g27649)&(~g26604));
assign g34255 = (g34120)|(g24302);
assign g10312 = ((~g5881)&(~g5873));
assign g28684 = (g27432)|(g16636);
assign g29774 = (g28287&g10233);
assign g25370 = ((~g22228));
assign g6800 = ((~g203));
assign g10157 = ((~g2036));
assign g24639 = (g6181&g23699);
assign g34989 = ((~II33267));
assign g27555 = (g26095)|(g24686);
assign g31300 = (g30148&g27858);
assign g26363 = (g2965)|(g24965);
assign g27255 = (g25936&g19689);
assign g22114 = (g6565&g19277);
assign II12728 = ((~g4291))|((~g4287));
assign g16969 = ((~g14262));
assign g16718 = ((~II17932));
assign II31292 = (g32877&g32878&g32879&g32880);
assign g31220 = (g30273&g25202);
assign g19483 = ((~g15969))|((~g10841))|((~g10922));
assign g31240 = (g14793&g30206);
assign g14330 = ((~II16486));
assign g26792 = ((~g25439));
assign g16582 = ((~g13915));
assign II31535 = ((~g33377));
assign g8964 = ((~g4269));
assign g15070 = ((~g6829)&(~g13416));
assign g20659 = ((~g17873));
assign g16523 = ((~g14041));
assign g16099 = ((~g13437));
assign g11666 = ((~g8172)&(~g8125));
assign g29669 = ((~II27941));
assign g12869 = ((~g10376));
assign g22171 = ((~g18882));
assign g18823 = (g6727&g15680);
assign g32999 = (g32337)|(g18401);
assign g21991 = (g5595&g19074);
assign g28430 = (g27229)|(g15914);
assign g6917 = ((~g3684));
assign g32596 = ((~g31070));
assign g24672 = (g19534&g22981);
assign g26248 = ((~II25220))|((~II25221));
assign II31196 = (g30825&g31830&g32738&g32739);
assign g23085 = ((~g19957));
assign g23822 = (g20218)|(g16929);
assign g29344 = (g29168&g18932);
assign II17989 = ((~g14173));
assign II14241 = ((~g8356));
assign g29717 = (g28200)|(g10883);
assign g34608 = (g34568)|(g15082);
assign g29286 = (g28542)|(g18759);
assign g31496 = (g2338&g30312);
assign g28492 = ((~g3857)&(~g7121)&(~g27635));
assign g16587 = ((~II17763));
assign g24657 = (g22644&g19730);
assign II13937 = (g7340&g7293&g7261);
assign g30508 = (g30199)|(g22029);
assign g18308 = (g6832&g16931);
assign gbuf141 = (g1576);
assign g30102 = ((~g29157));
assign g7673 = (g4153)|(g4172);
assign g14406 = ((~g12249));
assign g7436 = ((~g5276));
assign g33996 = (g33862)|(g18426);
assign g34189 = (g33801)|(g33808);
assign g29237 = (g28185)|(g18289);
assign II32929 = ((~g34649));
assign g27239 = (g25881)|(g24465);
assign g24047 = ((~g19919));
assign g21410 = ((~g15224));
assign g32866 = ((~g30614));
assign g28132 = (g27932)|(g27957);
assign g18411 = (g2093&g15373);
assign II32904 = ((~g34708));
assign II17098 = ((~g14336));
assign II27524 = (g28037&g24114&g24115&g24116);
assign g28142 = ((~II26649));
assign g34269 = (g34083)|(g18732);
assign g34214 = (g33772&g22689);
assign II30469 = (g31672)|(g31710)|(g31021)|(g30937);
assign g25193 = ((~g22763));
assign II32967 = ((~g34648));
assign g17249 = ((~II18265));
assign g29646 = (g1816&g28675);
assign g22654 = ((~g7733)&(~g19506));
assign g20132 = ((~g16931));
assign g7594 = ((~II12064));
assign g24977 = (g23209&g20232);
assign g8928 = ((~g4340));
assign g25848 = (g25539&g18977);
assign II31137 = (g32654&g32655&g32656&g32657);
assign g23929 = ((~g19147));
assign g33572 = (g33339)|(g18414);
assign g27177 = (g25997&g16651);
assign g19879 = (g15841)|(g13265);
assign g10531 = ((~g8925));
assign II12544 = ((~g191))|((~g194));
assign g24272 = (g23056)|(g18629);
assign g28428 = (g27227)|(g15912);
assign g23446 = ((~g21562));
assign g28556 = (g27431&g20374);
assign g34563 = (g34372&g17465);
assign g9372 = ((~g5080))|((~g5084));
assign II23961 = ((~g23184))|((~g13631));
assign g17764 = ((~II18758));
assign g12894 = ((~g10401));
assign g25881 = (g3821&g24685);
assign g14946 = ((~g6247))|((~g12173))|((~g6346))|((~g12672));
assign g20113 = ((~g16826));
assign g23751 = (g21415)|(g21402)|(II22880);
assign g25929 = (g24395)|(g22193);
assign g15741 = ((~g5244))|((~g14490))|((~g5320))|((~g14631));
assign g18635 = (g3808&g17096);
assign g16735 = (g6235&g15027);
assign II21976 = ((~g7680))|((~g19620));
assign g15978 = (g246&g14032);
assign g29230 = (g28107)|(g18202);
assign g9645 = ((~g2060))|((~g2028));
assign g14697 = ((~g12662))|((~g12824));
assign g24808 = ((~II23986))|((~II23987));
assign g27405 = (g24572)|(g25968);
assign g30188 = (g28644&g23841);
assign g21249 = ((~g15509));
assign g8906 = ((~g3530)&(~g3522));
assign g18574 = (g2882&g16349);
assign g32380 = (g29907)|(g31467);
assign g33709 = (g32414)|(g33441);
assign g22524 = ((~g19720)&(~g1361));
assign g32817 = ((~g31376));
assign g32392 = (g31513)|(g30000);
assign g21051 = ((~g15171));
assign g22594 = ((~II21934));
assign g18317 = (g12846&g17873);
assign g18478 = (g2445&g15426);
assign II22604 = ((~g21143));
assign g25974 = ((~g24576))|((~g22837));
assign g17515 = ((~g13221)&(~g10828));
assign II29254 = ((~g29482))|((~II29253));
assign gbuf131 = (g887);
assign g21764 = (g3227&g20785);
assign g30243 = (g28731&g23929);
assign g12721 = ((~g10061));
assign g28390 = (g27207)|(g15861);
assign g28300 = (g27771&g26605);
assign g25623 = (g24552)|(g18219);
assign g28389 = (g27206)|(g15860);
assign g34234 = (g32520)|(g33952);
assign g29203 = (g24095&II27513&II27514);
assign g27241 = (g24584)|(g25984);
assign g14678 = ((~g12432)&(~g9907));
assign II31121 = (g30614&g31817&g32629&g32630);
assign g24963 = ((~g22342));
assign g25875 = (g8390&g24809);
assign g22168 = ((~g19147));
assign g25211 = ((~g22763));
assign g26670 = (g13385&g24428);
assign g29854 = (g2197&g29092);
assign g30400 = (g29766)|(g21759);
assign g25450 = (g6888&g22497);
assign g16713 = ((~II17924))|((~II17925));
assign g30275 = (g28816&g23984);
assign g34624 = (g34509)|(g18592);
assign g6855 = ((~g2711));
assign g9924 = ((~g5644));
assign g17953 = ((~II18861));
assign g23574 = (g20093)|(g20108);
assign g25997 = ((~II25095));
assign g14357 = ((~g12181));
assign g20214 = ((~g16854))|((~g13993))|((~g16776))|((~g13967));
assign g28586 = (g27484&g20497);
assign g33945 = (g32430)|(g33455);
assign g15608 = ((~g11885)&(~g14212));
assign g34121 = ((~II32056));
assign g18784 = (g15155&g18065);
assign g16627 = ((~II17819));
assign g16172 = ((~g13584));
assign g17396 = ((~g7345))|((~g14272));
assign g21369 = ((~g16285));
assign II15821 = ((~g11143));
assign g22871 = (g9523&g20871);
assign g34710 = (g34553&g20903);
assign g17518 = ((~g14918));
assign g32705 = ((~g30614));
assign II13634 = ((~g79));
assign II14687 = ((~g7753));
assign gbuf81 = (g3654);
assign II20486 = ((~g16696))|((~g16757));
assign II15176 = ((~g2661))|((~II15174));
assign II26409 = ((~g26187));
assign g24070 = ((~g20014));
assign g29069 = ((~g9381)&(~g28010));
assign g32903 = ((~g31376));
assign g23540 = (g16866&g20622);
assign II20867 = ((~g16216));
assign g28830 = ((~g27886))|((~g7451))|((~g7369));
assign g19356 = (g17784)|(g14874);
assign g33614 = (g33249)|(g18650);
assign II32591 = ((~g34287));
assign g9003 = ((~g790));
assign g10382 = ((~g6958));
assign g34208 = ((~g33838));
assign g16228 = ((~II17569));
assign g19866 = ((~g16540));
assign II32775 = ((~g34512));
assign g26093 = ((~g24814));
assign g18294 = (g15072&g16449);
assign g32030 = (g4172&g30937);
assign g28494 = (g27973&g17741);
assign g29620 = (g2399&g29097);
assign g26547 = (g13283&g25027);
assign g7479 = ((~g1008));
assign g11119 = ((~g9180)&(~g9203));
assign II31336 = (g31672&g31855&g32940&g32941);
assign g12837 = ((~g10354));
assign g34079 = (g33703&g19532);
assign II17873 = ((~g15017));
assign g24151 = (g18088)|(g21661);
assign g21291 = ((~g16620));
assign g25684 = (g24983)|(g18643);
assign g17144 = ((~g14085));
assign g16621 = (g8278&g13821);
assign g12115 = ((~g1926))|((~g8249));
assign g33073 = (g32386&g18828);
assign g34918 = ((~II33146));
assign II14346 = ((~g10233));
assign g26397 = (g19475&g25563);
assign g22068 = (g6219&g19210);
assign g30443 = (g29808)|(g21852);
assign II32843 = ((~g34499));
assign g9601 = ((~g4005));
assign g19574 = ((~g16826));
assign g31259 = (g25992)|(g29554);
assign II15298 = ((~g10112))|((~g1982));
assign g32039 = (g31476&g20070);
assign g7765 = ((~g4165));
assign g27985 = ((~g26131));
assign g29961 = ((~g28892));
assign g28564 = (g27314)|(g26252);
assign g22866 = ((~g20330));
assign g25323 = (g6888&g22359);
assign II12064 = ((~g617));
assign g33691 = ((~II31528));
assign g34754 = (g34677&g19602);
assign g9967 = (g1178&g1157);
assign g25223 = (g22523&g10652);
assign g22651 = ((~g20114))|((~g2873));
assign II18574 = ((~g13075));
assign g29746 = (g28279&g20037);
assign II19799 = ((~g17817));
assign g23840 = ((~g19074));
assign g30258 = (g28751&g23953);
assign g19799 = ((~g17062));
assign g33537 = (g33244)|(g21716);
assign II17932 = ((~g3310));
assign g12227 = ((~g8418))|((~g8330));
assign g9631 = ((~g6573));
assign g9983 = ((~g4239));
assign g23902 = ((~g21468));
assign g22358 = ((~g19801));
assign g11936 = ((~g8241))|((~g1783));
assign g27665 = (g26872&g23519);
assign g32045 = (g31491&g16187);
assign g33730 = (g7202&g4621&g33127&g4633);
assign g15837 = (g3255&g14127);
assign g8480 = ((~g3147));
assign g22128 = (g6629&g19277);
assign g30397 = (g29747)|(g21756);
assign II17924 = ((~g13378))|((~II17923));
assign g34396 = (g34194&g21337);
assign g29339 = ((~g28274));
assign II18180 = ((~g13605));
assign g23518 = ((~g21070));
assign g33726 = ((~II31581));
assign g33588 = (g33334)|(g18468);
assign g12680 = ((~g9631)&(~g9576));
assign g18194 = (g843&g17821);
assign g21070 = ((~II20937));
assign g14258 = ((~g9203))|((~g11903));
assign g23299 = ((~II22400));
assign g13046 = (g6870&g11270);
assign g21160 = ((~g17508));
assign II26438 = ((~g26549))|((~g14271));
assign g23000 = ((~g20453));
assign g22845 = ((~g20682));
assign g25545 = (g23551)|(g20658);
assign g29219 = ((~II27573));
assign g14845 = ((~g12558))|((~g12798));
assign II31227 = (g32784&g32785&g32786&g32787);
assign g14867 = ((~g10191)&(~g12314));
assign g17773 = ((~g5965))|((~g14549))|((~g5976))|((~g9935));
assign g30112 = (g28566&g20919);
assign II22331 = ((~g19417));
assign g19442 = ((~g11431))|((~g17794));
assign g32986 = (g31996)|(g18280);
assign g23386 = (g20034&g20207);
assign g34229 = ((~g33936));
assign II31087 = (g32580&g32581&g32582&g32583);
assign g18148 = (g562&g17533);
assign g23541 = ((~g21514));
assign g18893 = (g16215&g16030);
assign g15714 = ((~II17228));
assign g17482 = ((~g9523)&(~g14434));
assign II16452 = ((~g11182));
assign g26781 = (g24913)|(g24921);
assign g21611 = ((~II21210));
assign g26313 = (g12645&g25326);
assign g31764 = (g30015)|(g30032);
assign g26236 = (g25357&g6856&g7586&g7558);
assign g27433 = (g26519&g17583);
assign g7995 = ((~g153));
assign g25551 = (g23822&g21511);
assign g14119 = (g10776)|(g8703);
assign g11618 = ((~g8114)&(~g8070));
assign g6983 = ((~g4698));
assign g32696 = ((~g30825));
assign g20231 = ((~g17821));
assign g12194 = ((~g8373))|((~g8273));
assign g33530 = (g32960&II31346&II31347);
assign g25285 = (g22152&g13061);
assign g27480 = (g26400&g17638);
assign g12153 = ((~g2610))|((~g8330));
assign g22494 = ((~g19801));
assign gbuf103 = (g4294);
assign g34881 = (g34866)|(g18187);
assign g30556 = (g30236)|(g22127);
assign II14883 = ((~g9500))|((~g5489));
assign g21935 = (g5196&g18997);
assign g25900 = (g24390&g19368);
assign g17476 = ((~g14665));
assign g16196 = ((~g13496))|((~g13513))|((~g13079))|((~g13476));
assign g25127 = (g13997&g23524);
assign g15903 = (g13796&g13223);
assign g9694 = ((~g1936)&(~g1862));
assign g24402 = (g4749&g22857);
assign g13257 = ((~g1389))|((~g10544));
assign g34414 = (g34206&g21457);
assign g21942 = (g5236&g18997);
assign g21251 = (g13969&g17470);
assign gbuf115 = (g4213);
assign g12553 = ((~g5170)&(~g9206));
assign g20660 = ((~g17873));
assign g23907 = ((~g19074));
assign g26648 = ((~g25115));
assign g20072 = ((~g17384));
assign II26643 = (g27073)|(g27058)|(g27045)|(g27040);
assign g19789 = ((~g17015));
assign g20196 = (g16207)|(g13497);
assign g30991 = ((~II28925));
assign g30438 = (g29890)|(g21847);
assign g27101 = ((~g26770));
assign g31226 = (g30282&g25218);
assign g24916 = ((~g19450))|((~g23154));
assign g12183 = ((~II15033));
assign II31201 = (g31672&g31831&g32745&g32746);
assign g14226 = ((~g11618));
assign g28417 = (g27219)|(g15881);
assign II18341 = ((~g14308));
assign g23520 = ((~g21468));
assign g24855 = (g3050&g23534&II24027);
assign II13852 = ((~g7397))|((~II13850));
assign g11951 = ((~g9166))|((~g847))|((~g703));
assign g34819 = (g34741)|(g34684);
assign g9626 = ((~g6466));
assign g33085 = ((~g31978)&(~g4311));
assign g21727 = ((~II21300));
assign g27204 = (g26026&g16689);
assign g9019 = ((~II12950));
assign g24712 = (g19592&g23001);
assign g23681 = ((~g21012));
assign g28218 = (g27768&g26645);
assign g34939 = ((~g34922));
assign II31607 = ((~g33164));
assign II32868 = ((~g34579));
assign g23361 = ((~II22464));
assign g29041 = ((~II27385));
assign g14110 = ((~g11692))|((~g8906));
assign II20468 = ((~g16663))|((~II20467));
assign g15595 = ((~II17173));
assign g31903 = (g31374)|(g21911);
assign g21830 = (g3774&g20453);
assign g31291 = (g29581)|(g29593);
assign g18630 = (g3689&g17226);
assign g14151 = ((~g11692))|((~g11483));
assign g25735 = (g25077)|(g18783);
assign g23404 = (g20063&g20247);
assign g16127 = ((~g13437));
assign g30474 = (g30208)|(g21945);
assign g34366 = (g26257)|(g34133);
assign g16540 = ((~II17744));
assign II15837 = ((~g1459));
assign g27993 = ((~II26503));
assign g28034 = ((~g26365));
assign II31262 = (g32833&g32834&g32835&g32836);
assign g28667 = (g27410)|(g16616);
assign g34222 = ((~II32195));
assign g9685 = ((~g6533));
assign g16923 = ((~II18089));
assign g32340 = (g31468&g23585);
assign g22708 = (g19266)|(g15711);
assign g18808 = (g6390&g15656);
assign g19587 = (g15700)|(g13046);
assign g34101 = (g33693)|(g33700);
assign g31478 = (g29764&g23410);
assign g24094 = ((~g21143));
assign g26342 = (g8407)|(g24591);
assign g32994 = (g32290)|(g18367);
assign g28530 = (g27383&g20240);
assign g19633 = ((~g16931));
assign g34575 = ((~II32651));
assign g17315 = ((~g9564))|((~g9516))|((~g14503));
assign g20238 = ((~g17096));
assign g24307 = (g4486&g22228);
assign II16217 = ((~g3632));
assign II27539 = (g28040&g24135&g24136&g24137);
assign g20595 = ((~g15877));
assign g34346 = ((~g34162));
assign g16757 = ((~g13911))|((~g13886))|((~g14120))|((~g11675));
assign g34607 = (g34567)|(g15081);
assign g23124 = ((~g8443)&(~g20011));
assign g28476 = ((~g27627)&(~g26547));
assign g30036 = ((~g29085));
assign g32479 = ((~g30735));
assign g30530 = (g30224)|(g22076);
assign g26296 = ((~g8287)&(~g24732));
assign g24750 = (g17662&g22472);
assign g7558 = ((~II12041));
assign g26973 = ((~g26105));
assign g20189 = ((~II20447));
assign g29999 = ((~g28973));
assign g34274 = (g27822)|(g34205);
assign g15104 = (g6955&g14454);
assign g23318 = (g19716)|(g16192);
assign II32231 = ((~g34123));
assign g11534 = ((~g7121))|((~g8958));
assign g8948 = ((~g785));
assign g21388 = ((~g11608))|((~g17157));
assign g27306 = ((~g24787))|((~g26235));
assign g11136 = ((~II14192));
assign g7557 = ((~g1500));
assign g23620 = ((~II22769));
assign g14385 = ((~II16541));
assign g24352 = (g22157)|(g18821);
assign g25660 = (g24726)|(g21785);
assign g12587 = ((~g7497))|((~g6315));
assign g30091 = (g28127&g20716);
assign II22745 = ((~g19458));
assign g32755 = ((~g31672));
assign g32236 = (g31152)|(g29664);
assign g22940 = ((~g18918))|((~g2860));
assign g21669 = ((~II21230));
assign g8571 = ((~g57));
assign g25042 = (g23262&g20496);
assign g25299 = ((~g22763));
assign g26281 = (g24688&g8812&g8778&g8757);
assign g24934 = ((~g21283))|((~g23462));
assign g32129 = (g31658&g29955);
assign g11561 = ((~II14517))|((~II14518));
assign g22758 = ((~g20330));
assign g18330 = (g1668&g17873);
assign g33276 = (g32128)|(g29566);
assign g11975 = ((~g8267))|((~g8316));
assign g26839 = (g2988&g24516);
assign g30379 = (g30089)|(g18491);
assign II16289 = ((~g12107));
assign II13236 = ((~g5452));
assign g30410 = (g29857)|(g21769);
assign II28913 = ((~g30322));
assign g30416 = (g29858)|(g21800);
assign g22073 = (g6235&g19210);
assign g23887 = ((~g18997));
assign g26865 = ((~g25328)&(~g25290));
assign g24227 = (g890&g22594);
assign g27284 = (g9908&g26631);
assign g34026 = (g33715)|(g18682);
assign g32876 = ((~g30735));
assign g13306 = (g441&g11048);
assign g18536 = (g2748&g15277);
assign g29568 = (g2571&g28950);
assign g8530 = (g2902&g2907);
assign g24374 = (g19345)|(g24004);
assign g30419 = (g29759)|(g21803);
assign g32404 = ((~II29936));
assign g21961 = (g5424&g21514);
assign g34423 = ((~g34222));
assign g28370 = ((~g27528));
assign gbuf6 = (g4414);
assign g19505 = ((~g16349));
assign II16606 = ((~g3649));
assign g33408 = (g32358&g21407);
assign g31827 = ((~g29385));
assign g22905 = ((~II22114));
assign g22716 = ((~g19795));
assign g33032 = (g32326)|(g21842);
assign g23462 = ((~II22589));
assign g10200 = ((~g2138));
assign g32240 = (g24757)|(g31182);
assign g24346 = (g23725)|(g18789);
assign g27137 = (g26026&g16606);
assign g28360 = (g27401&g19861);
assign g34035 = (g33721)|(g18714);
assign g34086 = (g20114&g33766&g9104);
assign g32321 = (g27613&g31376);
assign g26278 = (g24545)|(g24549);
assign g6874 = ((~g3143));
assign g24786 = (g661&g23654);
assign II16401 = ((~g869));
assign g20923 = ((~g15277));
assign g19773 = ((~g17615));
assign II16468 = ((~g12760));
assign g12738 = ((~g9374));
assign g14124 = ((~g8830)&(~g11083));
assign g26915 = (g25900)|(g18230);
assign g28623 = (g27361)|(g16520);
assign II15590 = ((~g11988));
assign g9640 = ((~g1802)&(~g1728));
assign g34911 = (g34909)|(g18188);
assign g28401 = (g27212)|(g15871);
assign II23363 = ((~g23385));
assign II31206 = (g31710&g31832&g32752&g32753);
assign g25778 = ((~g25459)&(~g25420));
assign II25555 = ((~g25241));
assign g9467 = ((~g6434));
assign g20583 = ((~g17873));
assign g8125 = ((~g3869));
assign g32223 = (g31142)|(g29637);
assign g23608 = ((~g21611));
assign g29843 = (g28373&g23289);
assign g27723 = (g26512&g21049);
assign g22639 = (g18950)|(g15612);
assign g32385 = (g31480)|(g29938);
assign g26912 = (g25946)|(g18209);
assign g31519 = (g29864&g23490);
assign g29598 = (g28823&g22342);
assign g32764 = ((~g30937));
assign g10874 = (g7791&g6219&g6227);
assign g7617 = ((~II12089));
assign g10665 = (g209&g8292);
assign g29365 = ((~g29067));
assign g25659 = (g24707)|(g21784);
assign g33059 = (g31987)|(g22021);
assign g14953 = ((~g12646))|((~g12405));
assign g10733 = (g3639&g6905&g3625&g8542);
assign II21230 = ((~g16540));
assign g10759 = ((~g7537))|((~g324));
assign g16897 = ((~II18083));
assign g17759 = ((~g14864));
assign g11473 = ((~g8107)&(~g8059));
assign II31167 = (g32696&g32697&g32698&g32699);
assign g25189 = ((~g6082)&(~g23726));
assign g29800 = ((~g28363));
assign g32936 = ((~g31710));
assign g32306 = (g31289&g23499);
assign g33698 = ((~II31539));
assign g9815 = ((~g6098));
assign g24030 = ((~g21127));
assign g31182 = (g30240&g20682);
assign g17291 = ((~II18276));
assign g27379 = ((~g8492)&(~g26636));
assign g24636 = ((~g23121));
assign II11617 = ((~g1));
assign g29903 = ((~g6928)&(~g28484));
assign g12207 = ((~g9887))|((~g5794));
assign g19265 = ((~g15721))|((~g15715))|((~g13091))|((~g15710));
assign g27587 = ((~g24917))|((~g25018))|((~g24918))|((~g26857));
assign II32837 = ((~g34498));
assign g29585 = (g1756&g28920);
assign g24423 = (g4950&g22897);
assign g33912 = ((~II31770));
assign gbuf16 = (g5290);
assign g24087 = ((~g21143));
assign g18061 = ((~g14800));
assign II30717 = (g31787)|(g32200)|(g31940)|(g31949);
assign g27041 = (g8519&g26330);
assign II18526 = ((~g13055));
assign II14079 = ((~g7231));
assign g27274 = (g15779)|(g25915);
assign g20915 = ((~II20882));
assign g27552 = (g26092)|(g24676);
assign g18584 = (g2950&g16349);
assign II17476 = ((~g1105))|((~II17474));
assign g14411 = ((~g9460)&(~g11160));
assign g21923 = (g5029&g21468);
assign g14723 = ((~g7704))|((~g12772));
assign g27440 = (g8046&g26314&g518&g504);
assign g30613 = ((~g4507)&(~g29365));
assign g10934 = (g9197&g7918);
assign g6836 = ((~g1322));
assign g32654 = ((~g31070));
assign g8591 = ((~g3763));
assign II22938 = ((~g21228))|((~II22936));
assign II12878 = ((~g4180))|((~II12876));
assign g24866 = ((~II24038));
assign g24686 = (g5485&g23630);
assign g34303 = (g25768)|(g34045);
assign II24689 = (g20841&g24040&g24041&g24042);
assign g32503 = ((~g31194));
assign g17509 = ((~II18446));
assign g18105 = (g417&g17015);
assign g12591 = ((~g504)&(~g9040));
assign g34090 = (g33676)|(g33680);
assign g26965 = (g26336)|(g24317);
assign g25851 = ((~g4311)&(~g24380)&(~g24369));
assign g25982 = (g2351&g25008);
assign II18682 = ((~g14752))|((~II18680));
assign g23590 = ((~g20682))|((~g11111));
assign g30307 = (g28256)|(g27260);
assign g30170 = ((~g28846)&(~g14615));
assign g29600 = (g1840&g29049);
assign g21424 = ((~g15426));
assign g20274 = ((~g17847));
assign g29506 = (g28148)|(g25880);
assign g19276 = ((~g17367));
assign g23321 = ((~II22422));
assign g12413 = ((~g7521))|((~g5654));
assign g30139 = (g28596&g21184);
assign g12066 = ((~II14924))|((~II14925));
assign II22754 = ((~g11937))|((~II22753));
assign g32718 = ((~g30825));
assign g9380 = ((~g5471));
assign g29384 = (g26424&g22763&g28179);
assign g12762 = (g4358&g8977);
assign g29752 = (g28516&g10233);
assign g31287 = (g29578)|(g28292);
assign g10820 = ((~g9985))|((~g9920))|((~g9843));
assign g29977 = ((~g28920));
assign g11223 = (g8281&g8505);
assign II17447 = ((~g13336))|((~II17446));
assign g27019 = (g26822)|(g14610);
assign g25206 = ((~g23613));
assign g29271 = (g28333)|(g18637);
assign g31745 = (g29959)|(g29973);
assign g34847 = ((~II33067));
assign g20916 = ((~g18008));
assign g18488 = (g2495&g15426);
assign g22020 = (g5863&g19147);
assign g24202 = (g22899)|(g18106);
assign g11705 = ((~II14576));
assign g21185 = ((~g15277));
assign g23067 = ((~g20887))|((~g10721));
assign g33160 = ((~g8672)&(~g32057));
assign g28489 = (g27010&g12417);
assign g27350 = (g10217&g26803);
assign II30992 = ((~g32445));
assign g12333 = ((~g1624)&(~g8139));
assign g9778 = ((~g5069));
assign g24311 = (g4498&g22228);
assign g28914 = ((~g27937))|((~g7462))|((~g2555));
assign g9568 = ((~g6181));
assign g30368 = (g30098)|(g18435);
assign II31097 = (g32596&g32597&g32598&g32599);
assign II32431 = ((~g34056))|((~g34051));
assign g17611 = ((~g14822));
assign g11772 = ((~II14623));
assign g27877 = ((~g9397)&(~g25839));
assign g33187 = (g32014)|(II30740)|(II30741);
assign g24417 = ((~g22171));
assign g25973 = (g2342&g24994);
assign g30116 = ((~II28349));
assign g20709 = ((~g15426));
assign II24461 = ((~g23796))|((~g14437));
assign g15572 = ((~g12969))|((~g7219));
assign g20203 = (g6195&g17789);
assign g20773 = ((~II20830));
assign II30959 = ((~g32021));
assign g24197 = (g347&g22722);
assign II12749 = ((~g4575));
assign g32823 = ((~g31327));
assign g32147 = (g31616&g29980);
assign g34992 = ((~II33276));
assign g26273 = (g2122&g25389);
assign g20654 = ((~II20750));
assign g27767 = ((~II26367))|((~II26368));
assign g24709 = (g16690&g23000);
assign g29231 = (g28301)|(g18229);
assign g34570 = ((~g34392));
assign g23493 = ((~g21611));
assign g30522 = (g29332)|(g22064);
assign II32203 = ((~g33937))|((~II32202));
assign II12811 = ((~g4340));
assign g29208 = (g24138&II27538&II27539);
assign II28419 = ((~g29195));
assign II11623 = ((~g28));
assign g7717 = ((~II12172));
assign II26309 = ((~g26825));
assign II24839 = ((~g24298));
assign g32155 = (g30935)|(g29475);
assign II25105 = ((~g25284));
assign g10487 = ((~g10233));
assign g29533 = (g28958&g22417);
assign g32518 = ((~g30614));
assign g33433 = (g32238&g29694);
assign g25961 = (g25199&g20682);
assign g14832 = (g1489&g10939);
assign g22059 = (g6148&g21611);
assign g23302 = ((~g20330));
assign g16161 = (g5841&g14297);
assign g18274 = (g1311&g16031);
assign g13057 = ((~g969))|((~g11294));
assign g34203 = (g33726&g24537);
assign g15705 = ((~g13217));
assign g24291 = (g18660&g22550);
assign II24038 = ((~g22202));
assign g10143 = ((~g568));
assign g29194 = ((~II27492));
assign II14213 = ((~g9295))|((~II14211));
assign g10707 = (g3787&g8561);
assign g11165 = ((~II14222));
assign II17814 = ((~g3274));
assign g18702 = (g15133&g16856);
assign g18359 = (g1825&g17955);
assign g29750 = (g28296&g23215);
assign g23397 = (g11154&g20239);
assign g34097 = (g33772&g9104&g18957);
assign g23924 = ((~g18997));
assign g28085 = (g27263)|(g18700);
assign g25764 = (g25551)|(g18819);
assign II32243 = ((~g34134));
assign II31047 = (g32524&g32525&g32526&g32527);
assign g27223 = ((~II25908))|((~II25909));
assign g28246 = (g8572&g27976);
assign g15110 = (g4245&g14454);
assign g24792 = ((~II23950))|((~II23951));
assign g15483 = ((~II17128));
assign g30573 = ((~g29355))|((~g19666));
assign g17646 = ((~II18609));
assign g29988 = (g29187&g12235);
assign g18883 = ((~g15938));
assign g28084 = (g27254)|(g18698);
assign II18485 = ((~g1677))|((~g14611));
assign g18554 = (g2831&g15277);
assign g22536 = ((~g1379)&(~g19720));
assign g32069 = (g10878&g30735);
assign g19610 = (g1141&g16069);
assign g9239 = ((~g5511));
assign g16745 = ((~g3594))|((~g13730))|((~g3661))|((~g11389));
assign g27353 = ((~g8097)&(~g26616));
assign g11969 = ((~g7252))|((~g1636));
assign g17768 = (g13325&g10741);
assign g35000 = (g34953)|(g34999);
assign g28931 = ((~g27886))|((~g2070))|((~g1996));
assign II15306 = ((~g10116))|((~g2407));
assign g12317 = ((~g10026))|((~g6486));
assign g17420 = ((~g9456)&(~g14408));
assign g9461 = ((~II13140))|((~II13141));
assign g24467 = (g13761&g23047);
assign g24268 = (g23025)|(g18612);
assign g20008 = ((~g16449));
assign g20499 = ((~g15483));
assign g23764 = ((~g21308));
assign g21139 = ((~g15634));
assign g12968 = ((~g11793));
assign g23426 = ((~II22539));
assign g20504 = ((~g18008));
assign g20147 = ((~g17328));
assign g21815 = (g3598&g20924);
assign g20067 = ((~g17328));
assign g25548 = ((~g22550));
assign g16286 = ((~II17615));
assign g17326 = ((~II18307));
assign g33652 = (g33393&g18889);
assign g28708 = (g27462)|(g16674);
assign g30173 = (g28118&g13082);
assign g28638 = (g27551&g20583);
assign II15448 = ((~g10877));
assign g21853 = (g3917&g21070);
assign gbuf88 = (g3672);
assign g27087 = (g13872&g26284);
assign II14955 = ((~g9620))|((~g6181));
assign g21885 = (g4122&g19801);
assign g26299 = (g24551)|(g22665);
assign g24318 = (g4555&g22228);
assign II16391 = ((~g859));
assign g9483 = (g1008)|(g969);
assign gbuf69 = (g6490);
assign g28576 = (g27325)|(g26271);
assign g25507 = (g6098&g23844&II24616);
assign g21756 = (g3211&g20785);
assign g29374 = ((~II27742));
assign gbuf90 = (g3443);
assign g7880 = ((~g1291));
assign g25435 = ((~g22432))|((~g2342))|((~g8316));
assign II31864 = (g33510)|(g33511)|(g33512)|(g33513);
assign gbuf13 = (g4812);
assign g34840 = ((~II33056));
assign II18460 = ((~g5276));
assign g15154 = ((~g13782)&(~g12898));
assign g10084 = ((~g2837));
assign g32890 = ((~g30735));
assign II26466 = ((~g26870));
assign g21698 = ((~g18562));
assign II24018 = (g8155&g8390&g3396);
assign g34654 = ((~II32766));
assign g30567 = ((~g29930));
assign g32486 = ((~g30735));
assign g31115 = (g29487&g22882);
assign g18156 = (g572&g17533);
assign g14448 = ((~g12192)&(~g9699));
assign II18785 = (g13156&g6767&g11498);
assign g30313 = ((~g28843));
assign g28127 = ((~g27102));
assign g24116 = ((~g21143));
assign g16206 = ((~g13437));
assign g34874 = (g34833&g20060);
assign g22007 = (g5770&g21562);
assign g21771 = (g3255&g20785);
assign g7322 = ((~g1862));
assign g13060 = (g8587&g11110);
assign g10572 = ((~g10233));
assign g25741 = (g25178)|(g22056);
assign g26052 = ((~g22714))|((~g24662))|((~g22921));
assign g30516 = (g30233)|(g22037);
assign g7564 = ((~g336));
assign g23937 = ((~g19277));
assign g29323 = (g28539&g6905&g3639);
assign II11655 = ((~g1246));
assign g18591 = (g2965&g16349);
assign g30218 = ((~g28918));
assign g22369 = (g9354&g7717&g20783);
assign g20104 = ((~g17433));
assign g32531 = ((~g31070));
assign g26512 = (g24786)|(g23130);
assign g22667 = ((~g21156));
assign g18627 = (g15093&g17093);
assign g33039 = (g32187)|(g24312);
assign II15166 = ((~g9904))|((~g9823));
assign g24161 = ((~II23327));
assign g8608 = ((~g278));
assign g25259 = ((~II24445));
assign g34791 = (g34771)|(g18184);
assign g14314 = ((~II16476));
assign II13094 = ((~g2724));
assign g18751 = (g5156&g17847);
assign g23606 = (g16927&g20679);
assign g21706 = (g222&g20283);
assign g9744 = ((~g6486));
assign g20702 = ((~g17955));
assign g23390 = ((~g21468));
assign g24102 = ((~g21143));
assign g25652 = (g24777)|(g21747);
assign g15753 = ((~g6239))|((~g14529))|((~g6351))|((~g10003));
assign g25917 = (g22524)|(g24518);
assign g23576 = ((~II22718))|((~II22719));
assign g29524 = (g2004&g28864);
assign g34431 = ((~II32464));
assign g32625 = ((~g31070));
assign g29878 = ((~g28421));
assign g15884 = (g3901&g14113);
assign g18933 = (g16237&g13597);
assign g11468 = ((~g7624));
assign g34585 = (g24705&g34316);
assign g19714 = ((~g16821));
assign g32875 = ((~g31376));
assign g21400 = ((~g17847));
assign g31910 = (g31471)|(g21957);
assign g16303 = (g4527&g12921);
assign g10803 = ((~g1384)&(~g7503));
assign II31504 = ((~g33164));
assign g23255 = (g19655)|(g16122);
assign g7805 = ((~g4366));
assign g9663 = ((~g128))|((~g4646));
assign II31322 = (g32921&g32922&g32923&g32924);
assign g12087 = ((~g7431))|((~g2599));
assign g23599 = (g19050&g9104);
assign g8769 = ((~g691))|((~g714));
assign g16615 = ((~II17801));
assign g21801 = (g3554&g20924);
assign g24339 = (g23690)|(g18756);
assign g34009 = (g33863)|(g18477);
assign II15287 = ((~g10061))|((~g6697));
assign g29647 = (g28934&g22457);
assign g16591 = (g5256&g14879);
assign g26843 = ((~II25567));
assign II18293 = ((~g1079));
assign g34732 = (g34686)|(g18593);
assign g34317 = ((~g34115));
assign g24995 = ((~g22763));
assign g24203 = (g22982)|(g18107);
assign g12640 = ((~II15382));
assign II26522 = (g19890)|(g19935)|(g19984)|(g26365);
assign g28673 = (g1373&g27122);
assign g21958 = (g5396&g21514);
assign g30920 = (g29889&g21024);
assign II18875 = ((~g13782));
assign II31172 = (g32703&g32704&g32705&g32706);
assign g14637 = ((~g12255))|((~g9815));
assign g30145 = (g28603&g21247);
assign g9761 = ((~g2445));
assign g6990 = ((~g4742));
assign II13497 = ((~g255))|((~g232));
assign II29969 = ((~g30991));
assign g19068 = ((~g16031));
assign g13580 = ((~g11849))|((~g7503))|((~g7922))|((~g10544));
assign g10622 = ((~g10178))|((~g9973));
assign g26181 = (g2652&g25157);
assign g18130 = (g528&g16971);
assign g7933 = ((~g907));
assign II31555 = ((~g33212));
assign II32103 = ((~g33661));
assign g12118 = ((~g8259))|((~g8150));
assign g27954 = ((~g10014)&(~g25856));
assign g23374 = (g19767)|(g13514);
assign g17504 = ((~g15021));
assign g7267 = ((~g1604));
assign g13522 = ((~g10981));
assign g13283 = ((~g12440))|((~g12399))|((~g9843));
assign g8733 = ((~g3698));
assign g13288 = ((~g10946))|((~g1442));
assign g16729 = (g5240&g14720);
assign g27210 = (g26218&g8373&g2476);
assign II24393 = ((~g23453));
assign g28504 = ((~g758))|((~g27528))|((~g11679));
assign g34715 = (g34570&g33375);
assign g20634 = ((~g15373));
assign g20432 = ((~g17847));
assign g17789 = ((~g14321));
assign g29981 = ((~g28942));
assign g34181 = ((~g33913));
assign II24546 = (g5046&g5052&g9716);
assign g28604 = ((~g27759));
assign g25025 = ((~g22498));
assign II11824 = ((~g4593))|((~g4601));
assign g9960 = ((~g6474));
assign g14583 = (g10685)|(g542);
assign II12176 = ((~g5523));
assign g27224 = (g25870)|(g15678);
assign II31463 = ((~g33318));
assign g31009 = ((~g27187))|((~g29503))|((~g19644));
assign g27563 = (g26104)|(g24704);
assign g34559 = ((~g34384));
assign g33548 = (g33327)|(g18336);
assign g10411 = ((~g7086));
assign g28780 = ((~g27742))|((~g7308))|((~g1636));
assign g20037 = ((~g17328));
assign g8218 = ((~g3490));
assign g15612 = (g3143&g13530);
assign g13036 = ((~g10981));
assign g32194 = (g30601&g28436);
assign g20714 = ((~g15277));
assign II17128 = ((~g13835));
assign g28329 = (g27128)|(g15813);
assign g22760 = (g9360&g20237);
assign II18700 = ((~g6027));
assign II12092 = ((~g790));
assign g34096 = (g22957&g9104&g33772);
assign II19818 = ((~g1056));
assign g22849 = (g1227&g19653);
assign g15805 = (g3243&g14041);
assign g13932 = ((~g11534));
assign g33509 = (g32809&II31241&II31242);
assign II24228 = ((~g22409));
assign g10352 = ((~g6804));
assign g32263 = (g31631&g30306);
assign II27349 = (g25534&g26424&g22698);
assign g18561 = (g2841&g15277);
assign g33014 = (g32305)|(g18499);
assign g18145 = (g582&g17533);
assign g24383 = ((~g22409)&(~g22360));
assign II17425 = ((~g13416));
assign g29893 = ((~g28755));
assign g21379 = ((~g17873));
assign g7624 = ((~II12106));
assign g23305 = ((~g20391));
assign g12919 = ((~II15536));
assign g18460 = (g2351&g15224);
assign II12074 = ((~g996))|((~g979));
assign g30162 = ((~g28880)&(~g7462));
assign g33354 = ((~g32329));
assign g15717 = ((~g10754))|((~g13092));
assign g22357 = ((~g1024)&(~g19699));
assign g26148 = (g25357&g11724&g11709&g11686);
assign g24646 = (g22640&g19711);
assign g12036 = ((~g9245));
assign g28852 = (g27559)|(g16871);
assign g24134 = ((~g19984));
assign g21278 = ((~II21013));
assign g29001 = ((~g27937))|((~g2599))|((~g7431));
assign II18518 = ((~g13835));
assign g23188 = (g13994&g20025);
assign g30318 = ((~g28274));
assign II24022 = ((~g22182));
assign g17602 = ((~g14962));
assign g26336 = (g10307&g25480);
assign g20606 = ((~g17955));
assign g30548 = (g30204)|(g22119);
assign g14419 = ((~g12152)&(~g9546));
assign g32800 = ((~g31021));
assign II23351 = ((~g23263));
assign g25867 = (g25449)|(g23884);
assign g34742 = (g9000&g34698);
assign g22101 = (g6474&g18833);
assign g28593 = ((~g27727));
assign g22136 = ((~g20277));
assign II16626 = ((~g11986));
assign g34927 = ((~II33173));
assign g28645 = (g27556&g20599);
assign g34335 = (g8461&g34197);
assign g32560 = ((~g31070));
assign g34590 = ((~II32678));
assign g33313 = (g29649)|(g32171);
assign g24549 = (g23162&g20887);
assign g8229 = ((~g3881));
assign g22014 = (g5805&g21562);
assign g24668 = (g11754&g22979);
assign g14176 = ((~g9044)&(~g12259));
assign g31835 = ((~g29385));
assign g24077 = ((~g20720));
assign g12358 = ((~g10019)&(~g10022));
assign g22305 = ((~g19801));
assign g31143 = (g29506&g22999);
assign g32647 = ((~g31154));
assign g6999 = ((~g86));
assign g17191 = (g1384&g13242);
assign g30917 = ((~II28897));
assign II31001 = (g29385&g32456&g32457&g32458);
assign g16699 = (g7134&g12933);
assign g28093 = (g27981)|(g21951);
assign g31638 = ((~g29689));
assign g21682 = ((~g16540));
assign g17086 = ((~g14297));
assign g10387 = ((~g6996));
assign g23250 = ((~g21070));
assign II31622 = ((~g33204));
assign g13634 = ((~g11797))|((~g11261));
assign II22946 = ((~g19620))|((~II22944));
assign g20014 = ((~g17096)&(~g11244));
assign g21787 = (g15091&g20391);
assign II13520 = ((~g2518))|((~II13518));
assign II23969 = ((~g22202))|((~g490));
assign g20443 = ((~g15171));
assign g27494 = (g8038&g26314&g518&g9077);
assign II33258 = ((~g34976));
assign g15589 = (g411&g13334);
assign g11355 = ((~g9551))|((~g3310));
assign g11679 = ((~g8836))|((~g802));
assign g32687 = ((~g31376));
assign g22854 = ((~g20330));
assign g14912 = ((~II16917));
assign g13527 = ((~g182))|((~g168))|((~g203))|((~g12812));
assign g28233 = (g27827&g23411);
assign g12467 = ((~g9472)&(~g9407));
assign g18446 = (g2279&g18008);
assign g33466 = (g32498&II31026&II31027);
assign g15080 = (g12855&g12983);
assign g31882 = (g31115)|(g21776);
assign g14677 = ((~II16779))|((~II16780));
assign g33338 = (g32220&g20633);
assign g11450 = ((~II14455));
assign g20552 = ((~g17847));
assign g21409 = ((~g18008));
assign g34558 = (g34353&g20578);
assign g31068 = ((~g4801)&(~g29540));
assign g34118 = ((~II32051));
assign g15087 = ((~g12860)&(~g13144));
assign g7516 = ((~II12003));
assign II18238 = ((~g13144));
assign g33255 = (g32106)|(g29514);
assign g16000 = ((~II17425));
assign g22207 = ((~II21787));
assign g16598 = (g6283&g14899);
assign g24215 = (g23484)|(g18196);
assign g18705 = (g4801&g16782);
assign g27658 = (g22491&g25786);
assign g25186 = ((~g5396))|((~g23602));
assign g10795 = ((~g7202));
assign g23191 = ((~II22289));
assign g29787 = (g28334&g23249);
assign II17612 = ((~g13250));
assign g8725 = ((~g739));
assign g16691 = ((~g14160));
assign g14610 = (g1484&g10935);
assign g13570 = (g9223)|(g11130);
assign II15893 = ((~g10430));
assign g14566 = (g10566&g10551);
assign g23897 = ((~g19210));
assign g28549 = (g27304)|(g26233);
assign g26360 = (g10589&g25533);
assign g34801 = (g34756)|(g18588);
assign g32179 = (g31748&g27907);
assign g9792 = ((~g5401));
assign g33135 = ((~g32090)&(~g8350));
assign II22760 = ((~g11939))|((~g21434));
assign g18609 = (g3147&g16987);
assign g25367 = (g6946&g22407);
assign g20010 = ((~g17226));
assign g12911 = (g10278)|(g12768);
assign g25466 = (g23574&g21346);
assign g8070 = ((~g3518));
assign g17124 = ((~g14051));
assign g24348 = (g22149)|(g18804);
assign g13349 = (g4933&g11780);
assign g26898 = (g26387)|(g18194);
assign g8404 = ((~g5005));
assign g15782 = ((~g6585))|((~g14556))|((~g6697))|((~g10061));
assign g32733 = ((~g31672));
assign g24214 = (g23471)|(g18195);
assign g9688 = ((~g113));
assign g30199 = (g28664&g23861);
assign gbuf153 = (g1056);
assign g9729 = ((~g5138));
assign g25888 = ((~g914))|((~g24439));
assign g22409 = ((~II21860));
assign g23015 = ((~g20391));
assign II24075 = (g3736&g3742&g8553);
assign II29214 = ((~g30300));
assign g14987 = ((~g6593))|((~g12211))|((~g6692))|((~g12721));
assign g33720 = (g33161&g19439);
assign g10150 = ((~g1700));
assign g19962 = ((~g11470))|((~g17794));
assign g21295 = ((~g17533));
assign g33061 = (g32334)|(g22050);
assign g24680 = (g16422&g22986);
assign g16234 = (g6772&g6782&g11640&II17575);
assign g24452 = ((~g22722));
assign g21430 = ((~g15608));
assign g14217 = ((~II16417));
assign g8841 = ((~II12823));
assign g13883 = ((~g4709)&(~g4785)&(~g11155));
assign g8848 = ((~g358));
assign g27262 = (g25997&g17092);
assign g18905 = ((~g16077));
assign g14719 = (g4392&g10830);
assign g25078 = (g23298&g20538);
assign g22035 = (g5933&g19147);
assign g34562 = (g34369&g17411);
assign g11990 = ((~g9166))|((~g703));
assign g26851 = ((~II25579));
assign g33557 = (g33331)|(g18363);
assign g15818 = (g3941&g14082);
assign g21994 = (g5607&g19074);
assign g17121 = ((~g14321));
assign II23756 = (g23457)|(g23480)|(g23494)|(g23511);
assign g14035 = (g699&g11048);
assign g14248 = ((~g6065)&(~g10578));
assign g34969 = (g34960&g19570);
assign g20513 = ((~g18065));
assign g20326 = ((~g18008));
assign g18248 = (g15067&g16897);
assign g28263 = (g23747&g27711);
assign g22146 = ((~g18997));
assign g16231 = ((~g13515)&(~g4771));
assign g31856 = ((~g29385));
assign g16514 = ((~g14139));
assign g24505 = ((~g22689));
assign g32255 = (g31248&g20381);
assign g28541 = (g27403&g20274);
assign g12296 = ((~g9860)&(~g9862));
assign g12462 = ((~g7051))|((~g7064))|((~g10190));
assign gbuf70 = (g3303);
assign g27217 = (g26236&g8418&g2610);
assign g13342 = ((~g10961)&(~g10935));
assign II12227 = ((~g34));
assign g23355 = ((~g21070));
assign g18513 = (g2575&g15509);
assign g21701 = (g153&g20283);
assign g31988 = (g31768&g22199);
assign g30078 = (g28526&g20667);
assign g30066 = (g28518&g20636);
assign g30003 = (g28149&g9021);
assign g30457 = (g29369)|(g21885);
assign g32898 = ((~g30825));
assign g29379 = ((~II27749));
assign g29839 = (g1728&g29045);
assign g24679 = (g13289&g22985);
assign g23439 = (g13771&g20452);
assign g27463 = ((~g287))|((~g26330))|((~g23204));
assign g17325 = ((~II18304));
assign g28386 = (g27202)|(g13277);
assign g34051 = ((~II31973))|((~II31974));
assign g28710 = (g27589&g20703);
assign g33963 = (g33830)|(g18124);
assign g25245 = ((~g22763));
assign II24527 = (g9672&g9264&g5401);
assign g32880 = ((~g30614));
assign g10357 = ((~g6825));
assign g32362 = (g29870)|(g31301);
assign g10179 = ((~g2098)&(~g1964)&(~g1830)&(~g1696));
assign g28666 = (g27567&g20625);
assign II28002 = ((~g28153));
assign g30183 = ((~g28880)&(~g14644));
assign g20451 = ((~g15277));
assign g9907 = ((~g1959));
assign g25170 = ((~g22498));
assign g34948 = (g16540&g34935);
assign g28130 = (g27353&g23063);
assign g22897 = ((~g21024));
assign g15651 = (g429&g13414);
assign g13794 = (g7396)|(g10684);
assign g21985 = (g5571&g19074);
assign g33057 = (g31968)|(g22019);
assign g24651 = (g2741&g23472);
assign g18315 = (g1548&g16931);
assign g23341 = ((~g21163));
assign g10917 = (g9174&g1087);
assign g13793 = ((~II16120));
assign g33519 = (g32881&II31291&II31292);
assign g26155 = (g1945&g25134);
assign g29214 = ((~II27558));
assign II17658 = ((~g13394));
assign g32012 = (g8297&g31233);
assign g19948 = (g17515&g16320);
assign g27510 = (g26576&g17687);
assign g17676 = ((~g12941));
assign g18062 = ((~II18872));
assign g30590 = (g18911&g29812);
assign g25759 = (g25166)|(g22106);
assign g17415 = ((~g14797));
assign g10042 = ((~g2671));
assign g24517 = (g22158)|(g18906);
assign g34511 = ((~g34419));
assign g14555 = (g12521&g12356&g12307&II16671);
assign II18221 = ((~g13605));
assign g27116 = (g26026&g16527);
assign g13431 = ((~II15932));
assign g12772 = ((~g5188)&(~g9300));
assign g14089 = ((~g11755))|((~g4717));
assign g19585 = (g17180&g14004);
assign g32576 = ((~g30614));
assign g7763 = (g2965&g2960);
assign g14851 = ((~g7738))|((~g12505));
assign g27773 = ((~II26378));
assign g15072 = ((~g13416)&(~g12843));
assign g19781 = ((~g16489));
assign g15722 = (g464&g13437);
assign g30357 = (g30107)|(g18366);
assign g28519 = ((~g8011)&(~g27602)&(~g10295));
assign g11249 = ((~g8405));
assign g34375 = (g13077&g34049);
assign g33031 = (g32315)|(g21841);
assign g29810 = (g28259&g11317);
assign g30141 = (g28499)|(g16844);
assign g28010 = (g23032&g26223&g26424&g25535);
assign g28871 = ((~g27858))|((~g7418))|((~g2331));
assign g34426 = ((~II32449));
assign II31317 = (g32914&g32915&g32916&g32917);
assign g18235 = (g1141&g16326);
assign g7352 = ((~g1526)&(~g1514));
assign g25716 = (g25088)|(g21967);
assign g18980 = ((~g16136));
assign g24884 = (g3401&g23555&II24051);
assign g7314 = ((~g1740));
assign g13971 = ((~g8938)&(~g4975)&(~g11173));
assign g16869 = (g6259&g14902);
assign g12811 = ((~g10319));
assign g10571 = ((~g10233));
assign II33020 = ((~g34781));
assign g18219 = (g969&g16100);
assign g34859 = (g16540&g34820);
assign g33358 = (g32249&g20778);
assign II23366 = ((~g23321));
assign g34506 = (g8833&g34354);
assign g25966 = (g9364&g24985);
assign g29477 = (g14090&g28441);
assign g7867 = ((~g1489));
assign g31242 = (g29373&g25409);
assign g10666 = ((~g8462)&(~g1171));
assign g33981 = (g33856)|(g18371);
assign g18567 = (g2894&g16349);
assign g33847 = (g33260&g20383);
assign g26123 = (g1696&g25382);
assign g7696 = (g2955&g2950);
assign g10561 = ((~g7157))|((~g5712));
assign g16427 = (g5216&g14876);
assign g11325 = ((~g7543));
assign g31829 = ((~g29385));
assign g8728 = ((~g3618))|((~g3661))|((~g3632))|((~g3654));
assign g16774 = ((~g14024));
assign g17585 = ((~g14974));
assign g10998 = (g8567&g8509&g8451&g7650);
assign g33256 = (g32107)|(g29517);
assign g15693 = (g269&g13474);
assign g9715 = ((~g5011))|((~g4836));
assign g20696 = ((~g17533));
assign g24587 = ((~g23112));
assign g8403 = ((~II12568));
assign g28261 = (g27878&g23695);
assign g16724 = ((~g14079));
assign g17473 = ((~g14841));
assign g13101 = ((~II15736));
assign g13593 = ((~g10556));
assign g19398 = ((~g16489));
assign g18747 = (g5138&g17847);
assign g28510 = ((~g3530)&(~g27617));
assign II32297 = ((~g34059));
assign g13140 = ((~g10632));
assign g33448 = ((~g7785)&(~g31950));
assign gbuf71 = (g3281);
assign g13604 = (g4495&g10487);
assign g28256 = (g11398&g27984);
assign g31879 = (g31475)|(g21745);
assign g19337 = (g17770)|(g17785);
assign II15106 = ((~g9780))|((~II15105));
assign g33525 = (g32925&II31321&II31322);
assign g20083 = (g2902)|(g17058);
assign g28077 = (g27120)|(g21879);
assign II14862 = ((~g8092));
assign II18832 = ((~g13782));
assign g7073 = ((~g6191));
assign g21804 = (g3542&g20924);
assign g11424 = ((~g9662))|((~g4012));
assign II22929 = ((~g12223))|((~g21228));
assign II16829 = ((~g6715));
assign g20776 = ((~g18008));
assign g34983 = ((~II33249));
assign II12144 = ((~g554));
assign g12085 = ((~g10082)&(~g9700));
assign II27271 = ((~g27998));
assign g7192 = ((~g6444)&(~g6404));
assign g13928 = ((~g3562))|((~g11238))|((~g3680))|((~g11576));
assign g29844 = (g28374&g23290);
assign g28266 = (g23748&g27714);
assign g13662 = (g10896)|(g10917);
assign g29762 = (g28298&g10233);
assign II12954 = ((~g4358));
assign g22839 = ((~g20114))|((~g2988));
assign g10176 = ((~g44));
assign g19491 = ((~g16349));
assign II12907 = ((~g4322));
assign g34887 = (g34865)|(g21670);
assign g26381 = (g4456&g25548);
assign g24944 = ((~g21354))|((~g23363));
assign g13700 = ((~g3288)&(~g11615));
assign g31526 = (g22521&g29342);
assign g29611 = (g28540&g14209);
assign g34617 = (g34526)|(g18579);
assign II12109 = ((~g749));
assign g12256 = ((~g10136)&(~g6105));
assign g28523 = (g27704&g15585);
assign g22213 = ((~g19147));
assign g8112 = ((~g3419));
assign g28721 = (g27488)|(g16705);
assign g29225 = (g28451)|(g18158);
assign g31120 = (g1700&g29976);
assign g34348 = (g34125&g20128);
assign g31964 = (g31654)|(g14544);
assign g32723 = ((~g31327));
assign g34007 = (g33640)|(g18467);
assign g19498 = ((~g16752));
assign g12173 = ((~g10050)&(~g7074));
assign g16200 = ((~g13584));
assign g13846 = ((~g1116))|((~g10649));
assign g19979 = ((~g17226));
assign g33716 = ((~II31569));
assign g7626 = ((~II12112));
assign g16424 = ((~g8064)&(~g13628));
assign g30599 = (g18911&g29863);
assign g30369 = (g30066)|(g18439);
assign g33508 = (g32802&II31236&II31237);
assign II17704 = ((~g13144));
assign g19947 = ((~g17226));
assign g34964 = (g34947&g23060);
assign g22132 = (g6645&g19277);
assign g26324 = (g2661&g25439);
assign g33693 = (g33145&g13594);
assign g20616 = ((~g15277));
assign g31798 = ((~g29385));
assign II14291 = ((~g3835))|((~II14289));
assign g19744 = ((~g15885));
assign g18760 = (g5462&g17929);
assign g30543 = (g29338)|(g22110);
assign g7523 = ((~g305));
assign g31127 = ((~g4966)&(~g29556));
assign g18220 = (g1002&g16100);
assign II15250 = ((~g9152));
assign g23882 = ((~g19277));
assign g32109 = (g31609&g29920);
assign g18792 = (g7051&g15634);
assign g26916 = (g25916)|(g18232);
assign g28671 = (g27413)|(g16619);
assign II27192 = ((~g27662));
assign II21734 = ((~g19268));
assign g28039 = ((~g26365));
assign g26947 = (g26394)|(g24285);
assign g31015 = (g29476&g22758);
assign g34319 = (g9535&g34156);
assign g17776 = ((~g14905));
assign g34995 = ((~II33285));
assign g28327 = (g27365&g19785);
assign II17653 = ((~g14276));
assign II17839 = ((~g13412));
assign g18677 = (g4639&g15758);
assign II22973 = ((~g9657))|((~II22972));
assign g28284 = (g11398&g27994);
assign g17748 = ((~g562))|((~g14708))|((~g12323));
assign g13709 = ((~g11755))|((~g11261));
assign g13946 = ((~g8651)&(~g11083));
assign II32645 = ((~g34367));
assign g27503 = (g26488&g14668);
assign g28735 = (g27510)|(g16737);
assign g33249 = (g32144&g20026);
assign g28060 = (g27616)|(g18532);
assign g27488 = (g26549&g17648);
assign g26853 = (g94&g24533);
assign g13736 = ((~g11313));
assign g28290 = (g23780&g27759);
assign g27127 = (g25997&g16582);
assign g24390 = (g23779)|(g21285);
assign g23675 = (g19050&g9104);
assign g32266 = (g30604)|(g29354);
assign g11034 = ((~g7611));
assign g17405 = (g1422&g13137);
assign g25389 = ((~g22457))|((~g12082));
assign g25470 = ((~g22457))|((~g2051))|((~g8365));
assign g24490 = ((~g22594));
assign g19554 = ((~g16861));
assign g10625 = (g3431&g7926);
assign g31706 = ((~II29270))|((~II29271));
assign g34243 = ((~II32228));
assign g25705 = (g25069)|(g18744);
assign II31032 = (g32501&g32502&g32503&g32504);
assign g28939 = (g17321&g25184&g26424&g27421);
assign II31849 = (g33483)|(g33484)|(g33485)|(g33486);
assign g27222 = (g26055&g13932);
assign g13074 = ((~II15702));
assign g32372 = (g29884)|(g31314);
assign g18520 = (g2661&g15509);
assign II15033 = ((~g10273));
assign g27259 = (g26755&g26725);
assign g20382 = ((~g15171));
assign g25800 = ((~g25518)&(~g25510));
assign g29484 = (g28124)|(g22191);
assign g17681 = ((~g14735));
assign g12797 = ((~g10275))|((~g7655))|((~g7643))|((~g7627));
assign g27515 = (g26051)|(g13431);
assign g23733 = ((~g20751))|((~g11178));
assign g24002 = (g19613&g10971);
assign II26679 = ((~g27773));
assign g34325 = ((~g34092));
assign g32111 = (g31616&g29922);
assign g25117 = ((~g22417));
assign g24168 = ((~II23348));
assign g7023 = ((~g5445));
assign g16680 = ((~g13223));
assign g31189 = ((~II29002));
assign II18048 = ((~g13638));
assign g12883 = ((~g10390));
assign g13517 = ((~g8541)&(~g12692));
assign g6989 = ((~g4575));
assign g33001 = (g32282)|(g18404);
assign g28817 = (g27548)|(g16845);
assign g24997 = (g22929&g10419);
assign g33340 = (g32222&g20639);
assign g24484 = (g16288&g23208);
assign g32095 = (g7619&g30825);
assign g8680 = ((~g686));
assign g10374 = ((~g6903));
assign g19510 = ((~g15969))|((~g10841))|((~g10899));
assign g29514 = (g1608&g28780);
assign g10366 = ((~g6895));
assign g25150 = (g17480&g23547);
assign g18687 = (g4664&g15885);
assign II15869 = ((~g11234));
assign g12979 = (g424&g11048);
assign g15123 = ((~g6975)&(~g13605));
assign g18501 = (g12854&g15509);
assign g32347 = (g29839)|(g31273);
assign g11913 = ((~g7197)&(~g9166));
assign II27481 = ((~g27928));
assign g26311 = (g2527&g25400);
assign g18549 = (g2799&g15277);
assign g9750 = ((~II13335))|((~II13336));
assign g18713 = (g4836&g15915);
assign g26845 = (g24391&g21426);
assign g23231 = ((~g20050));
assign g27400 = ((~g8553)&(~g26657));
assign g11706 = ((~II14579));
assign g10320 = ((~g817));
assign g19981 = ((~g3727)&(~g16316));
assign II25579 = ((~g25297));
assign g18974 = (g174&g16127);
assign g32186 = ((~II29720));
assign g8558 = ((~g3787));
assign g10410 = ((~g7069));
assign g28594 = (g27334)|(g26289);
assign g26050 = (g9630&g25047);
assign g33013 = (g32283)|(g18484);
assign g29284 = (g28554)|(g18747);
assign g13315 = ((~g1459))|((~g10715));
assign g12293 = ((~g7436))|((~g5283));
assign g24983 = (g23217&g20238);
assign g12893 = ((~g10391));
assign g20507 = ((~g15509));
assign g28665 = (g27409)|(g16614);
assign g10618 = ((~g10153))|((~g9913));
assign g21334 = ((~g14616))|((~g17596));
assign g27407 = (g26488&g17522);
assign g29631 = (g1682&g28656);
assign g22091 = (g6415&g18833);
assign g13176 = ((~g10715))|((~g7675))|((~g1322))|((~g1404));
assign g9951 = ((~g6133));
assign g34044 = ((~g33675));
assign II14370 = ((~g3303))|((~II14368));
assign gbuf60 = (g6675);
assign g33898 = (g33419&g15655);
assign II14964 = ((~g10230));
assign g16671 = (g6275&g14817);
assign II14230 = ((~g8055))|((~II14228));
assign g22157 = (g14608&g18892);
assign g16668 = (g5543&g14962);
assign g29042 = ((~II27388));
assign g9678 = ((~g5406));
assign g29322 = (g29192&g7074&g6336);
assign g19735 = (g9740&g17135);
assign II32809 = ((~g34586));
assign g28274 = ((~II26799));
assign g33038 = (g32184)|(g24311);
assign g23027 = ((~g20391));
assign g17756 = ((~g14858));
assign g12226 = ((~g2476)&(~g8373));
assign g12163 = ((~g5073)&(~g9989));
assign g13080 = (g6923&g11357);
assign g8186 = ((~g990));
assign g13108 = ((~g5551))|((~g12029))|((~g5685))|((~g9864));
assign g21357 = ((~g15736))|((~g13109))|((~g15726))|((~g13086));
assign g33114 = (g22139&g31945);
assign g24580 = (g22340)|(g13096);
assign g14180 = (g872&g10632);
assign g21355 = ((~g17821));
assign II29261 = ((~g29485))|((~g12046));
assign gbuf64 = (g6692);
assign gbuf139 = (g1426);
assign g8673 = ((~g4737));
assign II13287 = ((~g110));
assign g27335 = (g12087&g26776);
assign g27104 = (g25997&g16510);
assign g25018 = ((~g20107))|((~g23154));
assign g29596 = (g27823&g28620);
assign g17820 = ((~g5925))|((~g14549))|((~g6019))|((~g12614));
assign II24440 = ((~g14411))|((~II24438));
assign II31191 = (g30735&g31829&g32731&g32732);
assign g14825 = ((~g12806))|((~g12680));
assign g34012 = (g33886)|(g18480);
assign g16626 = ((~g14133));
assign g25790 = ((~g25027));
assign g31321 = (g30146&g27886);
assign g34126 = ((~II32067));
assign g14421 = ((~II16575));
assign g17521 = ((~g14727));
assign g34759 = ((~II32935));
assign II12709 = ((~g4284));
assign g14513 = ((~g12222)&(~g9754));
assign g30241 = (g28729&g23926);
assign II21250 = ((~g16540));
assign g32339 = (g31474&g20672);
assign g24316 = (g4527&g22228);
assign g14339 = ((~g12289)&(~g2735));
assign II30193 = (g31070)|(g30614)|(g30673)|(g31528);
assign II15906 = ((~g10430));
assign g10499 = ((~II13872));
assign g33043 = (g32195)|(g24325);
assign g24645 = (g22639&g19709);
assign g8340 = ((~g3050));
assign g30305 = ((~g28939));
assign g29144 = ((~g9518)&(~g26977));
assign g33122 = (g8859&g32192);
assign g19687 = ((~g17096));
assign g18161 = (g691&g17433);
assign g32154 = (g31277&g14184);
assign g24952 = (g21326)|(g21340)|(II24117);
assign g27031 = (g26213)|(g26190)|(g26166)|(g26148);
assign g24153 = ((~II23303));
assign g22921 = ((~g20219))|((~g2950));
assign II16077 = ((~g10430));
assign g32743 = ((~g30937));
assign g13085 = ((~II15717));
assign II12086 = ((~g622));
assign II14305 = ((~g8805));
assign g33563 = (g33361)|(g18383);
assign g23384 = ((~II22485));
assign g32773 = ((~g31376));
assign II24787 = ((~g24266));
assign g8033 = ((~g157));
assign g24023 = ((~g21127));
assign g32132 = (g31487)|(g31479);
assign g28579 = ((~g27714));
assign g19579 = ((~g16000));
assign g33146 = ((~g4669)&(~g32057));
assign g26545 = ((~g24881)&(~g24855));
assign g21732 = (g3004&g20330);
assign g14875 = (g1495&g10939);
assign II12546 = ((~g194))|((~II12544));
assign g31971 = ((~g30573))|((~g10511));
assign g29792 = (g28235)|(g28244);
assign g25080 = ((~g23742));
assign II12132 = ((~g577));
assign II19837 = ((~g1399));
assign g9644 = ((~g2016));
assign g31500 = (g29802&g23449);
assign g14101 = ((~g11653))|((~g11729));
assign g27237 = ((~g26162));
assign g23331 = ((~g20905));
assign g8876 = ((~II12855));
assign g7202 = ((~g4639));
assign g12946 = ((~II15564));
assign g19734 = ((~g16861));
assign g31133 = ((~g7953)&(~g29556));
assign g30146 = ((~g28833)&(~g7411));
assign II12469 = ((~g405))|((~II12468));
assign g8456 = ((~g56));
assign g28150 = (g10862&g11834&g11283&g27187);
assign g8064 = ((~g3376));
assign g32704 = ((~g31070));
assign g10395 = ((~g6995));
assign g34458 = (g34396)|(g18671);
assign g31748 = ((~II29303))|((~II29304));
assign g34389 = (g34170&g20715);
assign g17641 = ((~g14845));
assign g22541 = ((~II21911));
assign g25481 = ((~g22228));
assign g12023 = ((~g2453))|((~g8373));
assign g26085 = (g11906&g25070);
assign g32534 = ((~g30673));
assign g26084 = (g24926&g9602);
assign g12437 = ((~g2319)&(~g8267));
assign g22399 = ((~g1367)&(~g19720));
assign g25821 = (g25482)|(g25456)|(g25417)|(g25377);
assign g29622 = (g2579&g29001);
assign g24619 = ((~g23554)&(~g23581));
assign g20523 = ((~g17821));
assign g28032 = ((~g26365));
assign g33999 = (g33893)|(g18436);
assign g32342 = (g6545&g31579);
assign g25641 = ((~II24784));
assign g21408 = ((~g15373));
assign g16215 = ((~g1211)&(~g13545));
assign g15758 = ((~II17276));
assign g11273 = ((~g3061)&(~g8620));
assign g31670 = (g29937)|(g28573);
assign g12980 = ((~g7909)&(~g10741));
assign g18477 = (g2429&g15426);
assign g20046 = ((~g16540));
assign g11441 = ((~g9599))|((~g3267));
assign g12145 = ((~g8195))|((~g1760));
assign g10726 = ((~g7304))|((~g7661))|((~g979))|((~g1061));
assign g16531 = (g5232&g14656);
assign g21849 = (g3889&g21070);
assign g27263 = (g25940&g19713);
assign g32582 = ((~g31170));
assign g11419 = ((~II14428))|((~II14429));
assign g26162 = ((~g23052)&(~g24751));
assign II14331 = ((~g225))|((~II14330));
assign II31132 = (g32645&g32646&g32647&g32648);
assign II32446 = ((~g34127));
assign g9638 = ((~g1620));
assign g21694 = ((~g16540));
assign g10881 = ((~g7567));
assign g17093 = ((~II18165));
assign g25568 = (II24679&II24680);
assign g16155 = ((~II17495))|((~II17496));
assign g25633 = (g24420)|(g18282);
assign g12848 = ((~g6839)&(~g10430));
assign g22751 = (g19333)|(g15716);
assign g30329 = ((~II28588));
assign g18408 = (g2070&g15373);
assign g14015 = ((~g11658))|((~g11747));
assign g9808 = ((~g5827));
assign g34692 = ((~II32846));
assign g13241 = ((~g7503))|((~g10544));
assign g28289 = (g27734&g26575);
assign g25939 = (g24583&g19490);
assign g24601 = ((~g22957))|((~g2965));
assign g27014 = ((~g25888));
assign g19473 = ((~g16349));
assign g6767 = ((~II11626));
assign g33280 = (g32141)|(g29574);
assign g33366 = (g32268&g21010);
assign g32009 = (g31782&g22224);
assign g29228 = (g28426)|(g18173);
assign II15636 = ((~g12075));
assign g23586 = ((~g17284)&(~g20717));
assign g26962 = (g26295)|(g24307);
assign g34863 = (g16540&g34833);
assign gbuf123 = (g637);
assign g15734 = ((~g5228))|((~g12059))|((~g5290))|((~g14631));
assign g12515 = ((~g9511)&(~g5873));
assign g30169 = ((~g28833)&(~g14613));
assign g13064 = ((~g11705));
assign g29887 = (g28417&g23351);
assign g27646 = (g13094&g25773);
assign g28641 = (g27385)|(g16591);
assign g11609 = ((~g7660));
assign g34696 = (g34531&g20004);
assign g10231 = ((~g2661));
assign g22193 = (g19880&g20682);
assign g20162 = (g8737&g16750);
assign g19395 = ((~g16431));
assign g11185 = ((~g8038)&(~g8183)&(~g6804));
assign g26378 = (g19576&g25544);
assign g10158 = ((~g2461));
assign g13385 = (g11967)|(g9479);
assign g23246 = ((~g20785));
assign g15479 = ((~g14895));
assign g26350 = (g13087&g25517);
assign g25984 = ((~g24567))|((~g22668));
assign g11786 = ((~g7549));
assign g18948 = ((~g15800));
assign g24428 = ((~g22722));
assign g8068 = ((~g3457));
assign g26950 = (g26357)|(g24288);
assign g34384 = ((~II32391));
assign g12077 = ((~II14939));
assign g23819 = ((~g19147));
assign II13079 = ((~g5467))|((~II13077));
assign II12217 = ((~g1437))|((~g1478));
assign g7069 = ((~g6137));
assign g20386 = ((~g15224));
assign g9619 = ((~g5845));
assign g30214 = (g23424)|(g28572);
assign g29627 = (g28493&g11884);
assign g15680 = ((~II17207));
assign g9743 = ((~II13321));
assign g14091 = ((~g8854)&(~g12259));
assign g14688 = ((~g12604))|((~g12453));
assign g28888 = ((~g27738))|((~g8139));
assign g25969 = (g9310&g24987);
assign II24497 = ((~g22592));
assign g12037 = ((~II14893));
assign g14705 = ((~II16803));
assign g33600 = (g33418)|(g18501);
assign g34302 = ((~II32305));
assign g18423 = (g12851&g18008);
assign g21423 = ((~g15224));
assign g19691 = (g9614&g17085);
assign g33952 = (g33478)|(II31843)|(II31844);
assign g19614 = ((~g1542))|((~g16047));
assign g20910 = ((~g15171));
assign g18247 = (g1178&g16431);
assign g32794 = ((~g30937));
assign g13877 = ((~g11350));
assign g34802 = (g34757)|(g18589);
assign g28603 = (g27340)|(g26300);
assign g31996 = (g31779&g18979);
assign II20840 = ((~g17727));
assign II12262 = ((~g1454))|((~II12261));
assign g16653 = (g8343&g13850);
assign g14237 = ((~g11666));
assign g19268 = ((~g15979)&(~g962));
assign g18172 = (g15058&g17328);
assign g7003 = ((~g5152));
assign g23338 = ((~g20453));
assign g26844 = (g25261&g21418);
assign g23645 = ((~g20875));
assign g10878 = (g7858&g1135);
assign g26309 = ((~g8575)&(~g24825));
assign g32796 = ((~g31376));
assign g33891 = (g33264)|(g33269);
assign g25199 = ((~II24364))|((~II24365));
assign g23226 = ((~g20924));
assign g22085 = (g6295&g19210);
assign g29503 = ((~g22763)&(~g28250));
assign g13670 = ((~g8123)&(~g10756));
assign g23373 = (g13699&g20195);
assign g9708 = ((~g2741));
assign II32991 = ((~g34759));
assign g26899 = (g26844)|(g18199);
assign II20929 = ((~g17663));
assign g32289 = (g24796)|(g31230);
assign g33070 = (g32010)|(g22114);
assign g34676 = ((~II32812));
assign g27957 = (g25947&g15995);
assign g14190 = (g859&g10632);
assign g24242 = (g22834)|(g18253);
assign g26255 = ((~g8075))|((~g24779));
assign g25414 = (g5406&g22194&II24549);
assign g24905 = ((~g534))|((~g23088));
assign g29309 = (g28722)|(g18818);
assign g33471 = (g32535&II31051&II31052);
assign g25011 = ((~g22763));
assign g30039 = ((~g29134));
assign g32973 = ((~g31021));
assign g12432 = ((~g1894)&(~g8249));
assign g30059 = (g28106&g12467);
assign g23281 = ((~g18957))|((~g2898));
assign g32467 = ((~g31194));
assign g11658 = ((~g8021)&(~g3506));
assign g11810 = ((~g9664));
assign g26633 = (g24964&g20616);
assign g15969 = ((~II17416));
assign g29296 = (g28586)|(g18781);
assign g31855 = ((~g29385));
assign g9909 = ((~g1978));
assign g32460 = ((~g31194));
assign g22064 = (g15162&g19210);
assign II23309 = ((~g21677));
assign g25904 = (g14001&g24791);
assign g7635 = ((~g1002));
assign g33815 = (g33449&g12911);
assign g13997 = (g11029)|(g11036);
assign g24031 = ((~g21193));
assign g29104 = ((~g5188)&(~g27999));
assign g22979 = ((~g20453));
assign g24368 = ((~g22228));
assign g32126 = (g31601&g29948);
assign g25543 = (g23795&g21461);
assign g18931 = ((~g16031));
assign g9728 = ((~g5109));
assign g6828 = ((~g1300));
assign g14535 = ((~g12318));
assign g18625 = (g15092&g17062);
assign g24186 = (g18102&g22722);
assign g28920 = ((~g27779))|((~g1802))|((~g7315));
assign g11231 = ((~g7928)&(~g4801)&(~g4793));
assign g10518 = ((~g9311));
assign g26611 = (g24935&g20580);
assign g15632 = (g3494&g13555);
assign g18812 = (g6509&g15483);
assign g21562 = ((~II21199));
assign g14797 = ((~g12593))|((~g12405));
assign g29610 = (g28483&g8026);
assign g14545 = ((~g12768));
assign g18190 = (g822&g17821);
assign g20582 = ((~g17873));
assign g6817 = ((~g956));
assign g25585 = (g21674)|(g24155);
assign g21708 = (g15049&g20283);
assign g34023 = (g33796)|(g24320);
assign II14429 = ((~g4005))|((~II14427));
assign g34509 = (g34283&g19473);
assign g19207 = (g7803&g15992);
assign g11016 = (g4888&g8984);
assign II13875 = ((~g1233));
assign g27520 = (g26519&g17714);
assign gbuf142 = (g1500);
assign g30377 = (g30124)|(g18472);
assign II12487 = ((~g3443));
assign g14399 = ((~g5297)&(~g12598));
assign g34377 = (g26304)|(g34141);
assign g7943 = ((~g1395));
assign g24403 = (g4894&g22858);
assign g34246 = ((~II32237));
assign g23555 = ((~II22692));
assign g32545 = ((~g31070));
assign g16044 = ((~g10961)&(~g13861));
assign g31495 = (g1913&g30309);
assign g26654 = ((~g25275));
assign g34294 = (g26855)|(g34225);
assign g13092 = ((~g1061))|((~g10761));
assign II30330 = (g29385)|(g31376)|(g30735)|(g30825);
assign g12558 = ((~g7738)&(~g5517)&(~g5511));
assign g12929 = ((~g12550));
assign II29891 = ((~g31578));
assign g28051 = (g27699)|(g18166);
assign g17673 = ((~g14723));
assign II13740 = ((~g85));
assign g24353 = (g23682)|(g18822);
assign g16485 = (g5563&g14924);
assign g34537 = (g34324)|(g34084);
assign g25734 = (g25058)|(g18782);
assign g27995 = (g26809&g23985);
assign II26394 = ((~g26488))|((~II26393));
assign g34133 = (g33845&g23958);
assign g24858 = (g3361&g23223&II24030);
assign g31768 = (g30033)|(g30045);
assign II17633 = ((~g13258));
assign g7243 = ((~II11892));
assign g18616 = (g6875&g17200);
assign g8703 = ((~II12709));
assign g31255 = (g25982)|(g29536);
assign g28125 = (g27381&g26209);
assign g26349 = (g24630)|(g13409);
assign g22027 = (g5889&g19147);
assign g30502 = (g30232)|(g22023);
assign II26378 = ((~g26850));
assign g32698 = ((~g30614));
assign g7804 = (g2975&g2970);
assign g24249 = (g22624)|(g18294);
assign g9337 = ((~g1608));
assign g21432 = ((~g17790))|((~g14820))|((~g17761))|((~g14780));
assign g11215 = ((~g8285));
assign g18636 = (g3817&g17096);
assign g25789 = (g25285)|(g14543);
assign g32768 = ((~g30825));
assign g8651 = ((~g758));
assign II13672 = ((~g106));
assign g34102 = (g33912&g23599);
assign g22332 = ((~II21838));
assign II30751 = (g32042)|(g32161)|(g31943)|(g31959);
assign g30090 = ((~g29134));
assign g34477 = (g26344&g34328);
assign g21820 = (g3712&g20453);
assign g26710 = ((~g25349));
assign g33857 = (g33267&g20445);
assign g32225 = (g30576)|(g29336);
assign gbuf4 = (g4449);
assign g25932 = ((~g7680)&(~g24528));
assign g16509 = ((~g13873));
assign g28295 = (g27094)|(g15783);
assign g28091 = (g27665)|(g21913);
assign II33047 = ((~g34776));
assign g32490 = ((~g30673));
assign g9970 = ((~g1714));
assign g19766 = ((~g16449));
assign g16100 = ((~II17471));
assign II15364 = ((~g10182))|((~II15363));
assign g14033 = ((~g8808)&(~g12259));
assign g22856 = ((~g20453));
assign g32257 = (g31184)|(g29708);
assign g33485 = (g32635&II31121&II31122);
assign g32878 = ((~g30937));
assign g14221 = (g8686&g11823);
assign g31801 = ((~g29385));
assign g33742 = (g7828&g33142&II31600);
assign g34924 = ((~II33164));
assign g14437 = ((~g9527)&(~g11178));
assign g33274 = (g32126)|(g29563);
assign g18367 = (g1783&g17955);
assign II17462 = ((~g1300))|((~II17460));
assign g18798 = (g6177&g15348);
assign g30475 = (g30220)|(g21946);
assign II13462 = ((~g2380))|((~g2384));
assign g8287 = ((~g160));
assign g12486 = ((~g9055)&(~g9013)&(~g8957)&(~g8905));
assign g23965 = ((~g21611));
assign g25958 = ((~g7779)&(~g24609));
assign g11923 = ((~II14734))|((~II14735));
assign g30931 = ((~II28913));
assign g18260 = (g1252&g16000);
assign g28161 = ((~II26676));
assign g17478 = ((~g14996));
assign g20546 = ((~g18008));
assign g18357 = (g1816&g17955);
assign g15169 = ((~II17094));
assign g10951 = ((~g7845))|((~g7868));
assign g20453 = ((~II20584));
assign g32433 = ((~II29961));
assign g32556 = ((~g31554));
assign g8497 = ((~g3436));
assign g27185 = (g26190&g8302&g1917);
assign g22637 = (g19363&g19489);
assign g12123 = ((~g6856)&(~g2748));
assign g33889 = (g33303&g20641);
assign g25224 = ((~g22763));
assign g10406 = ((~g7046));
assign g26302 = (g2393&g25349);
assign g30295 = ((~II28540));
assign g29939 = ((~g28857));
assign g20497 = ((~g18065));
assign g16192 = (g6191&g14321);
assign II12855 = ((~g4311));
assign g20515 = ((~g15483));
assign g11031 = ((~g8609));
assign g33162 = ((~g4859)&(~g32072));
assign g29363 = (g8458&g28444);
assign g18695 = (g4737&g16053);
assign g23842 = ((~g19147));
assign g33946 = (g32434)|(g33456);
assign g20615 = ((~g15509));
assign g23908 = ((~g20739));
assign g24089 = ((~g19890));
assign II20433 = ((~g16234));
assign g27564 = (g26305&g23378);
assign g27272 = (g26055&g17144);
assign g13256 = ((~g11846))|((~g11294))|((~g11812));
assign g31754 = (g29989)|(g30006);
assign g20192 = ((~g17268));
assign g21795 = (g3506&g20924);
assign g29348 = ((~g28194));
assign g28874 = ((~g27907))|((~g7424))|((~g2421));
assign g33478 = (g32584&II31086&II31087);
assign g7228 = ((~g6398))|((~g6444));
assign g31231 = (g30290&g25239);
assign g23859 = ((~g19074));
assign II20529 = ((~g16309));
assign g30317 = (g29208)|(II28566)|(II28567);
assign g23475 = (g19070&g8971);
assign g22686 = (g19335&g19577);
assign g30559 = (g30269)|(g22130);
assign g12000 = ((~g8418))|((~g2610));
assign g8010 = ((~II12345))|((~II12346));
assign g19745 = ((~g16877));
assign II14369 = ((~g8481))|((~II14368));
assign g26303 = (g2685&g25439);
assign g10180 = ((~g2259));
assign g20182 = ((~g16897));
assign g12692 = (g10323&g3522&g3530);
assign g30211 = (g28685&g23878);
assign g12933 = ((~g7150))|((~g10515));
assign g23496 = ((~g20248));
assign g31765 = (g30128&g23968);
assign g28565 = (g27315)|(g26253);
assign g13048 = (g8558&g11043);
assign g7857 = ((~II12241))|((~II12242));
assign g10216 = ((~II13684));
assign g19696 = ((~g17015));
assign g26818 = ((~II25530));
assign g28846 = (g21434&g26424&g25399&g27474);
assign g25927 = (g25004&g20375);
assign g8172 = ((~g3873));
assign g32913 = ((~g30825));
assign g8138 = ((~g1500));
assign g32397 = (g31068&g15830);
assign II32517 = ((~g34424))|((~II32516));
assign g25214 = ((~g22228));
assign g33862 = (g33272&g20504);
assign g7536 = ((~g5976));
assign g16801 = (g5120&g14238);
assign g31317 = (g29611)|(g29626);
assign g27368 = ((~g8119)&(~g26657));
assign g31902 = (g31744)|(g21910);
assign g19798 = ((~g17200));
assign g21060 = ((~g15509));
assign g23001 = ((~g19801));
assign g33413 = ((~g31971));
assign g12345 = ((~g7158));
assign g17139 = (g8635&g12967);
assign g29033 = ((~g5511)&(~g7738)&(~g28010));
assign g14529 = ((~g6336)&(~g12749));
assign g16727 = ((~g14454));
assign g23519 = ((~g21468));
assign g17468 = ((~g3215))|((~g13700))|((~g3317))|((~g8481));
assign g15579 = ((~II17159));
assign g19441 = (g15507)|(g12931);
assign g9739 = ((~g5752));
assign g32662 = ((~g30614));
assign g21725 = ((~II21294));
assign g32778 = ((~g31021));
assign g21069 = ((~g15277));
assign g18758 = (g7004&g15595);
assign g28319 = (g27115)|(g15807);
assign II32071 = ((~g33665));
assign g32867 = ((~g30673));
assign g25638 = (g24977)|(g18316);
assign g8087 = ((~g1157));
assign g20781 = ((~II20840));
assign g24226 = (g446&g22594);
assign II16541 = ((~g11929));
assign g31791 = ((~II29363));
assign g12922 = ((~g12297));
assign g24131 = ((~g21209));
assign g34192 = ((~g33921));
assign g8500 = ((~g3431))|((~g3423));
assign g15857 = (g3199&g14038);
assign g22902 = ((~g18957))|((~g2848));
assign g22874 = ((~g18918))|((~g2844));
assign g23490 = ((~g21514));
assign g33801 = (g33437&g25327);
assign g27456 = (g25978)|(g24607);
assign g32313 = (g31303&g23515);
assign g10114 = ((~g2116));
assign g21269 = ((~g15506));
assign g31277 = (g29570)|(g28285);
assign g18280 = (g1367&g16136);
assign g24377 = ((~g22594));
assign g21719 = (g358&g21037);
assign g23267 = ((~g20097));
assign g32944 = ((~g31021));
assign g10490 = ((~g9274));
assign g16808 = (g6653&g14825);
assign g25558 = ((~g22594));
assign g33087 = (g32391&g18888);
assign g30151 = (g28607&g21249);
assign g27524 = (g26050)|(g24649);
assign g8679 = (g222)|(g199);
assign g30422 = (g29795)|(g21806);
assign g14146 = ((~g11020))|((~g691));
assign II23396 = ((~g23427));
assign g11906 = ((~II14713))|((~II14714));
assign g34545 = ((~g11679))|((~g794))|((~g34354));
assign g24058 = ((~g20982));
assign g18225 = (g1041&g16100);
assign g10334 = ((~g4420));
assign g31229 = (g30288&g23949);
assign g20641 = ((~g15509));
assign g33232 = (g32034)|(g30936);
assign g9913 = ((~g2403));
assign II29909 = ((~g31791));
assign g34689 = ((~II32837));
assign g23002 = ((~II22177));
assign g22000 = (g5727&g21562);
assign g28113 = (g8016&g27242);
assign g15912 = (g3562&g14018);
assign g10026 = ((~g6494));
assign g21412 = ((~g15758));
assign g23451 = (g13805&g20510);
assign g8211 = ((~g2319));
assign g32802 = ((~g31327));
assign g27903 = ((~g21228))|((~g25316))|((~g26424))|((~g26218));
assign g29245 = (g28676)|(g18384);
assign g16031 = ((~II17436));
assign g16987 = ((~II18135));
assign g32028 = (g30569&g29339);
assign g26398 = (g24946&g10474);
assign g18258 = (g1221&g16897);
assign g17847 = ((~II18839));
assign g18165 = (g650&g17433);
assign g21891 = (g19948)|(g15103);
assign II14289 = ((~g8282))|((~g3835));
assign g21869 = (g4087&g19801);
assign g24510 = (g22488)|(g7567);
assign g15155 = ((~g12899)&(~g13782));
assign II28866 = ((~g29730));
assign g33269 = (g31970&g15582);
assign g13960 = ((~g11669))|((~g11537));
assign g11492 = ((~g6928))|((~g6941))|((~g8756));
assign g31467 = (g30162&g27937);
assign g18426 = (g2177&g18008);
assign g32781 = ((~g31376));
assign g13478 = ((~g12511))|((~g12460))|((~g12414))|((~g12344));
assign g27598 = (g25899&g10475);
assign g16326 = ((~II17658));
assign g33930 = ((~g33394))|((~g12767))|((~g9848));
assign II14352 = ((~g8848))|((~II14350));
assign g30160 = ((~g28846)&(~g7387));
assign g27178 = (g25997&g16652);
assign g28185 = (g27026&g19435);
assign II15335 = ((~g2116))|((~II15333));
assign g17408 = ((~II18341));
assign g25035 = ((~g23699));
assign g34074 = (g33685&g19498);
assign g26207 = (g2638&g25170);
assign g13097 = ((~g5204))|((~g12002))|((~g5339))|((~g9780));
assign II15550 = ((~g10430));
assign g31898 = (g31707)|(g21906);
assign g32868 = ((~g31376));
assign g26166 = (g25357&g11724&g11709&g7558);
assign g20445 = ((~g15224));
assign g11116 = (g9960&g6466);
assign g33759 = (g33123&g22847);
assign g30601 = ((~g16279)&(~g29718));
assign g14695 = ((~g5583))|((~g12029))|((~g5637))|((~g12301));
assign g33321 = (g29712)|(g32182);
assign g7017 = ((~g128));
assign g33006 = (g32291)|(g18447);
assign II14475 = ((~g10175));
assign g18555 = (g2834&g15277);
assign g17657 = ((~g14751)&(~g12955));
assign g26053 = ((~g22875))|((~g24677))|((~g22941));
assign g31275 = (g30147&g27800);
assign g20589 = ((~g15224));
assign g16927 = (g13524)|(g11126);
assign g13416 = ((~II15929));
assign g32552 = ((~g30825));
assign g33103 = ((~g32176)&(~g31212));
assign g32386 = (g31488)|(g29949);
assign g33605 = (g33352)|(g18521);
assign g29165 = ((~g5881)&(~g28020));
assign g30527 = (g30192)|(g22073);
assign g22535 = ((~g19699)&(~g1030));
assign g15129 = ((~g6984)&(~g13638));
assign g33391 = ((~g32384));
assign g10278 = ((~g4628));
assign g23912 = ((~g19147));
assign g27299 = (g26546&g23028);
assign g28611 = (g27348)|(g16485);
assign g7462 = ((~g2599));
assign g19389 = ((~g17532));
assign g24662 = ((~g22957))|((~g2955));
assign g34629 = (g34495)|(g18654);
assign g21767 = (g3239&g20785);
assign g23032 = ((~II22211));
assign II31357 = (g32970&g32971&g32972&g32973);
assign g26146 = (g9892&g25334);
assign g23789 = ((~g21308));
assign g33653 = ((~II31486));
assign g31134 = ((~g8033)&(~g29679)&(~g24732));
assign g16173 = (g8796)|(g13464);
assign g13259 = ((~II15824));
assign g8890 = ((~g376));
assign g26200 = (g24688&g10678&g10658&g10627);
assign II18482 = ((~g13350));
assign g15932 = ((~II17395));
assign g23398 = ((~g21468));
assign g10223 = ((~g4561));
assign g33713 = ((~II31564));
assign g17794 = ((~g13350));
assign g19935 = ((~g17062)&(~g8113));
assign g27064 = ((~II25786));
assign g23013 = ((~g20330));
assign g11350 = ((~II14369))|((~II14370));
assign II32788 = ((~g34577));
assign g32667 = ((~g30825));
assign g7701 = ((~g4859))|((~g4849))|((~g4843));
assign II30734 = (g31790)|(g32191)|(g32086)|(g32095);
assign g28803 = ((~g27730)&(~g22763));
assign g9686 = ((~g73));
assign g34662 = (g34576&g18931);
assign g33027 = (g32314)|(g21796);
assign II12644 = ((~g3689));
assign g21245 = ((~II20982));
assign g14204 = ((~g12155));
assign g8363 = ((~g239));
assign g21914 = (g5077&g21468);
assign g7850 = ((~g554))|((~g807));
assign g9824 = ((~g1825));
assign g32173 = (g160&g31134);
assign g18659 = (g4366&g17183);
assign g34727 = (g34655)|(g18213);
assign g31504 = (g29370&g10553);
assign g14045 = ((~g11571))|((~g11747));
assign II17507 = ((~g13416));
assign g32294 = (g31231)|(g31232);
assign g23218 = (g20200&g16530);
assign g28754 = ((~II27238));
assign g25602 = (g24673)|(g18113);
assign g18896 = ((~g16031));
assign g22592 = ((~II21930));
assign g18291 = (g1437&g16449);
assign g24256 = (g22873)|(g18309);
assign g30338 = (g29613)|(g18240);
assign g16319 = ((~g8224))|((~g8170))|((~g13736));
assign II16671 = (g10185&g12461&g12415);
assign g28917 = ((~II27314));
assign g29940 = (g1740&g28758);
assign g25624 = (g24408)|(g18224);
assign g32434 = ((~g31189));
assign g12739 = ((~g9321)&(~g9274));
assign g11345 = ((~g8477)&(~g8479));
assign g28209 = (g27223)|(g27141);
assign g34036 = (g33722)|(g18715);
assign g18916 = ((~g16053));
assign g18459 = (g2331&g15224);
assign g15979 = ((~II17420));
assign g19650 = ((~g16971));
assign g32608 = ((~g31376));
assign g8616 = ((~g2803));
assign g11483 = ((~g8165)&(~g3522));
assign II23586 = ((~g22409))|((~II23585));
assign g15563 = ((~II17140));
assign g18911 = ((~g15169));
assign g18289 = (g1448&g16449);
assign g30351 = (g30084)|(g18339);
assign g29200 = ((~g7791)&(~g26977));
assign g11761 = ((~II14610))|((~II14611));
assign g12527 = (g8680&g667);
assign II18443 = ((~g13027));
assign g30569 = ((~II28838));
assign g33611 = (g33243)|(g18632);
assign g13551 = ((~g11812))|((~g7479))|((~g7903))|((~g10521));
assign II32963 = ((~g34650));
assign g12450 = ((~g7738))|((~g10281));
assign II26070 = ((~g26026))|((~g13517));
assign g18155 = (g15056&g17533);
assign g26875 = (g21652)|(g25575);
assign g34584 = (g24653&g34315);
assign g24080 = ((~g21143));
assign g17180 = ((~g1559)&(~g13574));
assign g12423 = ((~II15242))|((~II15243));
assign g32993 = (g32255)|(g18352);
assign g25136 = ((~g22457));
assign g18537 = (g6856&g15277);
assign g10082 = ((~g2375));
assign g21740 = (g3085&g20330);
assign g23564 = (g16882&g20648);
assign g27817 = (g22498&g25245&g26424&g26236);
assign II31497 = ((~g33187));
assign g8916 = ((~II12887));
assign g14947 = ((~g12785))|((~g10491));
assign g16874 = ((~II18066));
assign II32985 = ((~g34736));
assign II16795 = ((~g5637));
assign g34282 = (g26838)|(g34214);
assign g9326 = ((~g6203));
assign g15137 = ((~g6992)&(~g13680));
assign g14126 = (g881&g10632);
assign g23270 = ((~g20785));
assign II18758 = ((~g6719));
assign g29319 = (g28812)|(g14453);
assign g7167 = ((~g5360))|((~g5406));
assign g18180 = (g767&g17328);
assign g23825 = (g20705)|(g20781);
assign g34125 = (g33724)|(g33124);
assign g33906 = (g33084&g22311);
assign g32086 = (g7597&g30735);
assign g23353 = ((~g20924));
assign g30208 = (g28681&g23875);
assign g20527 = ((~g18008));
assign g23763 = ((~g2795)&(~g21276));
assign g30383 = (g30138)|(g18513);
assign g13715 = ((~g10573));
assign g23257 = ((~g20924));
assign II16695 = (g10207&g12523&g12463);
assign g8132 = ((~II12411));
assign g25532 = ((~g21360))|((~g23363));
assign g16924 = ((~II18092));
assign g23732 = ((~g18833));
assign g21754 = (g3195&g20785);
assign g20708 = ((~g15426));
assign g17791 = ((~g14950));
assign g9567 = ((~g6116))|((~g6120));
assign g31870 = (g30607)|(g18262);
assign g13497 = (g2724&g12155);
assign II17783 = ((~g13304));
assign g18412 = (g2098&g15373);
assign g29189 = ((~g9462)&(~g26977)&(~g7791));
assign g24148 = ((~g19268)&(~g19338));
assign g24474 = ((~g23620));
assign g23275 = (g19680)|(g16160);
assign g25168 = ((~II24334));
assign g34673 = ((~II32803));
assign II15626 = ((~g12041));
assign g13906 = ((~II16201));
assign g23481 = ((~II22604));
assign II26516 = ((~g26824));
assign g18938 = ((~g16053));
assign g23862 = ((~g19147));
assign g18778 = (g5817&g18065);
assign g32601 = ((~g31376));
assign g26573 = ((~g24897)&(~g24884));
assign g22106 = (g6497&g18833);
assign II22923 = ((~g21284))|((~II22921));
assign g17570 = (g14419)|(g14397)|(g11999)|(II18495);
assign g24289 = (g4427&g22550);
assign g30287 = (g28653)|(g27677);
assign g10587 = ((~g2421))|((~g7456));
assign g28402 = (g27213)|(g15873);
assign II16663 = ((~g10981));
assign II14579 = ((~g8792));
assign g29350 = (g4939&g28395);
assign g34258 = (g34211)|(g18675);
assign g19458 = ((~II19927));
assign g27709 = ((~II26337));
assign g26838 = (g2860&g24515);
assign g34138 = (g33929&g23828);
assign g19630 = ((~g16897));
assign g32335 = (g6199&g31566);
assign g34744 = (g34668&g19481);
assign g24556 = (g4035&g23341);
assign g17575 = ((~g14921));
assign II18635 = ((~g14713))|((~II18633));
assign g16310 = ((~g13223));
assign g23458 = ((~II22583));
assign II24400 = ((~g23954));
assign g12067 = ((~g5990)&(~g7051));
assign g6976 = ((~II11750));
assign g24385 = ((~g22908));
assign g19361 = ((~II19843));
assign g23692 = ((~g9501))|((~g20995));
assign g30990 = ((~g29676));
assign g12860 = ((~g10368));
assign g13938 = (g11213)|(g11191);
assign II16709 = ((~g10430));
assign g25818 = (g8124&g24605);
assign g32151 = (g31639&g29996);
assign g14753 = ((~g11317));
assign II33103 = ((~g34846));
assign II18028 = ((~g13638));
assign g23391 = ((~g20645));
assign g10141 = ((~II13634));
assign g21300 = ((~II21047));
assign g27025 = (g26334&g7917);
assign g19379 = ((~g17327));
assign g24238 = (g23254)|(g18248);
assign g10652 = ((~g7601));
assign g33795 = (g33138&g20782);
assign g33476 = (g32570&II31076&II31077);
assign g27038 = ((~g25932));
assign g33882 = (g33293&g20587);
assign g34866 = (g34819&g20106);
assign g14295 = (g1811&g11894);
assign g28088 = (g27264)|(g18729);
assign g30220 = (g28699&g23888);
assign g28976 = ((~g27903))|((~g8273));
assign g16185 = (g3263&g14011);
assign g25834 = (g25366)|(g23854);
assign g15570 = ((~g822)&(~g14279));
assign g26615 = ((~g25432));
assign II29255 = ((~g12017))|((~II29253));
assign g26901 = (g26362)|(g24218);
assign g15092 = ((~g12864)&(~g13177));
assign II22893 = ((~g12189))|((~II22892));
assign g32697 = ((~g31070));
assign II27235 = ((~g27320));
assign g16805 = (g7187&g12972);
assign g29883 = (g2465&g29152);
assign g31842 = ((~g29385));
assign g8566 = ((~g3831));
assign g18269 = (g15069&g16031);
assign g31923 = (g31763)|(g22048);
assign g25357 = (g23810&g23786);
assign g23509 = ((~g21611));
assign g24230 = (g901&g22594);
assign g17492 = ((~g8655))|((~g14367));
assign g25159 = (g4907&g22908);
assign g14504 = ((~g12361));
assign g8921 = (II12902)|(II12903);
assign g34339 = ((~g34077));
assign g6940 = ((~g4035));
assign g31820 = ((~g29385));
assign g30167 = (g28622&g23793);
assign g32884 = ((~g30825));
assign g14414 = ((~g12145)&(~g9639));
assign II13139 = ((~g6154))|((~g6159));
assign g34332 = (g34071)|(g33723);
assign g19210 = ((~II19796));
assign g27674 = (g26873&g23543);
assign g34553 = ((~II32621));
assign g32559 = ((~g30825));
assign g34601 = (g34488)|(g18211);
assign g30375 = (g30149)|(g18466);
assign II22966 = ((~g12288))|((~II22965));
assign g21274 = ((~g15373));
assign II18647 = ((~g5320));
assign g21280 = ((~g16601));
assign g21880 = (g4135&g19801);
assign g25087 = (g17307&g23489);
assign g15858 = (g3542&g14045);
assign g33544 = (g33392)|(g18317);
assign II25567 = ((~g25272));
assign g30925 = (g29908&g23309);
assign g34445 = (g34382)|(g18548);
assign g29215 = ((~II27561));
assign II14398 = ((~g8542))|((~g3654));
assign g17194 = ((~g11039)&(~g13480));
assign g34195 = ((~II32150));
assign g19446 = ((~II19917));
assign g20550 = ((~g15864));
assign g9417 = ((~II13124));
assign II18614 = ((~g6315));
assign g19330 = ((~g17326));
assign g16638 = (g6271&g14773);
assign g12614 = ((~g9935));
assign g13246 = ((~g10939));
assign g21299 = ((~g16600));
assign gbuf44 = (g6023);
assign g7781 = ((~g4064)&(~g4057));
assign g20559 = (g336&g15831);
assign g20603 = ((~g17873));
assign g18486 = (g2485&g15426);
assign II13402 = ((~g2246))|((~II13401));
assign g32870 = ((~g31021));
assign g19965 = ((~g3380))|((~g16424));
assign g14615 = (g10604&g10587);
assign g32197 = (g31144&g20088);
assign g25744 = (g25129)|(g22059);
assign g28655 = (g27561&g20603);
assign g24727 = (g13300&g23016);
assign g11512 = ((~g7634));
assign g17639 = ((~II18600));
assign g33082 = (g32389&g18877);
assign II13066 = ((~g4308))|((~II13065));
assign g20033 = ((~g16579));
assign II13202 = ((~g5105));
assign g31846 = ((~g29385));
assign g24113 = ((~g19984));
assign II25683 = ((~g25642));
assign g15824 = ((~II17324));
assign g24279 = (g23218)|(g15105);
assign g31146 = (g12285&g30053);
assign g29789 = (g28270&g10233);
assign g29733 = (g2675&g29157);
assign g23794 = ((~g19147));
assign g16696 = ((~g13871))|((~g13855))|((~g14682))|((~g12340));
assign g25921 = (g24936&g9664);
assign g21888 = (g4165&g19801);
assign g29984 = (g2567&g28877);
assign g10353 = ((~g6803));
assign g26190 = (g25357&g11724&g7586&g11686);
assign g33076 = (g32336)|(g32446);
assign g30580 = ((~g29335))|((~g19666));
assign g25476 = ((~g22472))|((~g2476))|((~g8373));
assign II24191 = ((~g22360));
assign II12840 = ((~g4222))|((~g4235));
assign g13078 = ((~g7446)&(~g10762));
assign g20674 = ((~g15277));
assign II12123 = ((~g758));
assign g25334 = ((~g21253))|((~g23756));
assign g14589 = (g10586&g10569);
assign g20568 = ((~g15509));
assign II32824 = ((~g34475));
assign gbuf36 = (g5452);
assign g16473 = ((~g13977));
assign g26754 = ((~g25300));
assign g22498 = (g7753&g7717&g21334);
assign g29490 = (g25832)|(g28136);
assign g22835 = (g15803&g19633);
assign g8357 = ((~II12538));
assign g7854 = ((~g1152));
assign g12999 = ((~g4392))|((~g10476))|((~g4401));
assign g32758 = ((~g31327));
assign g8139 = ((~g1648));
assign g22303 = ((~g19277));
assign g22119 = (g6581&g19277);
assign II15954 = ((~g12381));
assign g14030 = (g11037)|(g11046);
assign g22078 = (g6267&g19210);
assign g34794 = (g34746)|(g18571);
assign g12190 = ((~g8365))|((~g8255));
assign g31853 = ((~g29385));
assign g15507 = (g10970&g13305);
assign gbuf111 = (g4204);
assign g17472 = ((~g14656));
assign II17772 = ((~g14888));
assign II24619 = (g6423&g6428&g10014);
assign g27578 = (g26155)|(g24747);
assign g22011 = (g15154&g21562);
assign g9755 = ((~g2070)&(~g1996));
assign g20144 = ((~g17533));
assign g16090 = ((~g10961)&(~g13315));
assign g20734 = ((~g14408))|((~g17312));
assign g8789 = ((~II12779));
assign g34080 = (g22957&g9104&g33750);
assign g32482 = ((~g30614));
assign g18828 = ((~g17955));
assign g25006 = ((~g22417));
assign g25957 = (g17190&g24960);
assign g34067 = ((~g33859)&(~g11772));
assign g29757 = (g28305&g23221);
assign g17617 = (g7885&g13326);
assign g14365 = ((~g12084)&(~g9339));
assign II13360 = ((~g5343));
assign g26049 = (g9621&g25046);
assign g15713 = ((~g5571))|((~g14425))|((~g5673))|((~g9864));
assign g25331 = (g5366&g22194&II24508);
assign g18137 = (g538&g17249);
assign g32326 = (g31317&g23539);
assign g14509 = ((~II16626));
assign g18174 = (g739&g17328);
assign g27201 = (g25997&g16685);
assign g18189 = (g812&g17821);
assign g19620 = ((~g17296));
assign g18669 = (g4608&g17367);
assign II16898 = ((~g10615));
assign g22882 = ((~g20391));
assign g23063 = ((~g16313)&(~g19887));
assign g23975 = ((~II23119))|((~II23120));
assign g21834 = (g3752&g20453);
assign g30005 = (g28230&g24394);
assign g30027 = (g29104&g12550);
assign g8541 = ((~g3498));
assign g12644 = ((~g10233))|((~g4531));
assign g14800 = ((~g7704))|((~g12443));
assign g20329 = ((~g15277));
assign g21655 = ((~g17657)&(~g17700));
assign g9527 = ((~g6500));
assign g23086 = ((~g20283));
assign g9509 = ((~g5770))|((~g5774));
assign II30750 = (g31788)|(g32310)|(g32054)|(g32070);
assign II13352 = ((~g4146));
assign gbuf56 = (g6373);
assign g32389 = (g31496)|(g29966);
assign g25670 = (g24967)|(g18626);
assign g32957 = ((~g31672));
assign g18113 = (g405&g17015);
assign g34923 = ((~II33161));
assign gbuf9 = (g4999);
assign g17200 = ((~II18238));
assign g30501 = (g29327)|(g22018);
assign g27714 = (g22384&g25195&g26424&g26171);
assign g13524 = (g9995&g11910);
assign g32788 = ((~g31327));
assign g18231 = (g1105&g16326);
assign II18333 = ((~g1083));
assign g24282 = (g23407)|(g18657);
assign g32390 = (g31501)|(g29979);
assign g31206 = (g30260&g23890);
assign g34683 = ((~II32827));
assign g32827 = ((~g31672));
assign g16069 = ((~II17447))|((~II17448));
assign g15107 = (g4258&g14454);
assign g7778 = ((~g1339));
assign g31786 = (g30189&g24010);
assign g16519 = (g5591&g14804);
assign g21686 = ((~g16540));
assign g25462 = (g6404&g22300&II24585);
assign g15100 = ((~g13191)&(~g12870));
assign g29836 = (g28425&g26841);
assign g23198 = (g20214)|(g20199)|(II22298);
assign g30075 = (g28525&g20662);
assign II14823 = ((~g8056));
assign II25552 = ((~g25240));
assign g29912 = ((~g28827));
assign g34047 = ((~g33637));
assign g9889 = ((~g6128));
assign g21187 = ((~g14616))|((~g17364));
assign g30409 = (g29842)|(g21768);
assign g24509 = ((~g22689));
assign g27213 = (g26026&g16721);
assign g16235 = ((~g13437));
assign g24502 = (g23428&g13223);
assign II18825 = ((~g6019));
assign g29006 = ((~g5180)&(~g27999));
assign g28509 = ((~g8107)&(~g27602));
assign g15840 = (g3949&g14142);
assign g20670 = ((~g15426));
assign g18738 = (g15142&g16826);
assign g15779 = (g13909&g11214);
assign g33957 = (g33523)|(II31868)|(II31869);
assign g22003 = (g5736&g21562);
assign g21845 = (g3881&g21070);
assign II20412 = ((~g16213));
assign g33333 = (g32218&g20612);
assign II31067 = (g32552&g32553&g32554&g32555);
assign II25594 = ((~g25531));
assign g30464 = (g30152)|(g21935);
assign g16258 = (g13247)|(g10856);
assign II22580 = ((~g20982));
assign g13155 = (g11496)|(g11546);
assign g34952 = ((~g34942));
assign g18151 = (g617&g17533);
assign g20899 = ((~II20861));
assign g9820 = ((~g99));
assign g15817 = (g3921&g13929);
assign g28544 = (g27300)|(g26229);
assign g28692 = (g27578&g20661);
assign g23253 = ((~g21037));
assign g34461 = (g34291)|(g18681);
assign II15564 = ((~g11949));
assign g9933 = ((~g5759));
assign g20321 = ((~g17821));
assign g18242 = (g962&g16431);
assign g16510 = ((~g14008));
assign g24682 = (g22662&g19754);
assign g18091 = ((~II18879));
assign g34820 = ((~II33034));
assign g7212 = ((~g6411));
assign g13573 = ((~g8002))|((~g10544))|((~g7582))|((~g1351));
assign g27394 = (g25957)|(g24573);
assign g14700 = ((~g12512));
assign g25527 = ((~g21294))|((~g23462));
assign g29564 = (g1882&g28896);
assign g26310 = (g2102&g25389);
assign g10172 = ((~g6459));
assign g19763 = ((~g16431));
assign II20187 = ((~g16272))|((~g1333));
assign g30009 = (g29034&g10518);
assign g16288 = ((~g13794)&(~g417));
assign g34571 = (g27225&g34299);
assign g12901 = ((~g10404));
assign g27627 = (g13266&g25790);
assign g27560 = (g26299&g20191);
assign g34053 = ((~g33683));
assign g11944 = ((~II14765))|((~II14766));
assign g26515 = ((~g24843)&(~g24822));
assign g33510 = (g32816&II31246&II31247);
assign g34767 = ((~II32947));
assign g24217 = (g18200&g22594);
assign gbuf77 = (g3321);
assign g31874 = (g31016)|(g21729);
assign g23346 = (g19736)|(g16204);
assign g21704 = (g164&g20283);
assign g34611 = (g34508)|(g18565);
assign g22649 = ((~g19063));
assign g11729 = ((~g3179)&(~g8059));
assign g18571 = (g2856&g16349);
assign g25174 = ((~g23890));
assign g27381 = ((~g8075)&(~g26657));
assign g25328 = (g5022&g23764&II24505);
assign g18407 = (g2016&g15373);
assign g26881 = (g26629)|(g24187);
assign g16207 = (g9839&g14204);
assign g31802 = ((~g29385));
assign g19996 = ((~g17271));
assign g9339 = ((~g2295));
assign g33794 = (g33126)|(g32053);
assign g14193 = (g7178&g10590);
assign g10031 = ((~II13552));
assign g6830 = ((~g1389));
assign g13854 = ((~g4765))|((~g11797));
assign g13886 = ((~g11804))|((~g4922));
assign g12479 = ((~g2028)&(~g8310));
assign g10805 = ((~II14046));
assign g23767 = ((~g18997));
assign g15146 = ((~g13716)&(~g7003));
assign g33462 = (g32470&II31006&II31007);
assign g9086 = ((~g847));
assign g6839 = ((~g1858));
assign g12336 = ((~II15175))|((~II15176));
assign g26101 = (g1760&g25098);
assign g34647 = (g34558)|(g18820);
assign g8821 = ((~II12811));
assign g24677 = ((~g22957))|((~g2975));
assign g11964 = ((~g9154));
assign g23428 = ((~g13945))|((~g20522));
assign g34148 = (g33758)|(g19656);
assign g33251 = (g32096)|(g29509);
assign g27511 = ((~g22137)&(~g26866)&(~g20277));
assign g18304 = (g1542&g16489);
assign g27388 = (g26519&g17502);
assign g13494 = ((~g11912));
assign g33866 = (g33276&g20528);
assign g23760 = ((~II22889));
assign g32140 = (g31609&g29961);
assign g7197 = ((~g812));
assign g27720 = ((~g9253)&(~g25791));
assign g12834 = ((~g10349));
assign g10869 = (g7766&g5873&g5881);
assign g22644 = (g18981)|(g15632);
assign g24397 = ((~g22908));
assign g27010 = ((~g6052)&(~g25839));
assign g25693 = (g24627)|(g18707);
assign g29684 = (g1982&g29085);
assign g26251 = (g1988&g25341);
assign g15795 = (g3566&g14130);
assign II13252 = ((~g6751));
assign g27357 = (g26400&g17414);
assign g18662 = (g15126&g17367);
assign II18205 = ((~g14563));
assign g7670 = ((~g4104));
assign g33965 = (g33805)|(g18179);
assign g27250 = (g25901)|(g15738);
assign II24684 = (g20014&g24033&g24034&g24035);
assign g13296 = (g10626)|(g10657);
assign II31122 = (g32631&g32632&g32633&g32634);
assign II18379 = ((~g13012));
assign g26822 = (g24841&g13116);
assign II18894 = ((~g16708));
assign g29580 = (g28519&g14186);
assign g9551 = ((~g3281));
assign g14816 = ((~g10166)&(~g12252));
assign g34017 = (g33880)|(g18504);
assign II13744 = ((~g3518));
assign g22852 = ((~g18957))|((~g2856));
assign g28706 = (g27584&g20681);
assign g34306 = (g25782)|(g34054);
assign g20579 = ((~g17249));
assign g34298 = (g8679&g34132);
assign g13266 = ((~g12440))|((~g9920))|((~g9843));
assign g19475 = (g16930)|(g14126);
assign g32908 = ((~g31327));
assign g11626 = ((~g7121)&(~g3863)&(~g3857));
assign g15838 = (g3602&g14133);
assign g23874 = ((~g18997));
assign g8718 = ((~g3333));
assign II31838 = (g33461)|(g33462)|(g33463)|(g33464);
assign g24699 = ((~g23047));
assign g10275 = ((~g4584));
assign g32233 = (g31150)|(g29661);
assign g28906 = ((~g27796))|((~g8150));
assign g32628 = ((~g31542));
assign II28147 = (g2946)|(g24561)|(g28220);
assign II17154 = ((~g13605));
assign II17819 = ((~g3618));
assign g9310 = ((~II13078))|((~II13079));
assign g18492 = (g2523&g15426);
assign g17493 = ((~g8659))|((~g14367));
assign g11720 = ((~II14589));
assign g20101 = ((~g17533));
assign g24649 = (g6527&g23733);
assign g10414 = ((~g7092));
assign g15345 = ((~II17108));
assign g14168 = (g887&g10632);
assign g15060 = ((~g13350)&(~g6814));
assign g33010 = (g32301)|(g18473);
assign g22406 = ((~g19506));
assign II24482 = (g9364&g9607&g5057);
assign g15585 = ((~g11862)&(~g14194));
assign g29299 = (g28587)|(g18794);
assign g27584 = (g26165)|(g24758);
assign g9091 = ((~g1430));
assign g11961 = ((~g9777))|((~g5105));
assign g24121 = ((~g20720));
assign g12443 = ((~g9374)&(~g9300));
assign II17448 = ((~g956))|((~II17446));
assign g27684 = (g26386&g20657);
assign g16821 = ((~II18031));
assign g28173 = ((~II26693));
assign g23815 = ((~g19074));
assign g15030 = ((~g12716))|((~g12680));
assign g8764 = ((~g4826));
assign II24384 = ((~g23721))|((~II24383));
assign g27581 = (g26161)|(g24750);
assign g23745 = ((~g20900));
assign g34170 = (g33790)|(g19855);
assign g18516 = (g2638&g15509);
assign g7566 = ((~II12049));
assign g25185 = ((~g22228));
assign II15242 = ((~g10003))|((~II15241));
assign g19750 = ((~g16326));
assign g13131 = ((~g6243))|((~g12101))|((~g6377))|((~g10003));
assign g31483 = ((~g4899)&(~g29725));
assign g32592 = ((~g30673));
assign g30432 = (g29888)|(g21816);
assign g8240 = ((~g1333));
assign II12902 = (g4235)|(g4232)|(g4229)|(g4226);
assign g23666 = ((~g20875))|((~g11139));
assign g32963 = ((~g30825));
assign g29265 = (g28318)|(g18620);
assign II17181 = ((~g13745));
assign g19904 = (g17636)|(g14654);
assign II26461 = ((~g14306))|((~II26459));
assign g31185 = (g10114&g30087);
assign g26023 = (g9528&g25036);
assign g33295 = (g32153)|(g29605);
assign g31117 = ((~g4991)&(~g29556));
assign g32950 = ((~g31672));
assign g8449 = ((~g3752));
assign g16594 = ((~II17772));
assign g32160 = (g31001&g22995);
assign II15284 = ((~g6697));
assign g17591 = ((~II18526));
assign g33296 = (g32156)|(g29617);
assign g23263 = ((~II22366));
assign g32894 = ((~g30614));
assign g10611 = ((~g10115))|((~g9831));
assign g14915 = ((~g12553))|((~g10266));
assign II33235 = ((~g34957));
assign g25283 = ((~g22763));
assign g19887 = ((~g3025)&(~g16275));
assign g18935 = (g4322&g15574);
assign g32683 = ((~g30614));
assign g29725 = ((~g28349));
assign g18128 = (g504&g16971);
assign g14636 = ((~g5595))|((~g12029))|((~g5677))|((~g12563));
assign II14033 = ((~g8912));
assign II17695 = ((~g14330));
assign g14181 = ((~g9083)&(~g12259));
assign g29656 = (g28515&g11666);
assign g18335 = (g1687&g17873);
assign g15737 = ((~g13240))|((~g13115))|((~g7903))|((~g13210));
assign II12899 = ((~g4232));
assign g20993 = ((~g15615));
assign g33421 = (g32374&g21455);
assign II26049 = ((~g25997))|((~g13500));
assign g18419 = (g2051&g15373);
assign II16486 = ((~g11204));
assign g24988 = ((~g546))|((~g23088));
assign g12109 = ((~II14967));
assign g27880 = ((~II26427));
assign g18271 = (g1296&g16031);
assign g26486 = (g4423&g24358);
assign g17216 = ((~g14454));
assign g32981 = (g32425)|(g18206);
assign g34489 = (g34421&g19068);
assign g18740 = (g4572&g17384);
assign g34665 = (g34583&g19067);
assign g17503 = ((~g14892));
assign g31932 = (g31792)|(g22107);
assign g12563 = ((~g9864));
assign II29279 = ((~g12081))|((~II29277));
assign g8783 = ((~II12761));
assign g24625 = ((~g23135));
assign II25736 = (g12)|(g22150)|(g20277);
assign g27085 = (g25835&g22494);
assign g18474 = (g2287&g15224);
assign g27276 = (g9750&g26607);
assign g21811 = (g3582&g20924);
assign g32507 = ((~g30735));
assign g22663 = ((~II21977))|((~II21978));
assign II21722 = ((~g19264));
assign g28702 = (g27457)|(g16670);
assign g34186 = (g33705&g24396);
assign g26924 = (g26153)|(g18291);
assign g24084 = ((~g20720));
assign g31915 = (g31520)|(g22001);
assign g30046 = (g29108&g10564);
assign g6956 = ((~g4242));
assign g7224 = ((~g4601));
assign g23357 = ((~g20201))|((~g11231));
assign g32454 = (g30322)|(g31795);
assign g23799 = (g14911&g21279);
assign g7753 = ((~II12183));
assign g7835 = ((~g4125));
assign g17189 = ((~g14708));
assign II20385 = ((~g16194));
assign II12003 = ((~g767));
assign g24105 = ((~g19935));
assign g28745 = (g27519)|(g16760);
assign g15853 = ((~g14714))|((~g9417))|((~g12337));
assign g21929 = (g5176&g18997);
assign g29530 = (g1612&g28820);
assign g24035 = ((~g20841));
assign g23041 = ((~g19882));
assign g23379 = ((~g20216))|((~g11248));
assign g25970 = (g1792&g24991);
assign g21906 = (g5022&g21468);
assign g21824 = (g3706&g20453);
assign g18544 = (g2791&g15277);
assign g34482 = (g34405&g18917);
assign gbuf18 = (g5276);
assign g20026 = ((~g17271));
assign g10307 = ((~II13730))|((~II13731));
assign g22859 = (g9456&g20734);
assign II30986 = ((~g32437));
assign g24260 = (g23373)|(g18313);
assign g19350 = (g15968&g13505);
assign g26285 = (g1834&g25300);
assign g24295 = (g4434&g22550);
assign g12053 = ((~g2587))|((~g8418));
assign g24547 = ((~g22638))|((~g22643))|((~g22754));
assign g34470 = (g7834&g34325);
assign g14712 = ((~g12479)&(~g9971));
assign g31969 = (g31189&g22139);
assign g20563 = ((~g15171));
assign g18210 = (g936&g15938);
assign g27972 = (g26131)|(g26105);
assign g12411 = ((~g7393))|((~g5276));
assign g22023 = (g5881&g19147);
assign g34961 = (g34944&g23019);
assign g24399 = (g3133&g23067);
assign g31865 = (g31149)|(g21709);
assign g20009 = ((~g16349));
assign g21950 = (g5268&g18997);
assign g25243 = ((~g22763));
assign g12436 = ((~II15263))|((~II15264));
assign g31894 = (g30671)|(g21870);
assign g33582 = (g33351)|(g18444);
assign g19675 = ((~g16987));
assign II22502 = ((~g19376));
assign g32399 = (g31527)|(g30062);
assign g18121 = (g424&g17015);
assign II25790 = ((~g26424));
assign g26969 = (g26313)|(g24329);
assign g22009 = (g5782&g21562);
assign g13620 = ((~g10556));
assign g20593 = ((~g15277));
assign g27831 = ((~II26406));
assign g27091 = ((~g26725));
assign g22976 = ((~II22149));
assign g14608 = (g12638&g12476&g12429&II16721);
assign g18978 = ((~g16000));
assign g32205 = (g30922&g28463);
assign g19679 = ((~g16782));
assign g24333 = (g4512&g22228);
assign g31138 = ((~g29778));
assign g24220 = (g255&g22594);
assign II12782 = (g4188)|(g4194)|(g4197)|(g4200);
assign g25951 = (g24500&g19565);
assign g15372 = ((~g817)&(~g14279));
assign g25142 = (g4717&g22885);
assign g24054 = ((~g19919));
assign g13584 = ((~g12735));
assign g9234 = ((~g5170));
assign g25182 = ((~g22763));
assign g31812 = ((~g29385));
assign g18114 = (g452&g17015);
assign II32659 = ((~g34391));
assign g16746 = ((~g14258));
assign II23694 = ((~g23252));
assign g21287 = ((~g14616))|((~g17571));
assign g10347 = ((~II13759));
assign g8790 = (II12782)|(II12783);
assign g15745 = (g686&g13223);
assign g34844 = ((~g34737));
assign g11852 = ((~II14668));
assign g23020 = ((~g19869));
assign g23208 = ((~g20035)&(~g16324));
assign II32452 = ((~g34241));
assign g19532 = ((~g16821));
assign g16281 = ((~g4754))|((~g13937))|((~g12054));
assign g31974 = (g31760&g22176);
assign g11996 = ((~g7280))|((~g2197));
assign g23921 = (g19379&g4146);
assign g25979 = (g24517&g19650);
assign g22032 = (g5921&g19147);
assign II18626 = ((~g2079))|((~II18625));
assign g21338 = ((~g15741))|((~g15734))|((~g15728))|((~g13097));
assign g13474 = ((~g11048));
assign g23372 = (g16448&g20194);
assign g17062 = ((~II18154));
assign g18276 = (g1351&g16136);
assign II31331 = (g30825&g31854&g32933&g32934);
assign g16221 = (g5791&g14231);
assign g13897 = ((~g3211))|((~g11217))|((~g3329))|((~g11519));
assign g7327 = ((~g2165));
assign g28159 = (g8553&g27317);
assign g9649 = ((~g2227)&(~g2153));
assign g34403 = (g34180)|(g25085);
assign II20216 = ((~g15862));
assign g34435 = ((~II32476));
assign g31282 = (g30130&g27779);
assign g20135 = (g16258&g16695);
assign II33158 = ((~g34897));
assign g18550 = (g2819&g15277);
assign g18328 = (g1657&g17873);
assign g34320 = ((~g34119));
assign g15166 = ((~g13835)&(~g7096));
assign g28599 = (g27027&g8922);
assign II33053 = ((~g34778));
assign g29380 = (g28134&g19396);
assign II14277 = ((~g3484))|((~II14275));
assign II13166 = ((~g5101));
assign g34761 = (g34679)|(g34506);
assign gbuf110 = (g4200);
assign g21347 = (g1339&g15750);
assign g28049 = (g27684)|(g18164);
assign g25784 = ((~g25507)&(~g25485));
assign II20750 = ((~g16677));
assign g20233 = ((~g17873));
assign g12187 = ((~II15042))|((~II15043));
assign g33978 = (g33892)|(g18356);
assign g32273 = (g31255&g20446);
assign g32563 = ((~g31554));
assign g29653 = ((~II27927));
assign g27662 = ((~II26296));
assign g32170 = (g31671&g27779);
assign g24945 = (g23183&g20197);
assign g7520 = (g2704&g2697&g2689);
assign g12301 = ((~II15148))|((~II15149));
assign g26802 = ((~II25514));
assign g9546 = ((~g2437));
assign g27043 = (g26335&g8632);
assign II33064 = ((~g34784));
assign II32770 = ((~g34505));
assign g24195 = (g74&g22722);
assign g19431 = ((~g16249));
assign g18569 = (g94&g16349);
assign g33915 = (g33140&g7846);
assign g28774 = (g27536)|(g16804);
assign g24439 = ((~g7400)&(~g22312));
assign g16197 = ((~g13861));
assign II15843 = ((~g11181));
assign g18127 = (g499&g16971);
assign g21947 = (g5256&g18997);
assign g11708 = ((~g10147))|((~g10110));
assign g11955 = ((~g8302))|((~g1917));
assign g25559 = (g13004&g22649);
assign g24974 = ((~g21301))|((~g23363));
assign g33869 = (g33279&g20543);
assign g28534 = (g27292)|(g26204);
assign g22900 = (g17137&g19697);
assign g23312 = ((~g21070));
assign g25084 = (g4737&g22885);
assign g21404 = (g16069&g13569);
assign g22152 = (g21188)|(g17469);
assign g17500 = ((~g14573))|((~g14548));
assign g11972 = ((~g9591)&(~g7361));
assign g17485 = ((~II18408));
assign g32475 = ((~g30614));
assign g20235 = ((~g15277));
assign g30227 = (g28708&g23899);
assign g18532 = (g2724&g15277);
assign g12539 = ((~II15341))|((~II15342));
assign g24914 = (g8721&g23301);
assign g30301 = ((~II28548));
assign II16590 = ((~g11966));
assign g19603 = ((~g16349));
assign II31082 = (g32573&g32574&g32575&g32576);
assign g30494 = (g30209)|(g21990);
assign II21254 = ((~g16540));
assign g34185 = (g33702&g24389);
assign g12044 = ((~g1657))|((~g8139));
assign g10124 = ((~g5276))|((~g5320))|((~g5290))|((~g5313));
assign II12253 = ((~g1129))|((~II12251));
assign g33593 = (g33417)|(g18482);
assign g32105 = (g4922&g30673);
assign g34523 = (g9162&g34351);
assign g32923 = ((~g31021));
assign g20052 = ((~g17533));
assign g20536 = ((~g18065));
assign g21509 = ((~g17820))|((~g14898))|((~g17647))|((~g17608));
assign g16602 = ((~g14101));
assign g25645 = (g24679)|(g21738);
assign g27309 = (g26603&g23057);
assign g34686 = (g34494&g19494);
assign g18386 = (g1964&g15171);
assign g11038 = ((~g8632));
assign II27677 = ((~g28156));
assign II18852 = ((~g13716));
assign g18787 = (g15158&g15634);
assign g24387 = (g3457&g22761);
assign g33129 = ((~g8630)&(~g32072));
assign g32346 = (g29838)|(g31272);
assign g23523 = ((~g21514));
assign g29176 = (g27661)|(g17177);
assign g29642 = (g27954&g28669);
assign g9299 = ((~g5124));
assign g24306 = (g4483&g22228);
assign II26366 = ((~g26400))|((~g14211));
assign g17760 = ((~II18752));
assign g29354 = (g4961&g28421);
assign g32691 = ((~g30673));
assign g34364 = (g34048&g24366);
assign g23626 = ((~g17309)&(~g20854));
assign g26231 = (g1854&g25300);
assign g12735 = (g7121&g3873&g3881);
assign II13336 = ((~g1691))|((~II13334));
assign g17782 = ((~II18788));
assign g32048 = (g31498&g13869);
assign g17510 = (g14393)|(g14362)|(g11972)|(II18449);
assign g34642 = (g34482)|(g18725);
assign g7235 = ((~g4521));
assign II15981 = ((~g11290));
assign g24138 = ((~g21143));
assign II16564 = ((~g10429));
assign g24762 = (g655&g23573);
assign g28620 = ((~g27679));
assign g27208 = (g9037&g26598);
assign g15870 = (g3231&g13948);
assign g19502 = ((~g15674));
assign g24073 = ((~g21127));
assign g34827 = ((~II33041));
assign g28090 = (g27275)|(g18733);
assign g15710 = ((~g319))|((~g13385));
assign g7640 = ((~II12128));
assign g23955 = ((~g2823)&(~g18890));
assign II28572 = ((~g28274));
assign g8124 = ((~II12402))|((~II12403));
assign g27858 = (g17405)|(g26737);
assign g30547 = (g30194)|(g22118);
assign g33362 = (g32259&g20914);
assign g29964 = (g2008&g28830);
assign II12730 = ((~g4287))|((~II12728));
assign g32806 = ((~g31710));
assign g18583 = (g2936&g16349);
assign g34809 = (g33677)|(g34738);
assign g25610 = (g24923)|(g18127);
assign g30348 = (g30083)|(g18329);
assign g32329 = ((~g31522));
assign g12180 = ((~g9477));
assign II31983 = ((~g33653))|((~g33648));
assign g33706 = (g32412)|(g33440);
assign g32212 = ((~g8859)&(~g31262)&(~g11083));
assign II32973 = ((~g34714));
assign g27538 = (g26549&g14744);
assign g30385 = (g30172)|(g18518);
assign g27247 = (g2759&g26745);
assign g20218 = (g6541&g17815);
assign g29184 = ((~g9631)&(~g26994));
assign g32909 = ((~g30614));
assign g14157 = ((~g11715))|((~g11763));
assign g18641 = (g3841&g17096);
assign g24379 = ((~g22550));
assign g26934 = (g26845)|(g18556);
assign II12470 = ((~g392))|((~II12468));
assign g29539 = (g2864)|(g28220);
assign g28953 = ((~g5170)&(~g27999));
assign g13051 = ((~g11964));
assign g28435 = (g27234)|(g15967);
assign g27489 = (g24608)|(g26022);
assign g27326 = (g12048&g26731);
assign g8107 = ((~g3179));
assign g25563 = ((~g22594));
assign g9777 = ((~g5112));
assign g13304 = ((~II15872));
assign g34638 = (g34484)|(g18721);
assign g23870 = ((~g21293));
assign gbuf53 = (g6346);
assign g28270 = ((~g10504))|((~g26105))|((~g26987));
assign g33787 = (g33103&g20595);
assign g12113 = ((~g1648)&(~g8187));
assign g7170 = ((~g5719));
assign g20270 = ((~g15277));
assign g8903 = ((~g1075));
assign g23400 = ((~g20676));
assign g24566 = ((~g22755))|((~g22713));
assign g28528 = (g27187&g12730);
assign g21955 = (g5385&g21514);
assign g24320 = (g6973&g22228);
assign g14397 = ((~g12120)&(~g9416));
assign g25878 = (g25503)|(g23920);
assign g23571 = ((~g18833));
assign g18390 = (g1978&g15171);
assign g22513 = ((~g1002)&(~g19699));
assign g32033 = ((~g30929));
assign g29152 = ((~g27907));
assign g17607 = ((~II18560));
assign II19661 = ((~g17587));
assign II31237 = (g32798&g32799&g32800&g32801);
assign g29847 = ((~g28395));
assign II12030 = ((~g595));
assign g27963 = (g25952&g16047);
assign g9000 = ((~g632));
assign g27304 = (g2273&g26682);
assign g26977 = (g23032&g26261&g26424&g25550);
assign g15050 = ((~g12834)&(~g13350));
assign g18101 = ((~II18909));
assign g27267 = (g26026&g17124);
assign g33721 = (g33163&g19440);
assign g34029 = (g33798)|(g18703);
assign g9012 = (g2047)|(g2066);
assign g10502 = ((~g8876));
assign g32859 = ((~g30614));
assign g26177 = (g2079&g25154);
assign g21858 = (g3937&g21070);
assign g25040 = (g12738&g23443);
assign g34632 = (g34565)|(g15119);
assign g25201 = (g12346&g23665);
assign g16882 = (g13508)|(g11114);
assign g26949 = (g26356)|(g24287);
assign g9904 = ((~II13443))|((~II13444));
assign g31773 = (g30044)|(g30056);
assign g16845 = (g6593&g15011);
assign g14150 = ((~g12381));
assign g33805 = (g33232&g20079);
assign g7577 = ((~g1263));
assign g23407 = (g9295&g20273);
assign g20572 = ((~g15833));
assign II31266 = (g31327&g31843&g32838&g32839);
assign g17321 = (g1418&g13105);
assign g26650 = (g10796&g24424);
assign II29248 = ((~g29491));
assign g28660 = (g27824&g20623);
assign g12875 = ((~II15494));
assign g21973 = (g5511&g19074);
assign g18690 = (g15130&g16053);
assign g11017 = ((~g10289));
assign g18908 = ((~g16100));
assign g23019 = ((~g19866));
assign g9833 = ((~g2449));
assign g11930 = ((~g9281));
assign II32687 = ((~g34431));
assign II14450 = ((~g4191));
assign g26861 = (g25021&g25003);
assign g33369 = (g32277&g21060);
assign g13030 = (g429&g11048);
assign g17691 = ((~II18674));
assign II13280 = ((~g6140));
assign g20090 = ((~g17433));
assign g18804 = (g15163&g15656);
assign II18469 = ((~g13809));
assign g27280 = (g9825&g26614);
assign II17879 = ((~g14386));
assign g20064 = ((~g17533));
assign g12244 = ((~g7343))|((~g5320));
assign g20076 = ((~g13795))|((~g16521));
assign g30393 = (g29986)|(g21748);
assign g21666 = ((~g16540));
assign g32308 = (g31293&g23503);
assign g27931 = ((~g25425))|((~g25381))|((~g25780));
assign g7410 = ((~g2008));
assign g29735 = (g28202)|(g10898);
assign g18251 = (g996&g16897);
assign II13857 = ((~g9780));
assign g34167 = (g33786)|(g19768);
assign g25021 = ((~g21417))|((~g23363));
assign g10738 = ((~g6961))|((~g10308));
assign g33497 = (g32723&II31181&II31182);
assign g19570 = ((~g16349));
assign II32681 = ((~g34429));
assign g34587 = ((~II32671));
assign g9037 = ((~g164));
assign g18709 = (g59&g17302);
assign g30236 = (g28724&g23916);
assign g29865 = (g1802&g29115);
assign g25309 = ((~g22384))|((~g12021));
assign g24965 = (g22667)|(g23825);
assign g28910 = ((~g27854))|((~g14614));
assign g33834 = (g33095&g29172);
assign gbuf143 = (g1582);
assign g30033 = (g29189&g12937);
assign g26666 = ((~g9229))|((~g25144));
assign II17404 = ((~g13378))|((~g1472));
assign g32407 = ((~II29939));
assign g32243 = (g31166)|(g29683);
assign II12837 = ((~g4222));
assign g20664 = ((~g15373));
assign g31909 = (g31750)|(g21956);
assign g21326 = ((~II21058));
assign g26709 = ((~g25435));
assign g8509 = ((~g4141));
assign g29927 = ((~g28861));
assign g28193 = (g8851&g27629);
assign g28627 = (g27543&g20574);
assign g12073 = ((~g10058))|((~g6490));
assign g34454 = (g34414)|(g18667);
assign g20530 = ((~g15509));
assign g13009 = ((~II15617));
assign g22312 = ((~g907))|((~g19063));
assign g29193 = ((~g9529)&(~g26994)&(~g7812));
assign g16655 = ((~g14151));
assign g32087 = (g1291&g30825);
assign g31886 = (g31481)|(g21791);
assign g8644 = ((~g3352));
assign g26048 = (g5853&g25044);
assign g30485 = (g30166)|(g21981);
assign g17707 = ((~g14758));
assign g23056 = (g16052&g19860);
assign II15872 = ((~g11236));
assign g28714 = (g27591&g20711);
assign g7553 = ((~g1274));
assign g24496 = (g24008)|(g21557);
assign II25530 = ((~g25222));
assign II31017 = (g32480&g32481&g32482&g32483);
assign g10755 = ((~g7352))|((~g7675))|((~g1322))|((~g1404));
assign g17811 = ((~g12925));
assign g16027 = ((~g10929)&(~g13260));
assign g22089 = (g6311&g19210);
assign g25049 = ((~g21344))|((~g23462));
assign II32884 = ((~g34690));
assign g7175 = ((~g6098)&(~g6058));
assign g12588 = ((~g10169))|((~g6336))|((~g6386));
assign g18360 = (g1830&g17955);
assign g7834 = (g2886)|(g2946);
assign g31474 = (g29668)|(g13583);
assign g34369 = (g26279)|(g34136);
assign g22039 = (g5949&g19147);
assign g15113 = (g4291&g14454);
assign g34031 = (g33735)|(g18705);
assign g25195 = ((~g22763));
assign g21419 = (g16681&g13595);
assign g14687 = ((~g5352)&(~g12166));
assign g12700 = ((~g9321)&(~g5857));
assign g17489 = ((~g12955));
assign g11819 = ((~g7717));
assign II21067 = ((~g15573));
assign II17916 = ((~g13087));
assign g34273 = (g27765)|(g34203);
assign g25562 = ((~g22763));
assign g34739 = ((~II32909));
assign g34321 = (g25866)|(g34065);
assign g17577 = ((~II18504));
assign g20111 = ((~g17513))|((~g14517))|((~g17468))|((~g14422));
assign g28042 = (g24148)|(g26879);
assign II16231 = ((~g10520));
assign II23985 = ((~g22182))|((~g482));
assign g23449 = ((~g18833));
assign g10155 = ((~g2643));
assign g22493 = ((~g19801));
assign g29705 = ((~g28399)&(~g8284)&(~g8404));
assign g12872 = ((~g10379));
assign g16739 = ((~g13223));
assign g18438 = (g2236&g18008);
assign g26276 = (g2461&g25476);
assign g18429 = (g2193&g18008);
assign g32992 = (g32242)|(g18351);
assign g13272 = ((~II15837));
assign g29858 = (g28387&g23306);
assign g29864 = (g28272)|(g26086);
assign g25308 = ((~g22763));
assign g33550 = (g33342)|(g18338);
assign g21365 = ((~g15744))|((~g13119))|((~g15730))|((~g13100));
assign g21982 = (g5547&g19074);
assign g32634 = ((~g30673));
assign g21221 = ((~g15680));
assign g15045 = ((~g12716))|((~g7142));
assign g28213 = (g27720&g23380);
assign g25356 = ((~g22763));
assign g19469 = ((~g16326));
assign g33399 = (g32346&g21379);
assign g27711 = (g22369&g25193&g26424&g26166);
assign g22658 = ((~II21969));
assign g20655 = ((~II20753));
assign g7396 = (g392&g441);
assign g25267 = ((~g22228));
assign g32287 = (g2823&g30578);
assign g20391 = ((~II20562));
assign g31000 = ((~g29737));
assign g23651 = ((~g20655));
assign g15746 = ((~g13121));
assign g23121 = (g19128&g9104);
assign g34236 = (g32650)|(g33954);
assign II18897 = ((~g16738));
assign g30254 = (g28747&g23944);
assign g18579 = (g2984&g16349);
assign g30190 = (g28646&g23842);
assign g21989 = (g5587&g19074);
assign g15796 = (g3586&g14015);
assign g21909 = (g5041&g21468);
assign g28969 = ((~g27854))|((~g8267));
assign g7963 = ((~g4146));
assign g9946 = ((~g6093));
assign g14332 = ((~II16492));
assign g30732 = (g13778)|(g29762);
assign g22308 = (g1135&g19738);
assign II28883 = ((~g30105));
assign g12546 = ((~g8740));
assign II16688 = ((~g10981));
assign g21190 = ((~g6077))|((~g17420));
assign g19333 = (g464&g16223);
assign g25518 = (g6444&g23865&II24625);
assign g25068 = (g17574&g23477);
assign II13552 = ((~g121));
assign II18900 = ((~g16767));
assign g13541 = (g7069&g12308);
assign g11615 = ((~g6875));
assign g34289 = (g26847)|(g34218);
assign g7511 = (g2145&g2138&g2130);
assign g32753 = ((~g30735));
assign g31927 = (g31500)|(g22091);
assign g22118 = (g6605&g19277);
assign II19813 = ((~g17952));
assign g17784 = (g1152&g13215);
assign II18587 = ((~g2370))|((~g14679));
assign g16600 = ((~II17780));
assign II17763 = ((~g13191));
assign g21460 = ((~g15628));
assign g25911 = (g22514)|(g24510);
assign g16586 = ((~g13851))|((~g13823));
assign g15277 = ((~II17104));
assign g8431 = ((~g3085));
assign g21384 = ((~g17734))|((~g14686))|((~g17675))|((~g14663));
assign g17870 = ((~II18842));
assign g25054 = (g12778&g23452);
assign g32542 = ((~g31554));
assign g16607 = ((~g13960));
assign g15709 = ((~g5224))|((~g14399))|((~g5327))|((~g9780));
assign g34781 = (g33431)|(g34715);
assign g23639 = (g19050&g9104);
assign g29777 = (g28227)|(g28234);
assign II31829 = ((~g33454));
assign g7647 = ((~II12132));
assign II23300 = ((~g21665));
assign g29772 = (g28323&g23243);
assign II12497 = ((~g49));
assign g33641 = ((~II31474));
assign g34604 = (g34563)|(g15076);
assign g30250 = (g28744&g23939);
assign g21055 = ((~g15224));
assign g24849 = (g4165&g22227);
assign g12711 = ((~g6209)&(~g9326));
assign g23128 = ((~g20283));
assign g12013 = ((~II14866));
assign g22044 = (g6058&g21611);
assign g31776 = (g21329&g29385);
assign g27926 = ((~g9467)&(~g25856));
assign g30128 = (g28495)|(g11497);
assign II22794 = ((~g21434))|((~II22792));
assign g17391 = (g9556&g14378);
assign g10224 = ((~g6661))|((~g6704))|((~g6675))|((~g6697));
assign g11744 = ((~II14602));
assign g9875 = ((~g5747));
assign II24089 = ((~g22409));
assign g13250 = ((~II15811));
assign g27453 = (g25976)|(g24606);
assign g18764 = (g5485&g17929);
assign g13345 = (g4754&g11773);
assign II23979 = ((~g23198))|((~II23978));
assign g12288 = ((~g2610)&(~g8418));
assign g23855 = (g4112&g19455);
assign g20211 = ((~g16931));
assign g28717 = (g27482)|(g16701);
assign g34000 = (g33943)|(g18441);
assign g15066 = ((~g12841)&(~g13394));
assign g28497 = (g27267)|(g16199);
assign g24366 = ((~g22594));
assign g29995 = ((~g28955));
assign g25679 = (g24728)|(g21836);
assign g19777 = ((~g17015));
assign g32301 = (g31276&g20547);
assign g31490 = (g29786&g23429);
assign g32529 = ((~g30735));
assign g20763 = ((~II20816));
assign g29079 = ((~g27742));
assign II26925 = ((~g27015));
assign g9332 = ((~g64));
assign II18092 = ((~g3668));
assign g34806 = (g34763)|(g18595);
assign g23293 = (g9104&g19200);
assign g29013 = ((~II27368));
assign g17587 = ((~II18518));
assign g19873 = ((~g15755)&(~g1395));
assign g28688 = (g27435)|(g16639);
assign g34917 = ((~II33143));
assign g33786 = (g33130&g20572);
assign g34251 = (g34157)|(g18147);
assign g11193 = ((~II14258))|((~II14259));
assign gbuf109 = (g4197);
assign II23333 = ((~g22683));
assign g29713 = ((~II27970));
assign II32079 = ((~g33937));
assign II12346 = ((~g3111))|((~II12344));
assign g28238 = (g27133&g19658);
assign g12234 = ((~g9776)&(~g9778));
assign II20166 = ((~g16246))|((~II20165));
assign g26098 = ((~g9073)&(~g24732));
assign g7518 = ((~g1024));
assign g28139 = (g27337&g26054);
assign g19862 = ((~II20233));
assign II20910 = ((~g17197));
assign g29149 = ((~g27837));
assign g14306 = ((~g10060)&(~g10887));
assign g17178 = ((~II18214));
assign g25885 = (g25522)|(g23957);
assign g24042 = ((~g20014));
assign g11544 = ((~g8700))|((~g3990))|((~g4045));
assign g7885 = ((~II12270))|((~II12271));
assign g31002 = (g29362)|(g28154);
assign g10598 = ((~g7191))|((~g6404));
assign g28813 = (g4104&g27038);
assign g30553 = (g30205)|(g22124);
assign g21381 = ((~g18008));
assign g23755 = (g14821&g21204);
assign g34592 = ((~II32684));
assign g30278 = (g28818&g23988);
assign g33920 = ((~II31786));
assign g7142 = ((~g6573)&(~g6565));
assign g30914 = (g29873&g20887);
assign g9007 = ((~g1083));
assign g19504 = ((~g16349));
assign II13334 = ((~g1687))|((~g1691));
assign g32708 = ((~g31376));
assign g10385 = ((~II13805));
assign g31960 = (g31749&g22153);
assign g27438 = ((~II26130));
assign g29806 = (g28358&g23271);
assign g18298 = (g15073&g16489);
assign g30404 = (g29758)|(g21763);
assign g25663 = (g24666)|(g21788);
assign g20626 = ((~g15483));
assign g27404 = (g26400&g17518);
assign g17777 = ((~g14908));
assign g17424 = (g1426&g13176);
assign g34265 = (g34117)|(g18711);
assign g19717 = (g6527&g17122);
assign g10961 = ((~g1442))|((~g7876));
assign g22679 = (g19145)|(g15701);
assign g18466 = (g2389&g15224);
assign g28089 = (g27269)|(g18731);
assign g30449 = (g29845)|(g21858);
assign g16971 = ((~II18131));
assign g29944 = ((~g28911));
assign g25628 = (g24600)|(g18249);
assign g11170 = ((~g8476));
assign g16620 = ((~II17808));
assign II22889 = ((~g18926));
assign g28796 = ((~g27858))|((~g7418))|((~g7335));
assign g31267 = (g29548)|(g28263);
assign g12343 = ((~g7470))|((~g5630));
assign g28231 = (g27187&g22763&g27074);
assign g17653 = (g11547&g11592&g6789&II18620);
assign gbuf102 = (g3798);
assign g30435 = (g30025)|(g21840);
assign g18374 = (g1878&g15171);
assign g13023 = ((~g11897));
assign II28597 = ((~g29374));
assign g23618 = (g19388&g11917);
assign g32714 = ((~g31528));
assign g14452 = ((~g3538))|((~g11207))|((~g3649))|((~g8542));
assign g8836 = ((~g736));
assign g10604 = ((~g7424))|((~g7456));
assign g9740 = ((~g5821));
assign g16180 = ((~g13437));
assign II29286 = ((~g12085))|((~II29284));
assign II18034 = ((~g13680));
assign II31182 = (g32719&g32720&g32721&g32722);
assign g24618 = (g22625&g19672);
assign g13485 = ((~g10476));
assign g32113 = (g31601&g29925);
assign g27346 = (g26400&g17389);
assign II13519 = ((~g2514))|((~II13518));
assign g11020 = ((~g9187))|((~g9040));
assign g24277 = (g23188)|(g18647);
assign g26784 = ((~g25341));
assign g25260 = ((~II24448));
assign g33577 = (g33405)|(g18430);
assign gbuf138 = (g1422);
assign g13504 = ((~g11303));
assign g16126 = (g5495&g14262);
assign g18215 = (g943&g15979);
assign g18353 = (g1772&g17955);
assign g13321 = (g847&g11048);
assign g16768 = ((~g13223));
assign g32090 = ((~g31003));
assign g18450 = (g2299&g15224);
assign g19525 = (g7696)|(g16811);
assign g9379 = ((~g5424));
assign g25871 = (g8334&g24804);
assign g14218 = (g875&g10632);
assign g28698 = (g27451)|(g16666);
assign g28304 = (g27226&g19753);
assign g22842 = ((~g19875));
assign g22626 = ((~II21941));
assign g22545 = ((~g1373)&(~g19720));
assign g7345 = ((~g6415));
assign II20982 = ((~g16300));
assign g33622 = (g33366)|(g18791);
assign g30122 = (g28578&g21054);
assign g21837 = (g3719&g20453);
assign g11261 = ((~g7928)&(~g4801)&(~g9030));
assign II17101 = ((~g14338));
assign g29256 = (g28597)|(g18533);
assign g24157 = ((~II23315));
assign g29198 = ((~g7766)&(~g28020));
assign g23914 = ((~g19210));
assign g9030 = ((~g4793));
assign g22861 = (g19792&g19670);
assign g21857 = (g3933&g21070);
assign II11843 = ((~g111));
assign g7472 = ((~g6329));
assign II31341 = (g31710&g31856&g32947&g32948);
assign g8224 = ((~g3774));
assign II31141 = (g31376&g31820&g32659&g32660);
assign g29333 = ((~g28167));
assign g24177 = ((~II23375));
assign g11135 = ((~II14186))|((~II14187));
assign g11639 = ((~g8933))|((~g4722));
assign g10370 = ((~g7095));
assign g11917 = ((~II14727));
assign g28341 = (g27240&g19790);
assign g32820 = ((~g31672));
assign g24717 = (g22684&g19777);
assign g33975 = (g33860)|(g18346);
assign g14962 = ((~g12558))|((~g10281));
assign g13119 = ((~g6625))|((~g12211))|((~g6715))|((~g10061));
assign g12716 = ((~g7812)&(~g6555)&(~g6549));
assign g34315 = ((~g34085));
assign II22422 = ((~g19330));
assign g25063 = (g13078&g22325);
assign II32059 = ((~g33648));
assign g9414 = ((~g2004));
assign II13708 = ((~g136));
assign II16755 = ((~g12377));
assign g32747 = ((~g30825));
assign g25504 = ((~g22550)&(~g7222));
assign II17883 = ((~g13336))|((~g1135));
assign g31325 = (g29625)|(g29639);
assign g28980 = ((~g27933))|((~g14680));
assign g30578 = ((~g29956));
assign g13603 = ((~g8009)&(~g10721));
assign g24628 = (g5835&g23666);
assign II22816 = ((~g19862));
assign g24702 = (g17464&g22342);
assign g18795 = (g6163&g15348);
assign g34393 = (g34189&g21304);
assign g32053 = (g14176&g31509);
assign g34653 = ((~II32763));
assign g19549 = ((~g15969))|((~g10841))|((~g10899));
assign g28635 = (g27375)|(g16537);
assign g31807 = ((~g29385));
assign g32350 = (g2697&g31710);
assign g16578 = ((~II17750));
assign g32929 = ((~g31710));
assign g17522 = ((~g14927));
assign g30261 = (g28772&g23961);
assign g22145 = (g14555&g18832);
assign g29481 = (g28117)|(g28125);
assign g20503 = ((~g15373));
assign g30426 = (g29785)|(g21810);
assign g22028 = (g5893&g19147);
assign gbuf68 = (g6486);
assign g12897 = ((~g10400));
assign g25718 = (g25187)|(g21971);
assign g23533 = (g19436&g13015);
assign g25701 = (g25054)|(g21920);
assign II18486 = ((~g1677))|((~II18485));
assign g28245 = (g11367&g27975);
assign g32966 = ((~g31021));
assign g33345 = (g32229&g20671);
assign g26518 = ((~g25233));
assign g19538 = ((~g16100));
assign g21350 = ((~g15751))|((~g15742))|((~g15735))|((~g13108));
assign g24324 = (g4540&g22228);
assign g23962 = ((~g19147));
assign II32432 = ((~g34056))|((~II32431));
assign g14833 = ((~g11405));
assign II23387 = ((~g23394));
assign II24128 = ((~g23009));
assign g22052 = (g6113&g21611);
assign g23023 = (g650&g20248);
assign g24571 = ((~g22942));
assign g22709 = ((~g1193))|((~g19611));
assign g28895 = ((~g27775))|((~g8146));
assign g18754 = (g5339&g15595);
assign g14626 = ((~g12232))|((~g9852))|((~g12159))|((~g9715));
assign g30523 = (g30245)|(g22069);
assign g25014 = (g17474&g23420);
assign g14438 = (g1087&g10726);
assign g25582 = (g21662)|(g24152);
assign g16160 = (g5499&g14262);
assign g30088 = ((~g29094));
assign g9154 = ((~II12994));
assign g14683 = ((~g12553))|((~g12443));
assign gbuf135 = (g194);
assign g18200 = ((~II19012));
assign g34430 = ((~II32461));
assign g18895 = ((~g16000));
assign g13966 = ((~II16246));
assign g12892 = ((~g10398));
assign II31181 = (g29385&g32716&g32717&g32718);
assign g30340 = (g29377)|(g18245);
assign g12082 = ((~g9645));
assign g33317 = (g29688)|(g32179);
assign g34407 = (g34185)|(g25124);
assign g20095 = (g8873&g16632);
assign g27960 = ((~g7134)&(~g25791));
assign g11184 = ((~g513)&(~g9040));
assign g14505 = ((~g12073))|((~g9961));
assign II29295 = ((~g29495))|((~g12117));
assign g9679 = ((~g5475));
assign II30904 = ((~g32424));
assign g8872 = ((~g4258));
assign g15754 = ((~g341)&(~g7440)&(~g13385));
assign g11396 = ((~g8713))|((~g4688));
assign g13081 = (g8626&g11122);
assign II14708 = ((~g9417));
assign g11128 = ((~g7993));
assign g19355 = ((~g16027));
assign g33733 = (g33105)|(g32012);
assign II18083 = ((~g13394));
assign g25248 = ((~g22228));
assign II16492 = ((~g12430));
assign g17645 = ((~g15018));
assign g29922 = ((~g28837));
assign g25606 = (g24761)|(g18117);
assign g29987 = (g29197&g26424&g22763);
assign g31943 = (g4717&g30614);
assign II17692 = (g14988&g11450&g6756);
assign g9556 = ((~g5448));
assign g10391 = ((~g6988));
assign g27275 = (g25945&g19745);
assign II16917 = ((~g10582));
assign g33292 = (g32150)|(g29601);
assign g26422 = (g24774)|(g23104);
assign g6869 = ((~II11691));
assign g18689 = (g15129&g16752);
assign g15062 = ((~g6817)&(~g13394));
assign g26088 = (g6545&g25080);
assign g32874 = ((~g30673));
assign g30053 = ((~g29121));
assign g14786 = ((~g12471));
assign g27362 = (g26080&g20036);
assign g13319 = (g4076&g8812&g10658&g8757);
assign II27549 = ((~g28161));
assign II14248 = ((~g1322))|((~II14247));
assign g32530 = ((~g30825));
assign II26417 = ((~g26519))|((~g14247));
assign g24292 = (g4443&g22550);
assign g26223 = (g24688&g10678&g10658&g8757);
assign g9492 = ((~g2759));
assign g17496 = ((~g14683));
assign g24992 = ((~g22417));
assign g24771 = (g7028&g23605);
assign g31780 = (g30163&g23999);
assign g33562 = (g33414)|(g18379);
assign g9892 = ((~g6428));
assign g29229 = (g28532)|(g18191);
assign g33894 = ((~II31748));
assign II13043 = ((~g5115))|((~g5120));
assign g26744 = ((~g25400));
assign g18684 = (g4681&g15885);
assign g15083 = (g10362&g12983);
assign II24030 = (g8390&g8016&g3396);
assign g16520 = (g5909&g14965);
assign g22986 = ((~g20330));
assign g32375 = (g29896)|(g31324);
assign g27352 = ((~g7975)&(~g26616));
assign II32240 = ((~g34131));
assign g33186 = (g32037&g22830);
assign g22920 = (g19764&g19719);
assign g13830 = (g11543&g11424&g11395&II16143);
assign g33018 = (g32312)|(g18525);
assign g34485 = (g34411&g18952);
assign g31116 = ((~g7892)&(~g29540));
assign g15806 = ((~II17302));
assign g34385 = (g34168&g20642);
assign g25767 = (g25207)|(g12015);
assign g15151 = ((~g13745)&(~g7027));
assign g19953 = ((~g16220)&(~g13712));
assign g27311 = (g12431&g26693);
assign g19739 = ((~g16931));
assign g24026 = ((~g19919));
assign g28333 = (g27239&g19787);
assign g33111 = (g24005&g32421);
assign g31899 = (g31470)|(g21907);
assign g30564 = (g21358&g29385);
assign g17147 = ((~g14321));
assign II33044 = ((~g34775));
assign g31655 = ((~II29233));
assign g8344 = ((~II12523));
assign g25899 = ((~g24997));
assign g31744 = (g30092&g23902);
assign g21464 = (g16181&g10872);
assign g17367 = ((~II18320));
assign g12149 = ((~g8205))|((~g2185));
assign g20275 = ((~g17929));
assign g19366 = ((~g15885));
assign g13265 = (g9018&g11493);
assign g29976 = ((~g29018));
assign g15163 = ((~g13809)&(~g12905));
assign g27678 = (g947&g25830);
assign g29623 = (g28496&g11563);
assign g23542 = ((~g21514));
assign g26680 = ((~g25300));
assign g34620 = (g34529)|(g18582);
assign g14315 = ((~II16479));
assign g32905 = ((~g30825));
assign g31787 = (g21281&g29385);
assign g28575 = ((~g27711));
assign g34228 = (g33750&g22942);
assign g31318 = ((~g4785)&(~g29697));
assign g17594 = (g14450)|(g14420)|(g12025)|(II18543);
assign g18383 = (g1950&g15171);
assign g18207 = (g925&g15938);
assign g23961 = ((~g19074));
assign g20202 = (g16211)|(g13507);
assign g10584 = ((~g7362))|((~g7405));
assign g32513 = ((~g31376));
assign g19618 = ((~g16349));
assign g7451 = ((~g2070));
assign g21184 = ((~g15509));
assign g13872 = ((~g8745)&(~g11083));
assign II32550 = ((~g34398));
assign g13056 = ((~g7400)&(~g10741));
assign g32494 = ((~g30825));
assign II23393 = ((~g23414));
assign g28463 = ((~II26952));
assign II11626 = ((~g31));
assign g23472 = ((~g21062));
assign g25058 = (g23276&g20513);
assign g8607 = ((~g37));
assign g26894 = (g25979)|(g18129);
assign g26328 = (g1183)|(g24591);
assign II22009 = ((~g21269));
assign g29745 = ((~g28500));
assign g23506 = ((~g21514));
assign g28851 = (g27558)|(g16870);
assign g9523 = ((~g6419));
assign g18888 = ((~g15426));
assign g32519 = ((~g30673));
assign g18932 = ((~g16136));
assign g22102 = (g6479&g18833);
assign g23549 = ((~g18833));
assign g30136 = ((~g28799)&(~g7380));
assign g27975 = ((~g26694));
assign g19738 = ((~g15992));
assign II13383 = ((~g269))|((~II13382));
assign g28616 = (g27532&g20551);
assign g11448 = ((~g4191)&(~g8790));
assign g20914 = ((~g15373));
assign g16537 = (g5937&g14855);
assign g15654 = (g3845&g13584);
assign g18343 = (g12847&g17955);
assign g21722 = ((~II21285));
assign g28646 = (g27388)|(g16595);
assign g13764 = ((~g11252))|((~g3072));
assign g18106 = (g411&g17015);
assign g19411 = ((~g16489));
assign g13910 = ((~g4899)&(~g4975)&(~g11173));
assign g32571 = ((~g31376));
assign II15241 = ((~g10003))|((~g6351));
assign g19913 = ((~g11430))|((~g17794));
assign g33551 = (g33446)|(g18342);
assign g23898 = ((~g19277));
assign g27998 = ((~II26512));
assign II27758 = ((~g28119));
assign g26966 = (g26345)|(g24318);
assign g14749 = ((~II16829));
assign g12027 = (g9499&g9729);
assign II14623 = ((~g8925));
assign g33053 = (g31967)|(g21974);
assign g29383 = (g28138&g19412);
assign g23494 = ((~II22619));
assign g27008 = (g26866)|(g21370)|(II25736);
assign g23775 = (g14872&g21267);
assign g16534 = (g5575&g14665);
assign g23256 = ((~g20785));
assign g21818 = (g3610&g20924);
assign g31554 = (g19050&g29814);
assign g19367 = ((~II19851));
assign g23227 = ((~g20924));
assign g8592 = ((~g3805));
assign g12399 = ((~g9920));
assign g30451 = (g29877)|(g21860);
assign g25936 = (g24403)|(g22209);
assign II22211 = ((~g21463));
assign g33142 = ((~g32072));
assign g24637 = (g16586&g22884);
assign g34040 = (g33818)|(g18737);
assign g29796 = (g28345&g23258);
assign g15095 = ((~g13177)&(~g12866));
assign g22127 = (g6625&g19277);
assign g9804 = ((~g5456));
assign g8438 = ((~g3100));
assign g23220 = (g19417&g20067);
assign g17243 = ((~g7247))|((~g14212));
assign g31755 = (g29991)|(g30008);
assign g21908 = (g5037&g21468);
assign g11204 = ((~II14271));
assign g23968 = ((~g18833));
assign g34848 = ((~II33070));
assign g23320 = ((~II22419));
assign g28468 = ((~g3155)&(~g10295)&(~g27602));
assign II14498 = ((~g9020))|((~II14497));
assign gbuf127 = (g875);
assign g32549 = ((~g31554));
assign g23154 = ((~II22264));
assign g29904 = (g28312)|(g26146);
assign g11562 = ((~g7648));
assign g31299 = (g30123&g27800);
assign g12844 = ((~g10360));
assign g19429 = ((~g16489));
assign g30210 = (g28684&g23877);
assign g19264 = ((~II19802));
assign g12201 = ((~g5417)&(~g10047));
assign g19713 = ((~g16816));
assign g27378 = (g26089&g20052);
assign g30673 = (g20175&g29814);
assign g24424 = ((~g22722));
assign g29676 = ((~g28381))|((~g13676));
assign g33865 = (g33275&g20526);
assign g34134 = ((~II32079));
assign g16606 = ((~g14110));
assign g14829 = ((~g6621))|((~g12137))|((~g6675))|((~g12471));
assign II15620 = ((~g12038));
assign g9616 = ((~g5452));
assign II15123 = ((~g2102))|((~II15121));
assign II33252 = ((~g34974));
assign g31578 = ((~II29199));
assign g32775 = ((~g30825));
assign g34502 = (g26363&g34343);
assign g32016 = (g8522&g31138);
assign g24210 = (g22900)|(g18125);
assign g20645 = ((~g14344))|((~g17243));
assign g10565 = (g8182&g424);
assign II22458 = ((~g18954));
assign g27112 = ((~g26793));
assign g18431 = (g2185&g18008);
assign g9166 = ((~g837));
assign g34685 = (g14164&g34550);
assign g13282 = (g3546&g11480);
assign g24038 = ((~g21193));
assign g32734 = ((~g31710));
assign II12950 = ((~g4287));
assign II26395 = ((~g14227))|((~II26393));
assign g10191 = ((~g6386));
assign g18734 = (g4966&g16826);
assign g28126 = ((~g27122));
assign g14889 = ((~g12609))|((~g12824));
assign g31292 = (g29735&g23338);
assign g34740 = (g34664&g19414);
assign II14765 = ((~g9808))|((~II14764));
assign II31011 = (g30735&g31797&g32471&g32472);
assign g21964 = (g5441&g21514);
assign g26195 = (g25357&g6856&g11709&g7558);
assign g32897 = ((~g30735));
assign g28514 = ((~g8165)&(~g27617));
assign g30049 = (g13114&g28167);
assign g9044 = ((~g604));
assign g34625 = (g34532)|(g18610);
assign g34498 = (g13888&g34336);
assign g6972 = ((~II11740));
assign II13141 = ((~g6159))|((~II13139));
assign g33985 = (g33896)|(g18382);
assign gbuf152 = (g1239);
assign g20512 = ((~g18062));
assign II26334 = ((~g26834));
assign g25171 = ((~g22228));
assign g21827 = (g3759&g20453);
assign g13037 = ((~g10981));
assign g21774 = (g3361&g20391);
assign g29121 = ((~g9755))|((~g27886));
assign g21873 = (g6946&g19801);
assign II32284 = ((~g34052));
assign g13633 = (g4567&g10509);
assign g14864 = ((~g7791))|((~g10421));
assign g22622 = (g19336&g19469);
assign g18309 = (g1339&g16931);
assign g9499 = ((~g5152));
assign g15885 = ((~II17374));
assign g16630 = ((~g14142));
assign g21036 = ((~II20910));
assign g23166 = (g13959&g19979);
assign g34422 = ((~II32432))|((~II32433));
assign II27381 = (g25549&g26424&g22698);
assign g18628 = (g15095&g17226);
assign g30462 = (g30228)|(g21933);
assign g24244 = (g23349)|(g18255);
assign g21677 = ((~II21238));
assign g26126 = (g1959&g25118);
assign g6840 = ((~g1992));
assign gbuf146 = (g1075);
assign g32502 = ((~g31070));
assign g11189 = ((~II14248))|((~II14249));
assign g18319 = (g1600&g17873);
assign g32938 = ((~g30937));
assign g32161 = (g3151&g31154);
assign g26942 = ((~II25692));
assign g25547 = ((~g22550));
assign g34117 = (g33742&g19755);
assign g29852 = (g1772&g29080);
assign g28225 = (g27770&g23400);
assign g16529 = ((~g14055));
assign g33062 = (g31977)|(g22065);
assign g33378 = ((~II30904));
assign g30196 = (g28659&g23858);
assign g14512 = ((~g11955)&(~g9753));
assign g12482 = ((~II15307))|((~II15308));
assign g12823 = ((~g9206));
assign g33791 = (g33379)|(g32430);
assign g25680 = (g24794)|(g21839);
assign g8407 = ((~g1171));
assign g11663 = ((~g6905));
assign g11201 = ((~g4125)&(~g7765));
assign II31823 = ((~g33149));
assign g28728 = (g27501)|(g16730);
assign g34329 = (g14511&g34181);
assign II12519 = ((~g3447));
assign II25391 = ((~g24483));
assign g32862 = ((~g30825));
assign II17754 = ((~g13494));
assign g31021 = (g26025&g29814);
assign g30934 = ((~g29836)&(~g29850));
assign g26831 = ((~g24836));
assign g34427 = ((~II32452));
assign g33442 = ((~g31937));
assign g24481 = ((~II23684));
assign g31522 = ((~II29185));
assign g9704 = ((~g2575));
assign g28861 = ((~g27837))|((~g7405))|((~g1906));
assign g20448 = ((~g15509));
assign g32412 = (g4765&g30998);
assign g15844 = ((~g14714))|((~g9340))|((~g12378));
assign g8056 = ((~g1246));
assign g17401 = (g1083&g13143);
assign g32673 = ((~g31376));
assign g7565 = ((~II12046));
assign g20887 = (g16282&g4864);
assign g16641 = (g6613&g14782);
assign g24528 = ((~g4098))|((~g22654));
assign g31514 = (g20041&g29956);
assign g18525 = (g2610&g15509);
assign g24755 = (g16022&g23030);
assign g17514 = ((~g3917))|((~g13772))|((~g4019))|((~g8595));
assign g25178 = (g20241&g23608);
assign g11986 = ((~II14830));
assign g32262 = (g31186)|(g29710);
assign g16249 = ((~II17590));
assign g27227 = (g26026&g16771);
assign II14589 = ((~g8818));
assign g33252 = (g32155&g20064);
assign g17624 = ((~II18588))|((~II18589));
assign g26159 = (g2370&g25137);
assign g11590 = ((~g6928))|((~g3990))|((~g4049));
assign g28945 = ((~g27854))|((~g8211));
assign g16489 = ((~II17699));
assign g24140 = (g17663&g21654);
assign g25371 = (g5062&g22173&II24524);
assign g16928 = (g13525)|(g11127);
assign g24010 = ((~g21562));
assign g29766 = (g28316&g23235);
assign g29980 = ((~g28935));
assign g31067 = (g29484&g22868);
assign g18510 = (g2625&g15509);
assign g24940 = (g5011&g23971);
assign II20913 = ((~g16964));
assign g28315 = (g27232&g19769);
assign g31836 = ((~g29385));
assign g12297 = ((~g9269)&(~g9239));
assign g32041 = (g13913&g31262);
assign g16428 = ((~II17668));
assign g20152 = (g11545&g16727);
assign g30117 = ((~g28739)&(~g7252));
assign II14006 = ((~g9104));
assign g11245 = ((~g7636))|((~g7733))|((~g7697));
assign II12277 = ((~g1467))|((~g1472));
assign g20713 = ((~g15277));
assign g13221 = (g6946&g11425);
assign g33962 = (g33822)|(g18123);
assign g33645 = ((~II31477));
assign g7992 = ((~g5008));
assign g16244 = (g11547&g11592&g6789&II17585);
assign g32717 = ((~g30735));
assign g21303 = (g10120&g17625);
assign gbuf34 = (g5681);
assign II17801 = ((~g14936));
assign g27462 = (g26576&g17612);
assign g24821 = (g21404)|(g23990);
assign g18285 = (g1395&g16164);
assign g25696 = (g25012)|(g21915);
assign g28326 = ((~g27414));
assign g26871 = (g25038&g25020);
assign g34741 = (g8899&g34697);
assign II31217 = (g32768&g32769&g32770&g32771);
assign g29488 = (g28547)|(g27600);
assign g16474 = (g8280&g13666);
assign g6991 = ((~g4888));
assign g7863 = ((~g1249));
assign g24285 = (g4388&g22550);
assign g32727 = ((~g31710));
assign g10603 = ((~g10077))|((~g9751));
assign g23066 = ((~g20330));
assign g33475 = (g32563&II31071&II31072);
assign II27573 = ((~g28157));
assign g18505 = (g2583&g15509);
assign g8685 = ((~g1430));
assign II25220 = ((~g482))|((~II25219));
assign g29743 = (g28206&g10233);
assign II12098 = ((~g1322))|((~II12096));
assign g15726 = ((~g6263))|((~g14529))|((~g6365))|((~g10003));
assign g28262 = ((~II26785));
assign g16590 = (g5236&g14683);
assign g27034 = (g26328&g8609);
assign g16685 = ((~g14038));
assign II26741 = (g22881)|(g22905)|(g22928)|(g27402);
assign g28426 = (g27257&g20006);
assign g21800 = (g3546&g20924);
assign g9541 = ((~g2012));
assign g14090 = ((~g8851)&(~g12259));
assign g29378 = (g28137&g22493);
assign g28731 = (g27504)|(g16733);
assign g33457 = ((~II30989));
assign g22126 = (g6621&g19277);
assign g9908 = ((~II13453))|((~II13454));
assign g6895 = ((~g3288));
assign g23167 = ((~g8219))|((~g19981));
assign g33388 = ((~g32382));
assign g21024 = (g16306&g4871);
assign g30595 = (g18911&g29847);
assign g25830 = ((~g24485));
assign g21204 = ((~g15656));
assign g9931 = ((~g5763));
assign g25064 = ((~II24228));
assign g28590 = ((~g27724));
assign g34955 = (g34931&g34320);
assign g25763 = (g25113)|(g18817);
assign g33459 = ((~II30995));
assign g25687 = (g24729)|(g21882);
assign g11948 = ((~g10224));
assign g24312 = (g4501&g22228);
assign g33312 = (g29646)|(g32170);
assign II18537 = ((~g2236))|((~II18536));
assign g9664 = ((~g4878)&(~g4871)&(~g4864)&(~g4836));
assign g18718 = (g4854&g15915);
assign II13109 = ((~g5808))|((~g5813));
assign g31124 = (g2259&g29997);
assign g24017 = ((~g18833));
assign g7356 = ((~g1802));
assign gbuf120 = (g4229);
assign g19067 = ((~g15979));
assign g18481 = (g2461&g15426);
assign g25325 = ((~g22228));
assign g10113 = ((~g2084));
assign g9692 = ((~g1756));
assign g20170 = ((~g16741))|((~g13897))|((~g16687))|((~g13866));
assign g32171 = (g31706&g27800);
assign g15076 = (g2130&g12955);
assign g18728 = (g4939&g16821);
assign g19692 = (g12066&g17086);
assign g8201 = ((~g1894));
assign g10205 = ((~g2657)&(~g2523)&(~g2389)&(~g2255));
assign g15508 = ((~g10320)&(~g14279));
assign g28035 = (g24103&II26530&II26531);
assign g22137 = ((~g21370));
assign g21253 = ((~g6423))|((~g17482));
assign g22634 = (g18934)|(g15590);
assign g29517 = (g1870&g28827);
assign g9732 = ((~g5481));
assign II15697 = ((~g6000));
assign II16724 = ((~g12108));
assign II13566 = ((~g2652))|((~II13564));
assign g31845 = ((~g29385));
assign g10621 = ((~g7567));
assign g19445 = ((~g15915));
assign II16143 = (g8751&g11491&g11445);
assign g12088 = ((~g7701));
assign g18445 = (g2273&g18008);
assign g32568 = ((~g31170));
assign g31936 = (g31213&g24005);
assign g34991 = ((~II33273));
assign g10489 = ((~g9259));
assign g32976 = (g32207)|(g21704);
assign g34200 = ((~g33895));
assign II18449 = (g14512)|(g14445)|(g14415);
assign g32127 = (g31624&g29950);
assign g24506 = ((~II23711));
assign g31018 = (g29480&g22855);
assign g9760 = ((~g2315));
assign g31911 = (g31784)|(g21969);
assign g34968 = (g34952&g23203);
assign g9860 = ((~g5417));
assign g24164 = ((~II23336));
assign II14275 = ((~g8218))|((~g3484));
assign g33118 = (g32413)|(g32418);
assign g26750 = (g24514&g24474);
assign g28072 = (g27086)|(g21874);
assign g15128 = ((~g13638)&(~g12880));
assign II22267 = (g20236)|(g20133)|(g20111);
assign g10555 = ((~g7227)&(~g4601)&(~g4608));
assign g24145 = ((~g19402)&(~g19422));
assign g27142 = ((~g26105));
assign II15102 = ((~g5313));
assign g33533 = ((~II31361));
assign g16873 = ((~II18063));
assign II11708 = ((~g3703));
assign g18951 = (g3484&g16124);
assign g18984 = ((~g17486));
assign g12793 = ((~g10287));
assign g25987 = (g9501&g25015);
assign g13512 = ((~g9077)&(~g12527));
assign g10368 = ((~g6887));
assign g27528 = ((~g8770)&(~g26352)&(~g11083));
assign II14660 = ((~g9746));
assign g29853 = (g1862&g29081);
assign g24553 = (g22983&g19539);
assign g16322 = ((~II17650));
assign g25876 = (g3470&g24667);
assign g15002 = ((~g12609))|((~g10312));
assign g25102 = (g4727&g22885);
assign g10109 = ((~g135));
assign g12953 = (g411&g11048);
assign g11042 = ((~g8691));
assign g28414 = ((~g27467)&(~g26347));
assign g26380 = (g19572&g25547);
assign g18364 = (g1844&g17955);
assign II17136 = ((~g14398));
assign g21744 = (g3103&g20330);
assign g17605 = ((~g5559))|((~g14425))|((~g5630))|((~g12563));
assign g19416 = ((~g15885));
assign g32381 = ((~II29909));
assign g30282 = ((~g6336)&(~g29073));
assign g26297 = ((~g8519)&(~g24825));
assign g24922 = (g4831&g23931);
assign g18657 = (g4308&g17128);
assign g31508 = (g29813&g23459);
assign gbuf85 = (g3625);
assign g22870 = ((~g20887));
assign g31790 = (g21299&g29385);
assign g30292 = ((~g28736));
assign g30189 = (g23401)|(g28543);
assign g27339 = (g26400&g17308);
assign g12639 = ((~g10194))|((~g6682))|((~g6732));
assign g22111 = (g6549&g19277);
assign g13012 = ((~II15626));
assign II27970 = ((~g28803));
assign g17497 = ((~g14879));
assign g23926 = ((~g19074));
assign g21910 = (g5016&g21468);
assign g29169 = ((~g27886));
assign g10337 = ((~g5016));
assign g28991 = (g14438&g25209&g26424&g27469);
assign II17108 = ((~g13782));
assign g18770 = (g15153&g15615);
assign II16090 = ((~g10430));
assign g25887 = ((~g24984)&(~g11706));
assign g34078 = (g33699&g19531);
assign g15936 = (g475&g13999);
assign g23513 = (g19430&g13007);
assign g33873 = (g33291&g20549);
assign g27232 = (g25874)|(g24450);
assign g24252 = (g22518)|(g18299);
assign g15628 = ((~g11907)&(~g14228));
assign g7499 = ((~g333)&(~g355));
assign II18835 = ((~g6365));
assign g24532 = (g22331&g19478);
assign II24215 = ((~g22360));
assign g25424 = ((~g23800));
assign g29668 = (g28527&g14255);
assign g14691 = ((~g12695))|((~g12505));
assign g25429 = ((~g22417))|((~g1917))|((~g8302));
assign g28570 = (g27456&g20434);
assign II33170 = ((~g34890));
assign g33998 = (g33878)|(g18428);
assign II21246 = ((~g16540));
assign g24658 = (g22645&g19732);
assign g14731 = ((~g5698)&(~g12204));
assign g15875 = (g3961&g13963);
assign g12571 = ((~g9511)&(~g9451));
assign g18564 = (g2844&g16349);
assign g14541 = ((~g11405));
assign g22993 = ((~g1322)&(~g16292)&(~g19873));
assign g20166 = ((~g16886));
assign g27981 = (g26751&g23924);
assign g33615 = (g33113)|(g21871);
assign II19778 = ((~g17781));
assign II24709 = (g21256&g24068&g24069&g24070);
assign g20114 = ((~II20385));
assign g24048 = ((~g19968));
assign g13096 = ((~II15727));
assign gbuf61 = (g6704);
assign g22838 = ((~g20219))|((~g2960));
assign g25941 = (g24416)|(g22219);
assign g21864 = (g3961&g21070);
assign g24159 = ((~II23321));
assign g19741 = ((~g16987));
assign II13453 = ((~g1955))|((~II13452));
assign g19461 = (g11708&g16846);
assign g11142 = (g6381&g10207);
assign g17873 = ((~II18849));
assign g32969 = ((~g30735));
assign g31130 = (g12191&g30019);
assign g24576 = ((~g22957))|((~g2902));
assign g18295 = (g1489&g16449);
assign g28689 = (g27575&g20651);
assign g26813 = (g24940)|(g24949);
assign II16160 = ((~g11237));
assign II23978 = ((~g23198))|((~g13670));
assign g32137 = ((~g31134));
assign g28205 = (g27516&g16746);
assign II33137 = ((~g34884));
assign g33971 = (g33890)|(g18330);
assign g21155 = ((~g15656));
assign g32393 = ((~g30922));
assign g24798 = ((~II23962))|((~II23963));
assign II16618 = (g10124&g12341&g12293);
assign II20861 = ((~g16960));
assign g28750 = (g27525)|(g16765);
assign g27332 = (g12538&g26758);
assign g31477 = (g29763&g23409);
assign g25774 = (g25223)|(g12043);
assign g20667 = ((~g15224));
assign g7627 = ((~g4311));
assign g21763 = (g3223&g20785);
assign g14078 = (g10776)|(g8703);
assign II13699 = ((~g4581));
assign II16780 = ((~g12332))|((~II16778));
assign g22082 = (g6283&g19210);
assign g18214 = (g939&g15979);
assign g23416 = (g20082&g20321);
assign g14424 = ((~g11136));
assign g21608 = ((~g17955));
assign g26987 = ((~g26131));
assign II23162 = (g19919)|(g19968)|(g20014)|(g20841);
assign g14517 = ((~g3231))|((~g11217))|((~g3321))|((~g8481));
assign g16705 = (g6299&g15024);
assign II31854 = (g33492)|(g33493)|(g33494)|(g33495);
assign g25620 = ((~II24759));
assign II17529 = (g13156&g11450&g6756);
assign g12523 = ((~g7563))|((~g6346));
assign g17183 = ((~II18221));
assign g18300 = (g1306&g16489);
assign g7183 = ((~g4608));
assign II31972 = ((~g33641))|((~g33631));
assign gbuf147 = (g1079);
assign II25115 = ((~g25322));
assign g10041 = ((~II13565))|((~II13566));
assign g18473 = (g2342&g15224);
assign g34656 = ((~II32770));
assign II19734 = ((~g17725));
assign g30531 = (g30274)|(g22077);
assign g14450 = ((~g12195)&(~g9598));
assign g21917 = (g5092&g21468);
assign g28429 = (g27228)|(g15913);
assign g13666 = ((~g11190))|((~g8441));
assign g33598 = (g33364)|(g18496);
assign g23971 = ((~g20751));
assign g20109 = (g17954&g17616);
assign g24624 = (g16524&g22867);
assign g11367 = ((~II14381));
assign g13412 = ((~g11963));
assign g30203 = (g28668&g23864);
assign gbuf134 = (g802);
assign g21999 = (g5723&g21562);
assign g17686 = ((~g6251))|((~g14529))|((~g6322))|((~g12672));
assign g15569 = ((~II17148));
assign g31470 = (g29753&g23398);
assign g32953 = ((~g31327));
assign g29643 = (g28192)|(g27145);
assign gbuf25 = (g5105);
assign g25210 = ((~g23802));
assign g30482 = (g30230)|(g21978);
assign g23395 = ((~II22502));
assign g27616 = (g26349&g20449);
assign g34156 = ((~g33907));
assign g30142 = ((~g28754));
assign g34465 = (g34295)|(g18712);
assign g28375 = (g27183)|(g15851);
assign g32011 = (g8287&g31134);
assign g32082 = (g4917&g30673);
assign g17264 = (g7118)|(g14309);
assign g7335 = ((~g2287));
assign g34254 = (g34116)|(g24301);
assign g30401 = (g29782)|(g21760);
assign g33095 = ((~g31997)&(~g7236));
assign II14481 = ((~g10074))|((~II14480));
assign g33303 = (g32159)|(g29638);
assign g7231 = ((~g5));
assign g33418 = (g32372&g21425);
assign g17574 = (g9554&g14546);
assign g32331 = (g31322&g20637);
assign g13222 = ((~g10590));
assign g32586 = ((~g31376));
assign g10529 = ((~g1592))|((~g7308));
assign g14208 = ((~g11563));
assign g20737 = ((~g15656));
assign II31291 = (g31021&g31847&g32875&g32876);
assign g31920 = (g31493)|(g22045);
assign g20704 = ((~g15373));
assign II20221 = ((~g16272))|((~g11170));
assign g8330 = ((~g2587));
assign g25722 = (g25530)|(g18768);
assign g33926 = ((~II31796));
assign g29578 = (g2491&g28606);
assign g6801 = ((~g391));
assign g26776 = ((~g25498));
assign II13444 = ((~g239))|((~II13442));
assign g24606 = (g5489&g23630);
assign g33886 = (g33297&g20614);
assign g32605 = ((~g30614));
assign g12361 = ((~g6455)&(~g10172));
assign g23948 = ((~g21012));
assign II26512 = ((~g26817));
assign g23271 = ((~g20785));
assign g29615 = (g1844&g29049);
assign g25948 = ((~g7752)&(~g24609));
assign II21918 = ((~g21290));
assign g23130 = (g728&g20248);
assign g20769 = ((~g17955));
assign g24746 = (g22588)|(g19461);
assign g12850 = ((~g10430)&(~g6845));
assign II29352 = (g29322)|(g29315)|(g30315)|(g30308);
assign g18817 = (g6533&g15483);
assign g23412 = (g7297&g21510);
assign g16957 = (g13064&g10418);
assign g34159 = ((~II32116));
assign II14054 = ((~g10028));
assign g29204 = (g24110&II27518&II27519);
assign g23162 = (g20184)|(g20170)|(II22267);
assign g30065 = ((~g29049));
assign II31197 = (g32740&g32741&g32742&g32743);
assign g33612 = (g33247)|(g18633);
assign g9639 = ((~g1752));
assign g10213 = ((~g6732));
assign g33034 = (g32340)|(g21844);
assign g20449 = ((~g15277));
assign g9187 = ((~g518));
assign g22047 = (g6077&g21611);
assign g32998 = (g32300)|(g18393);
assign g23787 = ((~g18997));
assign II12563 = ((~g3798));
assign II17787 = ((~g3267));
assign g29248 = (g28677)|(g18434);
assign g8113 = ((~g3466));
assign g32098 = (g4732&g30614);
assign g22099 = (g6462&g18833);
assign g23568 = ((~g21611));
assign g26203 = (g1632&g25337);
assign II14684 = ((~g7717));
assign g11755 = ((~g4709)&(~g8796));
assign II32170 = ((~g33638));
assign g34776 = ((~II32970));
assign g34722 = (g34707)|(g18137);
assign g19376 = ((~g17509));
assign g7548 = ((~g1036));
assign II32106 = ((~g33653));
assign g16761 = (g7170&g12947);
assign II24558 = ((~g23777));
assign II18376 = ((~g14332));
assign g19659 = ((~g17062));
assign g28674 = (g27569&g20629);
assign g22755 = ((~g20136))|((~g18984));
assign g16826 = ((~II18034));
assign g9340 = ((~II13094));
assign g15078 = (g10361&g12955);
assign g19655 = (g2729&g16966);
assign g19454 = ((~g16349));
assign II24463 = ((~g14437))|((~II24461));
assign g9501 = ((~g5731));
assign g25572 = (II24699&II24700);
assign g9443 = ((~g5489));
assign g25536 = (g23770&g21431);
assign g20900 = ((~II20864));
assign g17736 = ((~g5563))|((~g14522))|((~g5659))|((~g12563));
assign II15253 = ((~g10078))|((~g1848));
assign g29838 = (g1636&g29044);
assign g10656 = (g3782&g7952);
assign II18160 = ((~g14441));
assign g27828 = ((~g9892)&(~g25856));
assign g26876 = (g21655)|(g25576);
assign g22997 = ((~g20391));
assign g29901 = (g28429&g23376);
assign g32526 = ((~g30614));
assign g25094 = (g23318&g20554);
assign g9974 = ((~g2518));
assign g18440 = (g2255&g18008);
assign g27393 = (g26099&g20066);
assign g31616 = ((~II29214));
assign g11292 = ((~II14331))|((~II14332));
assign g13027 = ((~II15647));
assign g12835 = ((~g10352));
assign g7666 = ((~g4076));
assign g17581 = ((~g5607))|((~g12029))|((~g5623))|((~g14669));
assign g18676 = (g4358&g15758);
assign g31211 = (g10156&g30102);
assign g25791 = (g25411)|(g25371)|(g25328)|(g25290);
assign g9689 = ((~g124));
assign g31608 = ((~g29653));
assign II26448 = ((~g26860));
assign g17744 = ((~g6303))|((~g14529))|((~g6373))|((~g12672));
assign g28149 = ((~g27598)&(~g27612));
assign g28136 = (g27382&g23135);
assign g29277 = (g28440)|(g18710);
assign g24358 = ((~g22550));
assign g16734 = (g5961&g14735);
assign g12730 = (g9024&g4349);
assign g32841 = ((~g31672));
assign II12333 = ((~g45));
assign g13350 = ((~II15906));
assign g30441 = (g29787)|(g21850);
assign g13902 = ((~g11389));
assign g30133 = (g28591&g21179);
assign g18265 = (g1270&g16000);
assign g21284 = ((~g16646)&(~g9690));
assign g7393 = ((~g5320));
assign II23600 = ((~g22360))|((~g4322));
assign II19345 = ((~g15083));
assign g14095 = ((~g11326));
assign g23885 = (g4132&g19513);
assign g8519 = ((~g287));
assign g11812 = ((~g7567));
assign g19629 = ((~g17015));
assign g30224 = (g28704&g23896);
assign g34027 = (g33718)|(g18683);
assign g29634 = (g2108&g29121);
assign g28889 = (g17292&g25169&g26424&g27395);
assign g11412 = ((~g8666))|((~g6918))|((~g8697));
assign II18868 = ((~g14315));
assign g24343 = (g23724)|(g18773);
assign g19740 = (g2783&g15907);
assign g29665 = (g2375&g28696);
assign g27617 = (g23032&g26264&g26424&g24982);
assign g29614 = (g28860&g22369);
assign g8387 = ((~g3080));
assign g20524 = ((~g17873));
assign g22717 = (g9291&g20212);
assign g8002 = ((~g1389));
assign g21610 = ((~g15615));
assign g33819 = (g23088&g33176&g9104);
assign g28711 = ((~g27886));
assign g28659 = (g27404)|(g16610);
assign g18612 = (g3329&g17200);
assign II18523 = ((~g14443));
assign II30755 = (g30564)|(g32303)|(g32049)|(g32055);
assign g27428 = (g26400&g17576);
assign II29315 = ((~g12154))|((~II29313));
assign g18397 = (g2004&g15373);
assign II11685 = ((~g117));
assign g14539 = ((~g11977)&(~g9833));
assign g30824 = (g13833)|(g29789);
assign g14085 = ((~g7121))|((~g11584));
assign g12581 = ((~g9569)&(~g6219));
assign g33134 = ((~g7686)&(~g32057));
assign g30106 = ((~g28739)&(~g7268));
assign g34380 = (g34158&g20571);
assign g18404 = (g2066&g15373);
assign II15736 = ((~g12322));
assign II31136 = (g29385&g32651&g32652&g32653);
assign g30388 = (g30023)|(g18534);
assign g28165 = (g27018&g22455);
assign g27073 = (g7121&g3873&g3881&g26281);
assign II11665 = ((~g1589));
assign g25118 = ((~g22417));
assign g29572 = (g1620&g28885);
assign g18502 = (g2567&g15509);
assign g34290 = (g26848)|(g34219);
assign II20469 = ((~g16728))|((~II20467));
assign g26858 = (g2970&g24540);
assign g16815 = ((~g3909))|((~g13824))|((~g4005))|((~g11631));
assign g25805 = (g25453)|(g25414)|(g25374)|(g25331);
assign g33279 = (g32140)|(g29573);
assign g28033 = ((~g26365));
assign g34539 = ((~g34354));
assign II12033 = ((~g776));
assign g29178 = (g27163&g12687);
assign II15921 = ((~g12381));
assign g31825 = ((~g29385));
assign g25658 = (g24635)|(g21783);
assign g8283 = ((~II12493));
assign g27334 = (g12539&g26769);
assign g22067 = (g6215&g19210);
assign g12838 = ((~g10353));
assign g22318 = (g21394)|(g17783);
assign II32476 = ((~g34277));
assign g7437 = ((~g5666));
assign II18795 = ((~g5327));
assign II14742 = ((~g9534));
assign g22518 = (g12982&g19398);
assign g10706 = (g3338&g8691);
assign g32253 = (g24771)|(g31207);
assign II24699 = (g21127&g24054&g24055&g24056);
assign g31152 = (g10039&g30067);
assign II20882 = ((~g17619));
assign g33481 = (g32607&II31101&II31102);
assign g33870 = (g33280&g20545);
assign g9724 = ((~g5092))|((~g5084));
assign g26713 = (g25447&g20714);
assign II14530 = ((~g8840))|((~g8873));
assign g15018 = ((~g12739))|((~g12515));
assign II15834 = ((~g11164));
assign g28973 = ((~g27907))|((~g2465))|((~g7387));
assign g28066 = (g27553)|(g21819);
assign g26703 = (g24447)|(g10705);
assign g23560 = ((~g9607)&(~g20838));
assign g21749 = (g3155&g20785);
assign g15143 = ((~g6998)&(~g13680));
assign g14121 = ((~g8891)&(~g12259));
assign g33498 = (g32730&II31186&II31187);
assign g31251 = (g25973)|(g29527);
assign g23988 = ((~g19277));
assign g17271 = ((~II18270));
assign g30094 = (g28544&g20767);
assign g33679 = ((~g33394))|((~g10737))|((~g10308));
assign g33589 = (g33340)|(g18469);
assign g34890 = (g34863)|(g21674);
assign g21796 = (g3512&g20924);
assign g8504 = ((~g3451));
assign g8183 = ((~g482));
assign g16268 = ((~g7913)&(~g13121));
assign g25250 = ((~II24434));
assign g18632 = (g3698&g17226);
assign g23559 = ((~g21070));
assign II32874 = ((~g34504));
assign g8088 = ((~g1554));
assign g28779 = ((~II27253));
assign II30727 = (g31759)|(g32196)|(g31933)|(g31941);
assign g27292 = (g1714&g26654);
assign g30471 = (g30175)|(g21942);
assign g10491 = ((~g6573)&(~g9576));
assign g25083 = ((~g23782));
assign g8917 = ((~II12890));
assign g24745 = (g650&g23550);
assign g9281 = ((~II13057));
assign g32246 = (g31246&g20326);
assign g33670 = ((~II31504));
assign g23430 = ((~II22547));
assign g11533 = ((~g6905))|((~g3639))|((~g3698));
assign g34493 = (g34273&g19360);
assign g28440 = (g27274&g20059);
assign g20543 = ((~g17955));
assign g17636 = (g10829&g13463);
assign g30325 = ((~II28576));
assign g19609 = ((~g16264));
assign g19762 = ((~g16326));
assign g34278 = (g26829)|(g34212);
assign g34225 = (g33744&g22942);
assign g33107 = ((~g32180)&(~g31223));
assign g30023 = (g28508&g20570);
assign II16010 = ((~g11148));
assign g14154 = ((~g11669))|((~g8958));
assign g7764 = (g2999)|(g2932);
assign g7247 = ((~g5377));
assign g23479 = ((~g21562));
assign g24430 = (g23151)|(g8234);
assign g32478 = ((~g31376));
assign g31256 = (g25983)|(g29537);
assign g32316 = (g31307&g23522);
assign g22341 = ((~g19801));
assign g22489 = (g12954&g19386);
assign g11027 = (g5097&g9724);
assign g19634 = ((~g16349));
assign II27538 = (g21209&g24132&g24133&g24134);
assign g24181 = ((~II23387));
assign g25728 = (g25076)|(g22011);
assign g18743 = (g5115&g17847);
assign g30097 = ((~g29118));
assign II29242 = ((~g29313));
assign g17700 = ((~g14792)&(~g12983));
assign g31304 = (g29594)|(g29608);
assign g11139 = (g5990&g7051&g5976&g9935);
assign g20186 = ((~g16926))|((~g8177));
assign g27732 = ((~g9364)&(~g25791));
assign g18990 = ((~g16136));
assign g32146 = (g31624&g29978);
assign g31769 = (g30141&g23986);
assign II12401 = ((~g3808))|((~g3813));
assign g32917 = ((~g30937));
assign g19908 = ((~g16540));
assign g31709 = ((~II29285))|((~II29286));
assign g31225 = (g30276&g21012);
assign g22224 = ((~g19277));
assign g30270 = (g28624)|(g27664);
assign g21451 = ((~II21162));
assign g21250 = ((~g9417)&(~g9340)&(~g17494));
assign g28675 = ((~g27779));
assign g21557 = (g12980&g15674);
assign g18892 = ((~g15680));
assign g21978 = (g5551&g19074);
assign g17119 = (g5272&g14800);
assign g23998 = (g19631&g10971);
assign g21934 = (g5220&g18997);
assign g32928 = ((~g31672));
assign II21959 = ((~g20242));
assign g12154 = ((~g10155)&(~g9835));
assign g22981 = ((~g20283));
assign g27432 = (g26519&g17582);
assign g24720 = ((~g1322)&(~g23051)&(~g19793));
assign g13019 = (g194&g11737);
assign g27459 = (g26549&g17609);
assign g14873 = ((~II16898));
assign g22906 = ((~g20453));
assign g23235 = ((~g20785));
assign g26732 = ((~g25389));
assign II18003 = ((~g13638));
assign g26636 = (g24897)|(g24884)|(g24858)|(g24846);
assign II31494 = ((~g33283));
assign g23997 = (g20602)|(g17191);
assign g21799 = (g3530&g20924);
assign g23515 = ((~g20785));
assign g7117 = ((~II11816));
assign g25619 = (g24961)|(g18193);
assign g10077 = ((~g1724));
assign II22799 = ((~g11960))|((~g21434));
assign g18691 = (g4727&g16053);
assign g31959 = (g4907&g30673);
assign g34150 = ((~II32103));
assign g19558 = ((~g15938));
assign g8880 = ((~II12861));
assign g15702 = ((~g13066))|((~g7293));
assign g20611 = ((~g18008));
assign g26362 = (g19557&g25538);
assign g25122 = (g23374&g20592);
assign g21792 = (g3396&g20391);
assign g10407 = ((~g7063));
assign g13865 = ((~II16168));
assign g32192 = ((~g31262));
assign g24373 = ((~g22908));
assign II17395 = ((~g12952));
assign g29116 = ((~g27837));
assign g16214 = ((~g13437));
assign g24854 = (g21453)|(g24002);
assign g13333 = (g4743&g11755);
assign g15862 = ((~II17355));
assign g14855 = ((~g12700))|((~g12824));
assign g29679 = ((~g153))|((~g28353))|((~g23042));
assign g11236 = ((~g8357));
assign g24941 = (g23171&g20190);
assign g7876 = ((~g1495));
assign g28101 = (g27691)|(g22062);
assign g12307 = ((~g7395))|((~g5983));
assign g16613 = (g5925&g14732);
assign g12048 = ((~g7369))|((~g2040));
assign g24663 = (g16621&g22974);
assign II13726 = ((~g4537));
assign g24063 = ((~g20014));
assign g24711 = ((~g23139));
assign g34061 = (g33800&g23076);
assign g31313 = (g30160&g27907);
assign g21952 = (g5366&g21514);
assign g29241 = (g28638)|(g18332);
assign g29345 = (g4749&g28376);
assign II25750 = ((~g26823));
assign g32948 = ((~g30735));
assign g33236 = (g32044)|(g32045);
assign g25893 = ((~g24541));
assign II24530 = (g9501&g9733&g5747);
assign g30155 = ((~II28390));
assign g23055 = ((~g20887));
assign g11444 = ((~g6905))|((~g6918))|((~g8733));
assign g25554 = ((~g22550));
assign g32419 = (g4955&g31000);
assign g23657 = (g19401&g11941);
assign II21815 = ((~g21308));
assign g32626 = ((~g30614));
assign g19436 = ((~g17176)&(~g14233));
assign g34906 = (g34857)|(g21694);
assign g34540 = ((~II32607));
assign g32270 = (g31254&g20444);
assign g25220 = ((~II24396));
assign g13070 = ((~g11984));
assign g33576 = (g33401)|(g18423);
assign g14261 = (g4507&g10738);
assign g34549 = ((~II32617));
assign g28180 = (g20242)|(g27511);
assign g34532 = (g34314&g19710);
assign g23005 = ((~g20283));
assign g27736 = ((~II26356));
assign g14772 = ((~g6044)&(~g12252));
assign g27956 = ((~II26466));
assign g18673 = (g4643&g15758);
assign g24569 = (g5115&g23382);
assign g20071 = ((~g16826));
assign g14255 = ((~g12381));
assign g20838 = ((~g5041))|((~g17284));
assign g12888 = ((~g10395));
assign g8879 = ((~II12858));
assign g33416 = (g32370&g21423);
assign g18195 = (g847&g17821);
assign g13941 = (g11019)|(g11023);
assign g12659 = ((~g9451)&(~g9392));
assign g26616 = (g24881)|(g24855)|(g24843)|(g24822);
assign g20632 = ((~g15171));
assign II31177 = (g32710&g32711&g32712&g32713);
assign g30035 = (g22539&g28120);
assign g25286 = ((~g22228));
assign g9912 = ((~II13463))|((~II13464));
assign g27134 = (g25997&g16602);
assign g30511 = (g30180)|(g22032);
assign II27519 = (g28036&g24107&g24108&g24109);
assign II22512 = ((~g19389));
assign g16840 = (g5467&g14262);
assign g25754 = (g25179)|(g22101);
assign g25651 = (g24680)|(g21744);
assign g28582 = (g27330)|(g26277);
assign II12799 = ((~g59));
assign g29553 = (g2437&g28911);
assign g25865 = (g25545&g18991);
assign g26953 = (g26486)|(g24291);
assign g16201 = ((~g13462)&(~g4704));
assign g32652 = ((~g30735));
assign g34784 = ((~II32982));
assign g28058 = (g27235)|(g18268);
assign g10218 = ((~g2527));
assign g25634 = (g24559)|(g18284);
assign g32110 = (g31639&g29921);
assign g23317 = (g19715)|(g16191);
assign g27568 = (g26576&g17791);
assign g30555 = (g30227)|(g22126);
assign g31308 = (g26101)|(g29614);
assign g23079 = ((~g8390)&(~g19965));
assign g34790 = (g34774)|(g18151);
assign g21926 = (g15147&g18997);
assign g33351 = (g32236&g20707);
assign g22941 = ((~g20219))|((~g2970));
assign g32067 = (g4727&g30614);
assign g33919 = (g33438&g10795);
assign g9898 = ((~g6444));
assign II22880 = (g21509)|(g21356)|(g21351);
assign g14051 = ((~g10323))|((~g11527));
assign g30178 = (g28632&g23815);
assign g8744 = ((~g691));
assign g31262 = ((~g767))|((~g29916))|((~g11679));
assign g31978 = ((~g30580))|((~g15591));
assign g32144 = (g30927)|(g30930);
assign g29916 = ((~g8681)&(~g28504)&(~g11083));
assign g33432 = ((~g31997)&(~g6978));
assign g8840 = ((~g4277));
assign g13870 = ((~g11773))|((~g4732));
assign g12332 = ((~II15167))|((~II15168));
assign g25646 = (g24706)|(g21739);
assign g17612 = ((~g15014));
assign g22338 = ((~g19801));
assign g33991 = (g33885)|(g18400);
assign g23905 = ((~g21514));
assign g34344 = (g34107&g20038);
assign II24680 = (g24029&g24030&g24031&g24032);
assign g11894 = ((~II14702));
assign g30306 = ((~g28796));
assign g24634 = (g22634&g19685);
assign g18589 = (g2902&g16349);
assign g23501 = ((~g20924));
assign g27724 = (g22417&g25208&g26424&g26190);
assign g12768 = (g7785)|(g7202);
assign g32643 = ((~g31376));
assign II31650 = ((~g33212));
assign g27876 = ((~II26418))|((~II26419));
assign II32607 = ((~g34358));
assign g11868 = ((~g9185));
assign g15117 = (g4300&g14454);
assign g29209 = ((~II27543));
assign II31327 = (g32928&g32929&g32930&g32931);
assign g11779 = ((~g9602));
assign g16709 = ((~II17919));
assign II17471 = ((~g13394));
assign g20922 = ((~II20891));
assign g24968 = (g22360)|(g22409)|(g23389);
assign g27011 = ((~g25917));
assign II33164 = ((~g34894));
assign II17699 = ((~g13416));
assign g26513 = (g19501&g24365);
assign II21181 = ((~g17413));
assign g13173 = ((~g10632));
assign g14572 = ((~g12169))|((~g9678));
assign g18666 = (g4593&g17367);
assign g11771 = ((~g8921)&(~g4185));
assign g30735 = (g29814&g22319);
assign g27327 = (g2116&g26732);
assign g26272 = (g2036&g25470);
assign II13321 = ((~g6486));
assign g17733 = ((~g14238));
assign g16136 = ((~II17491));
assign g34110 = (g33732&g22935);
assign g8822 = ((~g4975));
assign g31656 = ((~II29236));
assign II32202 = ((~g33937))|((~g33670));
assign g33045 = (g32206)|(g24328);
assign g11394 = ((~g9600))|((~g3661));
assign g29799 = (g28271&g10233);
assign g25114 = ((~II24278));
assign g25566 = ((~g22550));
assign g28229 = (g27345&g17213);
assign g26799 = (g25247&g21068);
assign g13068 = ((~II15697));
assign II31779 = ((~g33212));
assign g23662 = ((~g17393)&(~g20995));
assign g25540 = ((~g22409)&(~g22360));
assign g21711 = (g291&g20283);
assign g28456 = (g27290&g20104);
assign g26180 = (g2587&g25156);
assign g18701 = (g4771&g16856);
assign g28647 = (g27389)|(g16596);
assign g32524 = ((~g31070));
assign g31833 = ((~g29385));
assign g32083 = (g947&g30735);
assign g29534 = (g28965&g22457);
assign g9600 = ((~g3632));
assign g27216 = (g26055&g16725);
assign g15069 = ((~g6828)&(~g13416));
assign g7749 = ((~g996));
assign g14911 = ((~g10213)&(~g12364));
assign II15078 = ((~g9827))|((~g1968));
assign II22601 = ((~g21127));
assign g17389 = ((~g14915));
assign II23330 = ((~g22658));
assign g10615 = ((~g1636)&(~g7308));
assign g33953 = (g33487)|(II31848)|(II31849);
assign g30355 = (g30131)|(g18360);
assign g11432 = ((~g10295))|((~g8864));
assign g9071 = ((~g2831));
assign g25801 = (g8097&g24585);
assign g27042 = (g25774&g19343);
assign g13637 = ((~g10556));
assign g20266 = ((~g17873));
assign g12416 = ((~g10133))|((~g7064))|((~g10166));
assign g23811 = (g4087&g19364);
assign g27146 = (g26148&g8187&g1648);
assign g23647 = ((~g18833));
assign g28083 = (g27249)|(g18689);
assign g23839 = ((~g18997));
assign II25847 = ((~g24799))|((~II25845));
assign g10551 = ((~g1728))|((~g7356));
assign g26289 = (g2551&g25400);
assign g25039 = ((~g22498));
assign g29549 = (g2012&g28900);
assign g28155 = ((~II26664));
assign g11724 = ((~II14593));
assign g8146 = ((~g1760));
assign II18270 = ((~g13191));
assign g16776 = ((~g3945))|((~g13772))|((~g4012))|((~g11419));
assign g26341 = (g24746&g20105);
assign g35001 = ((~II33297));
assign g27358 = (g26400&g17415);
assign g13279 = ((~II15843));
assign g26956 = (g26487)|(g24294);
assign g22522 = ((~g19699)&(~g1024));
assign g6782 = ((~II11632));
assign g20435 = ((~g15348));
assign g14822 = ((~g12755))|((~g12632));
assign g19916 = ((~g3029))|((~g16313));
assign II26654 = ((~g27576));
assign g29593 = (g28470&g7985);
assign g34788 = ((~II32994));
assign g12159 = ((~g8765))|((~g4864));
assign g23202 = ((~II22302));
assign g29896 = (g2599&g29171);
assign g29366 = (g13738)|(g28439);
assign g18437 = (g2241&g18008);
assign g13043 = ((~g10521))|((~g969));
assign g18124 = (g102&g16886);
assign g34823 = ((~II33037));
assign g32720 = ((~g31710));
assign g24129 = ((~g20857));
assign g25465 = ((~g23824));
assign g29272 = (g28346)|(g18638);
assign II17381 = ((~g1129))|((~II17379));
assign g24453 = ((~g7446)&(~g22325));
assign g27585 = ((~g25994));
assign g32242 = (g31245&g20324);
assign g23425 = ((~g20751));
assign g12418 = ((~g9999)&(~g10001));
assign g30260 = ((~g7018)&(~g28982));
assign II18364 = ((~g13009));
assign g33521 = (g32895&II31301&II31302);
assign II17842 = ((~g13051));
assign g18144 = (g590&g17533);
assign g16728 = ((~g13884))|((~g13870))|((~g14089))|((~g11639));
assign g33212 = (g32328)|(II30755)|(II30756);
assign II31086 = (g31554&g31811&g32578&g32579);
assign g21699 = (g142&g20283);
assign g18878 = ((~g15426));
assign g8179 = ((~g4999));
assign g13105 = ((~g10671))|((~g7675))|((~g1322))|((~g1404));
assign g16732 = (g5555&g14882);
assign g16624 = ((~II17814));
assign g30312 = ((~g28970));
assign g10719 = (g6841&g2138&g2130);
assign g33933 = ((~g33394))|((~g12491))|((~g12819))|((~g12796));
assign g14449 = ((~g12194)&(~g9653));
assign g23881 = ((~g19277));
assign g11024 = (g5436&g9070);
assign g11547 = ((~II14505));
assign g13679 = ((~g10573));
assign g16954 = ((~II18104));
assign II18680 = ((~g2638))|((~g14752));
assign g24126 = ((~g19935));
assign g34708 = (g33381)|(g34572);
assign g24464 = (g3480&g23112);
assign g28387 = (g27203)|(g15858);
assign g7689 = ((~II12159));
assign gbuf98 = (g4019);
assign g7831 = ((~II12227));
assign g20105 = ((~g17433));
assign g12050 = ((~g10038)&(~g9649));
assign g30000 = (g23685&g29029);
assign g24701 = ((~g979)&(~g23024)&(~g19778));
assign g16205 = (g11547&g6782&g11640&II17542);
assign II31863 = (g33506)|(g33507)|(g33508)|(g33509);
assign g11897 = ((~II14705));
assign g19531 = ((~g16816));
assign g20701 = ((~g17955));
assign g31965 = ((~g30583)&(~g4358));
assign g18943 = (g269&g16099);
assign g21461 = ((~g15348));
assign g27287 = (g26545&g23011);
assign g16853 = ((~g13584));
assign II30998 = ((~g32453));
assign g19536 = (g518&g16768);
assign g30015 = (g29040&g10519);
assign g8847 = ((~g4831))|((~g4681));
assign g24301 = (g6961&g22228);
assign g23936 = ((~g19210));
assign g33547 = (g33349)|(g18331);
assign II13518 = ((~g2514))|((~g2518));
assign g27410 = (g26549&g17527);
assign g21604 = ((~g15938));
assign g22109 = (g6455&g18833);
assign II12360 = ((~g528));
assign II12000 = ((~g582));
assign g24101 = ((~g20998));
assign gbuf14 = (g4815);
assign g10083 = ((~g2407));
assign g26921 = (g25955)|(g18285);
assign g32701 = ((~g31376));
assign g25438 = ((~g22763));
assign g23262 = (g19661)|(g16126);
assign g8993 = ((~g385));
assign g29722 = ((~g28410))|((~g13742));
assign g33554 = (g33407)|(g18353);
assign g25492 = ((~g12479))|((~g22457));
assign g21048 = ((~g17533));
assign g34946 = ((~g34934));
assign g29694 = ((~g28391))|((~g13709));
assign II28872 = ((~g30072));
assign g29375 = (g13946&g28370);
assign II25908 = ((~g26256))|((~II25907));
assign II28585 = ((~g30217));
assign g10419 = ((~g8821));
assign II33056 = ((~g34778));
assign g33911 = (g33137&g10725);
assign g18275 = (g15070&g16136);
assign g11841 = ((~g9800));
assign g28345 = (g27137)|(g15821);
assign g8632 = ((~g1514))|((~g1500));
assign g16210 = ((~g13479)&(~g4894));
assign g11166 = (g8363&g269&g8296&II14225);
assign g23925 = ((~g21514));
assign g23204 = ((~g10685)&(~g19462)&(~g16488));
assign g7704 = ((~II12167));
assign g26911 = (g26612)|(g24230);
assign g8715 = ((~g4927));
assign II18138 = ((~g14277));
assign g20383 = ((~g15373));
assign II25695 = ((~g25690));
assign g19611 = ((~g1070))|((~g1199))|((~g15995));
assign g14197 = ((~g12160));
assign g24685 = ((~g23139));
assign g24793 = ((~g3742))|((~g23124));
assign g8259 = ((~g2217));
assign g12761 = (g969&g7567);
assign g25521 = ((~g23955)&(~g14645));
assign g21292 = ((~II21033));
assign g18882 = ((~II19674));
assign g25601 = (g24660)|(g18112);
assign g22432 = (g9354&g7717&g21187);
assign g22938 = (g19782&g19739);
assign g12150 = ((~g2208)&(~g8259));
assign g13624 = ((~g10951));
assign g18750 = (g15145&g17847);
assign g15992 = ((~g10929)&(~g13846));
assign g33568 = (g33409)|(g18395);
assign g23332 = ((~g20785));
assign g18425 = (g2161&g18008);
assign g22846 = (g9386&g20676);
assign g28758 = ((~g27779))|((~g7356))|((~g7275));
assign g30612 = (g26338&g29597);
assign g12969 = ((~g4388))|((~g7178))|((~g10476));
assign g29094 = ((~g27858))|((~g9700));
assign g10074 = ((~g718));
assign g32201 = ((~g31509));
assign g8080 = ((~g3863));
assign g19478 = ((~g16000));
assign g24020 = ((~g20014));
assign g25772 = (g24944&g24934);
assign g13831 = ((~g11245)&(~g7666));
assign g18324 = (g1644&g17873);
assign g19754 = ((~g17062));
assign g19882 = ((~g16540));
assign g21378 = (g7887&g16090);
assign g23209 = (g19585)|(g19601);
assign g34578 = (g24578&g34308);
assign g15573 = ((~II17154));
assign g33515 = (g32853&II31271&II31272);
assign g10819 = ((~g7479)&(~g1041));
assign g16742 = ((~g13983));
assign g19671 = (g1454&g16155);
assign g16285 = ((~II17612));
assign II18031 = ((~g13680));
assign g14656 = ((~g12553))|((~g12405));
assign g9484 = ((~g1612));
assign g25666 = (g24788)|(g21793);
assign g29584 = (g1706&g29018);
assign g27149 = (g25997&g16623);
assign g32237 = (g31153)|(g29667);
assign II22725 = ((~g21250));
assign g27163 = ((~II25869));
assign g24050 = ((~g20841));
assign g13015 = ((~g11875));
assign g24235 = (g22632)|(g18238);
assign g27371 = (g26400&g17473);
assign II18728 = ((~g6012));
assign g25501 = ((~g23918)&(~g14645));
assign g24213 = (g23220)|(g18186);
assign II20690 = ((~g15733));
assign g30561 = (g30284)|(g22132);
assign g14584 = ((~g11048));
assign g28724 = (g27491)|(g16707);
assign g8353 = ((~II12530));
assign g8217 = ((~g3143));
assign g11968 = ((~g837))|((~g9334))|((~g9086));
assign g9051 = ((~g1426));
assign II16646 = (g10160&g12413&g12343);
assign g24723 = (g17490&g22384);
assign g32193 = (g30732&g25410);
assign g24774 = (g718&g23614);
assign g24336 = (g24012)|(g18753);
assign g18560 = (g2837&g15277);
assign g29358 = ((~II27718));
assign g28061 = (g27287)|(g21735);
assign g33372 = (g32285&g21183);
assign g30148 = ((~g28799)&(~g7335));
assign g22169 = ((~g19147));
assign g13569 = ((~g10951));
assign g20633 = ((~g15171));
assign g32421 = ((~g31213));
assign g13141 = ((~g11374));
assign g18765 = (g5489&g17929);
assign g18461 = (g2307&g15224);
assign g7623 = ((~II12103));
assign g34569 = ((~II32639));
assign II16803 = ((~g6369));
assign g25868 = (g25450)|(g23885);
assign g15613 = (g3490&g13555);
assign g20596 = ((~II20690));
assign g24109 = ((~g21143));
assign II23312 = ((~g21681));
assign g27592 = ((~g26715));
assign g24076 = ((~g19984));
assign g28252 = (g27159&g19682);
assign g30217 = ((~II28458));
assign g27553 = (g26293&g23353);
assign g24621 = ((~g22957))|((~g2927));
assign g27534 = (g26488&g17735);
assign g23082 = ((~g21024));
assign g20607 = ((~g17955));
assign g18587 = (g2980&g16349);
assign g24514 = ((~g23619)&(~g23657));
assign g23187 = (g13989&g20010);
assign g34336 = ((~g34112));
assign g30163 = (g23381)|(g28523);
assign g23342 = ((~g6928))|((~g21163));
assign g29786 = (g22843)|(g28240);
assign II14630 = ((~g7717));
assign g12487 = ((~g9340));
assign II15316 = ((~g10087));
assign g34095 = (g33681)|(g33687);
assign g28561 = (g27312)|(g26250);
assign g22831 = (g19441&g19629);
assign g26885 = (g26541)|(g24191);
assign g13808 = (g4543&g10607);
assign II29363 = ((~g30218));
assign g21660 = ((~g17694));
assign g17599 = ((~g14794));
assign g19071 = ((~g15591));
assign g24817 = (g22929&g7235);
assign g13130 = ((~g1351))|((~g11815))|((~g11336));
assign g34084 = (g9214&g33851);
assign g34473 = ((~g34426));
assign g32836 = ((~g31021));
assign g27824 = ((~II26394))|((~II26395));
assign g29877 = (g28405&g23340);
assign g19999 = ((~g16232)&(~g13742));
assign g29589 = (g2575&g28977);
assign g10358 = ((~g6827));
assign g28094 = (g27673)|(g21959);
assign g31631 = ((~II29221));
assign g10476 = (g7244&g7259&II13862);
assign g34441 = (g34381)|(g18540);
assign g18989 = ((~g16000));
assign g30070 = (g29167&g9529);
assign g34637 = (g34478)|(g18694);
assign g20612 = ((~g18008));
assign g10804 = ((~g9772));
assign g18606 = (g3133&g16987);
assign g17308 = ((~g14876));
assign g20903 = ((~g17249));
assign g22217 = (g21302)|(g17617);
assign g28105 = (g27997)|(g22135);
assign g34798 = (g34754)|(g18575);
assign II28349 = ((~g28367));
assign g9759 = ((~g2265));
assign g32555 = ((~g30673));
assign gbuf91 = (g3447);
assign II18060 = ((~g14198));
assign g28589 = (g27331)|(g26285);
assign gbuf52 = (g6322);
assign g21959 = (g5413&g21514);
assign g30921 = (g29900&g24789);
assign g10371 = ((~g6918));
assign g34752 = (g34675&g19544);
assign g33503 = (g32765&II31211&II31212);
assign II31321 = (g31376&g31852&g32919&g32920);
assign g29753 = (g28213)|(g22720);
assign g34324 = (g14064&g34161);
assign II16150 = ((~g10430));
assign g20640 = ((~g15426));
assign g31142 = (g2527&g30039);
assign g22074 = (g6239&g19210);
assign g8440 = ((~g3431));
assign g14063 = ((~g11048));
assign g28783 = ((~g27779))|((~g7315))|((~g1728));
assign g24117 = ((~g21209));
assign g20148 = (g16128)|(g13393);
assign g32094 = (g30612)|(g29363);
assign g32710 = ((~g30825));
assign g20875 = (g16281&g4681);
assign g27667 = (g26361&g20601);
assign g17506 = (g9744&g14505);
assign II29239 = ((~g29498));
assign g21995 = (g5611&g19074);
assign g18774 = (g5698&g15615);
assign g9462 = ((~g6215));
assign g16616 = (g6267&g14741);
assign g28321 = ((~g27317));
assign g21270 = ((~II20999));
assign g34318 = (g25850)|(g34063);
assign g12350 = ((~II15190));
assign g23605 = ((~g20739));
assign g34557 = (g34352&g20555);
assign g13698 = ((~g528)&(~g12527)&(~g11185));
assign g21361 = (g7869&g16066);
assign g30589 = (g18898&g29811);
assign g19334 = ((~II19818));
assign g32272 = (g31639&g30310);
assign g24418 = ((~g22722));
assign g34019 = (g33889)|(g18506);
assign g9479 = (g305&g324);
assign II12805 = ((~g4098));
assign g15820 = (g3578&g13955);
assign g28391 = ((~g27064))|((~g13637));
assign II15341 = ((~g10154))|((~II15340));
assign g8734 = ((~g4045));
assign g32597 = ((~g31154));
assign g14366 = ((~II16526));
assign g11147 = ((~g8417));
assign g18229 = (g1099&g16326);
assign g22640 = (g18951)|(g15613);
assign g27120 = (g25878&g22543);
assign g11991 = ((~g9485));
assign g10118 = ((~g2541));
assign g34641 = (g34479)|(g18724);
assign g16663 = ((~g13854))|((~g13834))|((~g14655))|((~g12292));
assign g9220 = ((~g843));
assign II18313 = ((~g13350));
assign g26937 = ((~II25683));
assign g28520 = ((~g8229)&(~g27635));
assign g22202 = ((~II21784));
assign II26093 = ((~g26055))|((~g13539));
assign II27509 = (g24084&g24085&g24086&g24087);
assign g17057 = (g446&g13173);
assign g14034 = ((~g11048));
assign g34876 = (g34844&g20534);
assign g32256 = (g31249&g20382);
assign g30928 = ((~II28908));
assign g27230 = (g25906&g19558);
assign g30540 = (g30275)|(g22086);
assign g19517 = ((~g16777));
assign g25133 = ((~g23733));
assign g30267 = (g28776&g23967);
assign g28709 = ((~II27192));
assign g22623 = (g19337&g19470);
assign g26394 = (g22530&g25560);
assign g24135 = ((~g20720));
assign g21842 = (g3863&g21070);
assign g25368 = (g6946&g22408);
assign g7216 = ((~g822));
assign g27652 = ((~g3355)&(~g26636));
assign g17412 = ((~g14520))|((~g14489));
assign g21457 = ((~g17367));
assign g7490 = ((~g2629));
assign g34772 = ((~II32960));
assign g30470 = (g30165)|(g21941);
assign g33264 = (g31965&g21306);
assign g22408 = ((~g19483));
assign g33384 = (g32248)|(g29943);
assign II23755 = (g22904)|(g22927)|(g22980)|(g23444);
assign g28540 = ((~g8125)&(~g27635)&(~g7121));
assign g30079 = ((~g29097));
assign g14418 = ((~g12151)&(~g9594));
assign g33674 = (g33164&g10710&g22319);
assign g18095 = ((~II18891));
assign g32888 = ((~g30673));
assign g21700 = (g150&g20283);
assign g16515 = ((~g13486));
assign g24962 = (g23194&g20210);
assign g27768 = ((~g9264)&(~g25805));
assign g30456 = (g29378)|(g21869);
assign g13882 = ((~g3590))|((~g11207))|((~g3672))|((~g11576));
assign g17601 = (g9616&g14572);
assign g20127 = ((~II20388));
assign g30126 = (g28582&g21058);
assign g31918 = (g31786)|(g22015);
assign g24110 = ((~g21209));
assign g16224 = (g14583&g14232);
assign g34871 = (g34823&g19908);
assign g22034 = (g5929&g19147);
assign g22015 = (g5719&g21562);
assign g28431 = ((~II26925));
assign g21786 = (g3436&g20391);
assign g8686 = ((~g2819));
assign g27095 = (g25997&g16473);
assign g30299 = ((~g28765));
assign II12271 = ((~g956))|((~II12269));
assign II31186 = (g31376&g31828&g32724&g32725);
assign II12241 = ((~g1111))|((~II12240));
assign g19480 = ((~g16349));
assign II31012 = (g32473&g32474&g32475&g32476);
assign g26542 = (g13102&g24376);
assign g18877 = ((~g15224));
assign g33241 = (g32173&g23128);
assign g28558 = (g7301&g27046);
assign g6887 = ((~g3333));
assign g13858 = (g209)|(g10685);
assign g32646 = ((~g31070));
assign II22974 = ((~g19638))|((~II22972));
assign g18621 = (g3476&g17062);
assign g7405 = ((~g1936));
assign g20068 = ((~g11293))|((~g17794));
assign g25003 = ((~g21353))|((~g23462));
assign g21778 = (g3355&g20391);
assign g7970 = ((~g4688));
assign g21393 = ((~g17264));
assign g29525 = (g2169&g28837);
assign g28965 = ((~g27882))|((~g8255));
assign g18499 = (g2476&g15426);
assign II21769 = ((~g19402));
assign g25030 = (g23251&g20432);
assign g30468 = (g30238)|(g21939);
assign g18321 = (g1620&g17873);
assign g29648 = (g2112&g29121);
assign g25838 = ((~g25250));
assign g12076 = ((~g9280));
assign II32093 = ((~g33670));
assign g13920 = ((~g11621))|((~g11483));
assign g34734 = (g34681)|(g18652);
assign g24066 = ((~g21127));
assign g33848 = (g33261&g20384);
assign II22280 = (g20271)|(g20150)|(g20134);
assign g20555 = ((~g15480));
assign g31881 = (g31018)|(g21775);
assign g27491 = (g26576&g17652);
assign g13799 = ((~g8584)&(~g11663));
assign g23304 = ((~g20785));
assign g29876 = (g28404&g23339);
assign g34668 = ((~II32788));
assign g7116 = ((~g22));
assign g32428 = (g31133&g16261);
assign g18831 = ((~g15224));
assign g33467 = (g32505&II31031&II31032);
assign II32621 = ((~g34335));
assign g30538 = (g30256)|(g22084);
assign g27254 = (g25935&g19688);
assign II21994 = ((~g19638))|((~II21992));
assign g30515 = (g30223)|(g22036);
assign g23192 = ((~g20248));
assign g31168 = (g2241&g30077);
assign g20979 = ((~g5385))|((~g17309));
assign g30194 = (g28651&g23849);
assign g19385 = ((~g16326));
assign g25756 = (g25112)|(g22103);
assign g12995 = ((~g11820));
assign g11676 = ((~g358))|((~g8944))|((~g376))|((~g385));
assign g32493 = ((~g30735));
assign g28548 = (g27303)|(g26232);
assign g23193 = (g19556)|(g15937);
assign g22304 = (g21347)|(g17693);
assign g12923 = ((~II15542));
assign g22021 = (g5869&g19147);
assign g16631 = ((~g14454));
assign g10184 = ((~g4486));
assign g13242 = (g11336)|(g7601);
assign g19963 = ((~g16326));
assign g18706 = (g4785&g16782);
assign g10823 = (g7704&g5180&g5188);
assign g19755 = ((~g15915));
assign g27634 = (g26805&g26793);
assign g24349 = (g23646)|(g18805);
assign g13521 = ((~g11357));
assign g14611 = ((~g12333)&(~g9749));
assign g25880 = (g8443&g24814);
assign g18312 = (g1579&g16931);
assign g16692 = ((~g14170));
assign g29312 = ((~g28877));
assign g22763 = ((~II22046));
assign g28339 = (g9946&g27693);
assign g33558 = (g33350)|(g18364);
assign g11976 = ((~g9595)&(~g7379));
assign g28651 = (g27392)|(g16599);
assign g32881 = ((~g30673));
assign g20325 = ((~g15171));
assign g14331 = ((~II16489));
assign g34016 = (g33867)|(g18503);
assign g16449 = ((~II17679));
assign g14868 = ((~g12755))|((~g12680));
assign g33409 = (g32359&g21408);
assign g20651 = ((~g15483));
assign g24447 = (g10948)|(g22450);
assign gbuf37 = (g6005);
assign g34211 = (g33891&g21349);
assign g10509 = ((~g10233));
assign g21418 = ((~g17821));
assign g22497 = ((~g19513));
assign g34884 = (g34858)|(g21666);
assign g7674 = ((~II12151));
assign g29991 = (g29179&g12922);
assign g26358 = (g19522&g25528);
assign g25675 = (g24769)|(g21832);
assign g10266 = ((~g5188)&(~g5180));
assign g9439 = ((~g5428));
assign g22713 = ((~g20114))|((~g2890));
assign g23619 = (g19453&g13045);
assign g14676 = ((~II16775));
assign g19388 = ((~g17181)&(~g14256));
assign g21960 = (g5421&g21514);
assign g34615 = (g34516)|(g18576);
assign g26607 = ((~g25382));
assign II27504 = (g24077&g24078&g24079&g24080);
assign II25534 = ((~g25448));
assign g24803 = (g22901&g20005);
assign g9510 = ((~g5835));
assign g30398 = (g29749)|(g21757);
assign g13967 = ((~g3929))|((~g11225))|((~g3983))|((~g11419));
assign g15147 = ((~g13716)&(~g12892));
assign II21911 = ((~g21278));
assign g32099 = ((~g31009));
assign g8237 = ((~g255));
assign II24920 = ((~g25513));
assign g13005 = ((~g7939)&(~g10762));
assign II24416 = ((~g14382))|((~II24414));
assign II31251 = (g31710&g31840&g32817&g32818);
assign g32904 = ((~g30735));
assign g33995 = (g33848)|(g18425);
assign g29551 = (g2173&g28867);
assign g15142 = ((~g13680)&(~g12889));
assign g34609 = (g34503)|(g18563);
assign g12017 = ((~g9969)&(~g9586));
assign g24477 = ((~II23680));
assign g20444 = ((~g15373));
assign g28491 = ((~g8114)&(~g27617));
assign g30259 = ((~g28463));
assign g29238 = (g28178)|(g18292);
assign g34893 = ((~II33119));
assign II20793 = ((~g17694));
assign g29801 = (g25987)|(g28251);
assign g9699 = ((~g2311));
assign g23650 = ((~g20653));
assign g25091 = (g12830&g23492);
assign g18305 = (g1521&g16489);
assign g15749 = (g1454&g13273);
assign g26095 = (g11923&g25090);
assign II15494 = ((~g10385));
assign g6918 = ((~g3639));
assign II16129 = (g8728&g11443&g11411);
assign g21898 = (g20152)|(g15112);
assign g8411 = ((~II12577));
assign g31499 = (g29801&g23446);
assign g22752 = (g15792&g19612);
assign g28551 = (g27305)|(g26234);
assign g31906 = (g31477)|(g21953);
assign g25595 = (g24835)|(g21717);
assign g17197 = ((~II18233));
assign g20165 = (g5156&g17733);
assign g33283 = (g31995)|(g30318);
assign II15087 = ((~g9832))|((~g2393));
assign g28234 = (g27877&g26686);
assign g18168 = (g681&g17433);
assign II14905 = ((~g9822));
assign g33840 = (g33253&g20267);
assign g28679 = (g27572&g20638);
assign g25229 = (g7636&g22654);
assign II31356 = (g31327&g31859&g32968&g32969);
assign g25166 = (g17506&g23571);
assign g27966 = ((~g7153)&(~g25805));
assign g34670 = ((~II32794));
assign g9518 = ((~g6219));
assign g8805 = ((~II12799));
assign g33486 = (g32642&II31126&II31127);
assign g9682 = ((~II13280));
assign g27539 = (g26576&g17745);
assign g19452 = ((~g16326));
assign g32810 = ((~g31376));
assign II21162 = ((~g17292));
assign g13215 = ((~g10909));
assign g33969 = (g33864)|(g18321);
assign II12493 = ((~g5002));
assign g24141 = (g17657&g21656);
assign g21681 = ((~II21242));
assign g14164 = ((~g9000)&(~g12259));
assign g22160 = (g8005&g19795);
assign g13341 = ((~g7863)&(~g10762));
assign g17480 = (g9683&g14433);
assign g33921 = (g33187&g9104&g19200);
assign g34268 = (g34082)|(g18730);
assign II16246 = ((~g3983));
assign g15733 = ((~II17249));
assign g27469 = (g8046&g26314&g518&g9077);
assign g22040 = (g5953&g19147);
assign g34161 = ((~g33851));
assign II16778 = ((~g11292))|((~g12332));
assign g30362 = (g30120)|(g18392);
assign II18842 = ((~g13809));
assign g21054 = ((~g15373));
assign g32818 = ((~g30735));
assign II29225 = ((~g30311));
assign g29732 = (g2514&g29131);
assign g18575 = (g2878&g16349);
assign g32845 = ((~g30673)&(~II30399)&(~II30400));
assign g26904 = (g26393)|(g24221);
assign g20215 = (g16479&g10476);
assign g16597 = (g6263&g15021);
assign g21398 = ((~g18008));
assign g29605 = (g2445&g28973);
assign II24695 = (g24050&g24051&g24052&g24053);
assign g24174 = ((~II23366));
assign g33022 = (g32306)|(g21750);
assign g24761 = (g22751&g19852);
assign g24797 = (g22872&g19960);
assign II29585 = ((~g31655));
assign g7515 = ((~II12000));
assign g28143 = (g27344&g26083);
assign g12285 = ((~II15122))|((~II15123));
assign II31247 = (g32812&g32813&g32814&g32815);
assign g12857 = ((~II15474));
assign g8567 = ((~g4082));
assign g33009 = (g32273)|(g18458);
assign g34746 = (g34670&g19526);
assign g13209 = ((~g10632));
assign g19526 = ((~g16349));
assign g33697 = (g33160&g13330);
assign g27967 = ((~II26479));
assign g29969 = (g28121&g20509);
assign g10151 = ((~g1992));
assign g19606 = ((~g17614));
assign g18162 = (g686&g17433);
assign II32834 = ((~g34472));
assign II12746 = ((~g4087));
assign g18528 = ((~II19348));
assign g23548 = ((~g18833));
assign g9535 = (g209)|(g538);
assign II14939 = ((~g10216));
assign g8751 = ((~g3969))|((~g4012))|((~g3983))|((~g4005));
assign g25447 = ((~g23883)&(~g14645));
assign g9498 = ((~g5101));
assign g15132 = ((~g12882)&(~g13638));
assign g20372 = ((~g17847));
assign g13545 = ((~II16010));
assign II31791 = ((~g33354));
assign g29252 = (g28712)|(g18486);
assign g26094 = (g24936&g9664);
assign g32291 = (g31268&g20527);
assign g14037 = ((~g8748)&(~g11083));
assign g25787 = (g24792&g20887);
assign g25154 = ((~g22457));
assign II14679 = ((~g9332));
assign g13115 = ((~g1008))|((~g11786))|((~g11294));
assign g33626 = (g33374)|(g18825);
assign g11356 = ((~g9552))|((~g3632));
assign g16184 = (g9285&g14183);
assign g27242 = ((~g26183));
assign g29951 = (g1874&g28786);
assign g24130 = ((~g20998));
assign g19359 = (g17786)|(g14875);
assign g11173 = ((~g4966))|((~g7898))|((~g9064));
assign g19145 = (g8450&g16200);
assign g6856 = ((~II11682));
assign g17174 = ((~g9194)&(~g14279));
assign g31170 = (g19128&g29814);
assign g24329 = (g4462&g22228);
assign II22800 = ((~g11960))|((~II22799));
assign g14434 = ((~g6415))|((~g11945));
assign g34209 = ((~II32170));
assign g15730 = ((~g6609))|((~g14556))|((~g6711))|((~g10061));
assign g17430 = ((~II18373));
assign g21366 = ((~II21100));
assign g10381 = ((~g6957));
assign II20895 = ((~g16954));
assign g32031 = (g31372&g13464);
assign g26694 = (g24444)|(g10704);
assign g15049 = ((~g13350)&(~g6799));
assign g30408 = (g29806)|(g21767);
assign g28650 = (g27391)|(g16598);
assign II14158 = ((~g8806));
assign II25244 = ((~g24744))|((~II25242));
assign g24221 = (g232&g22594);
assign g16098 = (g5148&g14238);
assign g26546 = ((~g24858)&(~g24846));
assign g27382 = ((~g8219)&(~g26657));
assign g6831 = ((~g1413));
assign II17780 = ((~g13303));
assign g22865 = ((~g20330));
assign g11429 = ((~g7616));
assign g16764 = (g6307&g14776);
assign g25219 = ((~II24393));
assign g32368 = (g29881)|(g31310);
assign II13031 = ((~g6747));
assign g30274 = (g28815&g23983);
assign g32638 = ((~g30825));
assign g20173 = ((~g16696))|((~g13972));
assign g25264 = ((~g23828));
assign g15162 = ((~g13809)&(~g12904));
assign g34951 = ((~g34941));
assign g34261 = (g34074)|(g18688);
assign g11823 = ((~II14647));
assign g34841 = (g34761&g20080);
assign g28493 = ((~g3873)&(~g27635));
assign g7027 = ((~g5499));
assign g8398 = ((~II12563));
assign g10532 = ((~g10233));
assign g28188 = (g22535)|(g27108);
assign II18909 = ((~g16873));
assign g33941 = (g33380&g21560);
assign g21759 = (g3199&g20785);
assign II18822 = ((~g13745));
assign g12117 = ((~g10113)&(~g9755));
assign g14003 = ((~g9003)&(~g11083));
assign g16119 = ((~II17475))|((~II17476));
assign gbuf106 = (g4191);
assign g22659 = (g19062)|(g15673);
assign g34596 = ((~II32696));
assign g32388 = (g31495)|(g29962);
assign g24204 = (g22990)|(g18108);
assign g30180 = (g28635&g23820);
assign g23759 = ((~II22886));
assign g8279 = ((~II12487));
assign g13325 = ((~g7841)&(~g10741));
assign g32824 = ((~g31376));
assign g13868 = ((~g11493));
assign g29509 = (g1600&g28755);
assign g18769 = (g15151&g18062);
assign g21512 = (g16225&g10881);
assign g15139 = ((~g12886)&(~g13680));
assign g9373 = ((~g5142));
assign g26337 = ((~g24818));
assign g21382 = (g10086&g17625);
assign g32900 = ((~g30937));
assign g34867 = (g34826&g20145);
assign g25928 = (g25022&g23436);
assign g32789 = ((~g30735));
assign g18434 = (g2217&g18008);
assign II27523 = (g20857&g24111&g24112&g24113);
assign g18485 = (g2465&g15426);
assign g30997 = ((~g29702));
assign g10677 = (g4141&g7611);
assign g13500 = ((~g8480)&(~g12641));
assign g28308 = (g27105)|(g15795);
assign II14992 = ((~g9685))|((~II14991));
assign g10756 = (g3990&g6928&g3976&g8595);
assign g16960 = ((~II18114));
assign g22197 = ((~g19074));
assign g15042 = ((~g12806))|((~g10491));
assign g18944 = ((~g15938));
assign g22056 = (g6133&g21611);
assign II32195 = ((~g33628));
assign II18858 = ((~g13835));
assign g28202 = (g27659&g11413);
assign g18454 = (g2303&g15224);
assign g7471 = ((~g6012));
assign II21210 = ((~g17526));
assign g32450 = ((~g31591));
assign g18110 = (g441&g17015);
assign g23918 = ((~g2799)&(~g21382));
assign g32044 = (g31483&g20085);
assign g9472 = ((~g6555));
assign g24273 = (g23166)|(g18630);
assign g10057 = ((~g6455));
assign g17788 = ((~g5232))|((~g14490))|((~g5327))|((~g12497));
assign II22717 = ((~g11916))|((~g21434));
assign II22710 = ((~g11915))|((~g21434));
assign g22523 = ((~g1345)&(~g19720));
assign g27329 = (g12052&g26743);
assign g32784 = ((~g31672));
assign g32117 = (g24482)|(g30914);
assign g11797 = ((~g8883)&(~g8796));
assign g21902 = ((~II21477));
assign g27704 = ((~g7239)&(~g25791));
assign II21300 = ((~g18598));
assign g23612 = ((~II22745));
assign g18553 = (g2827&g15277);
assign II13684 = ((~g128));
assign g12238 = ((~II15102));
assign g14758 = ((~g7704))|((~g12405));
assign g28095 = (g27674)|(g21970);
assign II26051 = ((~g13500))|((~II26049));
assign g34413 = (g34094&g22670);
assign g26314 = ((~g24808)&(~g24802));
assign II24552 = (g9733&g9316&g5747);
assign g33688 = ((~II31523));
assign g34072 = (g33839&g24872);
assign II20460 = ((~g17515))|((~g14187));
assign g17532 = ((~II18479));
assign II20816 = ((~g17088));
assign g12160 = ((~g9721)&(~g9724));
assign g11959 = ((~g8316))|((~g2342));
assign g32657 = ((~g31528));
assign II14576 = ((~g8791));
assign g30498 = (g30251)|(g21994);
assign g6873 = ((~g3151));
assign g18723 = (g4922&g16077);
assign g32322 = (g31308&g20605);
assign g25417 = (g5712&g23816&II24552);
assign g18783 = (g5841&g18065);
assign g34217 = (g33736&g22876);
assign g7620 = ((~II12097))|((~II12098));
assign g12578 = ((~g7791))|((~g10341));
assign g18378 = (g1932&g15171);
assign g32183 = (g2795&g31653);
assign g22095 = (g6428&g18833);
assign g10946 = ((~g1489))|((~g7876));
assign g27341 = (g10203&g26788);
assign g29956 = ((~II28185));
assign g17481 = ((~g15005));
assign g30507 = (g30190)|(g22028);
assign II31126 = (g30673&g31818&g32636&g32637);
assign g18824 = (g6732&g15680);
assign g29949 = (g23575&g28924);
assign g21783 = (g3419&g20391);
assign g20532 = ((~g15277));
assign II20495 = ((~g16283));
assign g18255 = (g1087&g16897);
assign g15902 = (g441&g13975);
assign g28481 = ((~g3506)&(~g10323)&(~g27617));
assign g15582 = (g8977)|(g12925);
assign II31081 = (g30673&g31810&g32571&g32572);
assign g32277 = (g31211)|(g29733);
assign g12195 = ((~g2619))|((~g8381));
assign g16195 = ((~g13437));
assign II19851 = ((~g16615));
assign g26104 = (g2250&g25101);
assign g9434 = ((~g5385));
assign g26293 = (g24550)|(g24555);
assign g25901 = (g24853&g16290);
assign g28624 = (g22357&g27009);
assign g34434 = ((~II32473));
assign g33149 = (g32204)|(II30717)|(II30718);
assign g14790 = ((~II16855));
assign g21860 = (g3945&g21070);
assign g28219 = (g9316&g27573);
assign g24097 = ((~g19935));
assign g13020 = (g401&g11048);
assign II23949 = ((~g23162))|((~g13603));
assign g18595 = (g2927&g16349);
assign g14567 = (g10568&g10552);
assign g9575 = ((~g6509));
assign II14609 = ((~g8993))|((~g8678));
assign g27994 = ((~g26793));
assign II32797 = ((~g34581));
assign g30347 = (g29383)|(g18304);
assign g9416 = ((~g2429));
assign g24915 = (g23087&g20158);
assign g11653 = ((~g7980)&(~g7964));
assign g18338 = (g1710&g17873);
assign g32355 = (g29855)|(g31286);
assign g11740 = (g8769&g703);
assign g33808 = (g33109&g22161);
assign g31875 = (g31066)|(g21730);
assign g32985 = (g31963)|(g18266);
assign g26235 = ((~g8016))|((~g24766));
assign g25324 = ((~g22228));
assign g9291 = ((~g3021));
assign g26782 = ((~g9467))|((~g25203));
assign g33723 = (g14091&g33299);
assign g25238 = (g12466&g23732);
assign g34527 = (g34303&g19603);
assign g34974 = (g34870)|(g34963);
assign g10120 = ((~g1902));
assign g32893 = ((~g30937));
assign g33822 = (g33385&g20157);
assign g30321 = ((~II28572));
assign g30444 = (g29901)|(g21853);
assign II12067 = ((~g739));
assign II28185 = ((~g28803));
assign II15212 = ((~g10035))|((~g1714));
assign g31816 = ((~g29385));
assign g10139 = ((~g136));
assign g23526 = ((~g21611));
assign g27574 = (g26145)|(g24730);
assign g31486 = (g29777&g23422);
assign II24015 = (g8334&g7975&g3045);
assign g29716 = (g28199)|(g15856);
assign g25683 = (g24669)|(g18641);
assign g27300 = (g12370&g26672);
assign II31286 = (g30825&g31846&g32868&g32869);
assign g34400 = ((~g34142));
assign g34066 = (g33730&g19352);
assign g29960 = ((~g28885));
assign g34919 = ((~II33149));
assign II12618 = ((~g3338));
assign g27666 = (g26865&g23521);
assign g16871 = (g6597&g14908);
assign g30605 = (g29529)|(g29520);
assign g34990 = ((~II33270));
assign g14188 = ((~g9162)&(~g12259));
assign g26825 = ((~II25541));
assign II11892 = ((~g4408));
assign g20239 = ((~g17128));
assign g30431 = (g29875)|(g21815);
assign g19856 = ((~g13626))|((~g16278))|((~g8105));
assign g8696 = ((~g3347));
assign II16455 = ((~g11845));
assign g18592 = (g2994&g16349);
assign g17714 = ((~g14930));
assign g33690 = (g33146&g16280);
assign g21714 = (g278&g20283);
assign g29211 = ((~II27549));
assign g9780 = ((~II13360));
assign g24971 = ((~g23590));
assign g30084 = (g28534&g20700);
assign g19878 = ((~g17271));
assign II22177 = ((~g21366));
assign g10060 = ((~g6541));
assign g28749 = (g27523)|(g16764);
assign g34085 = (g33761&g9104&g18957);
assign g28812 = (g26972&g13037);
assign II24784 = ((~g24265));
assign g14599 = ((~g12207))|((~g9739));
assign g6905 = ((~II11708));
assign g27153 = (g26055&g16629);
assign g12322 = ((~II15162));
assign g32567 = ((~g31070));
assign g20180 = ((~g17533));
assign g32471 = ((~g31376));
assign g18645 = (g15100&g17271);
assign g24191 = (g319&g22722);
assign II18568 = (g13156&g11450&g11498);
assign g28658 = (g27563&g20611);
assign g20608 = ((~g15171));
assign g29180 = ((~g9569)&(~g26977));
assign II22684 = ((~g11893))|((~II22683));
assign g29328 = (g28553&g6928&g3990);
assign II13731 = ((~g4537))|((~II13729));
assign g18178 = (g758&g17328);
assign g11576 = ((~g8542));
assign g18393 = (g1917&g15171);
assign g20772 = ((~g15171));
assign g33736 = ((~II31597));
assign II14839 = ((~g9689));
assign g9552 = ((~g3654));
assign g31890 = (g31143)|(g21823);
assign g16129 = ((~II17488));
assign II14956 = ((~g9620))|((~II14955));
assign II11746 = ((~g4570));
assign g10488 = ((~g4616)&(~g7133)&(~g10336));
assign g24787 = ((~g3391))|((~g23079));
assign g13307 = ((~g1116))|((~g10695));
assign g15574 = (g4311&g13202);
assign g14548 = ((~g12208))|((~g5774));
assign g10683 = (g7289&g4438);
assign g34930 = ((~II33182));
assign II32820 = ((~g34474));
assign II29438 = ((~g30610));
assign g30417 = (g29874)|(g21801);
assign g22180 = ((~g19210));
assign g27320 = ((~II26004));
assign II14229 = ((~g979))|((~II14228));
assign g29635 = (g28910&g22432);
assign g14393 = ((~g12115)&(~g9488));
assign II32525 = ((~g34285));
assign g21661 = ((~II21222));
assign g7262 = ((~g5723));
assign g19402 = ((~g15979)&(~g13133));
assign g16966 = ((~g14291));
assign g24766 = ((~g3385)&(~g23132));
assign g7693 = ((~g4849));
assign g17156 = (g305&g13385);
assign g33608 = (g33322)|(g18537);
assign g30411 = (g29872)|(g21770);
assign II18421 = (g14447)|(g14417)|(g14395);
assign g12865 = ((~g10372));
assign g31221 = (g29494)|(g28204);
assign g17765 = ((~g6649))|((~g14556))|((~g6719))|((~g12721));
assign g16719 = ((~g3243))|((~g13700))|((~g3310))|((~g11350));
assign g17725 = (g11547&g11592&g6789&II18716);
assign g15054 = ((~g12837)&(~g13350));
assign g8956 = (g1913)|(g1932);
assign g20390 = ((~g17182)&(~g14257));
assign g33161 = ((~g32090)&(~g7806));
assign g32765 = ((~g31327));
assign g29106 = ((~g9451)&(~g28020));
assign g32614 = ((~g31542));
assign II26936 = ((~g27599));
assign g33125 = ((~g8606)&(~g32057));
assign II18101 = ((~g13416));
assign II31041 = (g31566&g31803&g32513&g32514);
assign g28621 = (g27359)|(g16518);
assign g10086 = ((~g2193));
assign g21943 = (g5240&g18997);
assign II14602 = ((~g9340));
assign g15789 = (g10819)|(g13211);
assign g29540 = ((~g28336))|((~g13464));
assign II21238 = ((~g16540));
assign g22317 = ((~g19801));
assign g31518 = (g20041&g29970);
assign g29172 = ((~g27020));
assign II22937 = ((~g12226))|((~II22936));
assign g18140 = (g559&g17533);
assign g17814 = ((~g5579))|((~g14522))|((~g5673))|((~g12563));
assign g32305 = (g31287&g20567);
assign g12135 = (g9684&g9959);
assign g7597 = ((~g952));
assign g28403 = (g27214)|(g13282);
assign g26387 = (g24813&g20231);
assign II18262 = ((~g13857));
assign g18331 = (g1682&g17873);
assign g7257 = ((~II11903));
assign II16489 = ((~g12793));
assign g21726 = ((~II21297));
assign g32216 = (g31128)|(g29615);
assign II29303 = ((~g29496))|((~II29302));
assign II16512 = ((~g12811));
assign g20056 = (g16291&g9007&g8954&g8903);
assign g12012 = ((~g9213));
assign g18800 = (g6187&g15348);
assign g33067 = (g31989)|(g22111);
assign g21831 = (g3782&g20453);
assign g10873 = (g3004&g9015);
assign g28048 = (g27362)|(g18163);
assign g9648 = ((~g2177));
assign g32167 = (g3853&g31194);
assign g23886 = ((~g21468));
assign g34108 = (g22957&g9104&g33766);
assign g33839 = ((~II31686));
assign g30024 = (g28497&g23501);
assign g9984 = (g4300)|(g4242);
assign g30489 = (g30250)|(g21985);
assign g12879 = ((~g10381));
assign g28538 = (g27294)|(g26206);
assign g27108 = (g22522)|(g25911);
assign g22868 = ((~g20453));
assign g8920 = ((~II12899));
assign g7716 = ((~g1199));
assign g34365 = (g34149&g20451);
assign g19588 = (g3849&g16853);
assign g19567 = ((~g16164));
assign g27415 = ((~g26382));
assign g30113 = ((~g29154));
assign g33493 = (g32693&II31161&II31162);
assign g25960 = (g24566)|(g24678);
assign g23879 = ((~g19210));
assign g24308 = (g4489&g22228);
assign g33429 = (g32231&g29676);
assign g11950 = ((~g9220)&(~g9166));
assign g20197 = ((~g16987));
assign g25615 = (g24803)|(g18162);
assign g16816 = ((~II18028));
assign II23917 = ((~g23975))|((~g9333));
assign g32854 = ((~g30735));
assign g27305 = (g10041&g26683);
assign g17316 = ((~II18293));
assign g28531 = (g27722&g15608);
assign II32364 = ((~g34208));
assign g18799 = (g6181&g15348);
assign g23488 = ((~g21468));
assign g27100 = ((~g26759));
assign g25113 = (g23346&g20577);
assign g23942 = ((~g21562));
assign II24334 = ((~g22976));
assign g7533 = ((~g1306));
assign g23403 = ((~II22512));
assign g34020 = (g33904)|(g18514);
assign g8515 = ((~II12631));
assign g34718 = ((~II32884));
assign g27367 = ((~g8155)&(~g26636));
assign g6845 = ((~g2126));
assign II17585 = (g14988&g11450&g11498);
assign g8481 = ((~II12618));
assign g20575 = ((~g17929));
assign g11937 = (g1936&g7362);
assign g25594 = (g24772)|(g21708);
assign g18403 = (g2028&g15373);
assign g25045 = (g17525&g23448);
assign g24393 = (g3808&g22844);
assign g25892 = ((~g24528));
assign g33400 = (g32347&g21380);
assign g16021 = (g13047)|(g10706);
assign g23006 = (g19575&g19776);
assign g9620 = ((~g6187));
assign g28775 = (g27537)|(g16806);
assign II32228 = ((~g34122));
assign II33261 = ((~g34977));
assign g29672 = ((~g28376))|((~g13672));
assign g24013 = ((~g21611));
assign g16278 = ((~g8102))|((~g8057))|((~g13664));
assign g21389 = ((~g10143)&(~g17748)&(~g12259));
assign g19792 = ((~II20204))|((~II20205));
assign g14201 = ((~II16401));
assign g34450 = (g34281)|(g18663);
assign g12905 = ((~g10408));
assign g30056 = (g29165&g12659);
assign g12856 = ((~g10430)&(~g6855));
assign g24933 = ((~g19466))|((~g23154));
assign g32036 = (g31469&g13486);
assign g25298 = ((~g23760));
assign g14336 = ((~II16498));
assign g21814 = (g3594&g20924);
assign g34912 = ((~g34883)&(~g20277)&(~g20242)&(~g21370));
assign II18782 = (g13156&g11450&g6756);
assign g29811 = ((~g28376));
assign g25852 = (g4593&g24411);
assign g21969 = (g5373&g21514);
assign g10569 = ((~g2287))|((~g7418));
assign II24555 = (g9559&g9809&g6093);
assign II22128 = ((~g19968));
assign g18380 = (g1926&g15171);
assign g22058 = (g6098&g21611);
assign g25172 = ((~g5052))|((~g23560));
assign g32851 = ((~g31327));
assign g11862 = ((~g7134)&(~g7150));
assign g33856 = (g33266&g20442);
assign II20499 = ((~g16224));
assign g24127 = ((~g19984));
assign g24354 = (g23775)|(g18823);
assign II32671 = ((~g34388));
assign g24765 = (g17699&g22498);
assign g13305 = ((~g11048));
assign g31668 = (g29924)|(g28558);
assign g31228 = (g20028&g29713);
assign g17410 = ((~g12955));
assign g16026 = (g854&g14065);
assign g15112 = (g4284&g14454);
assign g21770 = (g3251&g20785);
assign g32258 = (g31624&g30303);
assign g23406 = ((~g20330));
assign II31157 = (g32682&g32683&g32684&g32685);
assign g28235 = (g9467&g27592);
assign g9834 = ((~g2579));
assign g20531 = ((~g15907));
assign g25817 = (g24807&g21163);
assign g24433 = (g10878)|(g22400);
assign g24248 = (g22710)|(g18286);
assign g9621 = ((~g6423));
assign g16726 = ((~g14454));
assign g8278 = ((~g3096));
assign g34803 = (g34758)|(g18590);
assign g28628 = (g27370)|(g16531);
assign II12013 = ((~g590));
assign II14222 = ((~g8286));
assign II20233 = ((~g17487));
assign g21967 = (g5456&g21514);
assign g29232 = (g28183)|(g18231);
assign g28112 = (g27352&g26162);
assign g16925 = ((~g3574))|((~g13799))|((~g3668))|((~g11576));
assign g27492 = ((~g26598));
assign g24732 = ((~g23042));
assign g23809 = ((~II22966))|((~II22967));
assign g23047 = ((~g482))|((~g20000));
assign g14220 = (g8612&g11820);
assign g9338 = ((~g1870));
assign II14999 = ((~g10030));
assign g16740 = ((~g13980));
assign g10695 = ((~g8462)&(~g8407));
assign g28092 = (g27666)|(g21924);
assign g7246 = ((~g4446));
assign g11192 = ((~g8038));
assign g26788 = ((~g25349));
assign g32779 = ((~g30937));
assign g30476 = (g30229)|(g21947);
assign g18366 = (g1854&g17955);
assign g18538 = (g2759&g15277);
assign g18615 = (g3347&g17200);
assign g25959 = (g1648&g24963);
assign g25048 = ((~g542))|((~g23088));
assign g14337 = ((~g12049)&(~g9284));
assign II15587 = ((~g11985));
assign g17812 = ((~II18810));
assign g7440 = ((~g329));
assign II30995 = ((~g32449));
assign g30532 = (g30193)|(g22078);
assign g26603 = ((~g24908)&(~g24900));
assign g30458 = (g30005)|(g24330);
assign g7636 = ((~g4098));
assign g21124 = ((~g5731))|((~g17393));
assign g32180 = (g2791&g31638);
assign g25662 = (g24656)|(g21787);
assign g7115 = ((~g12));
assign g24911 = ((~II24078));
assign g8904 = (g1779)|(g1798);
assign g34478 = (g34402&g18904);
assign II16847 = ((~g6329));
assign g10947 = (g9200&g1430);
assign g21852 = (g3909&g21070);
assign g27301 = (g11992&g26679);
assign II27534 = (g28039&g24128&g24129&g24130);
assign g33428 = (g32230&g29672);
assign g23028 = ((~g20391));
assign g9901 = ((~g84));
assign g33401 = (g32349&g21381);
assign gbuf10 = (g5002);
assign II14069 = ((~g9104));
assign II21978 = ((~g19620))|((~II21976));
assign g18358 = (g1811&g17955);
assign g29856 = (g28385&g23303);
assign g31646 = ((~II29228));
assign g28436 = ((~II26929));
assign g25587 = (g21682)|(g24157);
assign g9969 = ((~g1682));
assign g21559 = (g16236&g10897);
assign g32300 = (g31274&g20544);
assign g9184 = ((~g6120));
assign II15542 = ((~g1570));
assign g22178 = ((~g19147));
assign g23280 = (g19417&g20146);
assign g22063 = (g6109&g21611);
assign g9830 = ((~II13402))|((~II13403));
assign g16186 = ((~g13555));
assign g18489 = (g2509&g15426);
assign g28138 = (g27964)|(g27968);
assign g32383 = ((~II29913));
assign g33290 = (g32149)|(g29589);
assign g16759 = (g5587&g14761);
assign g13326 = ((~g10929)&(~g10905));
assign g25873 = (g24854&g16197);
assign g34275 = ((~g34047));
assign g29868 = (g2227&g29128);
assign g24059 = ((~g21193));
assign g30414 = (g30002)|(g21794);
assign g10877 = ((~II14079));
assign II15174 = ((~g9977))|((~g2661));
assign g18339 = (g1714&g17873);
assign g10732 = (g6850&g2697&g2689);
assign g30038 = ((~g29097));
assign g9809 = ((~g6082));
assign g25605 = (g24743)|(g18116);
assign g29921 = ((~g28864));
assign g10872 = ((~g7567));
assign g11545 = ((~II14498))|((~II14499));
assign g27283 = (g25922)|(g25924);
assign II16040 = ((~g10430));
assign g26684 = (g25407&g20673);
assign g15876 = (g13512&g13223);
assign g34024 = (g33807)|(g24331);
assign g31188 = (g20028&g29653);
assign g11250 = ((~g7502));
assign g24340 = (g24016)|(g18770);
assign g6818 = ((~g976));
assign g20066 = ((~g17433));
assign g30445 = (g29772)|(g21854);
assign g10685 = ((~II13995));
assign g27685 = (g13032&g25895);
assign g15119 = (g4249&g14454);
assign II21285 = ((~g18215));
assign g26655 = ((~g25492));
assign g12874 = ((~g10383));
assign g25586 = (g21678)|(g24156);
assign II26700 = ((~g27956));
assign g14384 = ((~II16538));
assign g34260 = (g34113)|(g18680);
assign g32034 = (g14124&g31239);
assign g32426 = (g26105)|(g26131)|(g30613);
assign g30328 = ((~II28585));
assign g9962 = ((~g6519));
assign g11980 = ((~II14817))|((~II14818));
assign g32553 = ((~g31170));
assign g26721 = (g10776)|(g24444);
assign g32307 = (g31291&g23500);
assign g22514 = ((~g19699)&(~g1018));
assign g11472 = ((~g7918));
assign g32544 = ((~g30735));
assign g33585 = (g33411)|(g18456);
assign g27800 = (g17321)|(g26703);
assign g20571 = ((~g15277));
assign g19631 = (g1484&g16093);
assign g33851 = ((~g8854)&(~g33299)&(~g12259));
assign g30273 = ((~g5990)&(~g29036));
assign g15168 = ((~g13835)&(~g12909));
assign g13866 = ((~g3239))|((~g11194))|((~g3321))|((~g11519));
assign g31288 = (g2955)|(g29914);
assign g16844 = (g7212&g13000);
assign g22194 = ((~II21776));
assign g33242 = (g32123&g19931);
assign g33616 = (g33237)|(g24314);
assign g14544 = ((~II16663));
assign g27107 = (g26055&g16514);
assign II28908 = ((~g30182));
assign g14490 = ((~g9853)&(~g12598));
assign g26091 = (g1691&g25082);
assign g12116 = ((~g2051))|((~g8255));
assign g33800 = ((~II31642));
assign g18904 = ((~g16053));
assign g29145 = ((~g6549)&(~g7812)&(~g26994));
assign g29710 = (g2380&g29094);
assign g28380 = ((~g27064));
assign II32109 = ((~g33631));
assign g33714 = (g32419)|(g33450);
assign g32678 = ((~g31528));
assign g25126 = (g16839&g23523);
assign g30172 = (g28625&g21286);
assign g21511 = ((~g15483));
assign g34960 = ((~II33218));
assign g24936 = ((~g20186))|((~g20173))|((~g23379))|((~g14029));
assign g34082 = (g33709&g19554);
assign g22756 = ((~g20436));
assign g24376 = ((~g22722));
assign g33484 = (g32628&II31116&II31117);
assign II31026 = (g31194&g31800&g32492&g32493);
assign gbuf89 = (g3676);
assign g28318 = (g27233&g19770);
assign g32244 = (g31609&g30297);
assign g23445 = ((~II22564));
assign g29963 = ((~g28931));
assign g21896 = (g20084)|(g15110);
assign g22161 = (g13202&g19071);
assign g18786 = (g15156&g15345);
assign g8219 = ((~g3731));
assign g21928 = (g5170&g18997);
assign g29034 = ((~g5527)&(~g28010));
assign g31266 = (g30129&g27742);
assign II14705 = ((~g7717));
assign g27340 = (g10199&g26784);
assign g9246 = ((~g847))|((~g812));
assign g25321 = ((~g23835)&(~g14645));
assign g17739 = ((~II18728));
assign g33037 = (g32177)|(g24310);
assign g14398 = ((~II16555));
assign g12018 = ((~g9538));
assign g24132 = ((~g19890));
assign g20642 = ((~g15277));
assign II15288 = ((~g10061))|((~II15287));
assign g28625 = (g27363)|(g26324);
assign g19275 = (g7823&g16044);
assign g18257 = (g1205&g16897);
assign g17428 = ((~II18367));
assign g29683 = (g1821&g29046);
assign II22461 = ((~g21225));
assign g23362 = ((~II22467));
assign II20744 = ((~g17141));
assign g14642 = ((~g12374)&(~g9829));
assign g33743 = (g33119&g19574);
assign g11117 = ((~g8087))|((~g8186))|((~g8239));
assign g32037 = (g30566)|(g29329);
assign II20584 = ((~g16587));
assign II32274 = ((~g34195));
assign g29060 = ((~g9649))|((~g27800));
assign II16593 = ((~g10498));
assign g11829 = ((~II14653));
assign g34210 = ((~II32173));
assign g18196 = (g703&g17821);
assign g8669 = ((~g3767));
assign g22903 = ((~g20330));
assign g9451 = ((~g5873));
assign g18164 = (g699&g17433);
assign g28311 = (g9792&g27679);
assign g21944 = (g5244&g18997);
assign II18581 = ((~g14678))|((~II18579));
assign g14145 = ((~g8945)&(~g12259));
assign g17502 = ((~g14697));
assign g17753 = (g13281&g13175);
assign g29195 = ((~II27495));
assign g27826 = ((~g9501)&(~g25821));
assign II27368 = ((~g27881));
assign g29349 = (g4760&g28391);
assign g14804 = ((~g12651))|((~g12798));
assign g26656 = ((~g25495));
assign II26130 = ((~g26510));
assign g18993 = (g11224&g16172);
assign g27205 = (g25833)|(g24421);
assign g29652 = (g2667&g29157);
assign g22652 = (g18992)|(g15653);
assign g27932 = (g25944&g19369);
assign g18102 = ((~II18912));
assign g29938 = (g23552&g28889);
assign II26451 = ((~g26862));
assign g13996 = ((~g8938)&(~g8822)&(~g11173));
assign g31766 = (g30029)|(g30042);
assign g17488 = (g14361)|(g14335)|(g11954)|(II18417);
assign g22122 = (g6601&g19277);
assign g23363 = ((~II22470));
assign g22031 = (g5917&g19147);
assign g15716 = (g468&g13437);
assign II14271 = ((~g8456));
assign g28899 = ((~g27833))|((~g14612));
assign g20537 = ((~g15345));
assign g15058 = ((~g12838)&(~g13350));
assign g11954 = ((~g9538)&(~g7314));
assign g23522 = ((~g21514));
assign g11032 = (g9354&g7717);
assign g34633 = (g34481)|(g18690);
assign g23061 = ((~g20283));
assign g25116 = ((~g22369));
assign II15556 = ((~g11928));
assign II18839 = ((~g13716));
assign g22492 = ((~g19614));
assign g13462 = ((~g12449))|((~g12412))|((~g12342))|((~g12294));
assign g23909 = ((~g7028))|((~g20739));
assign g24622 = (g19856&g22866);
assign g26298 = ((~g8297)&(~g24825));
assign g14405 = ((~g12170));
assign g33863 = (g33273&g20505);
assign g8461 = (g301)|(g534);
assign g18594 = (g12858&g16349);
assign g20917 = ((~g15224));
assign g15633 = (g3841&g13584);
assign g34041 = (g33829)|(g18739);
assign g26909 = (g26543)|(g24227);
assign II28838 = ((~g29372));
assign g23529 = ((~g20558));
assign g32398 = (g31526)|(g30061);
assign g20183 = ((~g17152)&(~g14222));
assign II14186 = ((~g8442))|((~II14185));
assign g31901 = (g31516)|(g21909);
assign g18191 = (g827&g17821);
assign g30316 = (g29199&g7097&g6682);
assign II14351 = ((~g8890))|((~II14350));
assign g24919 = (g21606)|(g22143);
assign g28535 = (g11981&g27088);
assign g21431 = ((~g18065));
assign g18462 = (g2361&g15224);
assign II14830 = ((~g10141));
assign g12184 = ((~II15036));
assign II32518 = ((~g34422))|((~II32516));
assign II14518 = ((~g661))|((~II14516));
assign g23528 = ((~g18833));
assign g30558 = (g30258)|(g22129);
assign g12208 = ((~g10096)&(~g5759));
assign g26102 = (g1825&g25099);
assign g19544 = ((~g16349));
assign g32891 = ((~g30825));
assign g28020 = (g23032&g26241&g26424&g25542);
assign g11938 = ((~g8259))|((~g2208));
assign g11953 = ((~g8195))|((~g8241));
assign g9683 = ((~g6140));
assign II14855 = ((~g5142))|((~II14853));
assign II31523 = ((~g33187));
assign g33523 = (g32909&II31311&II31312);
assign g32295 = (g27931&g31376);
assign II22761 = ((~g11939))|((~II22760));
assign g10222 = ((~g4492));
assign g13383 = (g4765&g11797);
assign g27093 = ((~g26712)&(~g26749));
assign g31316 = (g29609)|(g29624);
assign g10081 = ((~g2279));
assign g34073 = (g8948&g33823);
assign g31498 = ((~g9030)&(~g29540));
assign g32187 = (g30672&g25287);
assign g8227 = ((~g3770))|((~g3774));
assign g23659 = ((~g9434))|((~g20854));
assign g11006 = ((~g7686)&(~g7836));
assign II31642 = ((~g33204));
assign g12344 = ((~g10093))|((~g7041))|((~g10130));
assign g17767 = (g6772&g11592&g6789&II18765);
assign g17513 = ((~g3247))|((~g13765))|((~g3325))|((~g8481));
assign g31940 = (g943&g30735);
assign g20236 = ((~g16875))|((~g14014))|((~g16625))|((~g16604));
assign g9374 = ((~g5188));
assign g24274 = (g23187)|(g18631);
assign II18151 = ((~g13144));
assign g20212 = ((~g17194));
assign g13484 = ((~g10981));
assign g34216 = (g33778&g22689);
assign g23577 = (g19444&g13033);
assign gbuf82 = (g3632);
assign II15042 = ((~g9752))|((~II15041));
assign g6961 = ((~II11734));
assign g21058 = ((~g15426));
assign g24096 = ((~g19890));
assign g10527 = ((~II13892));
assign II14854 = ((~g9433))|((~II14853));
assign g34439 = (g34344)|(g18181);
assign g22593 = ((~g19801));
assign g13505 = ((~g10981));
assign g13963 = ((~g11715))|((~g11584));
assign g20627 = ((~g17433));
assign g21810 = (g3578&g20924);
assign g9295 = ((~II13066))|((~II13067));
assign g28208 = (g27025)|(g27028);
assign g17181 = (g1945&g13014);
assign g11163 = (g6727&g10224);
assign g15036 = ((~g12780))|((~g12581));
assign g15067 = ((~g12842)&(~g13394));
assign g27244 = (g24652)|(g25995);
assign g16963 = ((~II18117));
assign g22860 = ((~g20000));
assign g29882 = (g2361&g29151);
assign g32821 = ((~g31021));
assign g33990 = (g33882)|(g18399);
assign g28415 = (g27250&g19963);
assign g16855 = (g4392&g13107);
assign g15882 = (g3554&g13986);
assign g18154 = (g622&g17533);
assign II31232 = (g32791&g32792&g32793&g32794);
assign g21178 = ((~g17955));
assign g33703 = (g32410)|(g33434);
assign II12861 = ((~g4372));
assign g13271 = ((~II15834));
assign g30916 = (g13853)|(g29799);
assign II24383 = ((~g23721))|((~g14347));
assign g24298 = (g4392&g22550);
assign g34583 = ((~II32665));
assign g30926 = (g29903&g21163);
assign g33079 = ((~II30641));
assign II17557 = ((~g14510));
assign g23756 = ((~g9621))|((~g21206));
assign II14745 = ((~g10029));
assign g32996 = (g32256)|(g18377);
assign g28207 = ((~g12546))|((~g26131))|((~g27977));
assign g22449 = ((~g19597));
assign g16124 = ((~g13555));
assign g11697 = ((~g8080)&(~g3857));
assign II32352 = ((~g34169));
assign g11491 = ((~g9982))|((~g4000));
assign g10152 = ((~g2122));
assign g30161 = (g28614&g21275);
assign g18112 = (g182&g17015);
assign g25005 = ((~g6811)&(~g23324));
assign g33175 = ((~g32099)&(~g7828));
assign g33931 = ((~II31807));
assign II32150 = ((~g33923));
assign g21741 = (g15086&g20330);
assign II14532 = ((~g8873))|((~II14530));
assign g26837 = ((~g24869));
assign g7593 = ((~II12061));
assign g24661 = ((~g23210))|((~g23195))|((~g22984));
assign II20487 = ((~g16696))|((~II20486));
assign g23913 = ((~g19147));
assign g25017 = ((~g23699));
assign g20588 = ((~g18008));
assign g10384 = ((~II13802));
assign g28682 = (g27430)|(g16635);
assign g33758 = (g33133&g20269);
assign g32869 = ((~g30735));
assign g21304 = ((~g17367));
assign g16164 = ((~II17507));
assign g19440 = ((~g15915));
assign g19503 = ((~g16349));
assign g20328 = ((~g15867));
assign g29250 = (g28695)|(g18460);
assign II26430 = ((~g26856));
assign g11820 = ((~II14644));
assign g17120 = ((~g14262));
assign g8891 = ((~g582));
assign g24706 = (g15910&g22996);
assign g11931 = ((~II14749));
assign g34180 = (g33716&g24373);
assign II31161 = (g30614&g31824&g32687&g32688);
assign g33631 = ((~II31459));
assign g25625 = (g24553)|(g18226);
assign g7018 = ((~g5297));
assign g29941 = ((~g28900));
assign g19501 = (g16986)|(g14168);
assign g13210 = ((~g7479))|((~g10521));
assign g31566 = (g19050&g29814);
assign g18556 = (g2823&g15277);
assign g28496 = ((~g3179)&(~g27602));
assign g34945 = ((~g34933));
assign g13258 = ((~II15821));
assign g28566 = (g27316)|(g26254);
assign g12839 = ((~g10350));
assign g15086 = ((~g13144)&(~g12859));
assign II16579 = ((~g10981));
assign g23724 = (g14767&g21123);
assign g19957 = ((~g16540));
assign g17747 = (g6772&g11592&g11640&II18740);
assign g24384 = ((~g22885));
assign g7461 = ((~g2567));
assign g29805 = (g28357&g23270);
assign g33005 = (g32260)|(g18432);
assign g25024 = ((~g22472));
assign g21296 = (g7879&g16072);
assign g33555 = (g33355)|(g18357);
assign g11224 = ((~II14290))|((~II14291));
assign g29342 = ((~g28188));
assign g16325 = ((~g13223));
assign g20051 = (g15936)|(g13306);
assign g28470 = ((~g8021)&(~g27617));
assign g27537 = (g26549&g17742);
assign g8565 = ((~g3802));
assign g29351 = (g4771&g28406);
assign g32901 = ((~g31327));
assign g34605 = (g34566)|(g15077);
assign g12136 = ((~II14992))|((~II14993));
assign g10841 = (g8509&g8567);
assign g22867 = ((~g20391));
assign g33660 = ((~II31494));
assign g9989 = ((~g5077));
assign g34845 = ((~g34773));
assign II22240 = ((~g20086));
assign g16093 = ((~II17461))|((~II17462));
assign g28453 = (g27582&g10233);
assign g12604 = ((~g5517)&(~g9239));
assign g30110 = (g28564&g20916);
assign II21757 = ((~g21308));
assign g23259 = ((~g21070));
assign g24185 = ((~II23399));
assign g25733 = (g25108)|(g18778);
assign g25196 = ((~g22763));
assign g26785 = (g10776)|(g24468);
assign g9574 = ((~g6462));
assign g15571 = ((~g13211));
assign g20082 = (g16026)|(g13321);
assign g17225 = ((~g8612))|((~g14367));
assign g20102 = ((~g17533));
assign g19600 = ((~g16164));
assign g31781 = (g30058)|(g30069);
assign g34204 = (g33832)|(g33833);
assign g13202 = ((~g8347)&(~g10511));
assign g22520 = ((~g19801));
assign II30746 = (g32047)|(g31985)|(g31991)|(g32309);
assign g34616 = (g34519)|(g18577);
assign g27474 = (g8038&g26314&g518&g504);
assign g7474 = ((~II11980));
assign g25244 = ((~g23802));
assign g10503 = ((~g8879));
assign g23856 = (g4116&g19483);
assign g14754 = ((~g12821)&(~g2988));
assign II31212 = (g32761&g32762&g32763&g32764);
assign g19362 = ((~g16072));
assign g33268 = (g32116)|(g29538);
assign g26993 = ((~g5360)&(~g25805));
assign II12876 = ((~g4200))|((~g4180));
assign g14203 = ((~g12381));
assign g21707 = (g191&g20283);
assign g29554 = (g28997&g22472);
assign g29706 = (g28198)|(g27208);
assign II31843 = (g33470)|(g33471)|(g33472)|(g33473);
assign g17268 = (g9220)|(g14387);
assign g32960 = ((~g31327));
assign g24652 = ((~g22712))|((~g22940))|((~g22757));
assign g23545 = ((~g21562));
assign g30251 = (g28745&g23940);
assign g19776 = ((~g17015));
assign g18640 = (g3835&g17096);
assign g32152 = (g31631&g29998);
assign II17461 = ((~g13378))|((~II17460));
assign g34239 = (g32845)|(g33957);
assign g17815 = ((~g14348));
assign g9060 = ((~g3355));
assign g15136 = ((~g13680)&(~g12885));
assign II14228 = ((~g979))|((~g8055));
assign g21364 = ((~g15787))|((~g15781))|((~g15753))|((~g13131));
assign g29239 = (g28427)|(g18297);
assign g17588 = ((~g14782));
assign g24996 = ((~g22763));
assign g25070 = ((~g23590));
assign II22866 = ((~g21228))|((~II22864));
assign g13507 = (g7023&g12198);
assign g34283 = (g26839)|(g34215);
assign g23824 = ((~g21271));
assign g20707 = ((~g18008));
assign g24802 = ((~II23970))|((~II23971));
assign g32760 = ((~g30735));
assign g14596 = ((~g12196))|((~g9775))|((~g12124))|((~g9663));
assign g21838 = (g3747&g20453);
assign g32635 = ((~g31542));
assign g15907 = ((~g14833))|((~g9417))|((~g12487));
assign g18138 = (g546&g17249);
assign g25213 = ((~g23293));
assign g33905 = (g33089&g15574);
assign g29188 = (g27163&g12762);
assign g23762 = ((~II22900))|((~II22901));
assign g32613 = ((~g30673));
assign g18572 = (g2864&g16349);
assign g10794 = ((~g8470));
assign g29664 = (g2273&g29060);
assign g15098 = ((~g13191)&(~g6927));
assign g27879 = ((~g9523)&(~g25856));
assign g33929 = ((~II31803));
assign g8854 = ((~g613));
assign g23480 = ((~II22601));
assign g21395 = ((~g17873));
assign II28014 = ((~g28158));
assign g23613 = ((~II22748));
assign g29318 = ((~g29029));
assign g25268 = ((~g21124))|((~g23692));
assign II31021 = (g31070&g31799&g32485&g32486);
assign g13003 = ((~II15609));
assign g32279 = (g31220)|(g31224);
assign g11869 = ((~g7649)&(~g7534)&(~g7581));
assign g32819 = ((~g30825));
assign g32812 = ((~g30825));
assign g16581 = ((~g13756)&(~g8086));
assign g34771 = (g34693&g20147);
assign g21277 = ((~g9417)&(~g9340)&(~g17467));
assign g21766 = (g3235&g20785);
assign g19336 = (g17769)|(g14831);
assign g11114 = (g5689&g10160);
assign g23779 = (g1105&g19355);
assign g8037 = ((~g405));
assign g16307 = ((~II17633));
assign g14044 = (g10776)|(g8703);
assign g16716 = ((~g13948));
assign g7268 = ((~g1636));
assign g31830 = ((~g29385));
assign g21981 = (g5543&g19074);
assign g19569 = ((~g16349));
assign g26395 = (g22547&g25561);
assign g30434 = (g30024)|(g21818);
assign g9158 = ((~g513));
assign g23615 = (g20109)|(g20131);
assign g29567 = (g2357&g28593);
assign g29773 = (g28203&g10233);
assign g18593 = (g2999&g16349);
assign g24404 = ((~g22908));
assign g25910 = (g25565)|(g22142);
assign g25169 = ((~g22763));
assign g18131 = (g482&g16971);
assign g28330 = (g27238&g19786);
assign g29166 = (g27653)|(g17153);
assign g27708 = ((~II26334));
assign g18413 = (g2089&g15373);
assign g16968 = ((~g14238));
assign g8540 = ((~g3408));
assign g31949 = (g1287&g30825);
assign g12909 = ((~g10412));
assign II17901 = ((~g3976));
assign g13937 = ((~g8883)&(~g4785)&(~g11155));
assign g18775 = (g7028&g15615);
assign g28547 = (g6821&g27091);
assign g18703 = (g4776&g16782);
assign g23990 = (g19610&g10951);
assign II28567 = (g29204)|(g29205)|(g29206)|(g29207);
assign g17640 = ((~g5264))|((~g14399))|((~g5335))|((~g12497));
assign g25188 = ((~g23909));
assign g7191 = ((~g6398));
assign g28257 = (g27179&g19686);
assign g14219 = ((~g12381));
assign g14581 = (g12587&g12428&g12357&II16695);
assign g17474 = ((~g14547))|((~g14521));
assign II17661 = ((~g13329));
assign g9716 = ((~g5057));
assign g13983 = ((~g11658))|((~g8906));
assign g20079 = ((~g17328));
assign g28664 = (g27408)|(g16613);
assign g20675 = ((~g14377))|((~g17246))|((~g9442));
assign g34109 = (g33918&g23708);
assign g12812 = (g518&g9158);
assign g14296 = (g2638&g11897);
assign g11046 = (g9889&g6120);
assign g24640 = (g6509&g23733);
assign II23951 = ((~g13603))|((~II23949));
assign g25043 = (g20733&g23447);
assign g32757 = ((~g30937));
assign g28328 = (g27127)|(g15812);
assign g29108 = ((~g6219)&(~g26977));
assign II13906 = ((~g7620));
assign II21766 = ((~g19620));
assign II15030 = ((~g10073));
assign g24978 = ((~g22342));
assign g23865 = ((~g21308));
assign g14032 = ((~g11048));
assign g34743 = (g8951&g34703);
assign II32909 = ((~g34712));
assign g16511 = ((~g14130));
assign g20569 = ((~g15277));
assign g14668 = ((~g12450));
assign g12449 = ((~g7004))|((~g5297))|((~g5352));
assign g35002 = ((~II33300));
assign g30272 = (g28814&g23982);
assign g10348 = ((~II13762));
assign g10177 = ((~g1834));
assign g28587 = (g27487&g20498);
assign g23877 = ((~g19147));
assign g31924 = (g31486)|(g22049);
assign g26389 = (g19949&g25553);
assign g28260 = (g27703&g26518);
assign gbuf108 = (g4194);
assign g20131 = (g15170&g14309);
assign g12086 = ((~g9654));
assign g27117 = (g26055&g16528);
assign g14256 = (g2079&g11872);
assign g23194 = (g19564)|(g19578);
assign g32485 = ((~g31376));
assign g18143 = (g586&g17533);
assign g33257 = (g32108)|(g29519);
assign II31166 = (g30673&g31825&g32694&g32695);
assign g28683 = (g27876&g20649);
assign g21848 = (g3913&g21070);
assign gbuf72 = (g3310);
assign g24683 = ((~g23112));
assign g23424 = (g7345&g21556);
assign g29599 = (g1710&g29018);
assign g23349 = (g13662&g20182);
assign g31987 = (g31767&g22198);
assign II26503 = ((~g26811));
assign g24990 = ((~g8898)&(~g23324));
assign g9595 = ((~g2351))|((~g2319));
assign g12465 = ((~g7192));
assign II14816 = ((~g9962))|((~g6513));
assign g20320 = ((~g17015));
assign g24216 = (g23416)|(g18197);
assign g13663 = ((~g10971));
assign g13795 = ((~g11216))|((~g401));
assign g32787 = ((~g30937));
assign g33058 = (g31976)|(g22020);
assign II31604 = ((~g33176));
assign g33844 = (g33257&g20327);
assign g24231 = (g22589)|(g18201);
assign g32259 = (g31185)|(g29709);
assign g23889 = ((~g20682));
assign g27659 = ((~g3706)&(~g26657));
assign g13885 = ((~g10862));
assign g34564 = (g34373&g17466);
assign g23646 = (g16959&g20737);
assign g18879 = (g17365)|(g14423);
assign g19709 = ((~g16987));
assign g19954 = ((~g16540));
assign g29213 = ((~II27555));
assign g8091 = ((~g1579));
assign g18400 = (g2012&g15373);
assign g11992 = ((~g7275))|((~g1772));
assign g30731 = (g11374&g29361);
assign II28548 = ((~g28147));
assign g7972 = ((~g1046));
assign g23686 = ((~g2767)&(~g21066));
assign g17190 = ((~g723)&(~g14279));
assign g26889 = (g26689)|(g24195);
assign II16821 = ((~g5983));
assign g19586 = ((~g16349));
assign g34345 = ((~II32352));
assign g34469 = ((~II32517))|((~II32518));
assign g14639 = ((~II16747));
assign g9095 = ((~g3368));
assign II31550 = ((~g33204));
assign g16232 = ((~g13516)&(~g4950));
assign g8418 = ((~g2619));
assign g20558 = ((~II20650));
assign g17328 = ((~II18313));
assign II11980 = ((~g66));
assign g18809 = (g7074&g15656);
assign g13102 = ((~g7523))|((~g10759));
assign g8883 = ((~g4709));
assign g20553 = ((~g17929));
assign g18981 = (g11206&g16158);
assign g19784 = (g2775&g15877);
assign g28595 = (g27335)|(g26290);
assign II23688 = ((~g23244));
assign g24167 = ((~II23345));
assign g8362 = ((~g194));
assign g18236 = (g15065&g16326);
assign g10194 = ((~g6741));
assign g21349 = ((~g15758));
assign g12169 = ((~g9804))|((~g5448));
assign g32951 = ((~g31021));
assign g16516 = (g5228&g14627);
assign g29269 = (g28249)|(g18634);
assign g34099 = (g33684)|(g33689);
assign g13945 = ((~g691))|((~g11740));
assign g7227 = ((~g4584))|((~g4593));
assign g20006 = ((~g17328));
assign g14908 = ((~g7812))|((~g10491));
assign g29526 = (g28938&g22384);
assign g30356 = (g30096)|(g18365);
assign g21984 = (g5563&g19074);
assign g17087 = ((~g14321));
assign g30076 = ((~g29085));
assign g24759 = ((~g23003));
assign g18730 = (g4950&g16861);
assign g11306 = ((~g3412)&(~g8647));
assign g24953 = ((~g10262)&(~g23978)&(~g12259));
assign g28697 = (g27581&g20669);
assign g17584 = ((~g14773));
assign g29898 = ((~g6895)&(~g28458));
assign II31466 = ((~g33318));
assign g32363 = ((~II29891));
assign g32541 = ((~g30673));
assign g34505 = ((~g34409));
assign g23385 = ((~II22488));
assign g21777 = (g3380&g20391);
assign g18487 = (g2441&g15426);
assign g31151 = (g10037&g30065);
assign g13109 = ((~g6279))|((~g12173))|((~g6369))|((~g10003));
assign g24869 = ((~II24041));
assign g26963 = (g26306)|(g24308);
assign g11155 = ((~g4776))|((~g7892))|((~g9030));
assign g34127 = (g33657)|(g32438);
assign g15105 = (g4235&g14454);
assign g18521 = (g2667&g15509);
assign g27258 = (g25905)|(g15749);
assign g32217 = (g31129)|(g29616);
assign g7791 = ((~II12199));
assign g25290 = (g5022&g22173&II24482);
assign II18752 = ((~g6358));
assign g29588 = (g2311&g28942);
assign g15819 = (g3251&g14101);
assign II17668 = ((~g13279));
assign g11960 = (g2495&g7424);
assign g13954 = ((~g8663)&(~g11276));
assign g32666 = ((~g31376));
assign g25337 = ((~g22342))|((~g1648))|((~g8187));
assign g22873 = (g19854&g19683);
assign g32265 = (g2799&g30567);
assign g18292 = (g1472&g16449);
assign g12910 = ((~g11002))|((~g10601));
assign g33390 = (g32276)|(g29968);
assign g10341 = ((~g6227)&(~g6219));
assign g25751 = (g25061)|(g22098);
assign g8788 = ((~II12776));
assign g10624 = (g8387&g3072);
assign g27556 = (g26097)|(g24687);
assign g16237 = ((~g8088)&(~g13574));
assign II32470 = ((~g34247));
assign g12080 = ((~g1917))|((~g8201));
assign g18094 = ((~II18888));
assign g17952 = ((~II18858));
assign II25680 = ((~g25641));
assign g33316 = (g29685)|(g32178);
assign g25034 = ((~g23695));
assign g24814 = ((~g20011))|((~g23167));
assign g13605 = ((~II16040));
assign g31933 = (g939&g30735);
assign g8681 = ((~g763));
assign g34712 = ((~II32868));
assign g11363 = ((~g8626)&(~g8751));
assign g23217 = (g19588)|(g16023);
assign g33526 = (g32932&II31326&II31327);
assign g18122 = (g15052&g17015);
assign II13499 = ((~g232))|((~II13497));
assign g31852 = ((~g29385));
assign g27092 = ((~g26737));
assign g28818 = (g27549)|(g13998);
assign g21956 = (g5360&g21514);
assign g34326 = ((~g34091));
assign g30366 = (g30122)|(g18417);
assign g20617 = ((~g15277));
assign g32371 = (g29883)|(g31313);
assign g14602 = ((~g10099)&(~g12790));
assign g32782 = ((~g30735));
assign g13861 = ((~g1459))|((~g10671));
assign g33636 = ((~II31463));
assign g18129 = (g518&g16971);
assign g23323 = ((~g20283));
assign g34071 = (g8854&g33799);
assign g27009 = ((~g25911));
assign g26629 = (g14173&g24418);
assign g27377 = ((~g10685))|((~g25930));
assign g16639 = (g6291&g14974);
assign gbuf30 = (g5630);
assign g9751 = ((~g1710));
assign g30103 = (g28477)|(g16731);
assign II17575 = (g13156&g11450&g6756);
assign g26312 = (g2704&g25264);
assign g20381 = ((~g17955));
assign g15848 = (g3259&g13892);
assign g27347 = (g26400&g17390);
assign g13240 = ((~g1046))|((~g10521));
assign g18891 = ((~g16053));
assign g30611 = (g13671)|(g29743);
assign g18548 = (g2807&g15277);
assign II25689 = ((~g25688));
assign g21662 = ((~g16540));
assign g9252 = ((~g4304));
assign g32724 = ((~g30735));
assign g26183 = ((~g23079)&(~g24766));
assign g27212 = (g25997&g16717);
assign g27597 = ((~g26745));
assign g12920 = (g1227&g10960);
assign g22942 = (g9104&g20219);
assign g16806 = (g6247&g14971);
assign g27126 = (g24378)|(g25787);
assign g33507 = (g32795&II31231&II31232);
assign II28301 = ((~g29042));
assign g10581 = ((~g9529));
assign g30286 = (g28191)|(g28186);
assign g28850 = (g27557)|(g16869);
assign II13067 = ((~g4304))|((~II13065));
assign g25137 = ((~g22432));
assign g32730 = ((~g31327));
assign g33692 = (g32400)|(g33428);
assign g22133 = (g6649&g19277);
assign g32497 = ((~g30673));
assign g28722 = (g27955&g20738);
assign II18713 = (g13156&g6767&g6756);
assign II24434 = ((~g22763));
assign g32234 = (g31601&g30292);
assign II18006 = ((~g13638));
assign g23307 = ((~g20924));
assign g33682 = ((~II31515));
assign g18119 = (g475&g17015);
assign g34602 = (g34489)|(g18269);
assign g26846 = (g37&g24524);
assign g25835 = (g25367)|(g23855);
assign g32885 = ((~g31021));
assign g30147 = ((~g28768)&(~g14567));
assign II11877 = ((~g4388))|((~g4430));
assign g30152 = (g28609&g23767);
assign g29293 = (g28570)|(g18777);
assign g7157 = ((~g5706));
assign g32598 = ((~g30614));
assign g14413 = ((~g11914)&(~g9638));
assign g27487 = (g25990)|(g24629);
assign g20190 = ((~g16971));
assign II12764 = ((~g4194));
assign g22219 = (g19953&g20887);
assign g25181 = (g23405&g20696);
assign g14359 = ((~II16515));
assign II23357 = ((~g23359));
assign g30528 = (g30202)|(g22074);
assign g33028 = (g32325)|(g21797);
assign g16280 = ((~g13330));
assign g21883 = (g4141&g19801);
assign g22012 = (g5752&g21562);
assign g26946 = (g26389)|(g24284);
assign g22103 = (g15164&g18833);
assign g23796 = (g21462)|(g21433)|(II22958);
assign g26930 = (g26799)|(g18544);
assign g23793 = ((~g19074));
assign g21733 = (g3034&g20330);
assign g16773 = ((~g14021));
assign g31849 = ((~g29385));
assign g31145 = (g9970&g30052);
assign g32512 = ((~g31566));
assign II20369 = ((~g17690));
assign g20671 = ((~g15509));
assign g30006 = (g29032&g9259);
assign g29498 = ((~II27784));
assign g26917 = (g26122)|(g18233);
assign g15740 = ((~g13342));
assign g22214 = ((~g19210));
assign g23261 = (g19660)|(g16125);
assign g28643 = (g27386)|(g16592);
assign g33989 = (g33870)|(g18398);
assign g21286 = ((~g15509));
assign g25975 = (g9434&g24999);
assign g28578 = (g27327)|(g26273);
assign g21821 = (g3723&g20453);
assign g28755 = ((~g27742))|((~g7268))|((~g1592));
assign g18329 = (g1612&g17873);
assign g24225 = (g246&g22594);
assign g10699 = ((~g8526)&(~g1514));
assign g25546 = ((~g22550));
assign g32153 = (g31646&g29999);
assign g25952 = ((~g1542)&(~g24609));
assign g18600 = (g3111&g16987);
assign g9598 = ((~g2571));
assign II22819 = ((~g19862));
assign g22209 = (g19907&g20751);
assign II14884 = ((~g9500))|((~II14883));
assign g10999 = (g7880&g1472);
assign g21407 = ((~g15171));
assign g22006 = (g5767&g21562);
assign g24630 = (g23255&g14149);
assign g23203 = ((~g20073));
assign g21884 = (g4104&g19801);
assign II12263 = ((~g1448))|((~II12261));
assign g24887 = (g3712&g23239&II24054);
assign g27243 = (g25884)|(g24475);
assign g8163 = ((~g3419))|((~g3423));
assign g18757 = (g5352&g15595);
assign g26379 = (g19904&g25546);
assign g34953 = (g34935&g19957);
assign II13762 = ((~g6755));
assign g22001 = (g5731&g21562);
assign g28418 = (g27220)|(g15882);
assign g34701 = (g34536&g20179);
assign g26230 = (g1768&g25385);
assign g31826 = ((~g29385));
assign g15224 = ((~II17101));
assign g25777 = ((~g25482)&(~g25456));
assign g31895 = (g31505)|(g24296);
assign g24794 = (g11414&g23138);
assign g31747 = ((~II29296))|((~II29297));
assign g31970 = ((~g9024)&(~g30583));
assign II33119 = ((~g34852));
assign g33042 = (g32193)|(g24324);
assign g28087 = (g27255)|(g18720);
assign g26130 = (g24890&g19772);
assign g25747 = (g25130)|(g18795);
assign g13267 = ((~II15831));
assign g7752 = ((~g1542));
assign g9742 = ((~g6144));
assign g14874 = (g1099&g10909);
assign g21561 = ((~g15595));
assign II29985 = (g29385)|(g31376)|(g30735)|(g30825);
assign g25081 = ((~g22342));
assign g13314 = ((~g10893));
assign II22886 = ((~g18926));
assign II22753 = ((~g11937))|((~g21434));
assign g22540 = ((~g19720)&(~g1373));
assign g33914 = (g33305)|(g33311);
assign g24465 = (g3827&g23139);
assign g11388 = ((~II14395));
assign g32731 = ((~g31376));
assign g16047 = (g13322&g1500&g10699);
assign g25640 = ((~II24781));
assign g18322 = (g1608&g17873);
assign g6799 = ((~g199));
assign g26892 = (g26719)|(g24198);
assign g14858 = ((~g7766))|((~g12515));
assign g11431 = ((~g7618));
assign g32533 = ((~g30614));
assign g7487 = ((~g1259));
assign g33086 = (g32390&g18887);
assign g7544 = ((~g918));
assign g23607 = ((~g21611));
assign g23750 = (g20174)|(g16840);
assign g27977 = ((~g26105));
assign g16287 = ((~g13622)&(~g11144));
assign g29504 = (g28143)|(g25875);
assign g25482 = (g5752&g23816&II24597);
assign II27558 = ((~g28155));
assign g16052 = (g13060)|(g10724);
assign g10727 = ((~II14016));
assign g32703 = ((~g30825));
assign g33540 = (g33099)|(g18207);
assign g28119 = ((~g27008));
assign g18277 = (g1312&g16136);
assign g19756 = (g9899&g17154);
assign g33518 = (g32874&II31286&II31287);
assign g14755 = ((~g12593))|((~g12772));
assign g23339 = ((~g21070));
assign g32684 = ((~g30673));
assign g33812 = (g23088&g33187&g9104);
assign g29364 = (g27400&g28321);
assign g18226 = (g15064&g16129);
assign g22989 = ((~g20453));
assign g28451 = (g27283&g20090);
assign g18663 = (g4311&g17367);
assign g8052 = ((~g1211));
assign g16877 = ((~II18071));
assign g29251 = (g28679)|(g18464);
assign g28703 = (g27925&g20680);
assign g15156 = ((~g13782)&(~g7050));
assign g13045 = ((~g11941));
assign g28352 = (g10014&g27705);
assign gbuf15 = (g5313);
assign g10287 = ((~II13715));
assign g28744 = (g27518)|(g16759);
assign II17198 = ((~g13809));
assign g17092 = ((~g14011));
assign g34471 = ((~g34423));
assign g33559 = (g33073)|(g18368);
assign g30311 = (g28265)|(g27265);
assign g12225 = ((~g8324))|((~g2453));
assign II18778 = ((~g6704));
assign g19573 = ((~g16877));
assign g31961 = (g31751&g22154);
assign g29043 = ((~II27391));
assign g34390 = (g34172&g21069);
assign g13761 = (g490)|(g12527);
assign g32958 = ((~g31710));
assign g22759 = ((~g19857));
assign II28199 = ((~g28803));
assign g6754 = ((~II11617));
assign g19127 = ((~II19775));
assign g33365 = (g32267&g20994);
assign g34963 = (g34946&g23041);
assign g10229 = ((~g6736));
assign g34910 = ((~g34864));
assign II25511 = ((~g25073));
assign g24118 = ((~g19890));
assign g28153 = (g26424&g22763&g27031);
assign g33465 = (g32491&II31021&II31022);
assign g19676 = ((~g17062));
assign g24108 = ((~g20998));
assign g26817 = ((~g25242));
assign g27762 = (g22472&g25226&g26424&g26218);
assign g20700 = ((~g17873));
assign II31569 = ((~g33197));
assign g34882 = (g34876)|(g18659);
assign g19358 = ((~g15723))|((~g1399));
assign g20594 = ((~g15277));
assign gbuf63 = (g6668);
assign g19684 = (g2735&g17297);
assign g30001 = (g28490&g23486);
assign g19666 = ((~g17188));
assign g13059 = (g6900&g11303);
assign g29321 = (g29033&g22148);
assign g34300 = (g26864)|(g34230);
assign II24710 = (g24071&g24072&g24073&g24074);
assign g32235 = (g31151)|(g29662);
assign II27546 = ((~g29041));
assign g26171 = (g25357&g6856&g11709&g11686);
assign g22721 = ((~II22028));
assign g24429 = ((~g22722));
assign II17723 = ((~g13177));
assign g18700 = (g15132&g16816);
assign g9092 = ((~g3004))|((~g3050));
assign g30542 = (g29337)|(g22088);
assign g23843 = ((~g19147));
assign g28483 = ((~g8080)&(~g27635));
assign g33583 = (g33074)|(g18448);
assign II33106 = ((~g34855));
assign II15942 = ((~g12381));
assign g11621 = ((~g3512)&(~g7985));
assign g7836 = ((~g4653))|((~g4688));
assign II15073 = ((~g10109));
assign II23339 = ((~g23232));
assign g22024 = (g5897&g19147);
assign g10181 = ((~g2551));
assign g16625 = ((~g3203))|((~g13700))|((~g3274))|((~g11519));
assign g19672 = ((~g16931));
assign g30486 = (g30177)|(g21982);
assign g26544 = (g7446&g24357);
assign g13631 = ((~g8068)&(~g10733));
assign g12318 = ((~g10172)&(~g6451));
assign g18318 = (g1604&g17873);
assign g14420 = ((~g12153)&(~g9490));
assign g34872 = (g34827&g19954);
assign g9298 = ((~g5080));
assign II16775 = ((~g12183));
assign g20534 = ((~g17183));
assign g34447 = (g34363)|(g18552);
assign g10308 = ((~g4459));
assign g27057 = (g7791&g6219&g6227&g26261);
assign g29583 = (g28182)|(g27099);
assign g9488 = ((~g1878));
assign g18416 = (g2112&g15373);
assign g32877 = ((~g30825));
assign II24603 = (g9892&g9467&g6439);
assign g27589 = (g26177)|(g24763);
assign gbuf5 = (g4446);
assign g20751 = (g16260&g4836);
assign II29207 = ((~g30293));
assign g6841 = ((~g2145));
assign g29618 = (g28870&g22384);
assign II17923 = ((~g13378))|((~g1478));
assign II16535 = ((~g11235));
assign g26247 = ((~g7995)&(~g24732));
assign II24385 = ((~g14347))|((~II24383));
assign g17292 = (g1075&g13093);
assign g14918 = ((~g12646))|((~g12772));
assign g11910 = ((~g10185));
assign g18498 = (g2547&g15426);
assign g7803 = ((~II12204))|((~II12205));
assign g21925 = (g5073&g21468);
assign g30230 = (g28717&g23906);
assign g19267 = (g17752)|(g17768);
assign g15735 = ((~g5547))|((~g14425))|((~g5659))|((~g9864));
assign g34301 = (g34064&g19415);
assign g24879 = (g21465)|(g24009);
assign g9776 = ((~g5073));
assign II31545 = ((~g33219));
assign g7400 = ((~g911));
assign g14830 = ((~g6605))|((~g12211))|((~g6723))|((~g12721));
assign g14828 = ((~II16875));
assign g30459 = (g29314)|(g21926);
assign g22957 = ((~II22143));
assign g27260 = (g26766&g26737);
assign gbuf116 = (g4216);
assign g20775 = ((~g18008));
assign g27013 = ((~II25743));
assign g29754 = (g28215)|(g28218);
assign II15365 = ((~g2675))|((~II15363));
assign g27141 = ((~II25846))|((~II25847));
assign g33099 = (g32395&g18944);
assign g15580 = ((~g13242));
assign g27004 = ((~g26131));
assign g24544 = ((~g22666))|((~g22661))|((~g22651));
assign g30509 = (g30210)|(g22030);
assign g29067 = ((~II27401));
assign g23201 = (g14027&g20040);
assign g25300 = ((~g22369))|((~g12018));
assign g9316 = ((~g5742));
assign II18078 = ((~g13350));
assign g28606 = ((~g27762));
assign g15371 = ((~II17114));
assign g18173 = (g736&g17328);
assign g19557 = (g17123)|(g14190);
assign g29895 = (g2495&g29170);
assign g13063 = (g8567&g10808);
assign g26574 = ((~g24887)&(~g24861));
assign II29278 = ((~g29488))|((~II29277));
assign g14937 = ((~g12667))|((~g10421));
assign g9602 = ((~g4688)&(~g4681)&(~g4674)&(~g4646));
assign g16654 = ((~g14136));
assign g24602 = (g16507&g22854);
assign g33951 = (g33469)|(II31838)|(II31839);
assign g8593 = ((~g3759));
assign g21426 = ((~g15277));
assign g26254 = (g2413&g25349);
assign g34677 = ((~II32815));
assign II32803 = ((~g34584));
assign g9177 = ((~g3355))|((~g3401));
assign g18495 = (g2533&g15426);
assign g17618 = ((~II18580))|((~II18581));
assign g18698 = (g15131&g16777);
assign II31272 = (g32849&g32850&g32851&g32852);
assign g13628 = ((~g3372))|((~g11107));
assign g6838 = ((~g1724));
assign g9449 = ((~g5770));
assign II22366 = ((~g19757));
assign g12940 = ((~g11744));
assign g18949 = (g10183&g17625);
assign g24775 = (g17594&g22498);
assign II14330 = ((~g225))|((~g9966));
assign g20506 = ((~g15426));
assign g10159 = ((~g4477));
assign g10350 = ((~g6800));
assign II29185 = ((~g30012));
assign II15667 = ((~g12143));
assign g32641 = ((~g30614));
assign g13177 = ((~II15782));
assign g23083 = (g16076&g19878);
assign g18422 = ((~II19238));
assign g9848 = ((~g4462));
assign g25673 = (g24727)|(g21830);
assign g13671 = (g4498&g10532);
assign II12823 = ((~g4311));
assign g32611 = ((~g31154));
assign g25567 = (II24674&II24675);
assign g15594 = ((~g10614)&(~g13026)&(~g7285));
assign g19439 = ((~g15885));
assign g12144 = ((~II15003))|((~II15004));
assign II19348 = ((~g15084));
assign g24120 = ((~g19984));
assign g15832 = ((~g7903))|((~g7479))|((~g13256));
assign g31503 = (g20041&g29945);
assign g13927 = ((~g3578))|((~g11207))|((~g3632))|((~g11389));
assign g22405 = ((~g18957)&(~g20136)&(~g20114));
assign g29875 = (g28403&g23337);
assign g11893 = (g1668&g7268);
assign II22852 = (g21459)|(g21350)|(g21339);
assign g31484 = (g29775&g23418);
assign g24982 = ((~g22763));
assign II31326 = (g30735&g31853&g32926&g32927);
assign g24790 = (g7074&g23681);
assign g27645 = (g26488&g15344);
assign g20163 = ((~g16663))|((~g13938));
assign g19343 = ((~g16136));
assign g27221 = (g26055&g16747);
assign g25632 = (g24558)|(g18277);
assign g28371 = (g27177)|(g15847);
assign g23931 = ((~g20875));
assign g33564 = (g33332)|(g18388);
assign g29334 = (g29148&g18908);
assign g25690 = (g24864)|(g21889);
assign g33431 = (g32364&g32377);
assign g30396 = (g29856)|(g21755);
assign g19472 = ((~g16349));
assign g23585 = ((~g21070));
assign g25207 = (g22513&g10621);
assign g28642 = (g27555&g20598);
assign g24540 = ((~g22942));
assign g12038 = ((~II14896));
assign g12414 = ((~g7028))|((~g7041))|((~g10165));
assign g23491 = ((~g21514));
assign II14428 = ((~g8595))|((~II14427));
assign g33994 = (g33841)|(g18424);
assign g34147 = ((~g33823));
assign g29531 = (g1664&g28559);
assign g29520 = (g28291)|(g28281)|(g28264)|(g28254);
assign g32239 = (g30595)|(g29350);
assign g30378 = (g30125)|(g18487);
assign g33696 = ((~II31535));
assign g34520 = (g34294&g19505);
assign g32989 = (g32241)|(g18326);
assign g28443 = ((~II26936));
assign g10472 = ((~II13851))|((~II13852));
assign II17442 = ((~g13638));
assign g34092 = (g33750&g9104&g18957);
assign g29998 = ((~g28966));
assign g33281 = (g32142)|(g29576);
assign g13889 = ((~g11566))|((~g11435));
assign g32832 = ((~g30735));
assign g33176 = (g32198)|(II30734)|(II30735);
assign g31252 = (g29643&g20101);
assign II16476 = ((~g10430));
assign g33750 = ((~II31607));
assign g29326 = (g29105&g22155);
assign g30213 = (g28688&g23880);
assign g7928 = ((~g4776));
assign g15995 = (g13314&g1157&g10666);
assign g8830 = ((~g767));
assign g19604 = (g15704)|(g13059);
assign g12378 = ((~g9417));
assign g16072 = ((~g10961)&(~g13273));
assign g24332 = (g4459&g22228);
assign g30421 = (g29784)|(g21805);
assign g7236 = ((~g4608));
assign g32916 = ((~g31021));
assign g32410 = (g4933&g30997);
assign g18533 = (g2729&g15277);
assign g34536 = ((~II32601));
assign g12577 = ((~g7051))|((~g5990))|((~g6044));
assign g23954 = ((~II23099));
assign g27827 = ((~g9456)&(~g25839));
assign g9517 = ((~g6163));
assign g33735 = (g33118&g19553);
assign g25598 = (g24904)|(g21720);
assign g26275 = (g2417&g25349);
assign g32029 = (g31318&g16482);
assign g29355 = ((~g24383))|((~g28109));
assign g17364 = ((~g8639))|((~g14367));
assign II31342 = (g32949&g32950&g32951&g32952);
assign g24072 = ((~g20982));
assign g24719 = (g681&g23530);
assign g6849 = ((~g2551));
assign g23219 = ((~II22316));
assign g22088 = (g6307&g19210);
assign g17138 = (g255&g13239);
assign g34191 = (g33713&g24404);
assign g20041 = ((~g15569));
assign II21810 = ((~g20596));
assign g24495 = (g6928&g23127);
assign g17477 = ((~g14848));
assign g32665 = ((~g31579));
assign g15706 = (g13296&g13484);
assign g16883 = (g13509)|(g11115);
assign g11268 = ((~g7515));
assign g11963 = ((~g9153));
assign g11039 = ((~g9056)&(~g9092));
assign g18387 = (g1955&g15171);
assign g23236 = ((~g20785));
assign g15591 = ((~g4332))|((~g4322))|((~g13202));
assign g27483 = (g26488&g17642);
assign g32805 = ((~g31672));
assign g31271 = (g29706&g23300);
assign g21068 = ((~g15277));
assign g25694 = (g24638)|(g18738);
assign g20271 = ((~g16925))|((~g14054))|((~g16657))|((~g16628));
assign g29244 = (g28692)|(g18380);
assign II14610 = ((~g8993))|((~II14609));
assign g18252 = (g990&g16897);
assign g34978 = (g34874)|(g34967);
assign g29153 = ((~g27937));
assign II19796 = ((~g17870));
assign g12483 = ((~g2453)&(~g8324));
assign g27565 = ((~g26645));
assign g23996 = (g19596&g10951);
assign II14749 = ((~g10031));
assign g32692 = ((~g31528));
assign II33288 = ((~g34989));
assign g18582 = (g2922&g16349);
assign g18198 = (g15059&g17821);
assign g23450 = ((~II22571));
assign g32345 = (g2138&g31672);
assign II11721 = ((~g4145));
assign g22199 = ((~g19210));
assign g9862 = ((~g5413));
assign g25104 = (g16800&g23504);
assign g30098 = (g28548&g20774);
assign g31854 = ((~g29385));
assign g27044 = (g7766&g5873&g5881&g26241);
assign g33092 = ((~g31978)&(~g4332));
assign g24043 = ((~g20982));
assign g33727 = (g33115&g19499);
assign g18568 = (g37&g16349);
assign g25012 = (g20644&g23419);
assign g11875 = ((~II14687));
assign g27338 = ((~g9291)&(~g26616));
assign II18885 = ((~g16643));
assign g18672 = (g15127&g15758);
assign g9916 = ((~g3625));
assign II25845 = ((~g26212))|((~g24799));
assign g32351 = (g29851)|(g31281);
assign g32882 = ((~g31376));
assign II31515 = ((~g33187));
assign g28654 = (g1030&g27108);
assign g27731 = ((~g9229)&(~g25791));
assign g30300 = (g28246)|(g27252);
assign g18288 = (g1454&g16449);
assign II22922 = ((~g14677))|((~II22921));
assign g8676 = ((~g4821));
assign g12886 = ((~g10393));
assign II13729 = ((~g4534))|((~g4537));
assign g28342 = (g27134)|(g15819);
assign g15913 = (g3933&g14021);
assign g20193 = (g15578&g17264);
assign g24169 = ((~II23351));
assign g7535 = ((~g1500));
assign II32473 = ((~g34248));
assign g34032 = (g33816)|(g18706);
assign II31236 = (g30735&g31837&g32796&g32797);
assign g15914 = (g3905&g14024);
assign g32474 = ((~g31194));
assign II12580 = ((~g1239));
assign g25783 = ((~g25250));
assign g27182 = (g25818)|(g24410);
assign g28529 = ((~g8070)&(~g27617)&(~g10323));
assign II14593 = ((~g9978));
assign g26803 = ((~g25389));
assign g12124 = ((~g8741))|((~g4674));
assign g26755 = (g10776)|(g24457);
assign g21798 = (g3522&g20924);
assign g30032 = (g29072&g9326);
assign g30331 = ((~II28594));
assign g14116 = ((~g11697))|((~g11584));
assign g23474 = (g13830&g20533);
assign II24781 = ((~g24264));
assign g31707 = (g30081&g23886);
assign g8281 = ((~g3494));
assign g30226 = (g28707&g23898);
assign g7960 = ((~g1404));
assign g34270 = ((~g34159));
assign II16111 = (g8691&g11409&g11381);
assign g11018 = (g7655&g7643&g7627);
assign g24360 = ((~g22228));
assign g28313 = (g27231&g19766);
assign g6975 = ((~g4507));
assign g22901 = (g19384)|(g15745);
assign g10160 = ((~g5623))|((~g5666))|((~g5637))|((~g5659));
assign g31666 = ((~II29248));
assign g32281 = (g31257&g20500);
assign g15871 = (g3203&g13951);
assign g33235 = (g32040)|(g30982);
assign g10402 = ((~g7023));
assign g32506 = ((~g31376));
assign g25613 = (g25181)|(g18140);
assign g12120 = ((~g2476))|((~g8273));
assign II33297 = ((~g35000));
assign g16802 = (g5567&g14807);
assign II12790 = ((~g4340));
assign g16856 = ((~II18048));
assign g19513 = ((~g15969))|((~g10841))|((~g10922));
assign g29579 = (g28457&g7964);
assign g12954 = (g12186)|(g9906);
assign g9364 = ((~g5041));
assign g9013 = (g2472)|(g2491);
assign g16191 = (g5475&g14262);
assign g17699 = ((~II18681))|((~II18682));
assign g26834 = ((~II25552));
assign g30493 = (g30198)|(g21989);
assign g7586 = ((~II12056));
assign g32430 = ((~g30984));
assign g17706 = ((~g3921))|((~g11255))|((~g3983))|((~g13933));
assign II21258 = ((~g16540));
assign g21951 = (g5272&g18997);
assign II30331 = (g31672)|(g31710)|(g31021)|(g30937);
assign g14343 = ((~g11961))|((~g9670));
assign g13330 = ((~g4664))|((~g11006));
assign g12043 = (g1345&g7601);
assign g17141 = ((~II18191));
assign II13805 = ((~g6976));
assign g32459 = ((~g31070));
assign g7777 = (g723&g822&g817);
assign g33833 = (g33093&g25852);
assign g10570 = ((~g9021));
assign g25377 = (g5712&g22210&II24530);
assign g33494 = (g32700&II31166&II31167);
assign g20091 = ((~g17328));
assign g20167 = ((~g16971));
assign II31242 = (g32805&g32806&g32807&g32808);
assign gbuf144 = (g1399);
assign II15572 = ((~g10499));
assign g32941 = ((~g30735));
assign g26874 = (II25612)|(II25613);
assign g27521 = (g26519&g14700);
assign g34925 = ((~II33167));
assign g12550 = ((~g9300)&(~g9259));
assign g9036 = ((~g5084));
assign g34508 = (g34282&g19472);
assign g23987 = ((~g19277));
assign g32455 = ((~g31566)&(~II29985)&(~II29986));
assign g23589 = ((~g21468));
assign g25561 = ((~g22550));
assign g32629 = ((~g31376));
assign II26393 = ((~g26488))|((~g14227));
assign g25725 = (g25127)|(g22008);
assign g28038 = ((~g26365));
assign g16722 = ((~II17938));
assign g21918 = (g5097&g21468);
assign g29360 = (g27364&g28294);
assign g28843 = ((~g27907))|((~g7456))|((~g7387));
assign g6992 = ((~g4899));
assign g12235 = ((~g9234)&(~g9206));
assign g23057 = ((~g20453));
assign g29926 = (g1604&g28736);
assign g25138 = ((~g22472));
assign g25531 = ((~g22763))|((~g2868));
assign g32769 = ((~g31672));
assign g9971 = ((~g2093));
assign g26711 = (g25446&g20713);
assign g10058 = ((~g6497));
assign g8643 = (g2927&g2922);
assign g31473 = (g26180)|(g29666);
assign g9547 = ((~g2735));
assign II16193 = ((~g3281));
assign g21456 = ((~g15509));
assign II22298 = (g20371)|(g20161)|(g20151);
assign g34130 = ((~II32071));
assign g18336 = (g1700&g17873);
assign g34372 = (g26287)|(g34137);
assign g30505 = (g30168)|(g22026);
assign g19716 = (g12100&g17121);
assign g24438 = ((~g22722));
assign g18642 = (g15097&g17096);
assign g17679 = ((~g5611))|((~g14425))|((~g5681))|((~g12563));
assign g13779 = ((~g11804))|((~g11283));
assign g14686 = ((~g5268))|((~g12059))|((~g5276))|((~g12239));
assign g16030 = ((~g13570));
assign g27612 = (g25887&g8844);
assign g9309 = ((~g5462));
assign g31800 = ((~g29385));
assign II26929 = ((~g27980));
assign g12889 = ((~g10396));
assign g17409 = ((~II18344));
assign g28054 = (g27723)|(g18170);
assign g17494 = ((~g14339));
assign g11686 = ((~II14567));
assign g23278 = ((~g20283));
assign g23558 = ((~g20924));
assign g19886 = ((~g11403))|((~g17794));
assign g32562 = ((~g30673));
assign g30012 = ((~II28241));
assign g32912 = ((~g30735));
assign g28162 = ((~II26679));
assign g16181 = ((~g13475))|((~g13495))|((~g13057))|((~g13459));
assign g21972 = (g15152&g19074);
assign II13872 = ((~g7474));
assign g23243 = ((~g21070));
assign g32858 = ((~g31327));
assign g28405 = (g27216)|(g15875);
assign g27929 = ((~II26448));
assign g33245 = (g32125&g19961);
assign g10232 = ((~g4527));
assign g34174 = ((~g617))|((~g33851))|((~g12323));
assign II15600 = ((~g10430));
assign g20178 = ((~g16971));
assign g29080 = ((~g27779));
assign g15051 = ((~g6801)&(~g13350));
assign g20065 = ((~g16846));
assign g31232 = (g30294&g23972);
assign g15170 = ((~g7118)&(~g14279));
assign II16163 = ((~g11930));
assign g14139 = ((~g11626))|((~g11584));
assign g14536 = ((~II16651));
assign g24398 = (g23801)|(g21296);
assign g26736 = ((~g25349));
assign g26651 = (g22707&g24425);
assign g11234 = ((~g8355));
assign g7616 = ((~II12086));
assign g10709 = ((~g7499)&(~g351));
assign g31774 = (g30046)|(g30057);
assign g14396 = ((~g12119)&(~g9489));
assign g29848 = (g28260)|(g26077);
assign g25202 = ((~g23932));
assign g25411 = (g5062&g23764&II24546);
assign g24060 = ((~g21256));
assign gbuf126 = (g869);
assign II22525 = ((~g19345));
assign II20609 = ((~g16539));
assign g13038 = (g8509&g11034);
assign g32770 = ((~g31710));
assign II18543 = (g14568)|(g14540)|(g14516);
assign g33604 = (g33345)|(g18520);
assign g19636 = ((~g16987));
assign g6829 = ((~g1319));
assign g32020 = (g4157&g30937);
assign g23487 = ((~g20924));
assign II30054 = (g29385)|(g31376)|(g30735)|(g30825);
assign g33594 = (g33421)|(g18485);
assign g32228 = (g31147)|(g29651);
assign g7163 = ((~g4593));
assign g26718 = ((~g25168));
assign g17692 = (g1124&g13307);
assign g17467 = ((~g14339));
assign g25884 = (g11153&g24711);
assign g23500 = ((~g20924));
assign g31373 = ((~g4975)&(~g29725));
assign II29271 = ((~g12050))|((~II29269));
assign g29177 = ((~g27937));
assign g23358 = (g19746)|(g16212);
assign II32309 = ((~g34210));
assign g25940 = (g24415)|(g22218);
assign g32949 = ((~g30825));
assign II32116 = ((~g33937));
assign g32752 = ((~g31376));
assign g23552 = ((~II22684))|((~II22685));
assign g33804 = ((~g33250));
assign g18354 = (g1792&g17955);
assign g28927 = ((~g27837))|((~g1906))|((~g7322));
assign II15932 = ((~g12381));
assign g32314 = (g31304&g23516);
assign g33578 = (g33410)|(g18433);
assign II14395 = ((~g3654));
assign II33264 = ((~g34978));
assign g22299 = (g19999&g21024);
assign g21724 = ((~II21291));
assign II22762 = ((~g21434))|((~II22760));
assign g23392 = (g7247&g21430);
assign g24557 = (g22308)|(g19207);
assign g18201 = (g15061&g15938);
assign g28526 = (g27285)|(g26178);
assign g23691 = (g14731&g20993);
assign g32849 = ((~g31021));
assign g34749 = ((~II32921));
assign g32828 = ((~g31710));
assign g33412 = (g32362&g21411);
assign g20036 = ((~g17433));
assign g16809 = ((~g14387));
assign g10760 = ((~g1046)&(~g7479));
assign g23399 = ((~g21514));
assign g9806 = ((~g5782));
assign g27063 = ((~g26485)&(~g26516));
assign g23457 = ((~II22580));
assign II23711 = ((~g23192));
assign g28718 = (g27483)|(g16702);
assign g8133 = ((~g4809));
assign g26828 = (g24919&g15756);
assign g28885 = ((~g27742))|((~g1668))|((~g7268));
assign g23538 = ((~g20924));
assign g29302 = (g28601)|(g18798);
assign g23569 = ((~g21611));
assign II31061 = (g30825&g31806&g32543&g32544);
assign II31672 = ((~g33149));
assign g12629 = ((~g7812))|((~g7142));
assign g29785 = (g28332&g23248);
assign g33355 = (g32243&g20769);
assign g8806 = ((~g358))|((~g370))|((~g376))|((~g385));
assign g11927 = ((~g10207));
assign g24239 = (g22752)|(g18250);
assign II15107 = ((~g5313))|((~II15105));
assign g20764 = ((~II20819));
assign g34297 = (g26858)|(g34228);
assign g28291 = (g7411&g2070&g27469);
assign g26900 = (g26819)|(g24217);
assign II26508 = ((~g26814));
assign g33479 = (g32593&II31091&II31092);
assign II21838 = ((~g19263));
assign g18467 = (g2380&g15224);
assign g29078 = (g27633)|(g26572);
assign g9489 = ((~g2303));
assign g26612 = (g901&g24407);
assign II26418 = ((~g26519))|((~II26417));
assign g29886 = ((~g3288)&(~g28458));
assign g23210 = ((~g18957))|((~g2882));
assign II17143 = ((~g14412));
assign g33204 = (g32317)|(II30750)|(II30751);
assign g25720 = (g25042)|(g18765);
assign g29619 = (g2269&g29060);
assign g11326 = ((~g8993))|((~g376))|((~g365))|((~g370));
assign g20656 = ((~g17249));
assign g30130 = ((~g28761)&(~g7275));
assign g17871 = ((~II18845));
assign g28363 = ((~g27064))|((~g13593));
assign g32584 = ((~g30673));
assign g30184 = ((~g28144));
assign g14968 = ((~g12739))|((~g10312));
assign g11290 = ((~II14326));
assign g34316 = ((~g34093));
assign g23901 = (g19606&g7963);
assign II32960 = ((~g34653));
assign g25731 = (g25128)|(g22014);
assign g24716 = (g15935&g23004);
assign II25161 = ((~g24920));
assign g24550 = (g3684&g23308);
assign g33659 = ((~II31491));
assign II16328 = ((~g878));
assign g29376 = (g14002&g28504);
assign g9748 = ((~g114));
assign g32991 = (g32322)|(g18349);
assign g34286 = (g26842)|(g34216);
assign g27429 = (g25969)|(g24589);
assign g32286 = (g31658&g29312);
assign g13542 = (g10053&g11927);
assign g11414 = ((~g8591)&(~g8593));
assign g29857 = (g28386&g23304);
assign g23431 = ((~g21514));
assign g17672 = ((~g14720));
assign g32338 = (g31466&g20668);
assign II31800 = ((~g33164));
assign g23623 = ((~g9364))|((~g20717));
assign g26634 = ((~g25317));
assign g27774 = ((~II26381));
assign g18779 = (g5821&g18065);
assign g25266 = ((~g22228));
assign g17792 = ((~g6601))|((~g14602))|((~g6697))|((~g12721));
assign g10212 = ((~g6390));
assign g28147 = ((~II26654));
assign II33249 = ((~g34971));
assign g7110 = ((~g6682));
assign g22982 = (g19535&g19747);
assign g12143 = ((~II14999));
assign g13809 = ((~II16135));
assign g14914 = ((~g12822)&(~g12797));
assign g29955 = ((~g28950));
assign g16482 = ((~g13464));
assign II22149 = ((~g21036));
assign g32209 = (g31122)|(g29599);
assign g16506 = (g13294)|(g10966);
assign g10115 = ((~g2283));
assign II18788 = ((~g13138));
assign II30756 = (g32088)|(g32163)|(g32098)|(g32105);
assign g7947 = ((~g1500));
assign g30386 = (g30139)|(g18523);
assign g25872 = (g3119&g24655);
assign g33094 = ((~g31950)&(~g4639));
assign g8310 = ((~g2051));
assign g19363 = (g17810)|(g14913);
assign g34726 = (g34665)|(g18212);
assign g12367 = ((~II15205));
assign II32237 = ((~g34130));
assign g33329 = (g32210&g20585);
assign g24288 = (g4417&g22550);
assign g12294 = ((~g10044))|((~g7018))|((~g10090));
assign g10720 = (g2704&g10219&g2689);
assign II11835 = ((~g101));
assign g28614 = (g27351)|(g26311);
assign g24872 = (g23088&g9104);
assign II12373 = ((~g3457))|((~II12372));
assign g32602 = ((~g30825));
assign g9927 = ((~g5689));
assign g28303 = (g7462&g2629&g27494);
assign g8623 = ((~g3990));
assign g34062 = ((~g33711));
assign g27219 = (g26026&g16742);
assign g34674 = ((~II32806));
assign g19788 = (g9983&g17216);
assign g27710 = (g26422&g20904);
assign g23861 = ((~g19147));
assign g34942 = ((~g34928));
assign g29835 = (g28326&g24866);
assign g15101 = ((~g12871)&(~g14591));
assign II15682 = ((~g12182));
assign g32114 = (g31624&g29927);
assign g19746 = (g9816&g17147);
assign g31750 = (g30103&g23925);
assign g14097 = (g878&g10632);
assign g34139 = (g33827&g23314);
assign g15674 = ((~g921))|((~g13110));
assign g31928 = (g31517)|(g22092);
assign II31277 = (g32856&g32857&g32858&g32859);
assign g7431 = ((~g2555));
assign II32678 = ((~g34428));
assign g7315 = ((~g1772));
assign g16608 = ((~g14116));
assign II31051 = (g31376&g31804&g32529&g32530);
assign g7497 = ((~g6358));
assign II22353 = ((~g19375));
assign II29211 = ((~g30298));
assign II27513 = (g19984&g24089&g24090&g28034);
assign g34250 = (g34111)|(g21713);
assign g7275 = ((~g1728));
assign g34483 = (g34406&g18938);
assign II29221 = ((~g30307));
assign g27577 = ((~g25019))|((~g25002))|((~g24988))|((~g25765));
assign g14075 = ((~g11658))|((~g11527));
assign g9021 = ((~II12954));
assign g16769 = ((~g13530));
assign g7957 = ((~g1252));
assign g21465 = (g16155&g13663);
assign g30191 = (g28647&g23843);
assign g18451 = (g2295&g15224);
assign II18350 = ((~g13716));
assign g12526 = ((~g10194))|((~g7110))|((~g10213));
assign g27525 = (g26576&g17720);
assign g22051 = (g6105&g21611);
assign g31795 = ((~II29371));
assign g30984 = (g29765)|(g29755);
assign g23283 = ((~g20785));
assign g24005 = ((~II23149));
assign g30983 = ((~g29657));
assign g27996 = ((~II26508));
assign g22019 = (g5857&g19147);
assign g11134 = ((~g8138))|((~g8240))|((~g8301));
assign g33976 = (g33869)|(g18347);
assign g34748 = (g34672&g19529);
assign g33036 = (g32168)|(g24309);
assign g30609 = (g13633)|(g29742);
assign g20229 = ((~g17015));
assign g7344 = ((~g5659));
assign g12830 = ((~g9995));
assign g25905 = (g24879&g16311);
assign g19140 = ((~g7939)&(~g15695));
assign g10967 = (g7880&g1448);
assign g24178 = ((~II23378));
assign g23652 = ((~II22785));
assign II17892 = ((~g3325));
assign g12841 = ((~g10357));
assign g24156 = ((~II23312));
assign gbuf137 = (g1418);
assign g33623 = (g33370)|(g18792);
assign g19651 = (g1111&g16119);
assign g23800 = ((~g21246));
assign g19522 = (g17057)|(g14180);
assign g14320 = ((~g9257)&(~g11111));
assign g16738 = ((~II17956));
assign g21803 = (g3538&g20924);
assign g34795 = (g34753)|(g18572);
assign II13637 = ((~g102));
assign g12422 = ((~II15238));
assign g19353 = ((~II19831));
assign g29255 = (g28714)|(g18516);
assign II11697 = ((~g3352));
assign II22785 = ((~g18940));
assign g31809 = ((~g29385));
assign g7362 = ((~g1906));
assign g27673 = (g25769&g23541);
assign g20110 = ((~g16897));
assign g26700 = ((~g25429));
assign g21066 = (g10043&g17625);
assign g22488 = ((~g19699)&(~g1002));
assign g11346 = ((~g7980)&(~g7964));
assign g23915 = ((~g19277));
assign g21703 = (g146&g20283);
assign II14714 = ((~g5128))|((~II14712));
assign g25539 = (g23531)|(g20628);
assign II16201 = ((~g4023));
assign g34446 = (g34390)|(g18550);
assign g28950 = ((~g27937))|((~g7490))|((~g2599));
assign g30264 = (g28774&g23963);
assign g25629 = (g24962)|(g18258);
assign g29945 = ((~II28174));
assign g26208 = ((~g7975))|((~g24751));
assign g13024 = ((~g11900));
assign g20528 = ((~g15224));
assign g34591 = ((~II32681));
assign II18154 = ((~g13177));
assign g16731 = (g7153&g12941);
assign g27437 = (g26576&g17589);
assign g14307 = ((~II16468));
assign g10272 = ((~II13705));
assign g27613 = ((~g24942))|((~g24933))|((~g25048))|((~g26871));
assign II12568 = ((~g5005));
assign g31507 = ((~g9064)&(~g29556));
assign II22499 = ((~g21160));
assign g31003 = ((~g27163))|((~g29497))|((~g19644));
assign g24744 = ((~g22202));
assign g25495 = ((~g12483))|((~g22472));
assign g20387 = ((~g15426));
assign II18177 = ((~g13191));
assign g20698 = ((~g17873));
assign g13716 = ((~II16090));
assign g21333 = (g1300&g15740);
assign g21915 = (g5080&g21468);
assign g12287 = ((~g8381))|((~g2587));
assign g23725 = (g14772&g21138);
assign g29850 = (g28340&g24893);
assign g25576 = (g24141)|(g24142);
assign g18658 = (g15121&g17183);
assign g7397 = ((~g890));
assign g10090 = ((~g5348));
assign g14519 = ((~g3889))|((~g11225))|((~g4000))|((~g8595));
assign g20446 = ((~g15224));
assign g21737 = (g3068&g20330);
assign g24603 = ((~g23108));
assign g30157 = ((~g28833)&(~g7369));
assign g30552 = (g30283)|(g22123);
assign g12342 = ((~g7004))|((~g7018))|((~g10129));
assign g29071 = ((~g5873)&(~g28020));
assign g34244 = ((~II32231));
assign g13410 = ((~II15921));
assign g7648 = ((~II12135));
assign g33332 = (g32217&g20608);
assign g18375 = (g1902&g15171);
assign g17392 = ((~g14924));
assign g8282 = ((~g3841));
assign g30294 = ((~g7110)&(~g29110));
assign II23601 = ((~g22360))|((~II23600));
assign g13415 = (g837&g11048);
assign g24255 = (g22835)|(g18308);
assign g14453 = ((~II16610));
assign II23120 = ((~g417))|((~II23118));
assign g17684 = ((~g15036));
assign II24448 = ((~g22923));
assign g12853 = ((~g6848)&(~g10430));
assign g33133 = ((~g32278)&(~g31503));
assign II27555 = ((~g28142));
assign g25453 = (g5406&g23789&II24576);
assign g34541 = (g34331&g20087);
assign g7139 = ((~g5406)&(~g5366));
assign g27925 = ((~II26439))|((~II26440));
assign g29573 = (g1752&g28892);
assign g24607 = (g5817&g23666);
assign g27964 = (g25956&g22492);
assign g17654 = (g962&g13284);
assign g18820 = (g15166&g15563);
assign g15968 = (g13038)|(g10677);
assign g25879 = (g11135&g24683);
assign g25425 = ((~g20081))|((~g23172));
assign II16762 = ((~g5290));
assign g33100 = ((~g32172)&(~g31188));
assign g12890 = ((~g10397));
assign g21246 = ((~II20985));
assign g34460 = (g34301)|(g18677);
assign II25146 = ((~g24911));
assign g9259 = ((~g5176));
assign g16861 = ((~II18051));
assign g19399 = ((~g16489));
assign II19775 = ((~g17780));
assign g9800 = ((~g5436))|((~g5428));
assign g13077 = (g11330)|(g943);
assign g9660 = ((~g3267));
assign g14048 = ((~g11658))|((~g11483));
assign g31944 = (g31745&g22146);
assign g18940 = ((~II19719));
assign g12188 = ((~g8249))|((~g1894));
assign g11878 = ((~II14690));
assign g30255 = (g28748&g23946);
assign g19139 = (g452&g16195);
assign g19801 = ((~II20216));
assign g32122 = (g31646&g29944);
assign g10827 = (g8914&g4258);
assign g28789 = (g21434&g26424&g25340&g27440);
assign g19063 = ((~g7909)&(~g15674));
assign g13516 = ((~g11533))|((~g11490))|((~g11444))|((~g11412));
assign g28441 = ((~g27629));
assign g25297 = ((~g23746));
assign g33377 = ((~II30901));
assign g20637 = ((~g15224));
assign g30534 = (g30213)|(g22080);
assign g12191 = ((~II15052))|((~II15053));
assign g28076 = (g27098)|(g21878);
assign g18134 = (g534&g17249);
assign g25407 = ((~g23871)&(~g14645));
assign g29763 = (g28217)|(g22762);
assign g18283 = (g1384&g16136);
assign II29571 = ((~g31783));
assign g18829 = ((~g15171));
assign g34857 = (g16540&g34813);
assign g18712 = (g4843&g15915);
assign g12862 = ((~g10370));
assign g29742 = (g28288&g10233);
assign II18446 = ((~g13028));
assign g27202 = (g25997&g13876);
assign g7456 = ((~g2495));
assign g24979 = ((~g22369));
assign II13140 = ((~g6154))|((~II13139));
assign g8356 = ((~g54));
assign g33110 = (g32404&g32415);
assign g12046 = ((~g10036)&(~g9640));
assign g17668 = ((~g3235))|((~g13765))|((~g3310))|((~g13877));
assign g33968 = (g33855)|(g18320);
assign g12651 = ((~g9269)&(~g5511));
assign g34869 = (g34816&g19869);
assign g34813 = ((~II33027));
assign g33902 = (g33085&g13202);
assign g33897 = (g33315&g20777);
assign g29712 = (g2643&g28726);
assign g33117 = ((~g31261)&(~g32205));
assign II22576 = ((~g21282));
assign II14368 = ((~g8481))|((~g3303));
assign g22079 = (g6271&g19210);
assign g33477 = (g32577&II31081&II31082);
assign g8296 = ((~g246));
assign g23062 = (g718&g20248);
assign g7522 = ((~g6661));
assign g10605 = ((~g2555))|((~g7490));
assign g31866 = (g31252)|(g18142);
assign g22456 = ((~g19801));
assign g29512 = (g2161&g28793);
assign g19662 = ((~g17432));
assign g23484 = (g20160&g20541);
assign g30080 = (g28121&g20674);
assign g32979 = (g32181)|(g18177);
assign g33004 = (g32246)|(g18431);
assign g29109 = ((~g9472)&(~g26994));
assign g34194 = (g33811)|(g33815);
assign g11126 = (g6035&g10185);
assign g12794 = (g1008&g7567);
assign g27209 = (g26213&g8365&g2051);
assign g26880 = (g26610)|(g24186);
assign g32176 = (g2779&g31623);
assign g34383 = ((~II32388));
assign g27145 = (g14121&g26382);
assign g10363 = ((~II13779));
assign g18299 = (g1526&g16489);
assign g9669 = ((~g5092));
assign g25175 = ((~g5736)&(~g23692));
assign g33030 = (g32166)|(g21826);
assign g24485 = (g10710&g22319);
assign g31995 = (g28274&g30569);
assign g18500 = (g2421&g15426);
assign g12511 = ((~g7028))|((~g5644))|((~g5698));
assign g26156 = (g2028&g25135);
assign g27403 = (g25962)|(g24581);
assign g31891 = (g31305)|(g21824);
assign g20151 = ((~g17598))|((~g14570))|((~g17514))|((~g14519));
assign g34420 = ((~g34152));
assign g13514 = ((~II15987));
assign g15014 = ((~g12785))|((~g12680));
assign g32583 = ((~g30614));
assign g31016 = (g29478&g22840);
assign II18531 = ((~g14640))|((~II18529));
assign g13125 = ((~g7863)&(~g10762));
assign II23324 = ((~g21697));
assign g21273 = ((~II21006));
assign g16637 = (g5949&g14968);
assign g34864 = ((~g34840));
assign g30045 = (g29200&g12419);
assign g23516 = ((~g20924));
assign g10597 = ((~g10233));
assign g31019 = (g29481&g22856);
assign g24579 = ((~g23067));
assign g9152 = ((~g2834));
assign g15712 = (g3791&g13521);
assign g26129 = (g2384&g25121);
assign g14528 = (g12459&g12306&g12245&II16646);
assign g8058 = ((~g3115));
assign II12167 = ((~g5176));
assign g18181 = (g772&g17328);
assign g32674 = ((~g30735));
assign g18768 = (g5503&g17929);
assign g28532 = (g27394&g20265);
assign g28100 = (g27690)|(g22051);
assign g26829 = (g2844&g24505);
assign g9934 = ((~g5849));
assign g12798 = ((~g5535)&(~g9381));
assign g25502 = (g6946&g22527);
assign g31821 = ((~g29385));
assign II23980 = ((~g13670))|((~II23978));
assign g13959 = ((~g3698)&(~g11309));
assign g23393 = ((~g20739));
assign g17720 = ((~g15045));
assign g15130 = ((~g13638)&(~g6985));
assign g33081 = (g32388&g18875);
assign g10588 = (g7004&g5297);
assign g15841 = (g4273&g13868);
assign g19499 = ((~g16782));
assign g23254 = (g20056&g20110);
assign g22836 = ((~g18918))|((~g2852));
assign g33717 = (g14092&g33306);
assign II16651 = ((~g10542));
assign g15825 = ((~g7666)&(~g13217));
assign II18529 = ((~g1811))|((~g14640));
assign g32713 = ((~g30673));
assign g11513 = ((~g7948));
assign g6984 = ((~g4709));
assign g12817 = (g1351&g7601);
assign g34425 = ((~II32446));
assign g34778 = ((~II32976));
assign II20188 = ((~g16272))|((~II20187));
assign g23711 = ((~g9892)&(~g21253));
assign II24585 = (g9621&g9892&g6439);
assign g26122 = (g24557&g19762);
assign g27561 = (g26100)|(g24702);
assign g24482 = (g6875&g23055);
assign g33261 = (g32111)|(g29525);
assign g19764 = ((~II20166))|((~II20167));
assign g15694 = (g457&g13437);
assign g11881 = ((~g9060))|((~g3361));
assign g9264 = ((~g5396));
assign g32465 = ((~g30825));
assign g34122 = ((~II32059));
assign g14701 = ((~g12351));
assign g14348 = ((~g10887));
assign g34766 = ((~g34703));
assign g33539 = (g33245)|(g18178);
assign g25055 = ((~g23590));
assign g28395 = ((~g27074))|((~g13655));
assign g27546 = (g26549&g17758);
assign gbuf78 = (g3325);
assign g18566 = (g2860&g16349);
assign g18449 = (g12852&g15224);
assign g30463 = (g30140)|(g21934);
assign g27628 = (g26400&g18061);
assign g29983 = ((~g28977));
assign II13111 = ((~g5813))|((~II13109));
assign II23342 = ((~g23299));
assign g12081 = ((~g10079)&(~g9694));
assign g34764 = (g34691&g20009);
assign g30121 = (g28577&g21052);
assign g6957 = ((~g2932));
assign g27468 = ((~g24951))|((~g24932))|((~g24925))|((~g26852));
assign g28511 = (g27272)|(g16208);
assign g31513 = (g2606&g29318);
assign g24991 = ((~g22369));
assign g28691 = (g27437)|(g16642);
assign g32112 = (g31646&g29923);
assign g14194 = ((~g5029)&(~g10515));
assign II18297 = ((~g1418));
assign g30020 = ((~g29097));
assign g28269 = (g27205&g19712);
assign g6926 = ((~g3853));
assign g34610 = (g34507)|(g18564);
assign g19980 = ((~g17226));
assign g7097 = ((~II11809));
assign g23221 = ((~g20785));
assign g17775 = ((~g6255))|((~g14575))|((~g6351))|((~g12672));
assign g24822 = (g3010&g23534&II24003);
assign g34621 = (g34517)|(g18583);
assign g15093 = ((~g13177)&(~g6904));
assign g18543 = (g2779&g15277);
assign g25060 = ((~g23708));
assign g25669 = (g24657)|(g18624);
assign g8742 = ((~g4035));
assign g29612 = (g27875&g28633);
assign g13031 = ((~g7301)&(~g10741));
assign g29483 = (g25801)|(g28130);
assign g12871 = ((~g10378));
assign g24670 = (g5138&g23590);
assign g33909 = (g33131&g10708);
assign g10375 = ((~g6941));
assign g16526 = ((~g13898));
assign g22149 = (g14581&g18880);
assign g29012 = ((~g5863)&(~g28020));
assign g23340 = ((~g21070));
assign g28516 = ((~g10857))|((~g26105))|((~g27155));
assign g13708 = ((~g11200))|((~g8507));
assign II22583 = ((~g20998));
assign g11945 = ((~g7212)&(~g7228));
assign g16311 = ((~g13273));
assign g20841 = ((~g17847)&(~g12027));
assign II17626 = ((~g14582));
assign g30350 = (g30118)|(g18334);
assign g17152 = (g8635&g12997);
assign g15145 = ((~g12891)&(~g13716));
assign g21385 = ((~g17736))|((~g14696))|((~g17679))|((~g14636));
assign g13855 = ((~g4944))|((~g11804));
assign g24524 = ((~g22876));
assign g18737 = (g4975&g16826);
assign g13940 = ((~g11426))|((~g8889))|((~g11707))|((~g8829));
assign g24283 = (g4411&g22550);
assign g28857 = ((~g27779))|((~g1802))|((~g1728));
assign g10369 = ((~g6873));
assign g33982 = (g33865)|(g18372);
assign g13676 = ((~g11834))|((~g11283));
assign g24943 = ((~g20068))|((~g23172));
assign g18602 = (g3115&g16987);
assign II22024 = ((~g19350));
assign g7625 = ((~II12109));
assign g33383 = (g32244)|(g29940);
assign g18232 = (g1124&g16326);
assign g32015 = ((~II29571));
assign g18637 = (g3821&g17096);
assign g34006 = (g33897)|(g18462);
assign II12242 = ((~g1105))|((~II12240));
assign g10887 = (g7812&g6565&g6573);
assign g29913 = ((~g28840));
assign g26344 = (g2927)|(g25010);
assign g15071 = ((~g6831)&(~g13416));
assign g31298 = (g30169&g27886);
assign g32521 = ((~g31376));
assign g33532 = (g32974&II31356&II31357);
assign g24570 = ((~g22957))|((~g2941));
assign II30989 = ((~g32441));
assign g16521 = ((~g13543));
assign II16721 = (g10224&g12589&g12525);
assign g21933 = (g5212&g18997);
assign g28946 = ((~g27907))|((~g2495))|((~g2421));
assign g32972 = ((~g31710));
assign g30519 = (g30264)|(g22040);
assign g17414 = ((~g14627));
assign g30500 = (g29326)|(g21996);
assign g31525 = (g29892&g23526);
assign g30063 = ((~g29015));
assign g27506 = (g26021)|(g24639);
assign g21844 = (g3873&g21070);
assign g20150 = ((~g17705))|((~g17669))|((~g17635))|((~g14590));
assign g18509 = (g2587&g15509);
assign g32896 = ((~g31376));
assign g32276 = (g31646&g30313);
assign g14247 = ((~g9934)&(~g10869));
assign g9888 = ((~g5831));
assign g21188 = (g7666&g15705);
assign g34682 = ((~II32824));
assign g27579 = (g26157)|(g24748);
assign g21825 = (g3736&g20453);
assign g18241 = (g1183&g16431);
assign g8898 = ((~g676));
assign g15816 = ((~II17314));
assign g24247 = (g22623)|(g18259);
assign g34512 = ((~g34420));
assign g28172 = (g27469)|(g27440)|(g27416)|(g27395);
assign g34353 = (g26088)|(g34114);
assign g34048 = ((~g33669))|((~g10583))|((~g7442));
assign g33447 = ((~g31978)&(~g7643));
assign g32737 = ((~g31327));
assign g25965 = (g2208&g24980);
assign g31811 = ((~g29385));
assign II31312 = (g32905&g32906&g32907&g32908);
assign g25069 = (g23296&g20535);
assign g17689 = ((~g6645))|((~g12137))|((~g6661))|((~g14786));
assign g15725 = ((~g5603))|((~g14522))|((~g5681))|((~g9864));
assign g14041 = ((~g11610))|((~g11473));
assign g15797 = (g3909&g14139);
assign g24503 = (g22225&g19409);
assign g23378 = ((~g21070));
assign g20681 = ((~g15483));
assign II12779 = ((~g4210));
assign g14514 = ((~g11959)&(~g9760));
assign g14996 = ((~g12662))|((~g10312));
assign g15962 = ((~g14833))|((~g9417))|((~g9340));
assign g24420 = (g23997&g18980);
assign g33450 = (g32266&g29737);
assign g33937 = ((~II31823));
assign g23814 = ((~g19074));
assign g18934 = (g3133&g16096);
assign g13086 = ((~g6235))|((~g12101))|((~g6346))|((~g10003));
assign g34455 = (g34284)|(g18668);
assign g13132 = ((~g10632));
assign g16593 = (g5599&g14885);
assign g20207 = ((~g17015));
assign g27583 = ((~g26686));
assign g33422 = (g32375&g21456);
assign g25242 = ((~g23684));
assign g29227 = (g28456)|(g18169);
assign II18600 = ((~g5335));
assign g18433 = (g2197&g18008);
assign g7567 = ((~g979)&(~g990));
assign g33790 = (g33108&g20643);
assign g34171 = (g33925&g24360);
assign II32699 = ((~g34569));
assign II14633 = ((~g9340));
assign II11629 = ((~g19));
assign g22547 = (g16855)|(g20215);
assign g11202 = ((~II14267));
assign g32939 = ((~g31327));
assign g31118 = (g29490&g22906);
assign g33145 = ((~g8677)&(~g32072));
assign g24241 = (g22920)|(g18252);
assign g27395 = (g8046&g26314&g9187&g9077);
assign g32088 = (g27241&g31070);
assign g20706 = ((~g18008));
assign g21685 = ((~II21246));
assign g12902 = ((~g10409));
assign g26859 = ((~II25591));
assign g26284 = ((~g24875));
assign g28864 = ((~g27886))|((~g7411))|((~g1996));
assign g25557 = ((~g22763));
assign g32096 = (g31601&g29893);
assign II27508 = (g19935&g24082&g24083&g28033);
assign g31885 = (g31017)|(g21779);
assign g30394 = (g29805)|(g21753);
assign g22038 = (g5945&g19147);
assign g23003 = ((~II22180));
assign g16656 = ((~II17852));
assign g28116 = (g27366&g26183);
assign g13458 = ((~g11048));
assign g23894 = ((~g19074));
assign g9538 = ((~g1792))|((~g1760));
assign g30177 = (g28631&g23814);
assign g29183 = ((~g9392)&(~g28020)&(~g7766));
assign g18688 = (g4704&g16752);
assign g16216 = ((~II17557));
assign g23572 = (g20230&g20656);
assign g26250 = (g1902&g25429);
assign g20994 = ((~g15615));
assign g32572 = ((~g30735));
assign g11709 = ((~II14584));
assign g20087 = ((~g17249));
assign g13040 = ((~g5196))|((~g12002))|((~g5308))|((~g9780));
assign g28158 = (g26424&g22763&g27037);
assign g10262 = ((~g586));
assign g10610 = ((~g7462))|((~g7490));
assign g14575 = ((~g10050)&(~g12749));
assign II27388 = ((~g27698));
assign g24987 = ((~g23630));
assign g7632 = ((~II12117));
assign g14210 = (g4392&g10590);
assign g13821 = ((~g11251))|((~g8340));
assign g20782 = ((~g15853));
assign g21428 = ((~g15758));
assign g21721 = (g385&g21037);
assign g29906 = ((~g28793));
assign g22927 = ((~II22128));
assign g18301 = (g1532&g16489);
assign g31753 = ((~II29314))|((~II29315));
assign g11182 = ((~II14241));
assign g23021 = ((~g20283));
assign g17649 = ((~II18614));
assign g8778 = ((~II12758));
assign g25225 = ((~g23802));
assign g14727 = ((~g12604))|((~g12505));
assign g13493 = (g9880&g11866);
assign g34699 = ((~II32855));
assign g25895 = ((~g1259))|((~g24453));
assign g24583 = ((~g22753))|((~g22711));
assign II33167 = ((~g34890));
assign g15061 = ((~g6815)&(~g13394));
assign g13898 = ((~g11621))|((~g11747));
assign g32930 = ((~g31021));
assign g21182 = ((~g15509));
assign II15732 = ((~g6692));
assign g25985 = ((~g24631))|((~g23956));
assign g11442 = ((~g8644))|((~g3288))|((~g3343));
assign II32690 = ((~g34432));
assign g24567 = ((~g22957))|((~g2917));
assign g34490 = ((~II32547));
assign g25931 = (g24574&g19477);
assign g26325 = (g12644&g25370);
assign g22643 = ((~g20136))|((~g18954));
assign g34695 = (g34523)|(g34322);
assign g17719 = (g9818&g14675);
assign g27970 = (g26514)|(g25050);
assign II21242 = ((~g16540));
assign g13249 = ((~g10590));
assign II31352 = (g32963&g32964&g32965&g32966);
assign II18625 = ((~g2079))|((~g14712));
assign g10413 = ((~g7110));
assign II16502 = ((~g10430));
assign g17246 = ((~g9439))|((~g9379))|((~g14405));
assign g27375 = (g26519&g17479);
assign g28288 = ((~g10533))|((~g26105))|((~g27004));
assign g34305 = (g25775)|(g34050);
assign g33049 = (g31966)|(g21929);
assign II15609 = ((~g12013));
assign g12368 = ((~II15208));
assign g18517 = (g2652&g15509);
assign g34136 = (g33850&g23293);
assign g17193 = (g2504&g13023);
assign II13443 = ((~g262))|((~II13442));
assign g18887 = ((~g15373));
assign II31776 = ((~g33204));
assign g21872 = (g4098&g19801);
assign g23497 = (g20169&g20569);
assign g15839 = (g3929&g13990);
assign II33210 = ((~g34943));
assign g12981 = (g12219)|(g9967);
assign g19697 = ((~g16886));
assign g14423 = ((~II16579));
assign g10038 = ((~g2241));
assign g30499 = (g30261)|(g21995);
assign g29261 = (g28247)|(g18605);
assign g19474 = ((~g11609))|((~g17794));
assign g33048 = (g31960)|(g21928);
assign g16535 = (g5595&g14848);
assign g20578 = ((~g15563));
assign g28056 = (g27230)|(g18210);
assign g27971 = ((~g26673));
assign g27029 = (g26327&g11031);
assign g33890 = (g33310&g20659);
assign g18340 = (g1720&g17873);
assign g12820 = ((~g10233));
assign g12435 = ((~g9012)&(~g8956)&(~g8904)&(~g8863));
assign II15079 = ((~g9827))|((~II15078));
assign g9429 = ((~g3723));
assign g29222 = (g28252)|(g18105);
assign g12204 = ((~g9927)&(~g10160));
assign II24033 = (g8219&g8443&g3747);
assign g22975 = ((~g20391));
assign g27832 = ((~II26409));
assign g10473 = ((~II13857));
assign g32791 = ((~g31672));
assign g10394 = ((~g6994));
assign II26649 = ((~g27675));
assign g14092 = ((~g8774)&(~g11083));
assign g24122 = ((~g20857));
assign II31482 = ((~g33204));
assign g12022 = ((~g7335))|((~g2331));
assign g33297 = (g32157)|(g29621);
assign II31077 = (g32566&g32567&g32568&g32569);
assign g9842 = ((~g3274));
assign g29190 = ((~g27046));
assign g34499 = (g31288&g34339);
assign g16686 = ((~II17892));
assign II12214 = ((~g6561));
assign g23514 = (g20149&g11829);
assign g21352 = ((~g16322));
assign g25657 = (g24624)|(g21782);
assign g33123 = (g31962)|(g30577);
assign g33344 = (g32228&g20670);
assign g15650 = (g8362&g13413);
assign g34037 = (g33803)|(g18734);
assign g23324 = ((~g703))|((~g20181));
assign g32052 = (g31507&g13885);
assign g25255 = ((~g20979))|((~g23659));
assign g32620 = ((~g30673));
assign II12451 = ((~g3092));
assign g19733 = ((~g16856));
assign g8343 = ((~g3447));
assign g29371 = ((~II27735));
assign g33569 = (g33415)|(g18402);
assign g19414 = ((~g16349));
assign g12938 = ((~II15556));
assign g12107 = ((~g9687));
assign g34404 = (g34182)|(g25102);
assign g20695 = ((~II20781));
assign II14276 = ((~g8218))|((~II14275));
assign g32358 = (g29866)|(g31297);
assign g31783 = (II29351)|(II29352);
assign g16220 = ((~g13499)&(~g4939));
assign g26081 = ((~g24619));
assign g23223 = ((~g21308));
assign g32699 = ((~g31528));
assign g32839 = ((~g30735));
assign II12289 = ((~g1300))|((~II12287));
assign II23381 = ((~g23322));
assign II16371 = ((~g887));
assign g23172 = ((~II22275));
assign g15150 = ((~g12895)&(~g13745));
assign g31283 = (g30156&g27837);
assign II20846 = ((~g16923));
assign g21346 = ((~g17821));
assign g13475 = ((~g1008))|((~g11294))|((~g11786));
assign g20669 = ((~g15426));
assign g31139 = (g12221&g30036);
assign g9670 = ((~g5022));
assign g32984 = (g31934)|(g18264);
assign g31916 = (g31756)|(g22002);
assign g16674 = (g6637&g15014);
assign g18347 = (g1756&g17955);
assign g30233 = (g28720&g23913);
assign g15750 = ((~g13291));
assign g17525 = ((~g14600))|((~g14574));
assign g34920 = ((~II33152));
assign g27356 = ((~g9429)&(~g26657));
assign II13184 = ((~g6505))|((~II13182));
assign g28633 = ((~g27687));
assign g24626 = ((~g23139));
assign g28820 = ((~g27742))|((~g1668))|((~g1592));
assign g19430 = ((~g17150)&(~g14220));
assign g20871 = ((~g14434))|((~g17396));
assign g18175 = (g744&g17328);
assign g12896 = ((~g10402));
assign II15846 = ((~g11183));
assign g22683 = ((~II22000));
assign g15937 = (g11950&g14387);
assign II31817 = ((~g33323));
assign II13326 = ((~g66));
assign g26925 = (g25939)|(g18301);
assign g34187 = (g33708&g24397);
assign g23103 = (g10143&g20765);
assign g9283 = ((~g1736));
assign g20160 = (g16163)|(g13415);
assign g22707 = (g20559)|(g17156);
assign g27989 = ((~g26759));
assign g9073 = ((~g150));
assign g27277 = (g26359&g14191);
assign g22090 = (g6404&g18833);
assign g9212 = ((~g6466));
assign g11446 = ((~g8700))|((~g6941))|((~g8734));
assign g11425 = ((~g7640));
assign g23665 = ((~g21562));
assign g25708 = (g25526)|(g18751);
assign g21607 = ((~g17873));
assign g14004 = ((~g11149));
assign g22922 = ((~g20330));
assign g29632 = (g28899&g22417);
assign g18717 = (g4849&g15915);
assign g31293 = (g29582)|(g28299);
assign II26460 = ((~g26576))|((~II26459));
assign g24024 = ((~g21193));
assign g29778 = ((~g294))|((~g28444))|((~g23204));
assign II31112 = (g32617&g32618&g32619&g32620);
assign g32206 = (g30609&g25524);
assign g21905 = ((~II21486));
assign g18370 = (g1874&g15171);
assign g25938 = (g8997&g24953);
assign II18819 = (g13156&g11450&g11498);
assign g24296 = (g4382&g22550);
assign g25446 = ((~g23686)&(~g14645));
assign g7051 = ((~II11793));
assign g27084 = ((~g26673));
assign g10206 = ((~g4489));
assign II32639 = ((~g34345));
assign g24321 = (g4558&g22228);
assign g20564 = ((~g15373));
assign g24085 = ((~g20857));
assign g25153 = ((~g23733));
assign g12686 = ((~g7097))|((~g6682))|((~g6736));
assign g16296 = ((~g9360))|((~g13501));
assign g11769 = ((~g8626));
assign g25644 = (g24622)|(g21737);
assign g19208 = ((~g17367));
assign g22666 = ((~g18957))|((~g2878));
assign II32187 = ((~g33661))|((~II32185));
assign g26089 = (g24501)|(g22534);
assign II12605 = ((~g1570));
assign g24265 = (g22316)|(g18560);
assign g17527 = ((~g14741));
assign gbuf94 = (g4012);
assign g13914 = (g8643)|(g11380);
assign g31466 = (g26160)|(g29650);
assign g32539 = ((~g31170));
assign g12638 = ((~g7514))|((~g6661));
assign g20171 = (g16479&g10476);
assign g22447 = (g21464)|(g12761);
assign g21758 = (g3191&g20785);
assign II32192 = ((~g33628));
assign g7686 = ((~g4659));
assign g21762 = (g3219&g20785);
assign gbuf133 = (g799);
assign g28204 = (g26098&g27654);
assign g25553 = ((~g22550));
assign g12371 = ((~g1760)&(~g8195));
assign g16762 = (g5901&g14930);
assign g14447 = ((~g11938)&(~g9698));
assign g27457 = (g26519&g17606);
assign II15811 = ((~g11128));
assign g17685 = ((~II18662));
assign II25677 = ((~g25640));
assign g27248 = (g24880)|(g25953);
assign g14978 = ((~g12716))|((~g10491));
assign g24799 = (g23901)|(g23921);
assign g32394 = ((~g30601));
assign g9197 = ((~g1221));
assign g16125 = (g5152&g14238);
assign g10533 = ((~g8795));
assign g28499 = (g27982&g17762);
assign g8397 = ((~g3470));
assign g34671 = ((~II32797));
assign g21879 = (g4132&g19801);
assign II18168 = ((~g13191));
assign g29199 = (g27187&g12687);
assign g16610 = (g5260&g14918);
assign g16596 = (g5941&g14892);
assign g10110 = ((~g661));
assign g21383 = ((~g17367));
assign II22289 = ((~g19446));
assign g32864 = ((~g30937));
assign g11143 = ((~g8032));
assign g25773 = ((~g24453));
assign g32746 = ((~g30735));
assign g20585 = ((~g17955));
assign g7596 = ((~II12070));
assign II23963 = ((~g13631))|((~II23961));
assign g9456 = ((~g6073));
assign g33700 = (g33148&g11012);
assign II32756 = ((~g34469))|((~g25779));
assign g11480 = ((~g10323))|((~g8906));
assign g10380 = ((~g6960));
assign g34267 = (g34079)|(g18728);
assign g24092 = ((~g20857));
assign g23927 = ((~g19074));
assign g11002 = ((~g7475))|((~g862));
assign g33707 = (g33174&g13346);
assign II14668 = ((~g7753));
assign gbuf148 = (g1083);
assign g20106 = ((~g17328));
assign g9534 = ((~g90));
assign II22028 = ((~g20204));
assign g14079 = ((~g11626))|((~g11763));
assign g7751 = ((~g1521));
assign g24270 = (g23165)|(g18614);
assign g32825 = ((~g30735));
assign II31581 = ((~g33164));
assign g25621 = (g24523)|(g18205);
assign g22714 = ((~g20436));
assign g29644 = (g28216&g19794);
assign g34842 = (g34762&g20168);
assign g32382 = ((~g31657));
assign g31141 = (g12224&g30038);
assign g25737 = (g25045)|(g22052);
assign g29793 = (g28237)|(g27247);
assign g32138 = ((~g31233));
assign gbuf86 = (g3649);
assign g33947 = (g32438)|(g33457);
assign g25020 = ((~g21377))|((~g23462));
assign g18472 = (g2413&g15224);
assign g24229 = (g896&g22594);
assign g29809 = (g28362&g23274);
assign g20216 = ((~II20487))|((~II20488));
assign g19580 = ((~g16164));
assign g10108 = ((~g120));
assign g19417 = ((~g17178));
assign g21689 = ((~II21250));
assign g25995 = ((~g24621))|((~g22853));
assign II26381 = ((~g26851));
assign II16028 = ((~g12381));
assign II14257 = ((~g8154))|((~g3133));
assign g7918 = (g1205&g1087);
assign II12300 = ((~g1157));
assign II16024 = ((~g11171));
assign g23939 = ((~g19074));
assign g8612 = ((~g2775));
assign g22526 = ((~g19801));
assign g24923 = (g23129&g20167);
assign g7543 = ((~II12033));
assign g34914 = ((~II33134));
assign g22539 = ((~g1030)&(~g19699));
assign g8290 = ((~g218));
assign g15021 = ((~g12711))|((~g10341));
assign g13480 = ((~g3017)&(~g11858));
assign g30399 = (g29757)|(g21758);
assign g28457 = ((~g7980)&(~g27602));
assign g16321 = ((~g4955))|((~g13996))|((~g12088));
assign g22071 = (g6251&g19210);
assign g19467 = (g16896)|(g14097);
assign II14170 = ((~g8389))|((~II14169));
assign g11291 = ((~g7526));
assign g34556 = (g34350&g20537);
assign g32954 = ((~g31376));
assign g14360 = ((~g12078)&(~g9484));
assign g18547 = (g121&g15277);
assign g16747 = ((~g14113));
assign g22098 = (g6459&g18833);
assign g24961 = (g23193&g20209);
assign g18599 = (g2955&g16349);
assign g25221 = ((~g23653));
assign g8655 = ((~g2787));
assign g27233 = (g25876)|(g24451);
assign g34206 = (g33834)|(g33836);
assign g7823 = ((~II12218))|((~II12219));
assign II13007 = ((~g65));
assign g8390 = ((~g3385));
assign g33816 = (g33234&g20096);
assign g16629 = ((~g13990));
assign II23336 = ((~g22721));
assign g31609 = ((~II29211));
assign g23658 = (g14687&g20852);
assign g22417 = (g7753&g9285&g21186);
assign g10890 = (g7858&g1105);
assign g20623 = ((~g17929));
assign g34077 = (g22957&g9104&g33736);
assign g34184 = (g33698&g24388);
assign II12203 = ((~g1094))|((~g1135));
assign g31921 = (g31508)|(g22046);
assign g8774 = ((~g781));
assign g9747 = ((~II13329));
assign g30825 = (g29814&g22332);
assign g12609 = ((~g7766)&(~g5863)&(~g5857));
assign II11785 = ((~g5703));
assign g26024 = (g2619&g25039);
assign g29073 = (g27163&g10290&g21012&II27409);
assign g26907 = (g26513)|(g24224);
assign g27159 = (g25814)|(g12953);
assign g13623 = (g482)|(g12527);
assign g14096 = ((~II16328));
assign g13216 = ((~g10939));
assign II24027 = (g3029&g3034&g8426);
assign g9415 = ((~g2169));
assign II20189 = ((~g1333))|((~II20187));
assign g33404 = (g32353&g21397);
assign g21283 = ((~g11291))|((~g17157));
assign g32221 = (g31140)|(g29634);
assign II12049 = ((~g781));
assign g23821 = ((~g19210));
assign g7259 = ((~g4375));
assign g26549 = ((~II25391));
assign II18344 = ((~g13003));
assign g14127 = ((~g11653))|((~g11435));
assign II20747 = ((~g17141));
assign g12497 = ((~g9780));
assign gbuf47 = (g5798);
assign g22864 = ((~g7780))|((~g21156));
assign g25571 = (II24694&II24695);
assign g9444 = ((~g5535));
assign II31271 = (g29385&g32846&g32847&g32848);
assign II14902 = ((~g9821));
assign g32886 = ((~g31327));
assign g19455 = ((~g15969))|((~g10841))|((~g7781));
assign g34756 = (g34680&g19618);
assign g24853 = (g21452)|(g24001);
assign g15615 = ((~II17181));
assign g27602 = (g23032&g26244&g26424&g24966);
assign g34033 = (g33821)|(g18708);
assign g12181 = ((~g9478));
assign II24415 = ((~g23751))|((~II24414));
assign g27387 = (g26488&g17499);
assign g21360 = ((~g11510))|((~g17157));
assign g20657 = ((~g17433));
assign g29278 = (g28626)|(g18740);
assign g24788 = (g11384&g23111);
assign g32997 = (g32269)|(g18378);
assign g13223 = ((~II15800));
assign g28837 = ((~g27800))|((~g7374))|((~g2197));
assign II21860 = ((~g19638));
assign g10190 = ((~g6044));
assign g26485 = (g24968&g10502);
assign g31222 = (g2643&g30113);
assign g17818 = ((~II18822));
assign g25077 = (g23297&g20536);
assign g17743 = ((~II18734));
assign g11148 = ((~g8052)&(~g9197)&(~g9174)&(~g9050));
assign g31261 = (g14754&g30259);
assign g33406 = (g32355&g21399);
assign g17573 = ((~g12911));
assign g25570 = (II24689&II24690);
assign g17655 = (g7897&g13342);
assign g22081 = (g6279&g19210);
assign II14204 = ((~g8508))|((~g3821));
assign II14653 = ((~g9417));
assign g32840 = ((~g30825));
assign g8626 = ((~g4040));
assign II25869 = ((~g25851));
assign g6802 = ((~g468));
assign g13116 = ((~g10935));
assign g18694 = (g4722&g16053);
assign g32815 = ((~g30937));
assign g25103 = (g4927&g22908);
assign g33785 = (g33100&g20550);
assign g22173 = ((~II21757));
assign g29959 = (g28953&g12823);
assign II22685 = ((~g21434))|((~II22683));
assign g34230 = (g33761&g22942);
assign g13255 = ((~g10632));
assign g19770 = ((~g17062));
assign II18259 = ((~g12946));
assign II18382 = ((~g13350));
assign g30989 = ((~g29672));
assign g30365 = (g30158)|(g18412);
assign g13277 = (g3195&g11432);
assign g20699 = ((~g17873));
assign g10566 = ((~g7315))|((~g7356));
assign g28715 = (g27480)|(g16700);
assign g33972 = (g33941)|(g18335);
assign g28793 = ((~g27800))|((~g7328))|((~g2153));
assign g34849 = (g34842)|(g18154);
assign II15129 = ((~g9914))|((~II15128));
assign g14888 = (g10776)|(g8703);
assign II18107 = ((~g4019));
assign g14207 = (g8639&g11793);
assign g18825 = (g6736&g15680);
assign II32970 = ((~g34716));
assign g29667 = (g2671&g29157);
assign g29235 = (g28110)|(g18260);
assign g25050 = (g13056&g22312);
assign g20187 = (g16202)|(g13491);
assign g8236 = ((~g4812));
assign g14184 = ((~g12381));
assign g27875 = ((~g9875)&(~g25821));
assign g33000 = (g32270)|(g18403);
assign g30309 = ((~g28959));
assign g22046 = (g6073&g21611);
assign g29205 = (g24117&II27523&II27524);
assign g14750 = ((~g6633))|((~g12137))|((~g6715))|((~g12721));
assign g10632 = (g7475&g7441&g890);
assign g33573 = (g33343)|(g18415);
assign g12239 = ((~II15106))|((~II15107));
assign II32455 = ((~g34242));
assign g29292 = (g28556)|(g18776);
assign g19435 = ((~g16449));
assign g7438 = ((~g5983));
assign II24048 = (g3034&g3040&g8426);
assign g10613 = ((~g10233));
assign g9433 = ((~g5148));
assign g23873 = (g21222&g10815);
assign II17420 = ((~g13394));
assign g26971 = (g26325)|(g24333);
assign II14119 = ((~g7824));
assign g28490 = (g27262)|(g16185);
assign g17533 = ((~II18482));
assign g31494 = (g29792&g23435);
assign g17872 = ((~g6617))|((~g14602))|((~g6711))|((~g12721));
assign g17781 = (g6772&g11592&g6789&II18785);
assign g34284 = (g34046&g19351);
assign g20703 = ((~g15373));
assign g11754 = ((~g8229));
assign g8359 = ((~II12545))|((~II12546));
assign g24355 = (g23799)|(g18824);
assign g20441 = ((~g17873));
assign g14838 = ((~g12492))|((~g12405));
assign g26096 = (g9733&g25268);
assign g23127 = ((~g21163));
assign g32639 = ((~g31070));
assign II18662 = ((~g6322));
assign g33613 = (g33248)|(g18649);
assign g34524 = (g9083&g34359);
assign g22491 = ((~g1361)&(~g19720));
assign g27982 = ((~g7212)&(~g25856));
assign g27991 = ((~g25852));
assign g23525 = ((~g21562));
assign g16585 = ((~g14075));
assign g19263 = ((~II19799));
assign g31476 = ((~g4709)&(~g29697));
assign g21901 = (g21251)|(g15115);
assign g12878 = ((~g10386));
assign g23539 = ((~g21070));
assign II29894 = ((~g31771));
assign g33665 = ((~II31500));
assign g11309 = ((~g8587)&(~g8728));
assign g20055 = ((~g11269))|((~g17794));
assign II30728 = (g32345)|(g32350)|(g32056)|(g32018);
assign g30034 = (g29077&g10541);
assign g33499 = (g32737&II31191&II31192);
assign g15703 = (g452&g13437);
assign II12159 = ((~g608));
assign g21459 = ((~g17814))|((~g14854))|((~g17605))|((~g17581));
assign g14984 = ((~g7812))|((~g12680));
assign g11891 = ((~g812)&(~g9166));
assign g27518 = (g26488&g17709);
assign II23306 = ((~g21673));
assign g25755 = (g25192)|(g22102);
assign g31869 = (g30592)|(g18221);
assign g24436 = (g3125&g23067);
assign g34661 = (g34575&g18907);
assign g30554 = (g30216)|(g22125);
assign g8439 = ((~g3129));
assign g25044 = ((~g23675));
assign g28955 = ((~g27837))|((~g1936))|((~g7362));
assign II13968 = ((~g7697));
assign g30472 = (g30186)|(g21943);
assign g28479 = ((~g27654));
assign II25882 = ((~g25776));
assign g24728 = (g16513&g23017);
assign g23899 = ((~g19277));
assign g11984 = ((~g9186));
assign g13772 = ((~g3990)&(~g11702));
assign g8195 = ((~g1783));
assign g29802 = (g28243)|(g22871);
assign g10121 = ((~g2327));
assign g16814 = ((~g14058));
assign g18581 = (g2912&g16349);
assign II31600 = (g31009&g8400&g7809);
assign II11632 = ((~g16));
assign g34368 = (g26274)|(g34135);
assign g16669 = (g5611&g14993);
assign g21963 = (g5436&g21514);
assign g26269 = ((~II25243))|((~II25244));
assign g9966 = ((~II13498))|((~II13499));
assign II12219 = ((~g1478))|((~II12217));
assign g24975 = ((~g21388))|((~g23363));
assign g32254 = (g31247&g20379);
assign g9864 = ((~II13424));
assign g23629 = ((~g21514));
assign g34010 = (g33872)|(g18478);
assign g12492 = ((~g7704)&(~g5170)&(~g5164));
assign g32408 = (g31541)|(g30073);
assign g29218 = ((~II27570));
assign gbuf97 = (g4000);
assign g21856 = (g3929&g21070);
assign g17470 = ((~g14454));
assign g24655 = ((~g23067));
assign g6875 = ((~II11697));
assign g34276 = ((~g34058));
assign g24309 = (g4480&g22228);
assign g26294 = (g4245&g25230);
assign II14766 = ((~g5821))|((~II14764));
assign g26812 = ((~g25439));
assign II31101 = (g30735&g31813&g32601&g32602);
assign g23409 = ((~g21514));
assign g23402 = ((~g20875));
assign g30389 = (g29969)|(g18554);
assign g30093 = (g28467)|(g11397);
assign g18611 = (g15090&g17200);
assign g30221 = (g28700&g23893);
assign g33480 = (g32600&II31096&II31097);
assign g24932 = ((~g19886))|((~g23172));
assign g18806 = (g6381&g15656);
assign g17635 = ((~g3542))|((~g13730))|((~g3654))|((~g8542));
assign g32402 = (g4888&g30990);
assign g20852 = ((~g15595));
assign g25307 = ((~g22763));
assign g29863 = ((~g28410));
assign g8466 = ((~g1514));
assign g23148 = (g19128&g9104);
assign g32548 = ((~g30673));
assign g18108 = (g433&g17015);
assign g32694 = ((~g31376));
assign g24344 = (g22145)|(g18787);
assign g31859 = ((~g29385));
assign g19589 = ((~g15969))|((~g10841))|((~g10884));
assign g34224 = (g33736&g22670);
assign II15193 = ((~g9935))|((~g6005));
assign g12767 = ((~g4467))|((~g6961));
assign g19872 = ((~g17015));
assign g34681 = (g34491&g19438);
assign II17552 = (g13156&g11450&g11498);
assign g14813 = ((~g7766))|((~g12824));
assign g28676 = (g27570&g20632);
assign g29975 = (g28986&g10420);
assign II20318 = ((~g16920));
assign g18405 = (g2040&g15373);
assign g23460 = ((~g21611));
assign II13759 = ((~g6754));
assign g26725 = (g24457)|(g10719);
assign g7232 = ((~g4411));
assign II22692 = ((~g21308));
assign g33278 = (g32139)|(g29572);
assign g27569 = (g26124)|(g24721);
assign g33273 = (g32122)|(g29553);
assign g30490 = (g30167)|(g21986);
assign g18707 = (g15134&g16782);
assign g9817 = ((~II13374));
assign g27135 = (g24387)|(g25803);
assign g18363 = (g1840&g17955);
assign g34646 = (g34557)|(g18803);
assign g28583 = (g12009&g27112);
assign g30402 = (g29871)|(g21761);
assign g31376 = (g24952&g29814);
assign g33607 = (g33091)|(g18526);
assign g11563 = ((~g8059)&(~g8011));
assign II33285 = ((~g34988));
assign g14872 = ((~g6736)&(~g12364));
assign g32304 = (g31284&g20564);
assign g18789 = (g6035&g15634);
assign g24769 = (g19619&g23058);
assign II31748 = ((~g33228));
assign g31184 = (g1950&g30085);
assign g8812 = ((~II12805));
assign g14981 = ((~g12785))|((~g12632));
assign II28832 = ((~g30301));
assign g18396 = (g2008&g15373);
assign g13028 = ((~II15650));
assign g21050 = ((~g17873));
assign II31973 = ((~g33641))|((~II31972));
assign g28712 = (g27590&g20708);
assign g17723 = ((~g6597))|((~g14556))|((~g6668))|((~g12721));
assign g26967 = (g26350)|(g24319);
assign g28554 = (g27426&g20372);
assign g23993 = ((~g19277));
assign g20511 = ((~g17929));
assign g18534 = (g2735&g15277);
assign g26994 = (g23032&g26226&g26424&g25557);
assign g12705 = ((~g7051));
assign g30506 = (g30179)|(g22027);
assign g24500 = (g24011)|(g21605);
assign g13301 = ((~g10862));
assign g28629 = (g27371)|(g16532);
assign g7619 = ((~g1296));
assign g30412 = (g29885)|(g21771);
assign g30466 = (g30174)|(g21937);
assign g14977 = (g10776)|(g8703);
assign g27344 = ((~g8390)&(~g26636));
assign g18296 = (g1495&g16449);
assign g21345 = ((~g11429))|((~g17157));
assign g30107 = (g28560&g20909);
assign g33068 = (g31994)|(g22112);
assign II26050 = ((~g25997))|((~II26049));
assign g12040 = ((~II14902));
assign g25583 = (g21666)|(g24153);
assign g29179 = ((~g9311)&(~g28010)&(~g7738));
assign g26857 = (g25062&g25049);
assign g30380 = (g30161)|(g18492);
assign g28539 = (g27187&g12762);
assign g30343 = (g29344)|(g18278);
assign g17146 = (g5965&g14895);
assign II15264 = ((~g2273))|((~II15262));
assign g19576 = (g17138)|(g14202);
assign g29315 = (g29188&g7051&g5990);
assign g25609 = (g24915)|(g18126);
assign g29925 = ((~g28820));
assign g34028 = (g33720)|(g18684);
assign g26229 = (g1724&g25275);
assign II15190 = ((~g6005));
assign II20035 = ((~g15706));
assign g22066 = (g6209&g19210);
assign g12941 = ((~g7167))|((~g10537));
assign g26077 = (g9607&g25233);
assign g10399 = ((~g7017));
assign g21940 = (g5228&g18997);
assign II27567 = ((~g28181));
assign g16614 = (g5945&g14933);
assign g22843 = (g9429&g20272);
assign g23380 = ((~g20619));
assign g11957 = ((~g8205))|((~g8259));
assign g21715 = (g160&g20283);
assign g7780 = ((~g2878));
assign g33910 = (g33134&g7836);
assign g26673 = (g24433)|(g10674);
assign g17423 = ((~II18360));
assign g34279 = (g34231&g19208);
assign g25097 = ((~g22342));
assign g27690 = (g25784&g23607);
assign g29537 = (g28976&g22472);
assign g33710 = (g14037&g33246);
assign g27961 = ((~g26816));
assign g15831 = ((~g13385));
assign g12593 = ((~g9234)&(~g5164));
assign g26329 = (g8526)|(g24609);
assign g21748 = (g15089&g20785);
assign g25866 = (g3853&g24648);
assign g31212 = (g20028&g29669);
assign g18384 = (g1945&g15171);
assign g27663 = (g26323)|(g24820);
assign g21413 = ((~g15585));
assign g28469 = ((~g3171)&(~g27602));
assign g24949 = (g23796&g20751);
assign g8505 = ((~g3480));
assign g14149 = ((~g12381));
assign g32047 = (g27248&g31070);
assign g29141 = ((~g9374)&(~g27999));
assign g24641 = (g22151)|(g22159);
assign g34928 = ((~II33176));
assign g21948 = (g5260&g18997);
assign g32516 = ((~g31070));
assign g13566 = (g7092&g12358);
assign g18192 = (g817&g17821);
assign g25287 = ((~g22228));
assign g34401 = (g34199&g21383);
assign g30510 = (g30263)|(g22031);
assign g33732 = (g33104)|(g32011);
assign g17757 = ((~g5909))|((~g14549))|((~g6005))|((~g12614));
assign g24184 = ((~II23396));
assign g20631 = ((~g15171));
assign g16204 = (g6537&g14348);
assign g17761 = ((~g6291))|((~g14529))|((~g6358))|((~g12423));
assign II14482 = ((~g655))|((~II14480));
assign g18428 = (g2169&g18008);
assign g11527 = ((~g8165)&(~g8114));
assign II15617 = ((~g12037));
assign g32630 = ((~g30735));
assign g32659 = ((~g30735));
assign II16357 = ((~g884));
assign g16737 = (g6645&g15042);
assign g29196 = ((~g27059));
assign g18782 = (g5835&g18065);
assign g27380 = ((~II26071))|((~II26072));
assign g13974 = (g6243&g12578);
assign g14854 = ((~g5555))|((~g12093))|((~g5654))|((~g12563));
assign g24918 = ((~g136))|((~g23088));
assign g22330 = ((~g19801));
assign g22181 = ((~g19277));
assign II24008 = ((~g22182));
assign g32184 = (g30611&g25249);
assign g12155 = ((~g7753))|((~g7717));
assign g7532 = ((~g1157));
assign g17615 = ((~II18574));
assign g9413 = ((~g1744));
assign g14383 = ((~II16535));
assign g20533 = ((~g17271));
assign g25902 = (g24398&g19373);
assign g16967 = ((~II18125));
assign g31224 = (g30280&g23932);
assign g9661 = ((~g3661));
assign g22223 = ((~g19210));
assign g12880 = ((~g10387));
assign g11413 = ((~g9100));
assign g23543 = ((~g21514));
assign g23714 = ((~g20751));
assign g28216 = (g27036)|(g27043);
assign g21729 = (g3021&g20330);
assign g20566 = ((~g15224));
assign g26234 = (g2657&g25514);
assign g17429 = ((~II18370));
assign g7394 = ((~g5637));
assign g26652 = (g10799&g24426);
assign g11973 = ((~g8365))|((~g2051));
assign g14451 = ((~II16606));
assign g34883 = ((~g34852));
assign II12577 = ((~g1227));
assign g21556 = ((~g15669));
assign g33597 = (g33344)|(g18495);
assign g32191 = (g27593&g31376);
assign g28622 = (g27360)|(g16519);
assign g26933 = (g26808)|(g18551);
assign g24400 = (g3466&g23112);
assign g9995 = ((~g6035));
assign II16438 = ((~g11165));
assign g27431 = (g24582)|(g25977);
assign g21053 = ((~g15373));
assign g25027 = ((~II24191));
assign g30390 = (g29985)|(g18555);
assign II13892 = ((~g1576));
assign g28853 = ((~g27742))|((~g1636))|((~g7252));
assign g17783 = (g7851&g13110);
assign g18125 = (g15053&g16886);
assign II31985 = ((~g33648))|((~II31983));
assign g19919 = ((~g16987)&(~g11205));
assign g26365 = (g25504)|(g25141);
assign g11934 = ((~g8139))|((~g8187));
assign g14238 = ((~g10823));
assign g18588 = (g2970&g16349);
assign g27983 = ((~g26725));
assign g23532 = (g19400&g11852);
assign g14540 = ((~g12287)&(~g9834));
assign g34257 = (g34226)|(g18674);
assign g12538 = ((~II15334))|((~II15335));
assign g20668 = ((~g15426));
assign g23683 = ((~II22816));
assign g32617 = ((~g30825));
assign g13189 = ((~g10762));
assign g9542 = ((~g2173));
assign g33075 = ((~g31997)&(~g7163));
assign g12047 = ((~g9591));
assign g24049 = ((~g20014));
assign g8388 = ((~g3010));
assign g25121 = ((~g22432));
assign g33685 = (g32396)|(g33423);
assign gbuf101 = (g3794);
assign g24666 = (g11753&g22975);
assign g13530 = ((~g12641));
assign II31152 = (g32675&g32676&g32677&g32678);
assign g23448 = ((~g21611));
assign g34416 = (g34191)|(g25159);
assign g25237 = ((~g6434))|((~g23711));
assign g8839 = ((~II12819));
assign II18888 = ((~g16644));
assign g21979 = (g5559&g19074);
assign g32558 = ((~g30735));
assign g21832 = (g3787&g20453);
assign g34973 = ((~II33235));
assign g25618 = (g25491)|(g18192);
assign g32210 = (g31123)|(g29600);
assign II17495 = ((~g13378))|((~II17494));
assign g11958 = ((~g9543)&(~g7327));
assign g24710 = (g22679&g19771);
assign II15831 = ((~g10416));
assign g7502 = ((~II11992));
assign g11949 = ((~II14773));
assign g29986 = (g28468&g23473);
assign g8714 = ((~g4859));
assign g27097 = (g25867&g22526);
assign g33017 = (g32292)|(g18510);
assign g13765 = ((~g8531)&(~g11615));
assign g11435 = ((~g8107)&(~g3171));
assign g34408 = ((~g34144));
assign g24293 = (g4438&g22550);
assign g21340 = ((~II21074));
assign g31480 = (g1644&g30296);
assign g18117 = (g464&g17015);
assign g21953 = (g5377&g21514);
assign g18325 = (g1624&g17873);
assign g28082 = (g27369)|(g24315);
assign g27411 = (g26549&g17528);
assign g11404 = ((~g7596));
assign II22931 = ((~g21228))|((~II22929));
assign g14564 = ((~II16679));
assign g25665 = (g24708)|(g21790);
assign g22538 = (g14035&g20248);
assign g34970 = (g34868)|(g34961);
assign g17625 = ((~g14541)&(~g12123));
assign g31312 = (g30136&g27858);
assign g12075 = ((~II14935));
assign II18086 = ((~g13856));
assign g20060 = ((~g16540));
assign g26340 = ((~g24953));
assign g28166 = ((~II26687));
assign g29280 = (g28530)|(g18742);
assign g13529 = ((~g11590))|((~g11544))|((~g11492))|((~g11446));
assign g15755 = ((~g13134));
assign g8895 = ((~g599));
assign g10520 = ((~g7195))|((~g7115));
assign g33063 = (g31988)|(g22066);
assign gbuf99 = (g4023);
assign g15063 = ((~g6818)&(~g13394));
assign g28244 = (g27926&g26715);
assign g33293 = (g32151)|(g29602);
assign g19354 = (g471&g16235);
assign g22698 = ((~II22009));
assign g26941 = ((~II25689));
assign g23922 = ((~g18997));
assign g17716 = ((~g5957))|((~g14497))|((~g6027))|((~g12614));
assign g25766 = ((~g24439));
assign g24263 = (g23497)|(g18529);
assign g27089 = ((~g26703));
assign g21887 = (g15101&g19801);
assign g11999 = ((~g9654)&(~g7423));
assign g32689 = ((~g30825));
assign g26025 = ((~g22405))|((~g24631));
assign g16308 = ((~II17636));
assign g27312 = (g12019&g26700);
assign g23309 = ((~g6905))|((~g21024));
assign II22096 = ((~g19890));
assign g20070 = ((~g16173));
assign g26681 = ((~g25396));
assign g18272 = (g1283&g16031);
assign g21377 = ((~g11560))|((~g17157));
assign g22985 = ((~g20330));
assign g23108 = ((~g16424)&(~g19932));
assign g7374 = ((~g2227));
assign g26896 = (g26341)|(g18171);
assign g21293 = ((~II21036));
assign g17366 = ((~g14454));
assign g19931 = ((~g17200));
assign g28574 = (g27324)|(g26270);
assign g28334 = (g27131)|(g15817);
assign g24779 = ((~g3736)&(~g23167));
assign g13923 = ((~g11692))|((~g11527));
assign II14249 = ((~g8091))|((~II14247));
assign g18633 = (g6905&g17226);
assign g15807 = (g3570&g13898);
assign g34394 = (g34190&g21305);
assign g20069 = (g16312&g9051&g9011&g8955);
assign g32680 = ((~g31376));
assign g18221 = (g1018&g16100);
assign g23749 = ((~g18997));
assign g29325 = (g28813)|(g27820);
assign II24439 = ((~g23771))|((~II24438));
assign g25650 = (g24663)|(g21743);
assign g6854 = ((~g2685));
assign g31806 = ((~g29385));
assign g32157 = (g31646&g30021);
assign g22669 = (g7763)|(g19525);
assign g22004 = (g5742&g21562);
assign g14655 = ((~g4743))|((~g11755));
assign g32145 = (g31609&g29977);
assign g18618 = (g3457&g17062);
assign g28748 = (g27522)|(g16763);
assign g13049 = ((~II15677));
assign g30565 = ((~II28832));
assign g30089 = (g28538&g20709);
assign g25505 = ((~g22228));
assign g11380 = (g8583)|(g8530);
assign g7153 = ((~g5373));
assign g34142 = ((~II32089));
assign g19546 = ((~g15969))|((~g10841))|((~g10884));
assign g34088 = (g33736&g9104&g18957);
assign g26510 = ((~II25369));
assign g24590 = (g6154&g23413);
assign g24676 = (g2748&g23782);
assign g21904 = ((~II21483));
assign g15152 = ((~g13745)&(~g12896));
assign II17852 = ((~g3625));
assign g18667 = (g4601&g17367);
assign g30315 = (g29182&g7028&g5644);
assign g23847 = ((~g19210));
assign g12405 = ((~g9374)&(~g5180));
assign g11967 = (g311&g7802);
assign II30124 = (g31070)|(g31154)|(g30614)|(g30673);
assign g6927 = ((~g3845));
assign g10359 = ((~g6830));
assign g22144 = ((~g18997));
assign g25144 = ((~g5046)&(~g23623));
assign g12314 = ((~g10053)&(~g10207));
assign g15756 = ((~g13315));
assign II18620 = (g13156&g11450&g11498);
assign II21042 = ((~g15824));
assign II29936 = ((~g30606));
assign g15116 = (g4297&g14454);
assign g19539 = ((~g16129));
assign g25743 = (g25110)|(g22058);
assign gbuf67 = (g6719);
assign II15041 = ((~g9752))|((~g1834));
assign g6850 = ((~g2704));
assign g34634 = (g34483)|(g18691);
assign g24460 = (g10967)|(g22450);
assign g7150 = ((~g5016))|((~g5062));
assign g32627 = ((~g30673));
assign g13742 = ((~g11780))|((~g11283));
assign g27365 = ((~II26050))|((~II26051));
assign g32501 = ((~g30825));
assign II31619 = ((~g33212));
assign g29759 = (g28308&g23226);
assign g12831 = ((~g9569));
assign gbuf11 = (g5005);
assign g24104 = ((~g19890));
assign g33461 = (g32463&II31001&II31002);
assign g32310 = (g27577&g31376);
assign g14506 = (g1430&g10755);
assign g18753 = (g15148&g15595);
assign g27215 = (g26055&g16724);
assign g7361 = ((~g1874));
assign g21817 = (g3606&g20924);
assign g20276 = (g16243)|(g13566);
assign g18491 = (g2518&g15426);
assign g19771 = ((~g17096));
assign g33054 = (g31975)|(g21975);
assign II17956 = ((~g14562));
assign g17742 = ((~g14971));
assign g9153 = ((~II12991));
assign g22342 = (g9354&g9285&g21287);
assign g29689 = ((~II27954));
assign g11770 = ((~II14619));
assign g17384 = ((~II18323));
assign g24864 = (g11201&g22305);
assign g12148 = ((~g2060))|((~g8310));
assign g29382 = (g26424&g22763&g28172);
assign g23046 = ((~g20283));
assign g20622 = ((~g15595));
assign g29602 = (g2020&g28962);
assign g22935 = ((~g20283));
assign g12415 = ((~g7496))|((~g5976));
assign g21922 = (g5112&g21468);
assign g19428 = ((~g16090));
assign g29860 = (g28389&g23312);
assign g24425 = ((~g22722));
assign g27017 = ((~g25895));
assign g25678 = (g24709)|(g21835);
assign g29994 = ((~g29049));
assign g24638 = (g22763&g19690);
assign II14508 = ((~g370))|((~g8721));
assign g32632 = ((~g31070));
assign g26259 = (g24430&g25232);
assign II17118 = ((~g14363));
assign g32980 = (g32254)|(g18198);
assign g29905 = ((~g28783));
assign g30137 = (g28594&g21181);
assign g16259 = ((~g4743))|((~g13908))|((~g12054));
assign g22061 = (g6065&g21611);
assign g26895 = (g26783)|(g18148);
assign g19660 = (g12001&g16968);
assign g29587 = (g2181&g28935);
assign g14122 = ((~g8895)&(~g12259));
assign g34713 = ((~II32871));
assign g33552 = (g33400)|(g18343);
assign g16211 = (g5445&g14215);
assign gbuf31 = (g5654);
assign g19914 = (g2815&g15853);
assign g16644 = ((~II17842));
assign g23153 = (g19521)|(g15876);
assign g14739 = ((~g5929))|((~g12067))|((~g5983))|((~g12351));
assign g34486 = (g34412&g18953);
assign g12760 = ((~g10272));
assign II16747 = ((~g12729));
assign g20771 = ((~g15171));
assign g27742 = (g17292)|(g26673);
assign g31487 = ((~II29149));
assign g12093 = ((~g9924)&(~g7028));
assign g18107 = (g429&g17015);
assign g25915 = (g24926&g9602);
assign g20050 = ((~II20321));
assign g28636 = (g27376)|(g16538);
assign II30262 = (g31672)|(g31710)|(g31021)|(g30937);
assign g34135 = (g33926&g23802);
assign g9282 = ((~g723));
assign g28279 = (g27087)|(g25909);
assign g8786 = ((~II12770));
assign g12417 = ((~g7175));
assign g28536 = (g27293)|(g26205);
assign g27289 = (g25925)|(g25927);
assign g24875 = ((~g8725)&(~g23850)&(~g11083));
assign g18746 = (g5134&g17847);
assign g10261 = ((~g4555));
assign g27355 = ((~g8443)&(~g26657));
assign g18526 = (g2555&g15509);
assign g19564 = (g17175&g13976);
assign g29548 = (g1798&g28575);
assign g24688 = (g22681&g22663);
assign g29966 = (g23617&g28970);
assign g18184 = (g785&g17328);
assign g9083 = ((~g626));
assign g14169 = ((~g12381));
assign g21422 = ((~g15373));
assign g18660 = ((~II19484));
assign g33016 = (g32284)|(g18509);
assign g24415 = (g4760&g22869);
assign g18208 = (g930&g15938);
assign g32477 = ((~g31566));
assign g15108 = (g4264&g14454);
assign g31788 = (g21352&g29385);
assign g18977 = ((~g16100));
assign g27677 = (g13021&g25888);
assign g29329 = (g7995&g28353);
assign g10899 = ((~g4064)&(~g8451));
assign g29840 = (g2153&g29056);
assign g19274 = (g17753)|(g14791);
assign II31127 = (g32638&g32639&g32640&g32641);
assign g32906 = ((~g31021));
assign g25980 = (g1926&g25006);
assign II32806 = ((~g34585));
assign g13873 = ((~g11566))|((~g11729));
assign g11914 = ((~g8187))|((~g1648));
assign g19500 = (g504&g16712);
assign g20502 = ((~g15373));
assign g33560 = (g33404)|(g18369);
assign II22153 = ((~g20014));
assign II22124 = ((~g21300));
assign g10922 = ((~g7650)&(~g4057));
assign g7404 = (g933)|(g939);
assign gbuf112 = (g4207);
assign g19683 = ((~g16931));
assign g23300 = ((~g20283));
assign g28669 = ((~g27705));
assign g15082 = (g2697&g12983);
assign II22944 = ((~g9492))|((~g19620));
assign g13055 = ((~II15682));
assign g23421 = ((~g21562));
assign g33435 = ((~II30959));
assign g9891 = ((~g6173));
assign g33546 = (g33402)|(g18327);
assign g15614 = ((~g14914));
assign g31066 = (g29483&g22865);
assign II21189 = ((~g17475));
assign g29529 = (g28303)|(g28293)|(g28283)|(g28267);
assign g17507 = ((~g15030));
assign g29535 = (g2303&g28871);
assign II17488 = ((~g13394));
assign g10014 = ((~g6439));
assign g22544 = ((~g19589));
assign g8476 = (g1399)|(g1459)|(II12611);
assign g34474 = (g20083&g34326);
assign g17393 = ((~g9386)&(~g14379));
assign g18471 = (g2407&g15224);
assign II26799 = ((~g27660));
assign g29607 = (g28509&g14208);
assign g29871 = (g28400&g23332);
assign g26484 = (g24946&g8841);
assign g19751 = ((~g16044));
assign g31007 = (g29364)|(g28159);
assign g31822 = ((~g29385));
assign g30430 = (g29859)|(g21814);
assign g11397 = (g5360&g7139);
assign g23505 = ((~g21514));
assign g31880 = (g31280)|(g21774);
assign g13464 = ((~g10831))|((~g4793))|((~g4776));
assign g16580 = ((~II17754));
assign g13632 = (g10232&g12228);
assign g31986 = (g31766&g22197);
assign g20738 = ((~g15483));
assign g9591 = ((~g1926))|((~g1894));
assign g19998 = ((~g15915));
assign g18576 = (g2868&g16349);
assign g11591 = ((~II14531))|((~II14532));
assign g19688 = ((~g16777));
assign g20679 = ((~g15634));
assign g12863 = ((~g10371));
assign g24055 = ((~g19968));
assign II15727 = ((~g10981));
assign g13600 = ((~g3021))|((~g11039));
assign g24644 = (g11714&g22903);
assign g32328 = (g5853&g31554);
assign g28962 = ((~g27886))|((~g2040))|((~g7369));
assign II18912 = ((~g15050));
assign g13881 = ((~II16181));
assign g25002 = ((~g19474))|((~g23154));
assign g29264 = (g28248)|(g18618);
assign II13206 = ((~g5448));
assign g16770 = ((~g3263))|((~g13765))|((~g3274))|((~g8481));
assign g34636 = (g34476)|(g18693);
assign g30919 = (g29898&g23286);
assign g32783 = ((~g30825));
assign g8406 = ((~g232));
assign g21789 = (g3451&g20391);
assign g34116 = (g33933&g25140);
assign g18874 = ((~g15938));
assign II25028 = ((~g24484));
assign g14662 = ((~II16762));
assign g32413 = (g31121&g19518);
assign g34515 = (g34288&g19491);
assign II22302 = ((~g19353));
assign g23958 = (g9104&g19200);
assign g10289 = ((~g1319));
assign g12464 = ((~g10169))|((~g7087))|((~g10191));
assign II13401 = ((~g2246))|((~g2250));
assign g33918 = ((~II31782));
assign g15744 = ((~g6641))|((~g14602))|((~g6719))|((~g10061));
assign g32889 = ((~g31376));
assign g24507 = (g22304&g19429);
assign g18952 = ((~g16053));
assign g15784 = (g3235&g13977);
assign g22182 = ((~II21766));
assign g30539 = (g30267)|(g22085);
assign g20145 = ((~g17533));
assign g25184 = ((~g22763));
assign g13820 = (g11184)|(g9187)|(g12527);
assign g31862 = ((~II29444));
assign g17411 = ((~g14454));
assign g11793 = ((~II14633));
assign g31912 = (g31752)|(g21998);
assign g34987 = ((~II33261));
assign II12783 = (g4204)|(g4207)|(g4210)|(g4180);
assign g33253 = (g32103)|(g29511);
assign g12996 = ((~g11823));
assign g25179 = (g16928&g23611);
assign II22131 = ((~g19984));
assign g24021 = ((~g20841));
assign g32873 = ((~g30614));
assign g31319 = (g29612)|(g28324);
assign g30929 = ((~g29803)&(~g29835));
assign g31517 = (g29849&g23482);
assign II31281 = (g30735&g31845&g32861&g32862);
assign g27717 = ((~g9492)&(~g26745));
assign II16120 = ((~g11868));
assign g18832 = ((~g15634));
assign g17580 = ((~II18509));
assign g28265 = (g11367&g27989);
assign g9823 = ((~II13383))|((~II13384));
assign g8092 = ((~g1589));
assign g30071 = (g29184&g12975);
assign g9762 = ((~g2495)&(~g2421));
assign g23972 = ((~g7097))|((~g20751));
assign g7898 = ((~g4991));
assign g22307 = (g20027&g21163);
assign g10884 = ((~g7650)&(~g8451));
assign g20554 = ((~g15348));
assign g25108 = (g23345&g20576);
assign g21996 = (g5615&g19074);
assign g30197 = (g28661&g23859);
assign g18511 = (g2599&g15509);
assign g10556 = ((~g7971))|((~g8133));
assign g10815 = ((~g9917));
assign g30935 = (g8808&g29745);
assign g24835 = (g8720&g23233);
assign g8958 = ((~g3881)&(~g3873));
assign g13975 = ((~g11048));
assign g32374 = (g29895)|(g31323);
assign g14036 = ((~g8725)&(~g11083));
assign g33722 = (g33175&g19445);
assign g16512 = ((~g14015));
assign g24212 = (g23280)|(g18155);
assign g23949 = ((~g7074))|((~g21012));
assign g31479 = ((~II29139));
assign g21397 = ((~g15171));
assign g14215 = ((~g12198));
assign g18733 = (g15141&g16877);
assign g13958 = ((~g3610))|((~g11238))|((~g3618))|((~g11389));
assign g9905 = ((~g802));
assign g13729 = ((~g10951));
assign g14107 = ((~g11571))|((~g11527));
assign g13120 = ((~g10632));
assign II19843 = ((~g16594));
assign g9805 = ((~g5485));
assign g34775 = ((~II32967));
assign II24616 = (g6082&g6088&g9946);
assign II28128 = ((~g28314));
assign g19767 = (g16810&g14203);
assign g34199 = (g33820)|(g33828);
assign g31020 = (g29375)|(g28164);
assign g23024 = ((~g7936)&(~g19407));
assign g30455 = (g30041)|(g21864);
assign g18246 = (g1199&g16431);
assign g18805 = (g6377&g15656);
assign g33925 = ((~g33394))|((~g4462))|((~g4467));
assign g11019 = (g5092&g9036);
assign g18586 = (g2886&g16349);
assign g27113 = (g25997&g16522);
assign g21835 = (g3802&g20453);
assign g29837 = (g28369&g20144);
assign g11225 = ((~g3990)&(~g6928));
assign II13317 = ((~g6144));
assign g29131 = ((~g27907))|((~g9762));
assign g21037 = ((~II20913));
assign g29899 = (g28428&g23375);
assign II18810 = ((~g13716));
assign g28543 = (g27735&g15628);
assign g20324 = ((~g17955));
assign g7948 = (g1548&g1430);
assign g30461 = (g30219)|(g21932);
assign g25954 = ((~g7750)&(~g24591));
assign gbuf151 = (g1157);
assign g8763 = ((~II12749));
assign g11826 = ((~II14650));
assign g18559 = (g12856&g15277);
assign g29892 = (g28300)|(g26120);
assign g18098 = ((~II18900));
assign g19780 = ((~g16449));
assign g30064 = (g28517&g20630);
assign g22992 = (g1227&g19765);
assign g24457 = (g10902)|(g22400);
assign g10372 = ((~g6900));
assign g27096 = (g26026&g16475);
assign II13847 = ((~g7266));
assign g16236 = ((~g13573))|((~g13554))|((~g13058));
assign g6971 = ((~II11737));
assign g18620 = (g3470&g17062);
assign g22125 = (g6617&g19277);
assign g6868 = ((~II11688));
assign g26758 = ((~g25389));
assign g16693 = ((~II17901));
assign g34560 = (g34366&g17366);
assign g32593 = ((~g31542));
assign g15881 = (g3582&g13983);
assign g17772 = ((~g14297));
assign g28121 = ((~g27093));
assign g8606 = ((~g4653));
assign g23031 = ((~g19801));
assign g16617 = (g6287&g14940);
assign g8441 = ((~g3361));
assign g18563 = (g2890&g16349);
assign g32106 = (g31601&g29911);
assign g19712 = ((~g17096));
assign g9654 = ((~g2485))|((~g2453));
assign g9752 = ((~g1840));
assign II19762 = ((~g15732));
assign g22633 = (g19359&g19479);
assign g14362 = ((~g12080)&(~g9338));
assign g25326 = ((~g22228));
assign g9557 = ((~g5499));
assign II17999 = ((~g4012));
assign II12887 = ((~g4216));
assign g34877 = ((~II33103));
assign g25831 = (g3151&g24623);
assign g10620 = ((~g10233));
assign g19693 = (g6181&g17087);
assign g17155 = ((~II18205));
assign g13006 = (g12284)|(g10034);
assign g26841 = ((~g24893));
assign g7527 = ((~II12016));
assign g34730 = (g34658)|(g18271);
assign g18237 = (g1146&g16326);
assign g20913 = ((~g15373));
assign g31937 = ((~g30991));
assign g23483 = ((~g18833));
assign II27503 = (g19890&g24075&g24076&g28032);
assign g18826 = (g7097&g15680);
assign II25562 = ((~g25250));
assign g24967 = (g23197&g20213);
assign g25971 = (g1917&g24992);
assign g31758 = (g30115&g23945);
assign g24200 = (g22831)|(g18103);
assign g30546 = (g30277)|(g22117);
assign g16640 = ((~II17834));
assign II19789 = ((~g17793));
assign g33543 = (g33106)|(g18281);
assign g33872 = (g33282&g20548);
assign g24627 = (g22763&g19679);
assign g7308 = ((~g1668));
assign g25340 = ((~g22763));
assign g32488 = ((~g31194));
assign g19960 = ((~g17433));
assign g30922 = ((~g16662)&(~g29810));
assign g13824 = ((~g8623)&(~g11702));
assign g21745 = (g3017&g20330);
assign g30143 = ((~g28761)&(~g14566));
assign g14612 = (g11971&g11993);
assign II23950 = ((~g23162))|((~II23949));
assign g25009 = ((~g22472));
assign g18132 = (g513&g16971);
assign II14517 = ((~g10147))|((~II14516));
assign g24163 = ((~II23333));
assign g34684 = (g14178&g34545);
assign g13730 = ((~g3639)&(~g11663));
assign g18147 = (g599&g17533);
assign II20951 = ((~g17782));
assign g17056 = ((~g13437));
assign g19386 = ((~g16431));
assign g27549 = (g26576&g14785);
assign g23345 = (g19735)|(g16203);
assign g22762 = (g9305&g20645);
assign g9853 = ((~g5297));
assign II12858 = ((~g4340));
assign g22496 = ((~g19510));
assign g14585 = (g1141&g10905);
assign II15070 = ((~g10108));
assign g24313 = (g4504&g22228);
assign g32642 = ((~g31542));
assign g8974 = ((~II12930));
assign g8989 = ((~II12935));
assign g14178 = ((~g8899)&(~g11083));
assign g26105 = ((~II25146));
assign g31837 = ((~g29385));
assign g24136 = ((~g20857));
assign g32177 = (g30608&g25214);
assign g33635 = ((~g33436));
assign g22112 = (g6555&g19277);
assign g24209 = (g23415)|(g18122);
assign g20712 = ((~g15509));
assign g15096 = ((~g13191)&(~g12867));
assign g27536 = (g26519&g17738);
assign g27390 = (g26549&g17504);
assign g32716 = ((~g31376));
assign g17604 = ((~II18555));
assign g9861 = ((~g5459));
assign g25686 = (g24712)|(g21881);
assign g25385 = ((~g22369))|((~g1783))|((~g8241));
assign g34994 = ((~II33282));
assign II23585 = ((~g22409))|((~g4332));
assign g33311 = (g31942&g12925);
assign g22847 = ((~g20283));
assign g20604 = ((~g17873));
assign g21895 = (g20135)|(g15108);
assign g32481 = ((~g31194));
assign g32728 = ((~g31021));
assign g13501 = ((~g3368)&(~g11881));
assign g10602 = ((~g7411))|((~g7451));
assign g24284 = (g4375&g22550);
assign g32196 = (g27587&g31376);
assign g28591 = (g27332)|(g26286);
assign g21370 = ((~g16323));
assign g30118 = (g28574&g21050);
assign g24818 = ((~g23191));
assign g14417 = ((~g12149)&(~g9648));
assign g20373 = ((~g17929));
assign g26870 = ((~II25606));
assign g27822 = (g4157&g25893);
assign II12097 = ((~g1339))|((~II12096));
assign g21386 = ((~g15798))|((~g15788))|((~g15782))|((~g13139));
assign g17224 = ((~II18248));
assign g18284 = (g15071&g16164);
assign g11940 = ((~g2712)&(~g10084));
assign g30048 = (g29193&g12945);
assign g27226 = (g25872)|(g24436);
assign II12252 = ((~g1124))|((~II12251));
assign g10801 = ((~g1041)&(~g7479));
assign g11519 = ((~g8481));
assign g32261 = (g31251&g20386);
assign g14316 = (g2370&g11920);
assign g21652 = ((~g17619)&(~g17663));
assign g27769 = ((~g9434)&(~g25805));
assign g25473 = ((~g12437))|((~g22432));
assign g34094 = ((~g33772));
assign g20716 = ((~g15277));
assign g25869 = ((~g25250));
assign g8160 = ((~g3423));
assign g34501 = ((~g34400));
assign g7993 = ((~II12333));
assign g30524 = (g30255)|(g22070);
assign g9477 = ((~II13149));
assign g32594 = ((~g30735));
assign g22016 = (g5747&g21562);
assign g29297 = (g28683)|(g18784);
assign g9932 = ((~g5805));
assign g34438 = (g34348)|(g18150);
assign g34574 = ((~II32648));
assign g24813 = (g22685)|(g19594);
assign g30734 = (g13808)|(g29774);
assign g20039 = ((~g11250))|((~g17794));
assign II15536 = ((~g1227));
assign g14179 = ((~g11048));
assign g19853 = ((~g15746)&(~g1052));
assign g22753 = ((~g1536))|((~g19632));
assign g25839 = (g25507)|(g25485)|(g25459)|(g25420);
assign g19453 = ((~g17199)&(~g14316));
assign g25945 = (g24427)|(g22307);
assign g23138 = ((~g20453));
assign g34178 = (g33712&g24361);
assign g28057 = (g27033)|(g18218);
assign II13010 = ((~g6749));
assign g28610 = (g27347)|(g16484);
assign g31792 = (g30214&g24017);
assign g31905 = (g31746)|(g21952);
assign g34247 = ((~II32240));
assign g26204 = (g1720&g25275);
assign g33772 = ((~II31622));
assign g28050 = (g27692)|(g18165);
assign g6996 = ((~g4955));
assign g19791 = (g14253&g17189);
assign g29606 = (g28480&g8011);
assign g25263 = ((~g22763));
assign g25167 = ((~II24331));
assign g19373 = ((~g16449));
assign g21179 = ((~g15373));
assign g14645 = ((~II16755));
assign g16486 = (g6772&g11592&g6789&II17692);
assign g12744 = ((~g9402)&(~g6203));
assign g34967 = (g34951&g23189);
assign g12232 = ((~g8804))|((~g4878));
assign g8216 = ((~g3092));
assign g28115 = (g27354&g22759);
assign g24142 = (g17700&g21657);
assign g22883 = ((~g20391));
assign g13712 = ((~g8984))|((~g11283));
assign g23152 = ((~g20283));
assign g34201 = ((~II32158));
assign g24008 = (g7909&g19502);
assign g30060 = (g29146&g10581);
assign g20540 = ((~g16646));
assign g16884 = (g6159&g14321);
assign g19372 = (g686&g16289);
assign g32606 = ((~g30673));
assign g23434 = ((~g21611));
assign g32844 = ((~g30937));
assign g30134 = ((~g28768)&(~g7280));
assign g29306 = (g28689)|(g18813);
assign g19527 = ((~g16349));
assign g10655 = (g8440&g3423);
assign g34521 = ((~g34270));
assign g18421 = ((~II19235));
assign II16779 = ((~g11292))|((~II16778));
assign g23471 = (g20148&g20523);
assign g28942 = ((~g27858))|((~g2331))|((~g7335));
assign g21415 = ((~g17773))|((~g14771))|((~g17740))|((~g14739));
assign g34688 = ((~II32834));
assign g33843 = (g33256&g20325);
assign g26290 = (g2595&g25498);
assign g27452 = (g26400&g17600);
assign g13834 = ((~g4754))|((~g11773));
assign g12284 = (g1532&g7557);
assign g13124 = ((~g10666))|((~g7661))|((~g979))|((~g1061));
assign g17650 = ((~g6299))|((~g12101))|((~g6315))|((~g14745));
assign g20581 = (g10801&g15571);
assign g20652 = ((~II20744));
assign g15679 = (g3470&g13555);
assign g19578 = (g16183&g11130);
assign g33137 = ((~g4849)&(~g32072));
assign g18818 = (g15165&g15483);
assign g28070 = (g27050)|(g21867);
assign g23828 = (g9104&g19128);
assign g26879 = (g25580)|(g25581);
assign g27231 = (g25873)|(g15699);
assign II26094 = ((~g26055))|((~II26093));
assign g33159 = (g32016)|(g30730);
assign g32123 = (g30915)|(g30919);
assign II18411 = ((~g13018));
assign g8700 = ((~g4054));
assign II25327 = ((~g24641));
assign g33961 = (g33789)|(g21712);
assign g15089 = ((~g13144)&(~g12861));
assign g25247 = ((~g23763)&(~g14645));
assign g23131 = (g13919&g19930);
assign II12103 = ((~g572));
assign g21791 = (g3368&g20391);
assign II26948 = (g24981&g26424&g22698);
assign g8334 = ((~g3034));
assign g25674 = (g24755)|(g21831);
assign g29990 = (g29007&g9239);
assign g25535 = ((~g22763));
assign II16168 = ((~g3321));
assign g24749 = (g17511&g22432);
assign g16958 = ((~g14238));
assign g20636 = ((~g18008));
assign g24554 = (g22490&g19541);
assign g27651 = (g22448&g25781);
assign g33680 = (g33128&g4688);
assign g13142 = ((~g10632));
assign II31147 = (g32668&g32669&g32670&g32671);
assign g12512 = ((~g7766))|((~g10312));
assign g15008 = ((~g12780))|((~g10341));
assign g15426 = ((~II17121));
assign g18801 = (g15160&g15348);
assign g12858 = ((~g10365)&(~g10430));
assign II33176 = ((~g34887));
assign g7092 = ((~g6483));
assign II32173 = ((~g33645));
assign g17662 = ((~II18634))|((~II18635));
assign g19656 = (g2807&g15844);
assign g23943 = ((~g19147));
assign g23415 = (g20077&g20320);
assign g24476 = (g18879&g22330);
assign g7380 = ((~g2331));
assign g23786 = ((~II22945))|((~II22946));
assign g29372 = ((~II27738));
assign II32950 = ((~g34713));
assign g33441 = (g32251&g29722);
assign g24079 = ((~g20998));
assign g27050 = (g25789&g22338);
assign g28226 = (g27825&g26667);
assign g27461 = (g26576&g17611);
assign g8154 = ((~g3139));
assign g15161 = ((~g13809)&(~g7073));
assign g8971 = ((~II12927));
assign g33033 = (g32333)|(g21843);
assign g25218 = ((~g23949));
assign g12402 = ((~g7704))|((~g10266));
assign g31777 = (g21343&g29385);
assign g30195 = ((~II28434));
assign g18211 = (g15062&g15979);
assign g16272 = ((~g13580)&(~g11189));
assign g28751 = (g27526)|(g16766);
assign g15748 = ((~g13257))|((~g13130))|((~g7922))|((~g13241));
assign g9497 = ((~II13166));
assign g34378 = (g13095&g34053);
assign g25514 = ((~g12540))|((~g22498));
assign II18280 = ((~g12951));
assign g11640 = ((~II14550));
assign II25095 = ((~g25265));
assign g27573 = ((~g26667));
assign g9827 = ((~g1974));
assign g7387 = ((~g2421));
assign II20321 = ((~g16920));
assign g20665 = ((~g15373));
assign g7953 = ((~g4966));
assign g20201 = ((~II20468))|((~II20469));
assign g29979 = (g23655&g28991);
assign g28331 = (g27129)|(g15814);
assign g31469 = ((~g8822)&(~g29725));
assign g10040 = ((~g2652));
assign g24515 = ((~g22689));
assign g34868 = (g34813&g19866);
assign g30181 = (g28636&g23821);
assign II16498 = ((~g10430));
assign gbuf62 = (g6661);
assign g19779 = ((~g16431));
assign II32791 = ((~g34578));
assign g12356 = ((~g7438))|((~g6012));
assign g8913 = ((~II12877))|((~II12878));
assign g21828 = (g3767&g20453);
assign g24499 = (g22217&g19394);
assign g14741 = ((~g12711))|((~g10421));
assign g22837 = ((~g20219))|((~g2907));
assign II22444 = ((~g19626));
assign g31919 = (g31758)|(g22044);
assign g30202 = (g28667&g23863);
assign g20902 = ((~II20870));
assign g26850 = ((~II25576));
assign g15821 = (g3598&g14110);
assign g32118 = ((~g31008));
assign g20081 = ((~g11325))|((~g17794));
assign g8492 = ((~g3396));
assign g16305 = ((~g13346));
assign II22275 = ((~g20127));
assign g13745 = ((~II16102));
assign g18670 = (g4621&g15758);
assign g10542 = ((~g7196));
assign g22722 = ((~II22031));
assign g34158 = (g33784)|(g19740);
assign g28148 = (g27355&g26093);
assign g10335 = ((~g4483));
assign g15861 = (g3957&g14170);
assign II14993 = ((~g6527))|((~II14991));
assign g23376 = ((~g21070));
assign g34659 = ((~II32775));
assign g28201 = (g27499&g16720);
assign g32360 = (g29868)|(g31299);
assign g25723 = (g25033)|(g22006);
assign g28296 = (g27095)|(g15784);
assign g20783 = ((~g14616))|((~g17225));
assign g21809 = (g3574&g20924);
assign g11110 = ((~g8728));
assign g23565 = ((~g21562));
assign g20501 = ((~g17955));
assign II12896 = ((~g4229));
assign g24001 = (g19651&g10951);
assign g25272 = ((~g23715));
assign g23748 = ((~II22872))|((~II22873));
assign g18814 = (g6519&g15483);
assign g21225 = ((~g17428));
assign g25155 = ((~g22472));
assign g24205 = (g23006)|(g18109);
assign II14537 = ((~g10106));
assign g12522 = ((~g10133))|((~g5990))|((~g6040));
assign g28307 = ((~g27306));
assign g21867 = (g4082&g19801);
assign g28135 = (g27959)|(g27963);
assign g28043 = (g27323)|(g21714);
assign g28096 = (g27988)|(g21997);
assign II22873 = ((~g21228))|((~II22871));
assign g18910 = (g16227&g16075);
assign g32334 = (g31375&g23568);
assign g33979 = (g33942)|(g18361);
assign g22055 = (g6128&g21611);
assign II14350 = ((~g8890))|((~g8848));
assign g34013 = (g33901)|(g18488);
assign g21337 = ((~g15758));
assign g18654 = (g4146&g16249);
assign g33468 = (g32512&II31036&II31037);
assign g34464 = (g34340)|(g18687);
assign g21899 = (g20162)|(g15113);
assign g11349 = ((~II14365));
assign II32461 = ((~g34244));
assign g21307 = ((~g15719))|((~g13067))|((~g15709))|((~g13040));
assign g32809 = ((~g31327));
assign g14251 = ((~g12308));
assign g34240 = (g32910)|(g33958);
assign g31276 = (g29567)|(g28282);
assign g27543 = (g26085)|(g24670);
assign g30291 = (g28672)|(g27685);
assign g30298 = (g28245)|(g27251);
assign g23396 = (g20051&g20229);
assign g34451 = (g34393)|(g18664);
assign g12431 = ((~II15254))|((~II15255));
assign g14706 = ((~g6287))|((~g12101))|((~g6369))|((~g12672));
assign g11804 = ((~g8938)&(~g4975));
assign g22996 = ((~g20330));
assign g23419 = ((~g21468));
assign g24039 = ((~g21256));
assign g34153 = (g33899)|(g33451);
assign g33638 = ((~II31469));
assign g28799 = (g21434&g26424&g25348&g27445);
assign g19144 = ((~g16031));
assign g16448 = (g13287)|(g10934);
assign g14233 = (g8639&g11855);
assign g33425 = (g32380&g21466);
assign g17217 = ((~g7239))|((~g14194));
assign g29950 = ((~g28896));
assign II21993 = ((~g7670))|((~II21992));
assign g27591 = (g26181)|(g24765);
assign g13968 = ((~g3913))|((~g11255))|((~g4031))|((~g11631));
assign g33130 = ((~g32265)&(~g31497));
assign II25779 = ((~g26424));
assign g14793 = ((~g2988)&(~g12228));
assign g34595 = ((~II32693));
assign II22892 = ((~g12189))|((~g21228));
assign II14192 = ((~g10233));
assign g18540 = (g2775&g15277);
assign g16279 = (g4512&g14424);
assign g18266 = (g1274&g16000);
assign g21911 = (g5046&g21468);
assign g24194 = (g106&g22722);
assign g27968 = (g25958&g19614);
assign g32649 = ((~g30673));
assign g32863 = ((~g31021));
assign g23016 = ((~g20453));
assign g12002 = ((~g5297)&(~g7004));
assign II31694 = ((~g33176));
assign g26241 = (g24688&g10678&g8778&g10627);
assign g24535 = ((~g22942));
assign g28045 = (g27378)|(g18141);
assign g15131 = ((~g12881)&(~g13638));
assign g27316 = (g2407&g26710);
assign g24251 = (g22637)|(g18296);
assign g11083 = (g8836&g802);
assign g16245 = (g14278&g14708);
assign g28184 = ((~II26705));
assign g13091 = (g329)|(g319)|(g10796);
assign g11652 = ((~g7674));
assign g18379 = (g1906&g15171);
assign g33472 = (g32542&II31056&II31057);
assign II24694 = (g20982&g24047&g24048&g24049);
assign g8178 = ((~II12437));
assign g33876 = (g33286&g20562);
assign g11043 = ((~g8561));
assign g10199 = ((~g1968));
assign g13411 = (g4955&g11834);
assign II33037 = ((~g34770));
assign g29105 = (g27645)|(g17134);
assign g25637 = (g24618)|(g18307);
assign g23290 = ((~g20924));
assign g29247 = (g28694)|(g18410);
assign g33893 = (g33313&g20706);
assign g18350 = (g1779&g17955);
assign g10497 = ((~g10102));
assign g14568 = ((~g12000)&(~g9915));
assign II14735 = ((~g5475))|((~II14733));
assign g33415 = (g32368&g21422);
assign g23495 = ((~II22622));
assign g30606 = ((~II28866));
assign g16870 = (g6625&g14905);
assign g20174 = (g5503&g17754);
assign g19855 = (g2787&g15962);
assign g26751 = (g24903)|(g24912);
assign II32305 = ((~g34209));
assign g27290 = (g25926)|(g25928);
assign g29173 = ((~g9259)&(~g27999)&(~g7704));
assign g31760 = (g30007)|(g30027);
assign g10705 = (g6850&g10219&g2689);
assign g24721 = (g17488&g22369);
assign g31122 = (g12144&g29993);
assign g11122 = ((~g8751));
assign g26304 = (g2697&g25246);
assign g16970 = (g13567)|(g11163);
assign g23774 = (g14867&g21252);
assign g24064 = ((~g20841));
assign g34998 = ((~g34981));
assign II22844 = ((~g12113))|((~g21228));
assign g8016 = ((~g3391));
assign g11035 = (g5441&g9800);
assign g18392 = (g1988&g15171);
assign g21183 = ((~g15509));
assign g7582 = ((~g1361))|((~g1373));
assign g19612 = ((~g16897));
assign g26938 = (g26186)|(g21883);
assign II27735 = ((~g28779));
assign g14392 = ((~g12114)&(~g9537));
assign g16843 = (g6251&g14864);
assign g25654 = (g24634)|(g18606);
assign g14187 = (g8871)|(g11771);
assign g8691 = ((~g3267))|((~g3310))|((~g3281))|((~g3303));
assign g12323 = ((~g9480))|((~g640));
assign II25598 = ((~g25424));
assign g32623 = ((~g30735));
assign II14957 = ((~g6181))|((~II14955));
assign g28346 = (g27243&g19800);
assign g21738 = (g3072&g20330);
assign g21773 = (g3263&g20785);
assign g17613 = (g11547&g11592&g11640&II18568);
assign g31307 = (g29596)|(g28311);
assign g30425 = (g29770)|(g21809);
assign II18252 = ((~g13177));
assign g30996 = ((~g29694));
assign g20609 = ((~g15373));
assign g12374 = ((~g2185)&(~g8205));
assign g10035 = ((~g1720));
assign g23478 = ((~g21514));
assign g29240 = (g28655)|(g18328);
assign g21752 = (g3171&g20785);
assign g9333 = ((~g417));
assign g14735 = ((~g12739))|((~g12571));
assign II33291 = ((~g34983));
assign g28448 = ((~g23975))|((~g27377));
assign g34630 = (g34560)|(g15117);
assign g23878 = ((~g19147));
assign g27735 = ((~g7262)&(~g25821));
assign g8864 = ((~g3179)&(~g3171));
assign II27954 = ((~g28803));
assign g17135 = ((~g14297));
assign g34931 = (g2984)|(g34912);
assign g18724 = (g4907&g16077);
assign g21868 = (g4076&g19801);
assign g29812 = ((~g28381));
assign g29273 = (g28269)|(g18639);
assign II18148 = ((~g13526));
assign g7964 = ((~g3155));
assign g10511 = ((~g4628))|((~g7202))|((~g4621));
assign g32927 = ((~g30825));
assign g34787 = ((~II32991));
assign g18256 = (g1242&g16897);
assign g31878 = (g31015)|(g21733);
assign g22515 = (g12981&g19395);
assign g21062 = ((~g9547)&(~g17297));
assign g8347 = ((~g4358))|((~g4349))|((~g4340));
assign g25148 = (g16867&g23545);
assign g32238 = (g30594)|(g29349);
assign g20600 = ((~g15348));
assign II16479 = ((~g10430));
assign g29909 = (g28435&g23388);
assign g22198 = ((~g19147));
assign g27186 = (g26195&g8316&g2342);
assign g17669 = ((~g3570))|((~g11238))|((~g3632))|((~g13902));
assign g29330 = (g29114&g18894);
assign g18926 = ((~II19707));
assign g33126 = (g9044&g32201);
assign g8155 = ((~g3380));
assign gbuf57 = (g6140);
assign g9162 = ((~g622));
assign g26733 = (g10776)|(g24447);
assign g20208 = ((~g17533));
assign g18455 = (g2327&g15224);
assign g7187 = ((~g6065));
assign g10323 = ((~II13744));
assign g17175 = ((~g1216)&(~g13545));
assign gbuf1 = (g4520);
assign g13944 = ((~g10262)&(~g12259));
assign g31303 = (g29592)|(g29606);
assign g24259 = (g23008)|(g18312);
assign g11235 = ((~II14301));
assign g9258 = ((~II13044))|((~II13045));
assign II26705 = ((~g27967));
assign g34382 = (g34167&g20618);
assign g7851 = ((~g921));
assign g21861 = (g3949&g21070);
assign g32354 = (g29854)|(g31285);
assign II28576 = ((~g28431));
assign g12806 = ((~g9472)&(~g9407));
assign g33489 = (g32665&II31141&II31142);
assign g10403 = ((~g7040));
assign g33239 = (g32117&g19902);
assign g25816 = (g8164&g24604);
assign g34909 = (g34856&g20130);
assign II15168 = ((~g9823))|((~II15166));
assign g16292 = ((~g7943)&(~g13134));
assign g21206 = ((~g6419)&(~g17396));
assign g26054 = ((~g24804));
assign g28824 = ((~g27779))|((~g7356))|((~g1772));
assign g22115 = (g6573&g19277);
assign g28183 = (g27024&g19421);
assign II15717 = ((~g6346));
assign g30497 = (g30242)|(g21993);
assign g8135 = ((~II12418));
assign g20380 = ((~g17955));
assign g19905 = ((~g15885));
assign g28248 = (g27150&g19676);
assign g30332 = ((~II28597));
assign g14591 = ((~II16709));
assign g32656 = ((~g30673));
assign g13336 = ((~g11330)&(~g11011));
assign g31129 = (g1968&g30017);
assign II15223 = ((~g10119));
assign g34723 = (g34710)|(g18139);
assign g17752 = (g7841&g13174);
assign g33104 = (g26296&g32137);
assign g25614 = (g24797)|(g18161);
assign g29930 = ((~II28162));
assign g28639 = (g27767&g20597);
assign g34376 = (g26301)|(g34140);
assign g33271 = (g32120)|(g29549);
assign g9917 = ((~II13473));
assign g23836 = (g4129&g19495);
assign g31274 = (g29565)|(g28280);
assign g27331 = (g10177&g26754);
assign g28632 = (g27373)|(g16535);
assign g13539 = ((~g8594)&(~g12735));
assign g26779 = (g24497&g23620);
assign g24012 = (g14496&g21561);
assign II33075 = ((~g34843));
assign g33052 = (g31961)|(g21973);
assign g27416 = (g8046&g26314&g9187&g504);
assign II14381 = ((~g8300));
assign g28776 = (g27538)|(g13974);
assign g33924 = (g33335&g33346);
assign g13437 = ((~II15937));
assign II31036 = (g30673&g31802&g32506&g32507);
assign g33983 = (g33877)|(g18373);
assign g29146 = ((~g6565)&(~g26994));
assign g34717 = ((~II32881));
assign g19626 = ((~g17409));
assign g32247 = (g31168)|(g29686);
assign g7134 = ((~g5029));
assign g26808 = (g25521&g21185);
assign g30164 = (g28618&g23787);
assign g29782 = (g28328&g23245);
assign g28482 = ((~g3522)&(~g27617));
assign II17104 = ((~g12932));
assign g28241 = ((~g27064));
assign g6814 = ((~g632));
assign II17249 = ((~g13605));
assign II27579 = ((~g28184));
assign g26359 = (g24651)|(g22939);
assign II18536 = ((~g2236))|((~g14642));
assign g18646 = (g4031&g17271);
assign g20590 = ((~g15426));
assign g29115 = ((~g27779));
assign g20181 = ((~g13252))|((~g16846));
assign g20547 = ((~g15224));
assign g17726 = (g1467&g13315);
assign g11026 = ((~g8434));
assign g24394 = ((~g22228));
assign II31246 = (g31672&g31839&g32810&g32811);
assign g7280 = ((~g2153));
assign g18813 = (g6513&g15483);
assign g17675 = ((~g5252))|((~g14399))|((~g5320))|((~g12239));
assign g32317 = (g5507&g31542);
assign g24825 = ((~g23204));
assign g33883 = (g33294&g20589);
assign g7261 = ((~g4449));
assign g18261 = (g1256&g16000);
assign g32945 = ((~g30937));
assign g25090 = ((~g23630));
assign g28410 = ((~g27074))|((~g13679));
assign g32653 = ((~g30825));
assign g34531 = ((~II32594));
assign g20544 = ((~g15171));
assign g33023 = (g32313)|(g21751);
assign g30057 = (g29144&g9462);
assign g25593 = (g24716)|(g21707);
assign II32878 = ((~g34501));
assign g26714 = ((~g9316))|((~g25175));
assign g13034 = ((~g11920));
assign g21782 = (g3416&g20391);
assign g33798 = (g33227&g20058);
assign g14547 = ((~g9439))|((~g12201));
assign g17713 = ((~g12947));
assign g30281 = (g28850&g23992);
assign g10085 = ((~g1768));
assign g9978 = ((~g2756));
assign g32661 = ((~g31070));
assign g10674 = (g6841&g10200&g2130);
assign g12695 = ((~g9269)&(~g9239));
assign II12336 = ((~g52));
assign II21006 = ((~g15579));
assign g24330 = (g18661&g22228);
assign g29311 = ((~g28998));
assign II23119 = ((~g20076))|((~II23118));
assign g22710 = (g19358&g19600);
assign g7660 = ((~II12144));
assign II11688 = ((~g70));
assign g30069 = (g29175&g12708);
assign g19543 = ((~g16349));
assign g19401 = ((~g17193)&(~g14296));
assign g28617 = (g27533&g20552);
assign g12211 = ((~g10099)&(~g7097));
assign II18504 = ((~g5283));
assign g9581 = ((~g91));
assign g24703 = (g17592&g22369);
assign g27293 = (g9972&g26655);
assign g9615 = ((~II13236));
assign II30641 = ((~g32024));
assign g27152 = (g24393)|(g25817);
assign g15781 = ((~g6267))|((~g12173))|((~g6329))|((~g14745));
assign II14365 = ((~g3303));
assign g17498 = ((~g14688));
assign g24527 = ((~g22670));
assign g24266 = (g22329)|(g18561);
assign g26271 = (g1992&g25341);
assign g32414 = (g4944&g30999);
assign g25565 = (g13013&g22660);
assign g18163 = (g79&g17433);
assign g9975 = ((~II13519))|((~II13520));
assign g34293 = (g26854)|(g34224);
assign g32566 = ((~g30825));
assign g17732 = ((~g3937))|((~g13824))|((~g4012))|((~g13933));
assign g30207 = (g28680&g23874);
assign g16284 = ((~II17609));
assign g33838 = ((~g33083))|((~g4369));
assign II15254 = ((~g10078))|((~II15253));
assign g24363 = (g7831)|(g22138);
assign g12866 = ((~g10369));
assign g31815 = ((~g29385));
assign g9490 = ((~g2563));
assign g28404 = (g27215)|(g15874);
assign g18204 = (g914&g15938);
assign g18444 = (g2269&g18008);
assign g22316 = (g2837&g20270);
assign g16316 = ((~g9429))|((~g13518));
assign g13782 = ((~II16117));
assign g27385 = (g26400&g17497);
assign g27270 = (g26805&g26793);
assign g30346 = (g29381)|(g18303);
assign g26153 = (g24565&g19780);
assign II24041 = ((~g22182));
assign g26388 = (g19595&g25552);
assign g29636 = (g2403&g29097);
assign g23983 = ((~g19210));
assign g15788 = ((~g6613))|((~g12211))|((~g6675))|((~g14786));
assign g24908 = (g3752&g23239&II24075);
assign g11815 = ((~g7582));
assign g18332 = (g1677&g17873);
assign g32168 = (g30597&g25185);
assign g25786 = ((~g24518));
assign II20647 = ((~g17010));
assign II29304 = ((~g12121))|((~II29302));
assign g20739 = (g16259&g4674);
assign g32462 = ((~g30673));
assign g18793 = (g6159&g15348);
assign g7715 = ((~g1178));
assign g29797 = (g28347&g23259);
assign g11447 = ((~II14450));
assign g23247 = ((~g20924));
assign g11205 = (g8217&g8439);
assign g22680 = (g19530&g7781);
assign g21429 = ((~g17788))|((~g14803))|((~g17578))|((~g17520));
assign g25038 = ((~g21331))|((~g23363));
assign g12887 = ((~g10394));
assign g34913 = ((~II33131));
assign g26922 = (g25902)|(g18288);
assign g34004 = (g33879)|(g18453);
assign g23387 = (g16506&g20211);
assign g9103 = ((~g5774));
assign g28154 = (g8492&g27306);
assign II25846 = ((~g26212))|((~II25845));
assign g32797 = ((~g30825));
assign g23007 = (g681&g20248);
assign g10614 = ((~g9024))|((~g8977))|((~g8928));
assign g32282 = (g31258&g20503);
assign g28736 = ((~g27742))|((~g7308))|((~g7252));
assign g14771 = ((~g5961))|((~g12129))|((~g5969))|((~g12351));
assign g9226 = ((~g1564));
assign g16775 = ((~II17999));
assign II13183 = ((~g6500))|((~II13182));
assign g25112 = (g10428&g23510);
assign g8871 = ((~II12841))|((~II12842));
assign g29337 = (g29166&g22180);
assign g16158 = ((~g13555));
assign II18891 = ((~g16676));
assign II14267 = ((~g7835));
assign g25935 = (g24402)|(g22208);
assign g27139 = (g26055&g16608);
assign g23810 = ((~II22973))|((~II22974));
assign g34113 = (g33734&g19744);
assign g16577 = ((~II17747));
assign g24958 = ((~g21330))|((~g23462));
assign g30450 = (g29861)|(g21859);
assign g7004 = ((~II11777));
assign g27037 = (g26236)|(g26218)|(g26195)|(g26171);
assign II25613 = (g25571)|(g25572)|(g25573)|(g25574);
assign g15509 = ((~II17136));
assign g34494 = (g26849)|(g34413);
assign g33141 = ((~g32099)&(~g8400));
assign g23648 = ((~g18833));
assign g25804 = (g8069&g24587);
assign g26218 = (g25357&g6856&g7586&g11686);
assign g22521 = ((~g1036)&(~g19699));
assign g27026 = (g26828)|(g17726);
assign g12906 = ((~g10413));
assign g27580 = (g26159)|(g24749);
assign g13278 = ((~g10738));
assign g28959 = (g17401&g25194&g26424&g27440);
assign g21761 = (g3215&g20785);
assign g14821 = ((~g6390)&(~g12314));
assign g32588 = ((~g30825));
assign g15055 = ((~g6808)&(~g13350));
assign g12780 = ((~g9402)&(~g9326));
assign g22585 = (g20915)|(g21061);
assign g11023 = (g9669&g5084);
assign g14275 = ((~g12358));
assign g29367 = (g8575&g28325);
assign g10862 = ((~g7701)&(~g7840));
assign g28884 = (g27568)|(g16885);
assign g32499 = ((~g31376));
assign g23890 = ((~g7004))|((~g20682));
assign g27370 = (g26400&g17472);
assign g26288 = (g2259&g25309);
assign g30405 = (g29767)|(g21764);
assign g34941 = ((~g34926));
assign g7922 = ((~g1312));
assign II12930 = ((~g4349));
assign II31459 = ((~g33219));
assign g28314 = (g27552&g14205);
assign g22648 = (g18987)|(g15652);
assign g26630 = (g7592&g24419);
assign g11858 = ((~g9014))|((~g3010));
assign g33490 = (g32672&II31146&II31147);
assign g33956 = (g33514)|(II31863)|(II31864);
assign g34220 = ((~II32186))|((~II32187));
assign g13707 = ((~g11360));
assign g31977 = (g31764&g22179);
assign g32934 = ((~g30735));
assign g32790 = ((~g30825));
assign g13871 = ((~g4955))|((~g11834));
assign g21938 = (g5216&g18997);
assign g29046 = ((~g27779))|((~g9640));
assign II31839 = (g33465)|(g33466)|(g33467)|(g33468);
assign g8743 = ((~g550));
assign II26337 = ((~g26835));
assign g19619 = (g15712)|(g13080);
assign II21033 = ((~g17221));
assign g11674 = ((~g8676))|((~g4674));
assign g16662 = (g4552&g14753);
assign g17595 = ((~g8616))|((~g14367));
assign II23390 = ((~g23395));
assign g18681 = (g4653&g15885);
assign g16538 = (g6255&g15005);
assign g12026 = ((~g9417)&(~g9340));
assign g10429 = ((~g7148));
assign g9070 = ((~g5428));
assign g29201 = (g24081&II27503&II27504);
assign g33603 = (g33372)|(g18515);
assign g13067 = ((~g5240))|((~g12059))|((~g5331))|((~g9780));
assign II32441 = ((~g34220))|((~II32439));
assign g7258 = ((~g4414));
assign g11395 = ((~g9601))|((~g3983));
assign g9959 = ((~g6177));
assign g25760 = (g25238)|(g22109);
assign g32835 = ((~g31710));
assign g32967 = ((~g31327));
assign g32143 = (g31646&g29967);
assign II23918 = ((~g23975))|((~II23917));
assign II15002 = ((~g9691))|((~g1700));
assign g27507 = (g26549&g17683);
assign g9528 = ((~II13183))|((~II13184));
assign g22043 = (g5965&g19147);
assign g8955 = ((~g1418));
assign g31889 = (g31118)|(g21822);
assign g24724 = (g17624&g22432);
assign g23228 = ((~g21070));
assign g29592 = (g28469&g11832);
assign g25697 = (g25086)|(g21916);
assign II14198 = (g225&g8237&g232&g8180);
assign g34649 = (g33111)|(g34492);
assign g22094 = (g6398&g18833);
assign g33148 = ((~g4854)&(~g32072));
assign II31346 = (g31021&g31857&g32954&g32955);
assign g20384 = ((~g18008));
assign g9899 = ((~g6513));
assign g18344 = (g1740&g17955);
assign g32323 = (g31311&g20610);
assign g31657 = ((~II29239));
assign g17307 = (g9498&g14343);
assign g30016 = ((~g29049));
assign g29841 = (g28371&g23283);
assign II24524 = (g5041&g5046&g9716);
assign g32084 = (g10948&g30825);
assign g8182 = ((~g405)&(~g392));
assign g10390 = ((~g6987));
assign g12891 = ((~g10399));
assign g27030 = (g26343&g7947);
assign g27333 = (g10180&g26765);
assign g30280 = ((~g7064)&(~g29036));
assign g20560 = ((~g17328));
assign g11129 = ((~g7994));
assign II31486 = ((~g33197));
assign g26910 = (g26571)|(g24228);
assign g10830 = ((~g10087));
assign g23510 = ((~g18833));
assign g24325 = (g4543&g22228);
assign g19737 = ((~g17015));
assign g13911 = ((~g11834))|((~g4917));
assign II33282 = ((~g34987));
assign g29630 = (g28212&g19781);
assign g9671 = ((~g5134));
assign g31257 = (g29531)|(g28253);
assign g34691 = ((~II32843));
assign II33279 = ((~g34986));
assign g24302 = (g15124&g22228);
assign g19368 = ((~g16326));
assign g33349 = (g32233&g20699);
assign g11608 = ((~g7659));
assign g14198 = ((~g12180));
assign g20267 = ((~g17955));
assign g19412 = ((~g16489));
assign g13050 = ((~g5543))|((~g12029))|((~g5654))|((~g9864));
assign g12192 = ((~g8267))|((~g2319));
assign g26745 = ((~g6856))|((~g25317));
assign g28987 = ((~g27886))|((~g2070))|((~g7411));
assign g25963 = (g1657&g24978);
assign g17680 = ((~g14889));
assign g24518 = (g22517)|(g7601);
assign g29748 = (g28210)|(g28214);
assign g34799 = (g34751)|(g18578);
assign g13082 = ((~g10981));
assign g25522 = (g6888&g22544);
assign g33098 = ((~g31997)&(~g4616));
assign g7788 = ((~g4674));
assign g9491 = ((~g2729));
assign g25991 = (g2060&g25023);
assign g34312 = ((~g34098));
assign g21734 = (g3040&g20330);
assign g7738 = ((~II12176));
assign g29289 = (g28642)|(g18763);
assign g26205 = (g2098&g25492);
assign g10608 = ((~g9155));
assign g33246 = ((~g32212));
assign g9553 = ((~II13202));
assign g16623 = ((~g14127));
assign g32470 = ((~g31566));
assign g19520 = ((~g16826));
assign g28562 = (g27313)|(g26251);
assign g9985 = ((~g4332));
assign g22687 = ((~g19560))|((~g7870));
assign g23333 = ((~g20785));
assign g34341 = (g34101&g19952);
assign g10073 = ((~g134));
assign g19635 = ((~g16349));
assign g33689 = (g33144&g11006);
assign g27148 = (g25997&g16622);
assign g27286 = (g6856&g26634);
assign g18179 = (g763&g17328);
assign g18424 = (g2165&g18008);
assign g29813 = (g26020)|(g28261);
assign II31564 = ((~g33204));
assign II31616 = ((~g33219));
assign g13016 = ((~g11878));
assign g20096 = ((~g16782));
assign g22400 = ((~g19345)&(~g15718));
assign g11849 = ((~g7601));
assign g30114 = (g28488)|(g16761);
assign g32056 = (g27271&g31021);
assign gbuf45 = (g6027);
assign g33565 = (g33338)|(g18389);
assign g21247 = ((~g15171));
assign g13087 = ((~g12012));
assign g16677 = ((~II17879));
assign g29224 = (g28919)|(g18156);
assign g30085 = ((~g29082));
assign g31805 = ((~g29385));
assign II24675 = (g24022&g24023&g24024&g24025);
assign g9077 = ((~g504));
assign II25909 = ((~g24782))|((~II25907));
assign g10418 = ((~g8818));
assign g9999 = ((~g6109));
assign g21351 = ((~g15729))|((~g13098))|((~g15720))|((~g13069));
assign g28648 = ((~g27693));
assign g32550 = ((~g31376));
assign II20461 = ((~g17515))|((~II20460));
assign g14571 = ((~II16688));
assign II12935 = ((~g6753));
assign g31326 = (g29627)|(g29640);
assign g11987 = ((~II14833));
assign g23969 = ((~g19277));
assign g15027 = ((~g12667))|((~g10341));
assign II26682 = ((~g27774));
assign g19949 = (g17671)|(g14681);
assign g20662 = ((~g15171));
assign g20597 = ((~g17847));
assign g22662 = (g19069)|(g15679);
assign g29693 = (g28207&g10233);
assign g32202 = (g31069)|(g13410);
assign g23880 = ((~g19210));
assign g29626 = (g28584&g11415);
assign g7340 = ((~g4443));
assign g31322 = (g26128)|(g29635);
assign g9247 = ((~g1559));
assign g14625 = ((~g3897))|((~g11225))|((~g4031))|((~g8595));
assign II14885 = ((~g5489))|((~II14883));
assign g10552 = ((~g2153))|((~g7374));
assign g25719 = (g25089)|(g18761);
assign g26391 = (g19593&g25555);
assign II33179 = ((~g34893));
assign g12849 = ((~g6840)&(~g10430));
assign g32741 = ((~g31710));
assign g23904 = ((~g18997));
assign g27130 = (g26026&g16585);
assign g27160 = (g14163&g26340);
assign g26519 = ((~II25380));
assign g17528 = ((~g14940));
assign g14556 = ((~g6682)&(~g12790));
assign g13106 = ((~g10981));
assign g33522 = (g32902&II31306&II31307);
assign g28419 = (g27221)|(g15884);
assign g21358 = ((~g16307));
assign II13384 = ((~g246))|((~II13382));
assign g19537 = ((~g15938));
assign g27103 = (g25997&g16509);
assign gbuf38 = (g5983);
assign g18456 = (g2338&g15224);
assign g14008 = ((~g11610))|((~g11435));
assign g23963 = ((~g19147));
assign g34442 = (g34380)|(g18542);
assign g21603 = ((~g17872))|((~g14987))|((~g17723))|((~g17689));
assign g16955 = ((~II18107));
assign g27886 = (g14438)|(g26759);
assign g25906 = (g25559)|(g24014);
assign g29513 = (g28448&g14095);
assign II12261 = ((~g1454))|((~g1448));
assign g25704 = (g25173)|(g21925);
assign g8458 = ((~g294));
assign g31992 = (g31773&g22213);
assign g28283 = (g7380&g2361&g27445);
assign II18408 = ((~g13017));
assign g31966 = (g31754&g22166);
assign g33821 = (g33238&g20153);
assign g32702 = ((~g30735));
assign g32988 = (g32232)|(g18325);
assign g24029 = ((~g20982));
assign g34352 = (g26079)|(g34109);
assign g14338 = ((~II16502));
assign g34049 = ((~g33678));
assign g15653 = (g3119&g13530);
assign g26955 = (g26391)|(g24293);
assign g15731 = ((~g13326));
assign g18605 = (g3129&g16987);
assign g34412 = (g34187)|(g25143);
assign g22075 = (g6247&g19210);
assign g13807 = (g4504&g10606);
assign gbuf40 = (g5969);
assign g7040 = ((~g4821));
assign g10916 = ((~g1146))|((~g7854));
assign II18009 = ((~g13680));
assign II12270 = ((~g1141))|((~II12269));
assign g34856 = (g34811)|(g34743);
assign g33755 = ((~II31610));
assign g33536 = (g33241)|(g21715);
assign g18482 = (g2472&g15426);
assign g20613 = ((~g15224));
assign g24409 = (g3484&g23112);
assign g12882 = ((~g10389));
assign g7946 = ((~II12314));
assign II22539 = ((~g19606));
assign g13129 = ((~g7553)&(~g10762));
assign g34735 = (g34709)|(g15116);
assign gbuf29 = (g5623);
assign g33648 = ((~II31482));
assign g34419 = ((~g34151));
assign g22218 = (g19951&g20875);
assign g33942 = (g33383&g21608);
assign g21256 = ((~g15483)&(~g12179));
assign g9771 = ((~g3969));
assign g21659 = ((~g17727));
assign g13918 = ((~g3259))|((~g11217))|((~g3267))|((~g11350));
assign II12666 = ((~g4040));
assign g20680 = ((~g15348));
assign g29790 = (g25975)|(g28242);
assign g25479 = (g22646&g9917);
assign g15738 = (g1111&g13260);
assign g33711 = (g33176&g10727&g22332);
assign g20874 = ((~g15680));
assign g16634 = (g5264&g14953);
assign g18311 = (g1554&g16931);
assign g29767 = (g28317&g23236);
assign g12170 = ((~g10047)&(~g5413));
assign g28525 = (g27284)|(g26176);
assign g24575 = ((~g23498)&(~g23514));
assign g15959 = ((~II17405))|((~II17406));
assign g27649 = (g10820&g25820);
assign II23149 = ((~g19061));
assign g9731 = ((~g5366));
assign gbuf22 = (g5331);
assign g18167 = (g718&g17433);
assign g28322 = (g27117)|(g15809);
assign g10360 = ((~g6836));
assign g23279 = ((~g21037));
assign g32554 = ((~g30614));
assign g18675 = (g4349&g15758);
assign g33373 = (g32288&g21205);
assign g11889 = ((~g9954));
assign g28071 = (g27085)|(g21873);
assign g12924 = (g1570&g10980);
assign g18476 = (g2433&g15426);
assign g34388 = (g10802&g34062);
assign II12903 = (g4222)|(g4219)|(g4216)|(g4213);
assign g28104 = (g27697)|(g22108);
assign g14062 = (g11047)|(g11116);
assign g30041 = (g28511&g23518);
assign II31117 = (g32624&g32625&g32626&g32627);
assign g18771 = (g5685&g15615);
assign g14496 = (g12411&g12244&g12197&II16618);
assign g18729 = (g15139&g16821);
assign g27502 = (g26488&g17677);
assign g8553 = ((~g3747));
assign g18945 = ((~g16100));
assign g31237 = (g29366&g25325);
assign II12842 = ((~g4235))|((~II12840));
assign II31686 = ((~g33164));
assign II15053 = ((~g2259))|((~II15051));
assign g17247 = ((~II18259));
assign II31858 = (g33497)|(g33498)|(g33499)|(g33500);
assign g30596 = (g30279&g18947);
assign g22151 = ((~II21734));
assign g14165 = ((~g8951)&(~g11083));
assign g34760 = ((~II32938));
assign g23729 = ((~g17482)&(~g21206));
assign g30372 = (g30110)|(g18446);
assign g22166 = ((~g18997));
assign g28376 = ((~g27064))|((~g13620));
assign g28786 = ((~g27837))|((~g7405))|((~g7322));
assign g34397 = (g7673&g34068);
assign g32042 = (g27244&g31070);
assign g28725 = (g27596&g20779);
assign g21875 = (g4116&g19801);
assign g31169 = (g10083&g30079);
assign g19516 = (g7824&g16097);
assign g6978 = ((~g4616));
assign g14943 = ((~g7791))|((~g12622));
assign g27668 = (g1367&g25917);
assign II25380 = ((~g24481));
assign g32587 = ((~g30735));
assign g26823 = (g24401&g13106);
assign g18504 = (g2579&g15509);
assign g12790 = ((~g7097));
assign g23919 = (g4122&g19546);
assign g30149 = (g28605&g21248);
assign g28062 = (g27288)|(g21746);
assign II19831 = ((~g16533));
assign g14442 = ((~II16593));
assign g13568 = ((~g8046)&(~g12527));
assign g10389 = ((~g6986));
assign g31315 = (g29607)|(g29623);
assign g31665 = ((~II29245));
assign g29487 = (g25815)|(g28133);
assign g28584 = ((~g7121)&(~g27635));
assign g16177 = (g5128&g14238);
assign g28573 = (g7349&g27059);
assign II14187 = ((~g3470))|((~II14185));
assign g7812 = ((~II12214));
assign g7827 = ((~g4688));
assign g25380 = ((~g23776));
assign g11498 = ((~II14475));
assign g30248 = (g28743&g23938);
assign II25399 = ((~g24489));
assign g21712 = (g294&g20283);
assign g24648 = ((~g23148));
assign g16603 = ((~II17787));
assign g19074 = ((~II19772));
assign g24335 = (g22165)|(g18678);
assign g19595 = (g17149)|(g14218);
assign g26604 = (g13248&g25051);
assign g22832 = (g19354)|(g15722);
assign g12950 = ((~g12708));
assign g27823 = ((~g9792)&(~g25805));
assign g26883 = (g26670)|(g24189);
assign g23242 = ((~g21070));
assign g20027 = ((~g16242)&(~g13779));
assign g10047 = ((~g5421));
assign g27519 = (g26488&g17710);
assign g33627 = (g33376)|(g18826);
assign g9050 = ((~g1087));
assign g34626 = (g34533)|(g18627);
assign g24820 = (g13944&g23978);
assign g6953 = ((~g4157));
assign g32721 = ((~g31021));
assign g25649 = (g24654)|(g21742);
assign g28353 = ((~g9073)&(~g27654)&(~g24732));
assign g34083 = (g33714&g19573);
assign g14344 = ((~g5377))|((~g11885));
assign g13393 = (g703&g11048);
assign g23050 = (g655&g20248);
assign g31540 = (g29904&g23548);
assign g34999 = (g34998&g23085);
assign g26884 = (g26511)|(g24190);
assign g13699 = (g10921)|(g10947);
assign g29769 = (g28319&g23237);
assign g27533 = (g26078)|(g24659);
assign g32051 = (g31506&g10831);
assign II18337 = ((~g1422));
assign II15342 = ((~g2541))|((~II15340));
assign g18622 = (g3480&g17062);
assign g19494 = ((~g16349));
assign g25713 = (g25147)|(g21964);
assign g27703 = ((~g9607)&(~g25791));
assign g32774 = ((~g30735));
assign g34421 = (g27686)|(g34198);
assign II21115 = ((~g15714));
assign g12822 = ((~g6978))|((~g7236))|((~g7224))|((~g7163));
assign II31301 = (g31327&g31849&g32889&g32890);
assign g19742 = ((~g17096));
assign g30363 = (g30121)|(g18407);
assign g24067 = ((~g21256));
assign g7209 = ((~g6052))|((~g6098));
assign g30354 = (g30064)|(g18359);
assign g29475 = (g14033&g28500);
assign g31844 = ((~g29385));
assign g28515 = ((~g3881)&(~g27635));
assign g11566 = ((~g3161)&(~g7964));
assign g10185 = ((~g5969))|((~g6012))|((~g5983))|((~g6005));
assign g24056 = ((~g20014));
assign g11426 = ((~g8742))|((~g4878));
assign g25033 = (g17500&g23433);
assign g34227 = ((~II32203))|((~II32204));
assign g24586 = ((~g23067));
assign g13511 = ((~g182))|((~g174))|((~g203))|((~g12812));
assign g13680 = ((~II16077));
assign g28253 = (g23719&g27700);
assign g30125 = (g28581&g21056);
assign g33387 = (g32263)|(g29954);
assign g25968 = (g25215&g20739);
assign II22769 = ((~g21277));
assign g31247 = (g29513)|(g13324);
assign g23216 = ((~g20924));
assign g28399 = ((~g27074));
assign II18398 = ((~g13745));
assign g25059 = (g20870&g23460);
assign g28729 = (g27502)|(g16732);
assign g31123 = (g1834&g29994);
assign g14518 = ((~II16639));
assign g12977 = ((~II15590));
assign g15126 = ((~g12878)&(~g13605));
assign II12089 = ((~g744));
assign g7074 = ((~II11801));
assign g26862 = ((~II25598));
assign g27421 = (g8038&g26314&g9187&g9077);
assign g19427 = ((~g16292));
assign g16525 = ((~II17723));
assign g18443 = (g2265&g18008);
assign g11675 = ((~g8984))|((~g4912));
assign g16645 = ((~g13756));
assign g26891 = (g26652)|(g24197);
assign g27633 = (g13076&g25766);
assign g12220 = (g1521&g7535);
assign g21308 = ((~g17485));
assign g33514 = (g32844&II31266&II31267);
assign g31209 = (g2084&g30097);
assign g32429 = (g30318)|(g31794);
assign g34669 = ((~II32791));
assign II15003 = ((~g9691))|((~II15002));
assign g33849 = (g33262&g20387);
assign g30467 = (g30185)|(g21938);
assign g7028 = ((~II11785));
assign g12351 = ((~II15194))|((~II15195));
assign II12183 = ((~g2719));
assign g31521 = ((~II29182));
assign g13756 = ((~g203))|((~g12812));
assign g26125 = (g1894&g25117);
assign g26903 = (g26388)|(g24220);
assign g15792 = (g12920)|(g10501);
assign g26348 = (g8466)|(g24609);
assign g14408 = ((~g6069))|((~g11924));
assign g34956 = ((~II33214));
assign g26020 = (g9559&g25034);
assign g19492 = ((~g16349));
assign II14510 = ((~g8721))|((~II14508));
assign g32019 = (g30579&g22358);
assign g34057 = (g33911)|(g33915);
assign g12218 = ((~II15073));
assign g32461 = ((~g30614));
assign g19760 = ((~g17015));
assign g27253 = (g24661)|(g26052);
assign g28550 = (g12009&g27092);
assign g30266 = (g28775&g23966);
assign g32468 = ((~g30614));
assign g11832 = ((~g8011));
assign g10119 = ((~g2841));
assign II21744 = ((~g19338));
assign g16429 = ((~II17671));
assign g7196 = ((~II11860));
assign g23504 = ((~g21468));
assign g32492 = ((~g31376));
assign II18829 = ((~g13350));
assign g11276 = ((~g8534)&(~g8691));
assign II18051 = ((~g13680));
assign g23274 = ((~g21070));
assign g24471 = (g10999)|(g22450);
assign g34614 = (g34518)|(g18568);
assign II15122 = ((~g9910))|((~II15121));
assign g34666 = (g34587&g19144);
assign g33265 = (g32113)|(g29530);
assign g13295 = (g10625)|(g10655);
assign g21892 = (g19788)|(g15104);
assign II12767 = ((~g4197));
assign g24236 = (g22489)|(g18241);
assign II32467 = ((~g34246));
assign g30100 = ((~g29131));
assign g15729 = ((~g5949))|((~g14549))|((~g6027))|((~g9935));
assign g10034 = (g1521&g1500);
assign g32369 = (g2130&g31672);
assign g26873 = ((~g25374)&(~g25331));
assign g13044 = ((~g7349)&(~g10762));
assign g9511 = ((~g5881));
assign g15141 = ((~g12888)&(~g13680));
assign g22228 = ((~II21810));
assign g16475 = ((~g14107));
assign g19881 = ((~g15915));
assign g7907 = ((~g3072));
assign g28860 = ((~g27775))|((~g14586));
assign g34745 = (g34669&g19482);
assign g11313 = ((~g8669)&(~g3759));
assign g8457 = ((~g225));
assign g16609 = ((~g14454));
assign g34103 = (g33701)|(g33707);
assign II25591 = ((~g25380));
assign g30454 = (g29909)|(g21863);
assign g19396 = ((~g16431));
assign g30672 = (g13737)|(g29752);
assign g21841 = (g3857&g21070);
assign g16659 = ((~II17857));
assign g33454 = ((~II30980));
assign g28670 = (g27412)|(g16618);
assign II19772 = ((~g17818));
assign g12166 = ((~g9856)&(~g10124));
assign g27770 = ((~g9386)&(~g25821));
assign g14682 = ((~g4933))|((~g11780));
assign g7498 = ((~g6675));
assign g13990 = ((~g11669))|((~g11584));
assign g27542 = (g16190)|(g26094);
assign g15813 = (g3247&g14069);
assign g34894 = (g34862)|(g21678);
assign g15075 = (g12850&g12955);
assign g29290 = (g28569)|(g18764);
assign g24674 = (g446&g23496);
assign g7675 = ((~g1554)&(~g1559)&(~g1564)&(~g1548));
assign II27742 = ((~g28819));
assign g25107 = (g17643&g23508);
assign II24597 = (g5736&g5742&g9875);
assign g16223 = ((~g13437));
assign g22029 = (g5901&g19147);
assign g19652 = ((~g16897));
assign g13627 = ((~g11172))|((~g8388));
assign g6819 = ((~g1046));
assign g29157 = ((~g9835))|((~g27937));
assign g27499 = ((~g9095)&(~g26636));
assign g13595 = ((~g10951));
assign g33262 = (g32112)|(g29528);
assign g25088 = (g17601&g23491);
assign g26543 = (g12910&g24377);
assign II13750 = ((~g4608))|((~II13749));
assign g25524 = ((~g22228));
assign g23869 = ((~g19277));
assign II14866 = ((~g9748));
assign g9900 = ((~g6));
assign g16075 = ((~g13597));
assign g33529 = (g32953&II31341&II31342);
assign g7892 = ((~g4801));
assign g25130 = (g23358&g20600);
assign g32975 = ((~II30537));
assign g28686 = (g27574&g20650);
assign g33986 = (g33639)|(g18387);
assign g31948 = (g30670&g18884);
assign II11860 = ((~g43));
assign g17317 = (g1079&g13124);
assign g7026 = ((~g5507));
assign g30206 = ((~g28436));
assign g18227 = (g1052&g16129);
assign g18601 = (g3106&g16987);
assign g29910 = ((~g3990)&(~g28484));
assign g21267 = ((~g15680));
assign g21968 = (g5459&g21514);
assign g25672 = (g24647)|(g21829);
assign g33266 = (g32114)|(g29532);
assign g18240 = (g15066&g16431);
assign g20529 = ((~g15509));
assign g33382 = ((~g32033));
assign g32712 = ((~g30614));
assign g20870 = ((~g14432))|((~g17315))|((~g9567));
assign II12128 = ((~g4253));
assign g28268 = (g8572&g27990);
assign g19757 = ((~g17224));
assign gbuf105 = (g4287);
assign g12667 = ((~g7791)&(~g6209)&(~g6203));
assign g30077 = ((~g29057));
assign g14971 = ((~g12667))|((~g12581));
assign g27118 = (g26055&g16529);
assign g21840 = (g15099&g21070);
assign g24450 = (g3129&g23067);
assign g18736 = (g4991&g16826);
assign g29268 = (g28343)|(g18625);
assign g15780 = ((~g5937))|((~g14549))|((~g6012))|((~g14701));
assign g20198 = ((~g16813))|((~g13958))|((~g16745))|((~g13927));
assign II20355 = ((~g17613));
assign g33487 = (g32649&II31131&II31132);
assign g26338 = ((~g8458)&(~g24825));
assign g28009 = ((~II26516));
assign g24090 = ((~g19935));
assign II31469 = ((~g33388));
assign g9569 = ((~g6227));
assign g31872 = (g31524)|(g18535);
assign g31208 = (g30262&g25188);
assign g20995 = ((~g5727)&(~g17287));
assign gbuf93 = (g3983);
assign g19486 = (g15589)|(g12979);
assign g29897 = ((~II28128));
assign gbuf117 = (g4219);
assign g17324 = ((~II18301));
assign g28634 = (g27374)|(g16536);
assign g23687 = (g21384)|(g21363)|(II22830);
assign g25525 = ((~g22550));
assign g32540 = ((~g30614));
assign g24760 = ((~II23918))|((~II23919));
assign g28243 = (g27879&g23423);
assign g11238 = ((~g8584)&(~g6905));
assign g27766 = ((~g9716)&(~g25791));
assign g16226 = ((~g8052)&(~g13545));
assign g21916 = (g5084&g21468);
assign g13806 = ((~g11245)&(~g4076));
assign g15099 = ((~g13191)&(~g12869));
assign g26400 = ((~II25351));
assign II31844 = (g33474)|(g33475)|(g33476)|(g33477);
assign g33227 = (g32029)|(g32031);
assign g30017 = ((~g29085));
assign g34586 = (g11025&g34317);
assign g10585 = ((~g1996))|((~g7451));
assign g11467 = ((~g7623));
assign g16517 = (g5248&g14797);
assign II13392 = ((~g1825))|((~II13390));
assign g11845 = ((~II14663));
assign g32959 = ((~g30937));
assign II12787 = ((~g4311));
assign g18111 = (g174&g17015);
assign g15787 = ((~g6283))|((~g14575))|((~g6358))|((~g14745));
assign II19704 = ((~g17653));
assign g33556 = (g33329)|(g18362);
assign II27552 = ((~g28162));
assign g18821 = (g15168&g15680);
assign g14598 = ((~g5248))|((~g12002))|((~g5331))|((~g12497));
assign II17121 = ((~g14366));
assign II32617 = ((~g34333));
assign g15842 = ((~g13469));
assign g15798 = ((~g6629))|((~g14602))|((~g6704))|((~g14786));
assign g28546 = (g27302)|(g26231);
assign g23251 = (g19637)|(g16098);
assign g24264 = (g22310)|(g18559);
assign g26990 = ((~g26105));
assign g31848 = ((~g29385));
assign g27974 = (g26544)|(g25063);
assign g29582 = (g27766&g28608);
assign g29107 = ((~g6203)&(~g7791)&(~g26977));
assign g28372 = (g27178)|(g15848);
assign g33512 = (g32830&II31256&II31257);
assign g18830 = ((~g18008));
assign g32650 = ((~g31579)&(~II30192)&(~II30193));
assign g31311 = (g26103)|(g29618);
assign g12870 = ((~g10374));
assign g27526 = (g26576&g17721);
assign g15811 = ((~g13125));
assign gbuf75 = (g3298);
assign g21189 = ((~g15634));
assign g10550 = ((~g7268))|((~g7308));
assign g15106 = ((~g12872)&(~g10430));
assign g18093 = ((~II18885));
assign g24222 = (g262&g22594);
assign g21702 = (g157&g20283);
assign g14669 = ((~g12301));
assign g34770 = ((~II32956));
assign II12355 = ((~g46));
assign g22018 = (g15157&g19147);
assign g34055 = (g33909)|(g33910);
assign g8119 = ((~g3727));
assign g33021 = (g32302)|(g21749);
assign g24791 = ((~g23850));
assign II21297 = ((~g18597));
assign g32599 = ((~g30673));
assign g14297 = ((~g10869));
assign g6958 = ((~g4372));
assign g31867 = (g31238)|(g18175);
assign g8170 = ((~g3770));
assign g32990 = (g32281)|(g18341);
assign g27545 = (g26519&g17756);
assign g28694 = (g27579&g20664);
assign g27383 = (g24569)|(g25961);
assign g29982 = (g23656&g28998);
assign g12918 = ((~II15533));
assign g27654 = ((~g164))|((~g26598))|((~g23042));
assign g23348 = (g15570&g21393);
assign g31249 = (g25971)|(g29523);
assign II30745 = (g31777)|(g32321)|(g32069)|(g32084);
assign g29834 = (g28368&g23278);
assign g10417 = ((~g7117));
assign g10349 = ((~g6956));
assign g18118 = (g471&g17015);
assign II12877 = ((~g4200))|((~II12876));
assign g28930 = ((~g27833))|((~g8201));
assign II31796 = ((~g33176));
assign g22148 = ((~g19074));
assign g24684 = (g11769&g22989);
assign g14358 = ((~II16512));
assign II12534 = ((~g50));
assign g30513 = (g30200)|(g22034);
assign g30520 = (g30272)|(g22041);
assign g16690 = (g8399&g13867);
assign g21750 = (g3161&g20785);
assign g9594 = ((~g2307));
assign g7064 = ((~g5990));
assign g18401 = (g2036&g15373);
assign g33331 = (g32216&g20607);
assign g13032 = ((~g7577)&(~g10762));
assign g12065 = (g9557&g9805);
assign g17766 = (g6772&g11592&g11640&II18762);
assign g34603 = (g34561)|(g15075);
assign g34950 = ((~g34940));
assign g31375 = (g29628)|(g28339);
assign g13884 = ((~g11797))|((~g4727));
assign g13294 = (g1564&g11513);
assign g16807 = (g6585&g14978);
assign II17131 = ((~g14384));
assign II22936 = ((~g12226))|((~g21228));
assign g13526 = (g209)|(g10685)|(g301);
assign g31989 = (g31770&g22200);
assign g14569 = ((~g3195))|((~g11194))|((~g3329))|((~g8481));
assign g18704 = (g4793&g16782);
assign II15205 = ((~g10139));
assign II29717 = ((~g30931));
assign g6837 = ((~g968));
assign g21276 = (g10157&g17625);
assign g20134 = ((~g17572))|((~g14542))|((~g17495))|((~g14452));
assign g20601 = ((~g17433));
assign g8075 = ((~g3742));
assign g31485 = (g29776&g23421);
assign g24338 = (g23658)|(g18755);
assign g14061 = (g8715&g11834);
assign g25923 = (g24443&g19443);
assign g33174 = ((~g8714)&(~g32072));
assign g20078 = ((~g16846));
assign g25149 = (g14030&g23546);
assign g29495 = (g28563)|(g27614);
assign g6923 = ((~g3791));
assign g33502 = (g32758&II31206&II31207);
assign g24776 = ((~g3040))|((~g23052));
assign II31116 = (g31154&g31816&g32622&g32623);
assign g15090 = ((~g13144)&(~g12862));
assign g30583 = (g19666&g29355);
assign g25004 = ((~g676)&(~g23324));
assign g13248 = ((~g9985))|((~g12399))|((~g9843));
assign g27676 = (g26377&g20627);
assign g30730 = (g26346&g29778);
assign g33374 = (g32289&g21221);
assign g6994 = ((~g4933));
assign g7450 = (g1277)|(g1283);
assign g32522 = ((~g30735));
assign g34443 = (g34385)|(g18545);
assign g23306 = ((~g20924));
assign g27999 = (g23032&g26200&g26424&g25529);
assign g23088 = ((~II22240));
assign g21297 = ((~II21042));
assign g26769 = ((~g25400));
assign g32181 = (g31020&g19912);
assign g17619 = ((~g10179)&(~g12955));
assign g32739 = ((~g30735));
assign g34737 = ((~g34706)&(~g30003));
assign g21882 = (g4057&g19801);
assign g23453 = ((~II22576));
assign g31144 = (g29477)|(g28193);
assign II12199 = ((~g6215));
assign g7158 = ((~g5752)&(~g5712));
assign g21417 = ((~g11677))|((~g17157));
assign g8757 = ((~II12746));
assign g30007 = (g29141&g12929);
assign g30062 = (g13129&g28174);
assign g12196 = ((~g8764))|((~g4688));
assign g14582 = ((~II16698));
assign g16238 = ((~g4698))|((~g13883))|((~g12054));
assign g21285 = (g7857&g16027);
assign g22833 = ((~g1193))|((~g19560))|((~g10666));
assign g26849 = (g2994&g24527);
assign g34792 = (g34750)|(g18569);
assign g28533 = (g27291)|(g26203);
assign g25648 = (g24644)|(g21741);
assign g18638 = (g3827&g17096);
assign g19857 = ((~g13628))|((~g16296));
assign II19012 = ((~g15060));
assign g18529 = (g2712&g15277);
assign g33724 = (g14145&g33258);
assign g24099 = ((~g20720));
assign g32655 = ((~g30614));
assign g28471 = (g27187&g12762&g21024&II26960);
assign g23195 = ((~g20136))|((~g37));
assign g9251 = ((~II13037));
assign g23795 = (g20203)|(g16884);
assign g25023 = ((~g22457));
assign g11514 = ((~g10295)&(~g3161)&(~g3155));
assign g14412 = ((~II16564));
assign g19488 = (g16965)|(g14148);
assign g34197 = ((~g33812));
assign g25180 = ((~g23529));
assign g17787 = ((~II18795));
assign g18448 = (g2153&g18008);
assign g29352 = (g4950&g28410);
assign g6985 = ((~g4669));
assign g16077 = ((~II17456));
assign II21969 = ((~g21370));
assign g13076 = ((~g7443)&(~g10741));
assign g7936 = ((~g1061));
assign g16194 = (g11547&g6782&g11640&II17529);
assign g20676 = ((~g14379))|((~g17287));
assign g21057 = ((~g15426));
assign g7991 = ((~g4878));
assign g16636 = (g5929&g14768);
assign g26752 = ((~g9397))|((~g25189));
assign II28458 = ((~g28443));
assign g10606 = ((~g10233));
assign g22013 = (g5802&g21562);
assign g7514 = ((~g6704));
assign g20054 = ((~g17328));
assign II29302 = ((~g29496))|((~g12121));
assign g8787 = ((~II12773));
assign g34098 = (g33744&g9104&g18957);
assign g32590 = ((~g31154));
assign g18585 = (g2960&g16349);
assign g29521 = (g1744&g28824);
assign g17508 = ((~II18443));
assign g28086 = (g27268)|(g18702);
assign g10828 = (g6888&g7640);
assign g20035 = ((~g16430));
assign g19387 = ((~g16431));
assign g8228 = ((~g3835));
assign g32952 = ((~g30937));
assign g32738 = ((~g31376));
assign g32926 = ((~g31376));
assign g11977 = ((~g8373))|((~g2476));
assign g34711 = ((~g34559));
assign g28103 = (g27696)|(g22097);
assign II24396 = ((~g23453));
assign g20628 = (g1046&g15789);
assign g27094 = (g25997&g16472);
assign g30043 = (g29106&g9392);
assign g33065 = (g32008)|(g22068);
assign II14650 = ((~g9340));
assign g29907 = (g2629&g29177);
assign II12808 = ((~g4322));
assign g11357 = ((~g8558)&(~g8561));
assign II28241 = ((~g28709));
assign II13498 = ((~g255))|((~II13497));
assign g18142 = (g577&g17533);
assign g14206 = (g8655&g11790);
assign g30044 = (g29174&g12944);
assign g9485 = ((~g1657))|((~g1624));
assign g25682 = (g24658)|(g18640);
assign g16123 = ((~g13530));
assign g8766 = ((~g572));
assign g34944 = ((~g34932));
assign g21957 = (g5390&g21514);
assign gbuf46 = (g5794);
assign g18306 = (g15074&g16931);
assign g28320 = (g27116)|(g15808);
assign g28527 = (g27286)|(g26182);
assign g20327 = ((~g15224));
assign g25916 = (g24432&g19434);
assign g26628 = ((~g8990)&(~g24732));
assign g33423 = (g32225&g29657);
assign g32484 = ((~g31566));
assign g11993 = ((~g1894))|((~g8302));
assign II13802 = ((~g6971));
assign g29890 = (g28419&g23355);
assign g34141 = (g33932&g23828);
assign g31804 = ((~g29385));
assign g30927 = (g29910&g24795);
assign g26392 = (g24745)|(g23050);
assign g7219 = ((~g4405));
assign g22937 = (g753&g20540);
assign g20129 = ((~g17328));
assign g31930 = (g31769)|(g22094);
assign g27162 = (g26171&g8259&g2208);
assign II29277 = ((~g29488))|((~g12081));
assign g28743 = (g27517)|(g16758);
assign g30310 = ((~g28830));
assign g18742 = (g5120&g17847);
assign g34405 = (g34183)|(g25103);
assign g27366 = ((~g8016)&(~g26636));
assign g23498 = (g20234&g12998);
assign g11401 = ((~g7593));
assign g28197 = (g27647&g11344);
assign g34812 = ((~II33024));
assign g30610 = ((~II28872));
assign II12288 = ((~g1484))|((~II12287));
assign g20565 = ((~g18008));
assign g9072 = ((~g2994));
assign II11691 = ((~g36));
assign g33050 = (g31974)|(g21930);
assign g30025 = (g28492&g23502);
assign g22030 = (g5909&g19147);
assign g24297 = (g4455&g22550);
assign g25953 = ((~g22756))|((~g24570))|((~g22688));
assign g18176 = (g732&g17328);
assign g11469 = ((~g650)&(~g9903)&(~g645));
assign g23423 = ((~g20871));
assign g32538 = ((~g31070));
assign g22057 = (g15159&g21611);
assign g19677 = ((~g17096));
assign g28140 = (II26643)|(II26644);
assign g26926 = (g26633)|(g18531);
assign g22025 = (g5905&g19147);
assign g19673 = ((~g16931));
assign g21813 = (g3590&g20924);
assign g24107 = ((~g20857));
assign g18153 = (g626&g17533);
assign g27765 = (g4146&g25886);
assign g8324 = ((~g2476));
assign g27278 = (g15786)|(g25921);
assign g28484 = (g27187&g10290&g21163&II26972);
assign II22400 = ((~g19620));
assign g34487 = (g34416&g18983);
assign g19670 = ((~g16897));
assign g21920 = (g5062&g21468);
assign g14820 = ((~g6307))|((~g12173))|((~g6315))|((~g12423));
assign g22857 = ((~g20739));
assign g9203 = ((~g3706))|((~g3752));
assign g18608 = (g15087&g16987);
assign g11833 = ((~g8026));
assign g30182 = ((~II28419));
assign II20985 = ((~g16300));
assign g7222 = ((~g4427));
assign g28700 = (g27454)|(g16668);
assign II13442 = ((~g262))|((~g239));
assign g19534 = (g15650)|(g13019);
assign g22720 = (g9253&g20619);
assign g34411 = (g34186)|(g25142);
assign g19407 = ((~g16268));
assign g34472 = ((~II32525));
assign g24537 = (g22626&g10851);
assign g24082 = ((~g19890));
assign g22665 = (g17174&g20905);
assign g24100 = ((~g20857));
assign g25746 = (g25217)|(g22063);
assign g25089 = (g23317&g20553);
assign g32472 = ((~g30825));
assign g27051 = ((~II25779));
assign g21560 = ((~g17873));
assign g31810 = ((~g29385));
assign g7680 = ((~g4108));
assign g8479 = ((~g3057));
assign g33566 = (g33356)|(g18390);
assign g18484 = (g2491&g15426);
assign g24731 = (g6519&g23733);
assign g25643 = (g24602)|(g21736);
assign g32207 = (g31221&g23323);
assign II32440 = ((~g34227))|((~II32439));
assign g25341 = ((~g22417))|((~g12047));
assign g30124 = (g28580&g21055);
assign g31896 = (g31242)|(g24305);
assign II26972 = (g25011&g26424&g22698);
assign g29507 = ((~g28353));
assign g21927 = (g5164&g18997);
assign g29035 = ((~g9321)&(~g28020));
assign g20161 = ((~g17732))|((~g17706))|((~g17670))|((~g14625));
assign II18479 = ((~g13041));
assign g16748 = ((~II17970));
assign II27941 = ((~g28803));
assign II15382 = ((~g9071));
assign g21331 = ((~g11402))|((~g17157));
assign g11430 = ((~g7617));
assign g9935 = ((~II13483));
assign g30370 = (g30135)|(g18440);
assign g22974 = ((~g20330));
assign II33149 = ((~g34900));
assign g10925 = (g7858&g956);
assign g22534 = (g8766&g21389);
assign g14627 = ((~g12553))|((~g12772));
assign II27570 = ((~g28262));
assign g23769 = ((~g19074));
assign II14827 = ((~g9686));
assign g34736 = ((~II32904));
assign g23511 = ((~II22640));
assign g32357 = (g29865)|(g31296);
assign g14659 = ((~g12646))|((~g12443));
assign g28118 = (g27821)|(g26815);
assign g27833 = ((~g21228))|((~g25282))|((~g26424))|((~g26190));
assign g33913 = (g23088&g33204&g9104);
assign g21851 = (g3901&g21070);
assign g28563 = (g11981&g27100);
assign g34433 = ((~II32470));
assign g7379 = ((~g2299));
assign g10609 = ((~g10111))|((~g9826));
assign g17327 = ((~II18310));
assign g8741 = ((~g4821));
assign g30936 = (g8830&g29916);
assign g17432 = ((~II18379));
assign g16633 = (g5196&g14921);
assign g18542 = (g2787&g15277);
assign g13476 = ((~g7503))|((~g11336))|((~g11869));
assign g23895 = ((~g19147));
assign g14191 = ((~g12381));
assign g24133 = ((~g19935));
assign g28047 = (g27676)|(g18160);
assign g10578 = ((~g7174))|((~g6058));
assign g16876 = (g14028)|(g11773)|(g11755);
assign g18310 = (g1333&g16931);
assign g13895 = ((~II16193));
assign g14791 = (g1146&g10909);
assign g27218 = (g25997&g16740);
assign g27058 = (g10323&g3522&g3530&g26264);
assign g29527 = (g28945&g22432);
assign g33330 = (g32211&g20588);
assign II18803 = (g13156&g11450&g6756);
assign g18494 = (g2527&g15426);
assign g24861 = (g3712&g23582&II24033);
assign g10831 = ((~g7690)&(~g7827));
assign g26598 = ((~g8990)&(~g13756)&(~g24732));
assign g11389 = ((~II14399))|((~II14400));
assign g33813 = ((~II31659));
assign g14211 = ((~g9779)&(~g10823));
assign g15149 = ((~g13745)&(~g12894));
assign II27385 = ((~g27438));
assign g14726 = ((~g10090)&(~g12166));
assign g20038 = ((~g17328));
assign g18664 = (g4332&g17367);
assign g23104 = (g661&g20248);
assign g7328 = ((~g2197));
assign g29702 = ((~g28395))|((~g13712));
assign g29855 = (g2287&g29093);
assign g30234 = (g28721&g23914);
assign g23930 = ((~g19147));
assign g8302 = ((~g1926));
assign g34146 = (g33788&g20091);
assign g17648 = ((~g15024));
assign g32640 = ((~g31154));
assign g33591 = (g33082)|(g18474);
assign g15611 = (g471&g13437);
assign g27374 = (g26519&g17478);
assign g34379 = (g26312)|(g34143);
assign g7424 = ((~g2465));
assign g18159 = (g671&g17433);
assign g16097 = ((~g13319))|((~g10998));
assign g19568 = (g1467&g15959);
assign g34645 = (g34556)|(g18786);
assign g17390 = ((~g14755));
assign g26103 = (g2185&g25100);
assign g12601 = ((~g9381)&(~g9311));
assign g29731 = (g2089&g29118);
assign g24986 = ((~g23590));
assign g34091 = (g22957&g9104&g33761);
assign g29085 = ((~g9694))|((~g27837));
assign II14773 = ((~g9581));
assign g11962 = ((~II14789))|((~II14790));
assign g22167 = ((~g19074));
assign g8355 = ((~II12534));
assign g22718 = ((~g20887));
assign II32161 = ((~g33791));
assign g18557 = (g2771&g15277);
assign g33430 = ((~g32421));
assign g30577 = (g26267&g29679);
assign II26989 = ((~g27277));
assign g19438 = ((~g16249));
assign II18487 = ((~g14611))|((~II18485));
assign g23876 = ((~g19074));
assign g14988 = ((~g10816)&(~g10812)&(~g10805));
assign g25874 = (g11118&g24665);
assign II12927 = ((~g4332));
assign g24541 = (g22626&g10851);
assign g10416 = ((~g10318));
assign g24647 = (g19903&g22907);
assign g28254 = (g7268&g1668&g27395);
assign g28657 = (g27562&g20606);
assign g11892 = ((~g7777))|((~g9086));
assign g34398 = (g7684&g34070);
assign g33464 = (g32484&II31016&II31017);
assign II13124 = ((~g2729));
assign g22550 = ((~II21922));
assign g33012 = (g32274)|(g18483);
assign g12818 = ((~g8792));
assign g34750 = (g34673&g19542);
assign g32139 = (g31601&g29960);
assign g12903 = ((~g10411));
assign g34308 = ((~g34088));
assign g25691 = (g24536)|(g21890);
assign g32280 = (g24790)|(g31225);
assign g22646 = ((~g19389));
assign II17675 = ((~g13394));
assign g7828 = ((~g4871));
assign g24190 = (g329&g22722);
assign g13852 = ((~g11320)&(~g8347));
assign g18497 = (g2541&g15426);
assign g27229 = (g26055&g16774);
assign II18414 = ((~g14359));
assign g24123 = ((~g21143));
assign g32722 = ((~g30937));
assign g17610 = ((~g15008));
assign g15751 = ((~g5591))|((~g14522))|((~g5666))|((~g14669));
assign g27445 = (g8038&g26314&g9187&g504);
assign g33695 = ((~g33187));
assign g25503 = (g6888&g22529);
assign g29617 = (g2024&g28987);
assign II21831 = ((~g19127));
assign g29335 = ((~g25540))|((~g28131));
assign g25467 = ((~g12432))|((~g22417));
assign g14574 = ((~g12256))|((~g6120));
assign g32961 = ((~g31376));
assign g29603 = (g2265&g29060);
assign g26824 = ((~g25298));
assign g13066 = ((~g4430))|((~g7178))|((~g10590));
assign g27359 = (g26488&g17416);
assign g16657 = ((~g3554))|((~g13730))|((~g3625))|((~g11576));
assign g9480 = ((~g559));
assign g29029 = (g14506&g25227&g26424&g27494);
assign g18697 = (g4749&g16777);
assign g13739 = ((~g11773))|((~g11261));
assign g33954 = (g33496)|(II31853)|(II31854);
assign g33298 = (g32158)|(g29622);
assign g22632 = (g19356&g19476);
assign g18123 = (g479&g16886);
assign g19477 = ((~g16431));
assign g19875 = ((~g13667))|((~g16316));
assign g34309 = (g13947&g34147);
assign g31752 = (g30104&g23928);
assign g25656 = (g24945)|(g18609);
assign g33959 = ((~II31878));
assign g19698 = ((~g16971));
assign g26602 = (g7487&g24453);
assign g28719 = (g27485)|(g16703);
assign g23813 = ((~g18997));
assign II22467 = ((~g19662));
assign g10474 = ((~g8841));
assign g32636 = ((~g31376));
assign g33936 = ((~II31820));
assign II12076 = ((~g979))|((~II12074));
assign g34172 = (g33795)|(g19914);
assign g17505 = ((~g14899));
assign g18514 = (g2629&g15509);
assign g7162 = ((~g4521));
assign g31759 = (g21291&g29385);
assign g30018 = ((~g28987));
assign g20184 = ((~g16770))|((~g13918))|((~g16719))|((~g13896));
assign g24545 = (g3333&g23285);
assign g31008 = ((~g30004)&(~g30026));
assign g31669 = ((~II29254))|((~II29255));
assign g27882 = ((~g21228))|((~g25307))|((~g26424))|((~g26213));
assign II18495 = (g14539)|(g14515)|(g14449);
assign g22850 = ((~g1536))|((~g19581))|((~g10699));
assign g26488 = ((~II25366));
assign g8470 = ((~II12605));
assign g32621 = ((~g31542));
assign g32892 = ((~g31021));
assign g32766 = ((~g31376));
assign g9460 = ((~g6154));
assign g12971 = ((~g9024))|((~g8977))|((~g10664));
assign g30290 = ((~g6682)&(~g29110));
assign II23998 = ((~g22182));
assign g29532 = (g1878&g28861);
assign g18665 = (g4584&g17367);
assign g33437 = ((~g31997)&(~g10275));
assign g33513 = (g32837&II31261&II31262);
assign g28827 = ((~g27837))|((~g7362))|((~g1862));
assign g31784 = (g30176&g24003);
assign g11773 = ((~g8883)&(~g4785));
assign g24840 = (g21419)|(g23996);
assign g28553 = (g27187&g10290);
assign g26890 = (g26630)|(g24196);
assign g19885 = ((~g17249));
assign g34528 = (g34305&g19617);
assign g34479 = (g34403&g18905);
assign g31119 = ((~g7898)&(~g29556));
assign g22298 = (g19997&g21012);
assign g23649 = ((~g18833));
assign g26292 = (g2689&g25228);
assign g16741 = ((~g3207))|((~g13765))|((~g3303))|((~g11519));
assign g17297 = ((~g2729))|((~g14291));
assign g18417 = (g2116&g15373);
assign g27557 = (g26549&g17774);
assign II16733 = ((~g12026));
assign g9797 = ((~g5441));
assign g33542 = (g33102)|(g18265);
assign II32800 = ((~g34582));
assign g26021 = (g9568&g25035);
assign g26685 = ((~g9264))|((~g25160));
assign g22037 = (g5941&g19147);
assign g27928 = ((~g26810));
assign g31884 = (g31290)|(g21778);
assign g15068 = ((~g6826)&(~g13416));
assign g34577 = (g24577&g34307);
assign II22114 = ((~g19935));
assign II24549 = (g5385&g5390&g9792);
assign g32250 = (g30598)|(g29351);
assign g28815 = (g27546)|(g16842);
assign g18643 = (g3849&g17096);
assign g15052 = ((~g12835)&(~g13350));
assign g10851 = ((~II14069));
assign g24051 = ((~g21127));
assign g29867 = (g1996&g29117);
assign g11191 = ((~g4776)&(~g4801)&(~g9030));
assign g13657 = (g7251)|(g10616);
assign g25105 = (g13973&g23505);
assign g33291 = (g32154)|(g13477);
assign g14454 = ((~II16613));
assign g32853 = ((~g30673));
assign g9831 = ((~g2269));
assign g28924 = (g17317&g25183&g26424&g27416);
assign g11471 = ((~g7626));
assign II21977 = ((~g7680))|((~II21976));
assign g23838 = ((~g18997));
assign g27509 = (g26023)|(g24640);
assign g10684 = (g7998&g411);
assign g30031 = (g29071&g10540);
assign g33364 = (g32264&g20921);
assign g28369 = (g27160)|(g25938);
assign g32035 = (g4176&g30937);
assign II31610 = ((~g33149));
assign g29845 = (g28375&g23291);
assign g28605 = (g27341)|(g26302);
assign g32169 = (g31014&g23046);
assign g19506 = ((~g4087))|((~g15825));
assign g27261 = (g24544)|(g25996);
assign g9636 = ((~g72));
assign g25612 = (g24941)|(g18132);
assign g21059 = ((~g15509));
assign g24410 = (g3817&g23139);
assign g27686 = (g1291&g25849);
assign g6848 = ((~g2417));
assign g24025 = ((~g21256));
assign g24350 = (g23755)|(g18806);
assign g20574 = ((~g17847));
assign g29874 = (g28402&g23336);
assign g12672 = ((~g10003));
assign g28662 = (g27407)|(g16612);
assign g17519 = ((~II18460));
assign g11546 = (g7289&g4375);
assign II31092 = (g32589&g32590&g32591&g32592);
assign g27282 = ((~g11192))|((~g26269))|((~g26248))|((~g479));
assign g33243 = (g32124&g19947);
assign g32838 = ((~g31376));
assign g29718 = (g28512&g11136);
assign g31771 = ((~II29337));
assign g19572 = (g17133)|(g14193);
assign g32427 = (g8928)|(g30583);
assign g22170 = ((~g19210));
assign g30415 = (g29843)|(g21799);
assign g18802 = (g6195&g15348);
assign g7650 = ((~g4064));
assign g24564 = (g23198&g21163);
assign g17693 = (g1306&g13291);
assign g9961 = ((~g6404));
assign g25771 = ((~II24920));
assign g21992 = (g5599&g19074);
assign g11111 = (g5297&g7004&g5283&g9780);
assign g26720 = ((~g25275));
assign g23184 = (g20198)|(g20185)|(II22280);
assign g12873 = ((~g10380));
assign g17711 = ((~II18694));
assign g19519 = ((~g16795));
assign g28833 = (g21434&g26424&g25388&g27469);
assign II18191 = ((~g14385));
assign g12867 = ((~g10375));
assign g8507 = ((~g3712));
assign g28037 = ((~g26365));
assign g18355 = (g1748&g17955);
assign g9354 = ((~g2719));
assign g10318 = ((~g25)&(~g22));
assign g25491 = (g23615&g21355);
assign g9245 = ((~II13031));
assign g10929 = ((~g1099))|((~g7854));
assign g31976 = (g31762&g22178);
assign g22226 = (g21333)|(g17655);
assign g30111 = (g28565&g20917);
assign g20666 = ((~g15224));
assign g33923 = ((~II31791));
assign g34804 = (g34740)|(g18591);
assign g13970 = ((~g8883)&(~g8796)&(~g11155));
assign g33832 = (g33088&g27991);
assign g14956 = ((~g12604))|((~g10281));
assign II18165 = ((~g13177));
assign g13291 = ((~g10715))|((~g1500));
assign g30483 = (g30241)|(g21979);
assign g22339 = ((~g19801));
assign g34589 = ((~II32675));
assign g32241 = (g31244&g20323);
assign g28198 = (g26649&g27492);
assign g17813 = ((~II18813));
assign g32751 = ((~g31327));
assign g11144 = (g239&g8136&g246&II14198);
assign g18530 = (g2715&g15277);
assign g26541 = (g319&g24375);
assign g25262 = ((~g22763));
assign g23405 = (g19791)|(g16245);
assign g15111 = (g4281&g14454);
assign g33661 = ((~II31497));
assign II12240 = ((~g1111))|((~g1105));
assign II31222 = (g32775&g32776&g32777&g32778);
assign g34081 = (g33706&g19552);
assign g13459 = ((~g7479))|((~g11294))|((~g11846));
assign g21931 = (g5188&g18997);
assign g32469 = ((~g30673));
assign g33807 = (g33112&g25452);
assign g23029 = ((~g20453));
assign g24494 = ((~g23513)&(~g23532));
assign g16199 = (g3614&g14051);
assign II24003 = (g8097&g8334&g3045);
assign g20784 = ((~g14616))|((~g17595));
assign g17418 = (g9618&g14407);
assign g12151 = ((~g8316))|((~g8211));
assign g16304 = ((~g4765))|((~g13970))|((~g12054));
assign g24839 = ((~g23436));
assign g15171 = ((~II17098));
assign g24395 = (g4704&g22845);
assign II17970 = ((~g4027));
assign g9902 = ((~g100));
assign g14395 = ((~g12118)&(~g9542));
assign g27450 = (g2917)|(g26483);
assign g17638 = ((~g14838));
assign g15581 = ((~g7232))|((~g12999));
assign g14113 = ((~g11626))|((~g11537));
assign g29929 = ((~g28914));
assign g20854 = ((~g5381)&(~g17243));
assign g7469 = (g4382&g4438);
assign g18104 = (g392&g17015);
assign g17727 = ((~g12486)&(~g12983));
assign g19433 = ((~g15915));
assign g29649 = (g2241&g28678);
assign g26099 = (g24506)|(g22538);
assign g33080 = ((~II30644));
assign g24929 = (g23751&g20875);
assign g13672 = ((~g8933))|((~g11261));
assign g23060 = ((~g19908));
assign g18103 = (g401&g17015);
assign g18447 = (g2208&g18008);
assign g18507 = (g2595&g15509);
assign g26863 = (g24974&g24957);
assign g8462 = ((~g1183));
assign g11790 = ((~II14630));
assign g24785 = (g7051&g23645);
assign g7251 = (g452&g392);
assign II17406 = ((~g1472))|((~II17404));
assign g24912 = (g23687&g20682);
assign g33495 = (g32707&II31171&II31172);
assign g31472 = (g29642)|(g28352);
assign g26339 = (g225&g24836);
assign g24206 = (g23386)|(g18110);
assign II12251 = ((~g1124))|((~g1129));
assign II18882 = ((~g16580));
assign g30446 = (g29788)|(g21855);
assign g10311 = ((~g4633));
assign g30303 = ((~g28786));
assign g15721 = ((~g7564))|((~g311))|((~g13385));
assign g31528 = (g19050&g29814);
assign g23521 = ((~g21468));
assign g34014 = (g33647)|(g18493);
assign g8863 = (g1644)|(g1664);
assign g24361 = ((~g22885));
assign g29212 = ((~II27552));
assign g17427 = ((~II18364));
assign g10133 = ((~g6049));
assign g14803 = ((~g5208))|((~g12059))|((~g5308))|((~g12497));
assign g26804 = ((~g25400));
assign g27206 = (g26055&g16691);
assign g21966 = (g5406&g21514);
assign g14407 = ((~g12008))|((~g9807));
assign g7149 = ((~g4564));
assign g22121 = (g6593&g19277);
assign g13461 = (g2719&g11819);
assign g27155 = ((~g26131));
assign II11701 = ((~g4164));
assign g33681 = (g33129&g7991);
assign g28343 = (g27380&g19799);
assign g22087 = (g6303&g19210);
assign g15039 = ((~g12755))|((~g7142));
assign g16854 = ((~g3965))|((~g13824))|((~g3976))|((~g8595));
assign g25115 = ((~II24281));
assign g23502 = ((~g21070));
assign g20918 = ((~g15224));
assign g30330 = ((~II28591));
assign II15289 = ((~g6697))|((~II15287));
assign g30492 = (g30188)|(g21988);
assign g32883 = ((~g30735));
assign g7289 = ((~g4382));
assign g13137 = ((~g10699))|((~g7675))|((~g1322))|((~g1404));
assign g8239 = ((~g1056));
assign g9629 = ((~g6462))|((~g6466));
assign g25322 = ((~II24497));
assign g23486 = ((~g20785));
assign II14505 = ((~g10140));
assign g15719 = ((~g5256))|((~g14490))|((~g5335))|((~g9780));
assign II31539 = ((~g33212));
assign g33041 = (g32189)|(g24323);
assign g27660 = (g24688&g26424&g22763);
assign g8164 = ((~g3484));
assign g25597 = (g24892)|(g21719);
assign g13313 = (g475&g11048);
assign II24704 = (g21193&g24061&g24062&g24063);
assign g18822 = (g6723&g15680);
assign g29174 = ((~g9511)&(~g28020));
assign g12185 = ((~g9905))|((~g799));
assign g12110 = ((~II14970));
assign g34042 = ((~g33674));
assign g22840 = ((~g20330));
assign g17363 = ((~g8635))|((~g14367));
assign g19545 = (g3147&g16769);
assign g24193 = (g336&g22722);
assign g11251 = ((~g8438))|((~g3092));
assign g23440 = ((~II22557));
assign g15140 = ((~g12887)&(~g13680));
assign g23527 = ((~g21611));
assign II17374 = ((~g13638));
assign g27106 = (g26026&g16512);
assign g12377 = ((~g6856)&(~g2748)&(~g9708));
assign g32442 = ((~g31213));
assign g28608 = ((~g27670));
assign II14185 = ((~g8442))|((~g3470));
assign g10037 = ((~g1848));
assign II14702 = ((~g7717));
assign g32561 = ((~g30614));
assign g11952 = ((~g1624))|((~g8187));
assign g27532 = (g16176)|(g26084);
assign g16628 = ((~g3602))|((~g11207))|((~g3618))|((~g13902));
assign g7513 = ((~g6315));
assign g25782 = (g2936&g24571);
assign g12049 = ((~g2208))|((~g8150));
assign g20535 = ((~g17847));
assign g28030 = (g24018)|(g26874);
assign II17542 = (g13156&g6767&g6756);
assign g11154 = ((~II14212))|((~II14213));
assign g23537 = ((~g20785));
assign II30861 = ((~g32383));
assign II13850 = ((~g862))|((~g7397));
assign g26780 = (g4098&g24437);
assign g19915 = ((~g16349));
assign II27529 = (g28038&g24121&g24122&g24123);
assign II20447 = ((~g16244));
assign II29270 = ((~g29486))|((~II29269));
assign g21052 = ((~g15373));
assign g23296 = (g19691)|(g16177);
assign g32107 = (g31624&g29912);
assign g30437 = (g29876)|(g21846);
assign g6755 = ((~II11620));
assign g26827 = ((~g24819));
assign II26368 = ((~g14211))|((~II26366));
assign g26092 = (g9766&g25083);
assign g30345 = (g29644)|(g18302);
assign g21658 = ((~g17694)&(~g17727));
assign g34757 = (g34682&g19635);
assign II31151 = (g30825&g31822&g32673&g32674);
assign g17598 = ((~g3949))|((~g13824))|((~g4027))|((~g8595));
assign g31761 = (g30009)|(g30028);
assign g21406 = ((~g17955));
assign g30607 = (g30291&g18989);
assign g17140 = (g8616&g12968);
assign g29150 = ((~g27886));
assign g26833 = (g2852&g24509);
assign g18333 = (g1691&g17873);
assign g27825 = ((~g9316)&(~g25821));
assign g33734 = (g7806&g33136&II31593);
assign g32220 = (g31139)|(g29633);
assign g15872 = (g9095&g14234);
assign g22076 = (g6255&g19210);
assign g8105 = ((~g3068))|((~g3072));
assign g20237 = ((~g17213));
assign g23444 = ((~II22561));
assign g24795 = ((~g23342));
assign g29962 = (g23616&g28959);
assign g18785 = (g5849&g18065);
assign g19601 = (g16198&g11149);
assign II16102 = ((~g10430));
assign g26131 = ((~II25161));
assign g7595 = ((~II12067));
assign g34418 = ((~g34150));
assign g30257 = (g28750&g23952);
assign g25689 = (g24849)|(g21888);
assign g21510 = ((~g15647));
assign g9680 = ((~II13276));
assign g24707 = (g13295&g22997);
assign g15707 = (g4082&g13506);
assign II14730 = ((~g7717));
assign g31187 = (g10118&g30090);
assign g30395 = (g29841)|(g21754);
assign g26805 = (g10776)|(g24478);
assign g21462 = ((~g17816))|((~g14871))|((~g17779))|((~g14829));
assign g9982 = ((~g3976));
assign g19715 = (g9679&g17120);
assign g8807 = ((~g79));
assign g28626 = (g27542&g20573);
assign g18348 = (g1744&g17955);
assign g27669 = (g26840&g13278);
assign g34333 = (g9984&g34192);
assign g32359 = (g29867)|(g31298);
assign g17220 = ((~g9369))|((~g9298))|((~g14376));
assign II12061 = ((~g562));
assign g8534 = ((~g3338));
assign g32344 = (g29804)|(g31266);
assign g12308 = ((~g9951)&(~g9954));
assign g32761 = ((~g30825));
assign g9964 = ((~g126));
assign g21877 = (g6888&g19801);
assign g26361 = (g24674)|(g22991);
assign g32685 = ((~g31528));
assign g16219 = ((~g13498)&(~g4760));
assign g30360 = (g30145)|(g18386);
assign g10893 = ((~g1189)&(~g7715)&(~g7749));
assign g21945 = (g5248&g18997);
assign g10793 = ((~g1389)&(~g7503));
assign g17600 = ((~g14659));
assign g16163 = (g14254&g14179);
assign g33789 = (g33159&g23022);
assign g18199 = (g832&g17821);
assign g34606 = (g34564)|(g15080);
assign g18388 = (g1968&g15171);
assign II31241 = (g30825&g31838&g32803&g32804);
assign g14631 = ((~g12239));
assign II32953 = ((~g34656));
assign g17176 = (g8616&g13008);
assign II22865 = ((~g12146))|((~II22864));
assign g33342 = (g32226&g20660);
assign g34594 = ((~II32690));
assign g25883 = (g13728&g24699);
assign g27211 = (g25997&g16716);
assign g27285 = (g9912&g26632);
assign g8663 = ((~g3343));
assign g7615 = ((~II12083));
assign g7592 = ((~g347));
assign g26945 = (g26379)|(g24283);
assign g34263 = (g34078)|(g18699);
assign g10273 = ((~II13708));
assign g24715 = (g22189)|(g22207);
assign g17712 = ((~g5599))|((~g14425))|((~g5666))|((~g12301));
assign g29258 = (g28238)|(g18601);
assign II30686 = ((~g32381));
assign g12598 = ((~g7004));
assign g33704 = (g33176&g10710&g22319);
assign g20272 = ((~g17239));
assign g29233 = (g28171)|(g18234);
assign g28236 = (g8515&g27971);
assign g29210 = ((~II27546));
assign g29287 = (g28555)|(g18760);
assign g23322 = ((~II22425));
assign II32654 = ((~g34378));
assign g25575 = (g24139)|(g24140);
assign g33639 = (g33386&g18829);
assign g19860 = ((~g17226));
assign g10504 = ((~g8763));
assign g31280 = (g29717&g23305);
assign g7971 = ((~g4818));
assign g12341 = ((~g7512))|((~g5308));
assign II22464 = ((~g21222));
assign g28388 = (g27204)|(g15859);
assign g28588 = (g27489&g20499);
assign g28495 = (g27012&g12465);
assign g26914 = (g25949)|(g18227);
assign II32464 = ((~g34245));
assign g25661 = (g24754)|(g21786);
assign g21305 = ((~g15758));
assign g12967 = ((~g11790));
assign g18139 = (g542&g17249);
assign g8905 = (g2204)|(g2223);
assign g8630 = ((~g4843));
assign g7148 = ((~II11835));
assign g34579 = ((~II32659));
assign g28596 = (g27336)|(g26291);
assign g29640 = (g28498&g8125);
assign II11740 = ((~g4519));
assign g25626 = (g24499)|(g18235);
assign g29942 = ((~g28867));
assign g23578 = ((~II22725));
assign II18609 = ((~g5976));
assign g33127 = ((~g31950));
assign g21513 = (g16196&g10882);
assign g28302 = (g23809&g27817);
assign g26913 = (g25848)|(g18225);
assign g20672 = ((~g15277));
assign II32158 = ((~g33791));
assign g10383 = ((~g6978));
assign g34253 = (g34171)|(g24300);
assign II18765 = (g13156&g11450&g11498);
assign g21839 = (g3763&g20453);
assign g22670 = (g20114&g9104);
assign g28723 = (g27490)|(g16706);
assign g16743 = ((~g13986));
assign g18885 = ((~g15979));
assign g8277 = ((~II12483));
assign g7913 = ((~g1052));
assign g27436 = (g26576&g17588);
assign g25976 = (g9443&g25000);
assign g18372 = (g1886&g15171);
assign g13021 = ((~g7544)&(~g10741));
assign g20909 = ((~g17955));
assign II32388 = ((~g34153));
assign g29804 = (g1592&g29014);
assign g29070 = ((~g5857)&(~g7766)&(~g28020));
assign g32115 = (g31631&g29928);
assign g24150 = ((~g19268));
assign g17609 = ((~g14817));
assign g11939 = (g2361&g7380);
assign g10544 = ((~II13906));
assign g24171 = ((~II23357));
assign g16730 = (g5212&g14723);
assign g14377 = ((~g12201));
assign g14675 = ((~g12317))|((~g9898));
assign g25993 = (g2610&g25025);
assign g17651 = ((~g14868));
assign g6803 = ((~g496));
assign g25164 = (g16883&g23569);
assign g22201 = ((~g19277));
assign g14367 = ((~g9547)&(~g12289));
assign g11172 = ((~g8478))|((~g3096));
assign g18464 = (g2370&g15224);
assign II22901 = ((~g21228))|((~II22899));
assign g33524 = (g32918&II31316&II31317);
assign g8399 = ((~g3798));
assign g7441 = ((~g862));
assign g30246 = (g28734&g23936);
assign g32188 = (g27586&g31376);
assign g20375 = (g671&g16846);
assign g24275 = (g23474)|(g18645);
assign g23282 = ((~g20330));
assign II17392 = ((~g13680));
assign g23940 = ((~g19074));
assign II31311 = (g30673&g31851&g32903&g32904);
assign g29566 = (g2307&g28907);
assign g23616 = ((~II22754))|((~II22755));
assign II31027 = (g32494&g32495&g32496&g32497);
assign g10528 = (g1576&g9051);
assign g13869 = ((~g10831));
assign g8925 = ((~II12910));
assign g10197 = ((~g31));
assign II31062 = (g32545&g32546&g32547&g32548);
assign g16765 = (g6581&g15045);
assign g32813 = ((~g31710));
assign g17123 = (g225&g13209);
assign g21907 = (g5033&g21468);
assign g23935 = ((~g19210));
assign g20000 = ((~g13661)&(~g16264));
assign g26908 = (g26358)|(g24225);
assign g22624 = (g19344&g19471);
assign II19719 = ((~g17431));
assign g33624 = (g33371)|(g18808);
assign g16622 = ((~g14104));
assign II14853 = ((~g9433))|((~g5142));
assign II20891 = ((~g17700));
assign g13483 = ((~g11270));
assign g27132 = (g26055&g16589);
assign g19413 = ((~g17151)&(~g14221));
assign g12628 = ((~g7074))|((~g6336))|((~g6390));
assign II18671 = (g13156&g11450&g6756);
assign g25197 = ((~g23958));
assign g7733 = ((~g4093));
assign g25452 = ((~g22228));
assign g33973 = (g33840)|(g18344);
assign g13506 = ((~g10808));
assign g33579 = (g33357)|(g18437);
assign g23530 = ((~g20248));
assign g25061 = (g17586&g23461);
assign g33427 = ((~g10278)&(~g31950));
assign g10971 = ((~g7867))|((~g7886));
assign g33402 = (g32351&g21395);
assign g17955 = ((~II18865));
assign g13281 = ((~g10916))|((~g1099));
assign II27253 = ((~g27996));
assign g27554 = ((~g26625));
assign g6982 = ((~g4531));
assign g28478 = (g27007&g12345);
assign g12842 = ((~g10355));
assign g16751 = (g13155&g13065);
assign g34565 = (g34374&g17471);
assign g21177 = ((~II20957));
assign II18245 = ((~g14676));
assign II22748 = ((~g19458));
assign g20591 = ((~g15509));
assign II15214 = ((~g1714))|((~II15212));
assign g19400 = ((~g17139)&(~g14206));
assign g31917 = (g31478)|(g22003);
assign II13564 = ((~g2648))|((~g2652));
assign g30999 = ((~g29722));
assign g21900 = (g20977)|(g15114);
assign g24044 = ((~g21127));
assign II31192 = (g32733&g32734&g32735&g32736);
assign g14334 = ((~g12044)&(~g9337));
assign g34205 = (g33729&g24541);
assign g17487 = ((~II18414));
assign g27402 = ((~II26100));
assign g23916 = ((~g19277));
assign g14072 = ((~g11571))|((~g11483));
assign g28200 = (g27652&g11383);
assign g25668 = (g24646)|(g18623);
assign II15862 = ((~g11215));
assign g12854 = ((~g6849)&(~g10430));
assign g16750 = ((~g14454));
assign g22448 = ((~g1018)&(~g19699));
assign g27348 = (g26488&g17392);
assign g16721 = ((~g14072));
assign g13778 = (g4540&g10597);
assign g19790 = ((~g16971));
assign II22846 = ((~g21228))|((~II22844));
assign g34213 = (g33766&g22689);
assign II33267 = ((~g34979));
assign g31782 = (g30060)|(g30070);
assign g32473 = ((~g31070));
assign g21394 = (g13335&g15799);
assign g13508 = (g9927&g11888);
assign g12286 = ((~II15129))|((~II15130));
assign g28191 = (g27217)|(g27210)|(g27186)|(g27162);
assign g29711 = (g2541&g29134);
assign II31593 = (g31003&g8350&g7788);
assign gbuf107 = (g4188);
assign g30592 = (g30270&g18929);
assign g31877 = (g31278)|(g21732);
assign g29310 = ((~g28991));
assign II19671 = ((~g15932));
assign g17589 = ((~g14981));
assign g22495 = ((~g19801));
assign g20653 = ((~II20747));
assign g10948 = (g7880&g1478);
assign g14974 = ((~g12744))|((~g12622));
assign g17475 = ((~II18398));
assign g29954 = (g2299&g28796);
assign g21980 = (g5567&g19074);
assign g29207 = (g24131&II27533&II27534);
assign g32612 = ((~g30614));
assign II17747 = ((~g13298));
assign II31257 = (g32826&g32827&g32828&g32829);
assign II18071 = ((~g13680));
assign II24625 = (g6428&g6434&g10014);
assign g25296 = ((~g23745));
assign g18597 = (g2975&g16349);
assign g33618 = (g33353)|(g18757);
assign g34972 = ((~II33232));
assign g27074 = ((~II25790));
assign g34747 = (g34671&g19527);
assign g7655 = ((~g4332));
assign g29707 = ((~g28504));
assign II17474 = ((~g13336))|((~g1105));
assign g18573 = (g2898&g16349);
assign gbuf2 = (g4537);
assign g23076 = (g19128&g9104);
assign g9835 = ((~g2629)&(~g2555));
assign g30439 = (g29761)|(g21848);
assign g34238 = (g32780)|(g33956);
assign g18436 = (g2227&g18008);
assign g17929 = ((~II18855));
assign II23680 = ((~g23219));
assign II15162 = ((~g10176));
assign g22050 = (g6088&g21611);
assign g16717 = ((~g13951));
assign g32968 = ((~g31376));
assign g22116 = (g6589&g19277);
assign g27924 = ((~g9946)&(~g25839));
assign g30560 = (g30278)|(g22131);
assign g28040 = ((~g26365));
assign g31831 = ((~g29385));
assign g25757 = (g25132)|(g22104);
assign g26270 = (g1700&g25275);
assign g11970 = ((~g1760))|((~g8241));
assign g23614 = ((~g20248));
assign g31925 = (g31789)|(g22061);
assign g16584 = ((~g13920));
assign II32119 = ((~g33648));
assign II18589 = ((~g14679))|((~II18587));
assign g33352 = (g32237&g20712);
assign g9049 = ((~g640));
assign g17786 = (g1489&g13216);
assign g24972 = ((~g19962))|((~g23172));
assign g14308 = ((~II16471));
assign g13004 = ((~g7933)&(~g10741));
assign g27965 = (g25834&g13117);
assign g16931 = ((~II18101));
assign g30514 = (g30211)|(g22035);
assign g29662 = (g1848&g29049);
assign II23602 = ((~g4322))|((~II23600));
assign g32271 = (g31209)|(g29731);
assign g24419 = ((~g22722));
assign g31289 = (g29580)|(g29591);
assign g27629 = ((~g8891)&(~g26382)&(~g12259));
assign g29590 = (g2625&g28615);
assign II23987 = ((~g482))|((~II23985));
assign II27514 = (g24091&g24092&g24093&g24094);
assign g33339 = (g32221&g20634);
assign g13888 = (g2941)|(g11691);
assign g28454 = (g26976&g12233);
assign g30256 = (g28749&g23947);
assign g32902 = ((~g30673));
assign g29479 = (g28113)|(g28116);
assign g30271 = ((~g7041)&(~g29008));
assign g32420 = (g31127&g19533);
assign g23903 = ((~g18997));
assign II32594 = ((~g34298));
assign II22547 = ((~g20720));
assign II19484 = ((~g15122));
assign g18767 = (g15150&g17929);
assign g13211 = (g11294)|(g7567);
assign g12137 = ((~g6682)&(~g7097));
assign g10537 = ((~g7138))|((~g5366));
assign II18580 = ((~g1945))|((~II18579));
assign g34232 = (g33451)|(g33944);
assign g22042 = (g5961&g19147);
assign g18907 = ((~g15979));
assign g34343 = ((~g34089));
assign g17512 = ((~g12983));
assign g16920 = ((~II18086));
assign g13926 = ((~II16217));
assign II25514 = ((~g25073));
assign g29077 = ((~g6555)&(~g26994));
assign g27576 = ((~g26081));
assign g34640 = (g34487)|(g18723);
assign g27245 = ((~g26209));
assign II26419 = ((~g14247))|((~II26417));
assign g20580 = ((~g17328));
assign g21710 = (g287&g20283);
assign g27302 = (g1848&g26680);
assign g16589 = ((~g14082));
assign g30185 = (g28640&g23838);
assign g19481 = ((~g16349));
assign g9206 = ((~g5164));
assign g32574 = ((~g31070));
assign g29377 = (g28132&g19387);
assign g27409 = (g26519&g17524);
assign g20149 = ((~g17091)&(~g14185));
assign II14932 = ((~g9901));
assign g10153 = ((~g2417));
assign g9599 = ((~g3310));
assign g7868 = ((~g1099));
assign g28109 = ((~g27051))|((~g25783));
assign g13114 = ((~g7528)&(~g10741));
assign g23801 = (g1448&g19362);
assign g34002 = (g33857)|(g18451);
assign g26356 = (g15581&g25523);
assign g24155 = ((~II23309));
assign g29359 = ((~g7528)&(~g28167));
assign g10530 = ((~g8922));
assign g18762 = (g5475&g17929);
assign g23546 = ((~g21611));
assign g30252 = ((~g7028)&(~g29008));
assign g29997 = ((~g29060));
assign g26212 = ((~g23837)&(~g25408));
assign II22031 = ((~g21387));
assign II33273 = ((~g34984));
assign II25576 = ((~g25296));
assign g31900 = (g31484)|(g21908);
assign g31017 = (g29479&g22841);
assign II33300 = ((~g35001));
assign g34932 = ((~g34914));
assign g12982 = (g12220)|(g9968);
assign g28067 = (g27309)|(g21827);
assign g11885 = ((~g7153)&(~g7167));
assign g31131 = (g2393&g30020);
assign g10582 = ((~g7116));
assign g26343 = (g1514)|(g24609);
assign g7975 = ((~g3040));
assign g34313 = ((~g34086));
assign II21291 = ((~g18273));
assign g26847 = (g2873&g24525);
assign g22138 = ((~g21370));
assign g12930 = ((~g12347));
assign g32377 = ((~g30984));
assign g20204 = ((~g16578));
assign g10376 = ((~g6923));
assign II19674 = ((~g15932));
assign g33520 = (g32888&II31296&II31297);
assign g16242 = ((~g13529)&(~g4961));
assign g32349 = (g29840)|(g31275);
assign g13284 = ((~g10695))|((~g1157));
assign g29516 = (g28895&g22369);
assign g7873 = ((~g1266));
assign II22872 = ((~g12150))|((~II22871));
assign g20618 = ((~g15277));
assign g32496 = ((~g30614));
assign II23360 = ((~g23360));
assign g26928 = (g26713)|(g18541);
assign g21971 = (g5417&g21514);
assign g18976 = ((~g16100));
assign g31502 = (g2472&g29311);
assign g27505 = (g26519&g17681);
assign g13513 = ((~g1351))|((~g11815))|((~g8002));
assign g32675 = ((~g31070));
assign g33718 = (g33147&g19432);
assign g28444 = ((~g8575)&(~g27463)&(~g24825));
assign g8954 = ((~g1079));
assign g32536 = ((~g31376));
assign g15079 = (g2151&g12955);
assign II16135 = ((~g10430));
assign g25707 = (g25041)|(g18749);
assign g32010 = (g31785&g22303);
assign g33451 = ((~g32132));
assign g31166 = (g1816&g30074);
assign g28568 = ((~g10323)&(~g27617));
assign II14584 = ((~g9766));
assign g28325 = ((~g27463));
assign g27220 = (g26026&g16743);
assign g20158 = ((~g16971));
assign g32669 = ((~g30614));
assign g22455 = ((~g19801));
assign g33446 = (g32385&g21607);
assign g29497 = ((~g22763)&(~g28241));
assign II31347 = (g32956&g32957&g32958&g32959);
assign g26888 = (g26671)|(g24194);
assign II29284 = ((~g29489))|((~g12085));
assign gbuf100 = (g4027);
assign g31941 = (g1283&g30825);
assign g33506 = (g32788&II31226&II31227);
assign II26296 = ((~g26820));
assign g8977 = ((~g4349));
assign g21976 = (g5527&g19074);
assign II11777 = ((~g5357));
assign g33393 = (g32286)|(g29984);
assign g14058 = ((~g7121))|((~g11537));
assign g13948 = ((~g11610))|((~g8864));
assign g30545 = (g30268)|(g22116);
assign g15833 = ((~g14714))|((~g12378))|((~g12337));
assign g20191 = ((~g17821));
assign g27698 = ((~g26648));
assign g33144 = ((~g4664)&(~g32057));
assign g16213 = (g6772&g6782&g11640&II17552);
assign g33855 = (g33265&g20441);
assign g26931 = (g26778)|(g18547);
assign II22823 = ((~g11978))|((~II22822));
assign g26918 = (g25931)|(g18243);
assign g17013 = ((~g14262));
assign g27691 = (g25778&g23609);
assign II12849 = ((~g4281))|((~II12848));
assign g34861 = (g16540&g34827);
assign g10905 = ((~g1116))|((~g7304));
assign II18813 = ((~g5673));
assign g15849 = (g3538&g14136);
assign II20222 = ((~g16272))|((~II20221));
assign II12279 = ((~g1472))|((~II12277));
assign g30447 = (g29798)|(g21856);
assign g34169 = (g33804&g31227);
assign g9386 = ((~g5727));
assign g22636 = (g18943)|(g15611);
assign g27550 = ((~g24943))|((~g25772));
assign g22457 = (g7753&g7717&g21288);
assign g13951 = ((~g10295))|((~g11729));
assign g14537 = (g10550&g10529);
assign g32097 = (g25960&g31021);
assign g20277 = ((~g16487));
assign g24015 = (g19540&g10951);
assign g34005 = (g33883)|(g18454);
assign g34359 = ((~g9162)&(~g34174)&(~g12259));
assign II23970 = ((~g22202))|((~II23969));
assign g12470 = ((~II15284));
assign g19069 = (g8397&g16186);
assign g31838 = ((~g29385));
assign g19694 = ((~g16429));
assign g31934 = (g31670&g18827);
assign II16521 = ((~g10430));
assign g33003 = (g32323)|(g18429);
assign g22124 = (g6613&g19277);
assign g30535 = (g30225)|(g22081);
assign g34327 = ((~g34108));
assign g34496 = ((~g34370)&(~g27648));
assign g20912 = ((~g15171));
assign g33960 = (g33759)|(g21701);
assign g18249 = (g1216&g16897);
assign g17302 = ((~II18285));
assign g29741 = (g28205)|(g15883);
assign g21454 = ((~g15373));
assign g34966 = (g34950&g23170);
assign g32268 = (g24785)|(g31219);
assign g7903 = ((~g969));
assign g27257 = (g25904)|(g24498);
assign g25456 = (g5752&g22210&II24579);
assign II26742 = (g23430)|(g23445)|(g23458)|(g23481);
assign g20159 = ((~g17533));
assign II18849 = ((~g14290));
assign g33040 = (g32164)|(g24313);
assign g9500 = ((~g5495));
assign g33637 = ((~II31466));
assign g32175 = (g31709&g27858);
assign g33531 = (g32967&II31351&II31352);
assign g33887 = (g33298&g20615);
assign g14601 = ((~g12318))|((~g6466));
assign g22155 = ((~g19074));
assign g19800 = ((~g17096));
assign g24166 = ((~II23342));
assign g7096 = ((~g6537));
assign g33527 = (g32939&II31331&II31332);
assign g10364 = ((~g6869));
assign g32619 = ((~g30614));
assign g6987 = ((~g4754));
assign g9061 = ((~g3401)&(~g3361));
assign g23685 = ((~II22823))|((~II22824));
assign g26836 = ((~g24866));
assign g29482 = (g28524)|(g27588);
assign g20494 = ((~g17847));
assign g34852 = ((~g34845));
assign II14817 = ((~g9962))|((~II14816));
assign g13762 = (g499)|(g12527);
assign g12045 = ((~g1783))|((~g8146));
assign II15633 = ((~g12074));
assign g25925 = (g24990&g23234);
assign g18522 = (g2671&g15509);
assign g13323 = ((~g11048));
assign g31013 = ((~g29679));
assign g12795 = (g1312&g7601);
assign II28566 = (g29201)|(g29202)|(g29203)|(g28035);
assign g24653 = (g2848)|(g22585);
assign g32725 = ((~g30825));
assign g11047 = (g6474&g9212);
assign II27713 = ((~g28224));
assign g18711 = (g15136&g15915);
assign g27460 = (g26549&g17610);
assign g33219 = (g32335)|(II30760)|(II30761);
assign g32014 = (g8715&g30673);
assign II33024 = ((~g34783));
assign g18982 = (g3835&g16159);
assign g27700 = (g22342&g25182&g26424&g26148);
assign g33683 = (g33149&g10727&g22332);
assign g34619 = (g34528)|(g18581);
assign II14690 = ((~g9340));
assign g31823 = ((~g29385));
assign II13020 = ((~g6750));
assign g24232 = (g22686)|(g18228);
assign g27114 = (g25997&g16523);
assign g14257 = (g8612&g11878);
assign II17636 = ((~g14252));
assign g31492 = (g29790&g23431);
assign g30028 = (g29069&g9311);
assign II31102 = (g32603&g32604&g32605&g32606);
assign g27830 = ((~g26802));
assign g11214 = ((~g9602));
assign g18217 = (g15063&g16100);
assign g10627 = ((~II13968));
assign g18508 = (g2606&g15509);
assign g12453 = ((~g9444)&(~g5527));
assign g33379 = (g30984&g32364);
assign g18233 = (g1094&g16326);
assign g17413 = ((~II18350));
assign g33901 = (g33317&g20920);
assign g29633 = (g1978&g29085);
assign g25037 = (g23103)|(g19911);
assign g20434 = ((~g18065));
assign g28696 = ((~g27858));
assign g13667 = ((~g3723))|((~g11119));
assign g34504 = ((~g34408));
assign g28297 = (g27096)|(g15785);
assign g14768 = ((~g12662))|((~g12571));
assign g34468 = (g34342)|(g18718);
assign g14066 = ((~g11514))|((~g11473));
assign g32511 = ((~g30614));
assign g30518 = (g30254)|(g22039);
assign g29294 = (g28645)|(g18779);
assign g25908 = (g24782&g22520);
assign g20587 = ((~g15373));
assign g15724 = ((~g13858)&(~g11374));
assign g13796 = ((~g9158)&(~g12527));
assign II31306 = (g30614&g31850&g32896&g32897);
assign g8899 = ((~g807));
assign g25399 = ((~g22763));
assign g17583 = ((~g14968));
assign g28258 = (g27182&g19687);
assign g31294 = ((~g11326)&(~g29660));
assign II14788 = ((~g9891))|((~g6167));
assign g24246 = (g23372)|(g18257);
assign g16689 = ((~g13923));
assign g12490 = ((~II15316));
assign g29004 = ((~g27933))|((~g8330));
assign g33089 = ((~g31978)&(~g4322));
assign g7138 = ((~g5360));
assign g18732 = (g4961&g16877);
assign g21209 = ((~g15483)&(~g9575));
assign II18233 = ((~g14639));
assign g10361 = ((~g6841));
assign g32275 = (g31210)|(g29732);
assign II12776 = ((~g4207));
assign g19344 = (g17771)|(g14832);
assign g25964 = (g1783&g24979);
assign g16772 = ((~g3558))|((~g13799))|((~g3654))|((~g11576));
assign g11270 = ((~g8431)&(~g8434));
assign g34354 = ((~g9003)&(~g34162)&(~g11083));
assign g11978 = (g2629&g7462);
assign g14562 = ((~g12036));
assign g21987 = (g5579&g19074);
assign II26427 = ((~g26859));
assign II17228 = ((~g13350));
assign g29279 = (g28442)|(g18741);
assign g33020 = (g32160)|(g21734);
assign II25356 = ((~g24374));
assign g10829 = (g7289&g4375);
assign gbuf73 = (g3267);
assign II29368 = ((~g30321));
assign II22822 = ((~g11978))|((~g21434));
assign g33356 = (g32245&g20772);
assign g10761 = ((~g8411));
assign g13515 = ((~g12628))|((~g12588))|((~g12524))|((~g12464));
assign g10122 = ((~II13623));
assign g28880 = (g21434&g26424&g25438&g27494);
assign II31491 = ((~g33283));
assign g31150 = (g1682&g30063);
assign g26121 = (g6167&g25111);
assign g29613 = (g28208&g19763);
assign g21806 = (g3558&g20924);
assign g15122 = ((~g6959)&(~g13605));
assign g17213 = ((~g11107)&(~g13501));
assign g28075 = (g27083)|(g21877);
assign g14522 = ((~g9924)&(~g12656));
assign g18725 = (g4912&g16077);
assign g7897 = ((~II12288))|((~II12289));
assign g31244 = (g25963)|(g29515);
assign g18244 = (g1171&g16431);
assign g28663 = (g27566&g20624);
assign g34106 = (g33917&g23675);
assign g13660 = (g8183)|(g12527);
assign g20213 = ((~g17062));
assign g29885 = (g28416&g23350);
assign g32251 = (g30599)|(g29352);
assign g34783 = (g33110)|(g34667);
assign g33997 = (g33871)|(g18427);
assign g12015 = (g1002&g7567);
assign g25134 = ((~g22417));
assign g21716 = (g301&g20283);
assign g16312 = ((~g13580))|((~g13574));
assign g13039 = ((~II15663));
assign g21674 = ((~g16540));
assign g34060 = ((~g33704));
assign g24578 = (g2882)|(g23825);
assign g34694 = (g34530&g19885);
assign g16706 = (g6621&g14868);
assign g12900 = ((~g10406));
assign g31653 = ((~g29713));
assign g11715 = ((~g8080)&(~g8026));
assign g30359 = (g30075)|(g18385);
assign g13850 = ((~g11279))|((~g8396));
assign g33517 = (g32867&II31281&II31282);
assign g24262 = (g23387)|(g18315);
assign g13728 = (g6804)|(g12527);
assign II13045 = ((~g5120))|((~II13043));
assign g12147 = ((~g8302))|((~g8201));
assign g16687 = ((~g3255))|((~g13700))|((~g3325))|((~g11519));
assign g32872 = ((~g31327));
assign g27517 = (g26400&g17707);
assign g6815 = ((~g929));
assign g21847 = (g3905&g21070);
assign g25549 = ((~g22763));
assign II28390 = ((~g29185));
assign g26119 = (g11944&g25109);
assign g24483 = ((~II23688));
assign II11866 = ((~g4401))|((~II11864));
assign g9713 = ((~g3618));
assign g19422 = ((~g16031)&(~g13141));
assign II31751 = ((~g33228));
assign g16527 = ((~g14048));
assign g12466 = ((~g10057)&(~g10059));
assign g28949 = ((~g27903))|((~g14643));
assign g13999 = ((~g11048));
assign g33258 = ((~g32296));
assign g28994 = ((~g27907))|((~g2495))|((~g7424));
assign II32693 = ((~g34433));
assign g13117 = ((~g10981));
assign II29236 = ((~g29498));
assign g26682 = ((~g25309));
assign g24568 = ((~g22942));
assign g29262 = (g28327)|(g18608);
assign g25769 = ((~g25453)&(~g25414));
assign g8114 = ((~g3522));
assign g23884 = (g4119&g19510);
assign II27314 = ((~g28009));
assign g25894 = (g24817)|(g23229);
assign g22340 = (g19605&g13522);
assign g22684 = (g19206)|(g15703);
assign II21222 = ((~g18091));
assign II31561 = ((~g33197));
assign g22100 = (g6466&g18833);
assign g11181 = ((~g8134));
assign g28053 = (g27393)|(g18168);
assign g31962 = (g8033&g31013);
assign g34777 = ((~II32973));
assign g19471 = ((~g16449));
assign II13979 = ((~g7733));
assign g22642 = ((~g7870))|((~g19560));
assign g26326 = ((~g24872));
assign g32149 = (g31658&g29983);
assign g34698 = ((~g34550));
assign g27490 = (g26576&g17651);
assign g25986 = (g5160&g25013);
assign g25930 = ((~II25028));
assign g22325 = ((~g1252))|((~g19140));
assign g23244 = ((~II22343));
assign g16422 = (g8216&g13627);
assign g17705 = ((~g3586))|((~g13799))|((~g3661))|((~g13902));
assign g23844 = ((~g21308));
assign g28287 = ((~g10504))|((~g26131))|((~g26973));
assign II31351 = (g30937&g31858&g32961&g32962);
assign g22928 = ((~II22131));
assign g14054 = ((~g3550))|((~g11238))|((~g3649))|((~g11576));
assign g10182 = ((~g2681));
assign g29182 = (g27163&g12730);
assign II31586 = ((~g33149));
assign g30440 = (g29771)|(g21849);
assign gbuf125 = (g859);
assign g24421 = (g3835&g23139);
assign g30175 = (g28629&g23813);
assign g16159 = ((~g13584));
assign II14400 = ((~g3654))|((~II14398));
assign g34709 = (g34549&g17242);
assign g10724 = (g3689&g8728);
assign g15695 = ((~g1266))|((~g13125));
assign g28373 = (g27180)|(g15849);
assign II33270 = ((~g34982));
assign g33315 = (g29665)|(g32175);
assign g34491 = ((~II32550));
assign g18886 = ((~g16000));
assign g32610 = ((~g31070));
assign g10981 = ((~II14119));
assign g27821 = (g7680&g25892);
assign g9906 = (g996&g1157);
assign II17380 = ((~g13336))|((~II17379));
assign g13217 = ((~g4082))|((~g10808));
assign g18341 = (g1648&g17873);
assign g16202 = (g86&g14197);
assign g17091 = (g8659&g12940);
assign g29036 = (g27163&g12762&g20875&II27381);
assign g24426 = ((~g22722));
assign g32527 = ((~g30673));
assign g32931 = ((~g30937));
assign II31814 = ((~g33149));
assign II22899 = ((~g12193))|((~g21228));
assign g32831 = ((~g31376));
assign g13915 = ((~g11566))|((~g11473));
assign II26785 = ((~g27013));
assign g13320 = (g417&g11048);
assign g28264 = (g7315&g1802&g27416);
assign II14211 = ((~g9252))|((~g9295));
assign g12039 = ((~II14899));
assign g18432 = (g2223&g18008);
assign g29629 = (g28211&g19779);
assign g32445 = ((~II29973));
assign g16651 = ((~g14005));
assign g34456 = (g34395)|(g18669);
assign g33343 = (g32227&g20665);
assign g8945 = ((~g608));
assign g30216 = (g28691&g23882);
assign g22757 = ((~g20114))|((~g7891));
assign g12079 = ((~g1792))|((~g8195));
assign g21420 = (g16093&g13596);
assign g21425 = ((~g15509));
assign II21019 = ((~g17325));
assign g26749 = (g24494&g23578);
assign II13077 = ((~g5462))|((~g5467));
assign g23642 = ((~g9733)&(~g21124));
assign g20168 = ((~g17533));
assign g34985 = ((~II33255));
assign g18692 = (g4732&g16053);
assign II32067 = ((~g33661));
assign g24664 = (g22652&g19741);
assign g20705 = ((~II20793));
assign g23229 = (g18994&g4521);
assign g26258 = (g12875&g25231);
assign g10059 = ((~g6451));
assign g26952 = (g26360)|(g24290);
assign g28074 = (g27119)|(g21876);
assign g33072 = ((~g31945));
assign g28462 = ((~g3512)&(~g27617));
assign g26960 = (g26258)|(g24304);
assign g10428 = ((~g9631));
assign g31888 = (g31067)|(g21821);
assign g24240 = (g22861)|(g18251);
assign g33950 = (g32450)|(g33460);
assign g26257 = (g4253&g25197);
assign g25802 = (g8106&g24586);
assign II11816 = ((~g93));
assign g27522 = (g26549&g17717);
assign II24054 = (g8443&g8075&g3747);
assign g11911 = ((~g10022));
assign g23004 = ((~g20283));
assign g17644 = ((~g15002));
assign II12910 = ((~g4340));
assign g16182 = ((~g13846));
assign g18680 = (g15128&g15885);
assign g18503 = (g2563&g15509);
assign g34678 = (g34490&g19431);
assign g28282 = (g23762&g27727);
assign g23336 = ((~g20924));
assign g18685 = (g4688&g15885);
assign g27976 = ((~g26703));
assign g10050 = ((~g6336));
assign g23222 = ((~g20785));
assign g26307 = (g13070&g25288);
assign II24679 = (g19968&g24026&g24027&g24028);
assign g12029 = ((~g5644)&(~g7028));
assign g13062 = ((~g10981));
assign g27140 = (g25885&g22593);
assign g26893 = (g26753)|(g24199);
assign g28310 = (g27107)|(g15797);
assign g7633 = ((~II12120));
assign g32573 = ((~g30825));
assign g33116 = (g32403)|(g32411);
assign g19711 = ((~g17062));
assign g27955 = ((~II26460))|((~II26461));
assign g15085 = ((~II17008));
assign g21176 = ((~II20954));
assign g25163 = (g20217&g23566);
assign g24573 = (g17198&g23716);
assign II15300 = ((~g1982))|((~II15298));
assign g31465 = (g26156)|(g29647);
assign g27354 = ((~g8064)&(~g26636));
assign g14936 = (g10776)|(g8703);
assign g20086 = ((~II20355));
assign g15157 = ((~g13782)&(~g12900));
assign g18170 = (g661&g17433);
assign g8639 = ((~g2807));
assign II29297 = ((~g12117))|((~II29295));
assign g24488 = (g6905&g23082);
assign II18734 = ((~g6373));
assign g33845 = ((~II31694));
assign g23966 = ((~g19210));
assign g34391 = ((~g34200));
assign g29044 = ((~g27742));
assign g28120 = ((~g27108));
assign g20643 = ((~g15962));
assign g33019 = (g32339)|(g18536);
assign g19649 = ((~g17015));
assign g25208 = ((~g22763));
assign g10281 = ((~g5535)&(~g5527));
assign g8539 = ((~g3454));
assign g27268 = (g25942&g19733);
assign g11872 = ((~II14684));
assign II33140 = ((~g34884));
assign g12895 = ((~g10403));
assign g8984 = ((~g4899)&(~g4975));
assign II12890 = ((~g4219));
assign II11820 = ((~g3869));
assign g22899 = (g19486&g19695);
assign g16673 = (g6617&g14822);
assign g12224 = ((~II15088))|((~II15089));
assign g26082 = (g2898)|(g24561);
assign g28272 = (g27721&g26548);
assign g23690 = (g14726&g20978);
assign g13174 = ((~g10741));
assign g11445 = ((~g9771))|((~g3976));
assign g33896 = (g33314&g20771);
assign g34038 = (g33731)|(g18735);
assign g20509 = ((~g15277));
assign gbuf49 = (g6329);
assign g24322 = (g4423&g22228);
assign II18530 = ((~g1811))|((~II18529));
assign g32500 = ((~g30735));
assign g32804 = ((~g30735));
assign g18065 = ((~II18875));
assign g24314 = (g4515&g22228);
assign g10203 = ((~g2393));
assign g9213 = ((~II13020));
assign g16666 = (g5200&g14794);
assign II17401 = ((~g13394));
assign g14441 = ((~II16590));
assign g33306 = ((~g776))|((~g32212))|((~g11679));
assign g34702 = (g34537&g20208);
assign g21163 = (g16321&g4878);
assign g19685 = ((~g16987));
assign g32364 = ((~II29894));
assign II32766 = ((~g34522));
assign g14005 = ((~g11514))|((~g11729));
assign g27324 = (g10150&g26720);
assign g32200 = (g27468&g31376);
assign II19756 = ((~g17812));
assign g22384 = (g9354&g9285&g20784);
assign II17188 = ((~g13782));
assign g8918 = ((~II12893));
assign g8396 = ((~g3401));
assign g25152 = (g23383&g20626);
assign II26406 = ((~g26187));
assign II13329 = ((~g86));
assign g17524 = ((~g14933));
assign g12687 = (g9024&g8977);
assign g10430 = ((~II13847));
assign g23991 = (g19209&g21428);
assign g18631 = (g3694&g17226);
assign II14925 = ((~g5835))|((~II14923));
assign II30735 = (g32369)|(g32376)|(g32089)|(g32035);
assign g33234 = (g32039)|(g32043);
assign g18756 = (g5348&g15595);
assign II23315 = ((~g21685));
assign g20108 = (g15508&g11048);
assign g21776 = (g3376&g20391);
assign g34525 = (g34297&g19528);
assign g12021 = ((~g9543));
assign II26356 = ((~g26843));
assign g13912 = (g5551&g12450);
assign g21434 = ((~g17248));
assign g12246 = ((~g9880)&(~g9883));
assign g13083 = ((~g4392))|((~g10590))|((~g4434));
assign g14885 = ((~g12651))|((~g12505));
assign g19462 = (g7850&g14182&g14177&g16646);
assign g14446 = ((~g12190)&(~g9644));
assign g27361 = (g26519&g17419);
assign g29794 = (g28342&g23256);
assign g28420 = (g27222)|(g13290);
assign g11371 = ((~g7565));
assign g17526 = ((~II18469));
assign g29221 = ((~II27579));
assign g28452 = ((~g3161)&(~g27602));
assign g32771 = ((~g31021));
assign g28335 = (g27132)|(g15818);
assign g10393 = ((~g6991));
assign II12135 = ((~g807));
assign g12100 = ((~II14956))|((~II14957));
assign gbuf66 = (g6715);
assign g29320 = (g29068&g22147);
assign II29986 = (g31070)|(g31194)|(g30614)|(g30673);
assign g32327 = (g31319&g23544);
assign g9775 = ((~g4831))|((~g4681));
assign g20525 = ((~g17955));
assign g8342 = ((~II12519));
assign g18565 = (g2852&g16349);
assign g34219 = (g33736&g22942);
assign g9558 = ((~g5841));
assign g7998 = ((~g392));
assign g26186 = (g24580&g23031);
assign g11691 = ((~II14570));
assign g32745 = ((~g31376));
assign g27016 = (g26821)|(g14585);
assign g24128 = ((~g20720));
assign g20092 = ((~g11373))|((~g17794));
assign g30231 = (g28718&g23907);
assign II19863 = ((~g16675));
assign g18223 = (g1030&g16100);
assign g32120 = (g31639&g29941);
assign g22919 = ((~g21163));
assign g10521 = ((~II13889));
assign g29259 = (g28304)|(g18603);
assign g15808 = (g3590&g14048);
assign II32433 = ((~g34051))|((~II32431));
assign g21140 = ((~g6073)&(~g17312));
assign g21730 = (g3025&g20330);
assign II25005 = ((~g24417));
assign g19732 = ((~g17096));
assign g14807 = ((~g7738))|((~g12453));
assign g27183 = (g26055&g16658);
assign II18131 = ((~g13350));
assign II23369 = ((~g23347));
assign II18674 = ((~g13101));
assign II14247 = ((~g1322))|((~g8091));
assign g20778 = ((~g15224));
assign II16057 = ((~g10430));
assign g24589 = (g5471&g23630);
assign g34409 = ((~g34145));
assign g33561 = (g33408)|(g18376);
assign II29314 = ((~g29501))|((~II29313));
assign g24942 = ((~g20039))|((~g23172));
assign g11127 = (g6479&g10022);
assign g24764 = (g17570&g22472);
assign g10816 = ((~II14054));
assign g23171 = (g19536)|(g15903);
assign g22988 = ((~g20391));
assign II24281 = ((~g23440));
assign g19415 = ((~g15758));
assign g32715 = ((~g31327)&(~II30261)&(~II30262));
assign g16532 = (g5252&g14841);
assign II25541 = ((~g25180));
assign g25996 = ((~g24601))|((~g22838));
assign g22589 = (g19267&g19451);
assign g24896 = (g22863)|(g19684);
assign g13013 = ((~g7957)&(~g10762));
assign g29937 = (g13044&g29196);
assign g15634 = ((~II17188));
assign g31233 = ((~g8522)&(~g29778)&(~g24825));
assign g16190 = (g14626&g11810);
assign g18992 = (g8341&g16171);
assign II11750 = ((~g4474));
assign g9585 = ((~g1616));
assign II31072 = (g32559&g32560&g32561&g32562);
assign g26809 = (g24930)|(g24939);
assign g27730 = ((~g26424));
assign g17770 = (g7863&g13189);
assign g25710 = (g25031)|(g21961);
assign g26300 = (g1968&g25341);
assign g30327 = ((~II28582));
assign II12403 = ((~g3813))|((~II12401));
assign g10408 = ((~g7049));
assign g27430 = (g26488&g17579);
assign g24224 = (g269&g22594);
assign g8677 = ((~g4854));
assign g26608 = ((~g25334));
assign g24287 = (g4401&g22550);
assign g22528 = ((~g19801));
assign g13329 = ((~II15893));
assign II13464 = ((~g2384))|((~II13462));
assign g18671 = (g4628&g15758);
assign g27294 = (g9975&g26656);
assign g15915 = ((~II17392));
assign g34256 = (g34173)|(g24303);
assign g15135 = ((~g6990)&(~g13638));
assign g26176 = (g1964&g25467);
assign g28677 = (g27571&g20635);
assign g12121 = ((~g10117)&(~g9762));
assign g30099 = (g28549&g20776);
assign g29243 = (g28657)|(g18358);
assign g23778 = ((~II22922))|((~II22923));
assign g32292 = (g31269&g20530);
assign g32395 = (g31523)|(g30049);
assign g24146 = ((~g19422));
assign g32505 = ((~g31566));
assign g13867 = ((~g11312))|((~g8449));
assign g31756 = (g30114&g23942);
assign g26959 = (g26381)|(g24299);
assign g25226 = ((~g22763));
assign g7534 = ((~g1367));
assign g10233 = ((~II13699));
assign g28400 = (g27211)|(g15870);
assign g19409 = ((~g16431));
assign g9185 = ((~II13007));
assign g22191 = (g8119&g19875);
assign g11981 = ((~II14823));
assign g12125 = ((~g9728))|((~g5101));
assign g24068 = ((~g19919));
assign g20711 = ((~g15509));
assign g29346 = (g4894&g28381);
assign g33860 = (g33270&g20501);
assign g33091 = (g32392&g18897);
assign g16872 = ((~II18060));
assign II27784 = ((~g29013));
assign g26571 = (g10472&g24386);
assign g28187 = ((~II26710));
assign g16803 = (g5933&g14810);
assign g9915 = ((~g2583));
assign g24770 = ((~g22763));
assign g24061 = ((~g19919));
assign g19869 = ((~g16540));
assign g14730 = ((~g5615))|((~g12093))|((~g5623))|((~g12301));
assign g17149 = (g232&g13255);
assign g7840 = ((~g4878));
assign g25125 = (g20187&g23520);
assign g33328 = (g32209&g20584);
assign g18650 = (g6928&g17271);
assign g29501 = (g28583)|(g27634);
assign g34900 = (g34860)|(g21686);
assign g30284 = (g28852&g23994);
assign g10377 = ((~g6940));
assign g32850 = ((~g30937));
assign g34190 = (g33802)|(g33810);
assign g22876 = (g20136&g9104);
assign g22907 = ((~g20453));
assign g23708 = (g19050&g9104);
assign g26816 = ((~g25260));
assign g11509 = ((~g7632));
assign g7296 = ((~g5313));
assign g34543 = ((~g34359));
assign g32915 = ((~g31710));
assign II30644 = ((~g32024));
assign g17738 = ((~g14813));
assign g30367 = (g30133)|(g18418);
assign II27409 = (g25556&g26424&g22698);
assign g17466 = ((~g12983));
assign II18214 = ((~g12918));
assign g8381 = ((~g2610));
assign g16611 = (g5583&g14727);
assign g30477 = (g30239)|(g21948);
assign g12931 = (g392&g11048);
assign g28919 = (g27663&g21295);
assign g17226 = ((~II18252));
assign g34542 = (g34332&g20089);
assign g15864 = ((~g14833))|((~g12543))|((~g12487));
assign g24331 = (g6977&g22228);
assign g28362 = (g27154)|(g15840);
assign g18371 = (g1870&g15171);
assign g34507 = (g34280&g19454);
assign g11160 = (g6336&g7074&g6322&g10003);
assign II17808 = ((~g13311));
assign g20248 = ((~g17056))|((~g14146))|((~g14123));
assign g9843 = ((~g4311));
assign II27718 = ((~g28231));
assign g11994 = ((~g8310))|((~g8365));
assign II17569 = ((~g14564));
assign g33108 = ((~g32183)&(~g31228));
assign g23782 = ((~g2741))|((~g21062));
assign g32411 = (g31119&g13469);
assign g12836 = ((~g10351));
assign g33676 = (g33125&g7970);
assign g24207 = (g23396)|(g18119);
assign g29480 = (g28115)|(g22172);
assign g25556 = ((~g22763));
assign g6974 = ((~II11746));
assign II19384 = ((~g15085));
assign g32547 = ((~g30614));
assign g27482 = (g26488&g17641);
assign g28111 = (g27343&g22716);
assign g28580 = (g27328)|(g26275);
assign g25752 = (g25079)|(g22099);
assign II18276 = ((~g1075));
assign g8055 = ((~g1236));
assign g28309 = (g27106)|(g15796);
assign II30761 = (g32071)|(g32167)|(g32067)|(g32082);
assign II16471 = ((~g12367));
assign g8280 = ((~g3443));
assign g24372 = ((~g22885));
assign g9863 = ((~g5503));
assign g11330 = ((~g9483))|((~g1193));
assign g25096 = (g23778&g20560);
assign g23550 = ((~g20248));
assign g14133 = ((~g11692))|((~g11747));
assign g25288 = ((~g22228));
assign g20921 = ((~g15426));
assign g14148 = (g884&g10632);
assign g33411 = (g32361&g21410);
assign g31126 = ((~g7928)&(~g29540));
assign g10295 = ((~II13723));
assign g32664 = ((~g31528));
assign g17469 = (g4076&g13217);
assign g27386 = (g26488&g17498);
assign g27566 = (g26119)|(g24713);
assign g31270 = (g29692&g23282);
assign g8756 = ((~g4049));
assign g13025 = (g8431&g11026);
assign g23857 = (g19626&g7908);
assign g34934 = ((~g34918));
assign g18614 = (g3343&g17200);
assign g21067 = (g10085&g17625);
assign II26459 = ((~g26576))|((~g14306));
assign g21723 = ((~II21288));
assign g10028 = ((~g8));
assign g10708 = ((~g7836));
assign g24052 = ((~g21193));
assign g29574 = (g2016&g28931);
assign g8316 = ((~g2351));
assign g22319 = ((~II21831));
assign g34021 = (g33652)|(g18519);
assign II32846 = ((~g34502));
assign g30420 = (g29769)|(g21804);
assign g27997 = (g26813&g23995);
assign g12622 = ((~g9569)&(~g9518));
assign g21558 = (g15904&g13729);
assign g24582 = (g5808&g23402);
assign g30104 = (g28478)|(g11427);
assign g14231 = ((~g12246));
assign g21822 = (g3727&g20453);
assign g33272 = (g32121)|(g29551);
assign g28704 = (g27459)|(g16671);
assign g33932 = ((~II31810));
assign g9705 = ((~g2619))|((~g2587));
assign g21467 = ((~g15758));
assign g28044 = (g27256)|(g18130);
assign g33586 = (g33416)|(g18459);
assign g32027 = ((~II29585));
assign II21002 = ((~g16709));
assign g26737 = (g24460)|(g10720);
assign g23551 = (g10793&g18948);
assign g11233 = ((~g9664));
assign g15059 = ((~g12839)&(~g13350));
assign g34534 = (g34321&g19743);
assign g13995 = ((~g11261));
assign g9285 = ((~g2715));
assign g17671 = (g7685&g13485);
assign g17495 = ((~g3566))|((~g13730))|((~g3668))|((~g8542));
assign II24600 = (g6077&g6082&g9946);
assign g26856 = ((~II25586));
assign g32162 = (g31002&g23014);
assign g17721 = ((~g12915));
assign g21897 = (g20095)|(g15111);
assign g33132 = ((~g4843)&(~g32072));
assign g23277 = ((~II22380));
assign g26128 = (g2319&g25120);
assign g32670 = ((~g30673));
assign g19209 = ((~g12971)&(~g15614)&(~g11320));
assign II30055 = (g31070)|(g31170)|(g30614)|(g30673);
assign g12430 = ((~II15250));
assign g29675 = ((~g28380)&(~g8236)&(~g8354));
assign g21871 = (g4108&g19801);
assign g24523 = (g22318&g19468);
assign g17718 = ((~g14776));
assign g14183 = ((~g12381));
assign g33875 = ((~II31727));
assign II26670 = ((~g27709));
assign g8205 = ((~g2208));
assign g18399 = (g2024&g15373);
assign g26157 = (g2093&g25136);
assign g23872 = (g19389&g4157);
assign g29300 = (g28666)|(g18796);
assign g24341 = (g23564)|(g18771);
assign g31372 = ((~g8796)&(~g29697));
assign g34535 = (g34309)|(g34073);
assign g26645 = ((~g23602)&(~g25160));
assign g25588 = (g21686)|(g24158);
assign g24754 = (g19604&g23027);
assign II32547 = ((~g34397));
assign g9972 = ((~II13510))|((~II13511));
assign g7879 = ((~II12262))|((~II12263));
assign g32021 = ((~II29579));
assign g26719 = (g10709&g24438);
assign g30308 = (g29178&g7004&g5297);
assign II21288 = ((~g18216));
assign g29025 = ((~g27937))|((~g2629))|((~g7462));
assign g29686 = (g2246&g29057);
assign g29097 = ((~g9700))|((~g27858));
assign g14543 = ((~II16660));
assign g11010 = (g4698&g8933);
assign g24880 = ((~g23281))|((~g23266))|((~g22839));
assign g32911 = ((~g31376));
assign II29351 = (g29328)|(g29323)|(g29316)|(g30316);
assign g20447 = ((~g15426));
assign g10030 = ((~g116));
assign II33255 = ((~g34975));
assign g23359 = ((~II22458));
assign II26667 = ((~g27585));
assign II32871 = ((~g34521));
assign g20570 = ((~g15277));
assign g20241 = (g16233)|(g13541);
assign g20548 = ((~g15426));
assign g14387 = (g9086)|(g11048);
assign g14431 = ((~g12208));
assign g30504 = (g30253)|(g22025);
assign g30072 = ((~II28301));
assign g34248 = ((~II32243));
assign g34104 = (g33916&g23639);
assign g9684 = ((~g6191));
assign g19902 = ((~g17200));
assign g32055 = (g10999&g30825);
assign II27391 = ((~g27929));
assign g24432 = (g23900)|(g21361);
assign g6810 = ((~g723));
assign g34131 = ((~II32074));
assign g32227 = (g31146)|(g29648);
assign g34115 = (g20516&g9104&g33750);
assign g21123 = ((~g15615));
assign g33987 = (g33847)|(g18396);
assign g31579 = (g19128&g29814);
assign g11865 = ((~g10124));
assign g31819 = ((~g29385));
assign g32072 = ((~g31009))|((~g13301));
assign II15043 = ((~g1834))|((~II15041));
assign g26657 = (g24908)|(g24900)|(g24887)|(g24861);
assign g13977 = ((~g11610))|((~g11729));
assign g31253 = (g25980)|(g29533);
assign g14898 = ((~g5901))|((~g12129))|((~g6000))|((~g12614));
assign g18369 = (g12848&g15171);
assign g6993 = ((~g4859));
assign II28162 = ((~g28803));
assign g33829 = (g33240&g20164);
assign g14223 = ((~g9092))|((~g11858));
assign g21878 = (g4129&g19801);
assign II26072 = ((~g13517))|((~II26070));
assign II28174 = ((~g28803));
assign g23985 = ((~g19210));
assign g25726 = (g25148)|(g22009);
assign g24405 = ((~g22722));
assign II12712 = ((~g59));
assign g16507 = ((~g13797))|((~g13764));
assign g24656 = (g11736&g22926);
assign II14836 = ((~g9688));
assign g14641 = (g11994&g12020);
assign II20204 = ((~g16246))|((~II20203));
assign II22327 = ((~g19367));
assign g23986 = ((~g18833));
assign g24904 = (g11761&g23279);
assign g27548 = (g26576&g17763);
assign g23953 = ((~g19277));
assign II31156 = (g31070&g31823&g32680&g32681);
assign g21455 = ((~g15426));
assign g11410 = ((~g6875))|((~g6895))|((~g8696));
assign g25233 = ((~g20838))|((~g23623));
assign g15883 = (g9180&g14258);
assign g33483 = (g32621&II31111&II31112);
assign II32056 = ((~g33641));
assign g29142 = ((~g5535)&(~g28010));
assign g22080 = (g6275&g19210);
assign g33139 = ((~g8650)&(~g32057));
assign g25013 = ((~g23599));
assign II18452 = (g14514)|(g14448)|(g14418);
assign g34977 = (g34873)|(g34966);
assign g11737 = (g8359)|(g8292);
assign g32995 = (g32330)|(g18375);
assign g28163 = ((~II26682));
assign II22918 = ((~g21451));
assign g23995 = ((~g19277));
assign II13995 = ((~g8744));
assign g15877 = ((~g14833))|((~g9340))|((~g12543));
assign g10678 = ((~II13990));
assign g12370 = ((~II15213))|((~II15214));
assign g20059 = ((~g17302));
assign II12997 = ((~g351));
assign g29361 = ((~g7553)&(~g28174));
assign g18796 = (g6167&g15348);
assign g33831 = (g23088&g33149&g9104);
assign g26635 = (g25321&g20617);
assign g29755 = ((~II28002));
assign g29609 = (g28482&g11861);
assign g28174 = ((~g1270))|((~g27059));
assign g27614 = (g26785&g26759);
assign g25400 = ((~g22472))|((~g12086));
assign g16264 = ((~g518))|((~g9158))|((~g13223));
assign g11374 = ((~g9536))|((~g1536));
assign g29317 = ((~II27677));
assign g11115 = (g6133&g9954);
assign g32337 = (g31465&g20663);
assign g7304 = ((~g1183)&(~g1171));
assign g18209 = (g921&g15938);
assign g26613 = (g1361&g24518);
assign g30285 = ((~g7097)&(~g29110));
assign g10053 = ((~g6381));
assign g34675 = ((~II32809));
assign g33439 = ((~g31950)&(~g4633));
assign II28579 = ((~g29474));
assign II24117 = (g23088)|(g23154)|(g23172);
assign g27033 = (g25767&g19273);
assign g17290 = ((~g9506))|((~g9449))|((~g14431));
assign g24170 = ((~II23354));
assign g34720 = (g34694)|(g18134);
assign g14028 = (g8673&g11797);
assign g33093 = ((~g31997)&(~g4601));
assign g31524 = (g29897&g20593);
assign II14206 = ((~g3821))|((~II14204));
assign g28223 = (g27338&g17194);
assign II31297 = (g32884&g32885&g32886&g32887);
assign g10510 = ((~g7183)&(~g4593)&(~g4584));
assign g24443 = (g23917)|(g21378);
assign g21932 = (g5204&g18997);
assign g32843 = ((~g31021));
assign g13463 = ((~g10476));
assign g27962 = (g25954&g19597);
assign g23860 = ((~g19074));
assign g17572 = ((~g3598))|((~g13799))|((~g3676))|((~g8542));
assign II26676 = ((~g27736));
assign II12374 = ((~g3462))|((~II12372));
assign g13908 = ((~g4709)&(~g8796)&(~g11155));
assign g30293 = (g28236)|(g27246);
assign g20085 = ((~g16187));
assign g16483 = (g5224&g14915);
assign g34517 = (g34290&g19493);
assign II32988 = ((~g34755));
assign II22921 = ((~g14677))|((~g21284));
assign g14021 = ((~g11697))|((~g8958));
assign g8796 = ((~g4785));
assign g24629 = (g6163&g23699);
assign II31202 = (g32747&g32748&g32749&g32750);
assign g25732 = (g25201)|(g22017);
assign g25513 = ((~g23870));
assign g32603 = ((~g31070));
assign g23010 = ((~g20516))|((~g2984));
assign g33908 = (g33092&g18935);
assign g15094 = ((~g13177)&(~g12865));
assign g33549 = (g33328)|(g18337);
assign g17284 = ((~g9253)&(~g14317));
assign g17151 = (g8659&g12996);
assign g22999 = ((~g20453));
assign g34660 = ((~g34473));
assign g10721 = (g3288&g6875&g3274&g8481);
assign g18414 = (g2102&g15373);
assign g13499 = ((~g11479))|((~g11442))|((~g11410))|((~g11382));
assign g29281 = (g28541)|(g18743);
assign g28567 = (g6832&g27101);
assign g25538 = ((~g22594));
assign g23900 = (g1129&g19408);
assign g28340 = ((~g27439)&(~g26339));
assign g18202 = (g907&g15938);
assign g31279 = (g29571)|(g29579);
assign g27759 = (g22457&g25224&g26424&g26213);
assign g32942 = ((~g30825));
assign g32199 = (g30916&g25506);
assign g23699 = ((~g21012))|((~g11160));
assign g20767 = ((~g17873));
assign g6821 = ((~II11655));
assign g33474 = (g32556&II31066&II31067);
assign g8134 = ((~II12415));
assign g33880 = (g33290&g20568);
assign g24558 = (g22516&g19566);
assign g19787 = ((~g17096));
assign g22139 = ((~II21722));
assign g24016 = (g14528&g21610);
assign II31211 = (g31021&g31833&g32759&g32760);
assign g18186 = (g753&g17328);
assign II12269 = ((~g1141))|((~g956));
assign g32829 = ((~g30937));
assign g23456 = ((~g21514));
assign g33025 = (g32162)|(g21780);
assign g12592 = ((~II15364))|((~II15365));
assign g34245 = ((~II32234));
assign gbuf83 = (g3661);
assign g29303 = (g28703)|(g18801);
assign g26396 = (g24762)|(g23062);
assign II18694 = ((~g5666));
assign g34123 = ((~II32062));
assign g24004 = (g37&g21225);
assign g24188 = (g316&g22722);
assign II26523 = (g20720)|(g20857)|(g20998)|(g21143);
assign g9392 = ((~g5869));
assign g23411 = ((~g20734));
assign g10044 = ((~g5357));
assign g19370 = ((~g15915));
assign g25739 = (g25149)|(g22054);
assign II15333 = ((~g10152))|((~g2116));
assign g12851 = ((~g6846)&(~g10430));
assign g24604 = ((~g23112));
assign II22264 = ((~g20100));
assign II31807 = ((~g33149));
assign g30131 = (g28589&g21178);
assign g17845 = ((~II18835));
assign g25530 = (g23750&g21414);
assign g16702 = (g5615&g14691);
assign g24551 = (g17148&g23331);
assign g23233 = ((~g21037));
assign g14844 = (g10776)|(g8703);
assign g21332 = (g996&g15739);
assign g29881 = (g2040&g29150);
assign g29555 = (g29004&g22498);
assign g12008 = ((~g9932))|((~g5798));
assign g24280 = (g23292)|(g15109);
assign g8951 = ((~g554));
assign g33678 = (g33149&g10710&g22319);
assign g28416 = (g27218)|(g15880);
assign g25139 = ((~g22472));
assign II23399 = ((~g23450));
assign g21414 = ((~g17929));
assign g16187 = (g8822)|(g13486);
assign g14751 = ((~g10622)&(~g10617)&(~g10609)&(~g10603));
assign II32458 = ((~g34243));
assign II22683 = ((~g11893))|((~g21434));
assign g31506 = ((~g4793)&(~g29540));
assign g25073 = ((~II24237));
assign g30263 = (g28773&g23962);
assign g8654 = ((~g1087));
assign g13095 = (g11374)|(g1287);
assign g20710 = ((~g15509));
assign II14171 = ((~g3119))|((~II14169));
assign g10166 = ((~g6040));
assign II23345 = ((~g23320));
assign g10001 = ((~g6105));
assign g18720 = (g15137&g16795);
assign g23771 = (g21432)|(g21416)|(II22912);
assign g29974 = (g29173&g12914);
assign II14050 = ((~g9963));
assign g27775 = ((~g21228))|((~g25262))|((~g26424))|((~g26166));
assign II17460 = ((~g13378))|((~g1300));
assign g24960 = ((~g23716));
assign g27413 = (g26576&g17530);
assign g28681 = (g27428)|(g16634);
assign g30158 = (g28613&g21274);
assign g34076 = (g33694&g19519);
assign g29851 = (g1668&g29079);
assign g21769 = (g3247&g20785);
assign g18362 = (g1834&g17955);
assign g34725 = (g34700)|(g18183);
assign g12429 = ((~g7473))|((~g6675));
assign II11793 = ((~g6049));
assign g33008 = (g32261)|(g18457);
assign II13565 = ((~g2648))|((~II13564));
assign gbuf24 = (g5101);
assign g26295 = (g13070&g25266);
assign g11382 = ((~g8644))|((~g6895))|((~g8663));
assign g10617 = ((~g10151))|((~g9909));
assign g29663 = (g1950&g28693);
assign g33055 = (g31986)|(g21976);
assign g33101 = (g32398&g18976);
assign g23726 = ((~g9559))|((~g21140));
assign g25426 = ((~g12371))|((~g22369));
assign g24704 = (g17593&g22384);
assign g24254 = (g23265)|(g18306);
assign g18655 = (g15106&g14454);
assign g23655 = ((~II22793))|((~II22794));
assign g25776 = ((~g7166)&(~g24380)&(~g24369));
assign g25480 = ((~g22228));
assign g20388 = ((~g17297));
assign g15127 = ((~g12879)&(~g13605));
assign g26386 = (g24719)|(g23023);
assign II16544 = ((~g11931));
assign g23432 = ((~g21514));
assign g12347 = ((~g9321)&(~g9274));
assign g34296 = ((~II32297));
assign g7766 = ((~II12189));
assign II13152 = ((~g6746));
assign g10107 = ((~II13606));
assign g16306 = ((~g4944))|((~g13971))|((~g12088));
assign g12955 = ((~II15577));
assign g23531 = (g10760&g18930);
assign II32938 = ((~g34663));
assign g32384 = ((~g31666));
assign g11402 = ((~g7594));
assign g16707 = (g6641&g15033);
assign g18810 = (g6505&g15483);
assign g22177 = ((~g19074));
assign g32128 = (g31631&g29953);
assign g16929 = (g6505&g14348);
assign g28934 = ((~g27882))|((~g14641));
assign g11763 = ((~g3881)&(~g8172));
assign g17433 = ((~II18382));
assign g10112 = ((~g1988));
assign g24608 = (g6500&g23425);
assign g24743 = (g22708&g19789);
assign II12503 = ((~g215));
assign g14779 = ((~II16847));
assign g27878 = ((~g9559)&(~g25839));
assign g25580 = (g19268&g24149);
assign g27458 = (g24590)|(g25989);
assign II27401 = ((~g27051));
assign g15965 = (g13035)|(g10675);
assign g33286 = (g32145)|(g29585);
assign g30336 = (g29324)|(g18203);
assign II15773 = ((~g10430));
assign g9807 = ((~g5712));
assign II31057 = (g32538&g32539&g32540&g32541);
assign g19747 = ((~g17015));
assign g30050 = (g22545&g28126);
assign g16324 = (g13657&g182);
assign g15005 = ((~g12667))|((~g12622));
assign g10338 = ((~g5062)&(~g5022));
assign g15167 = ((~g13835)&(~g12908));
assign II18066 = ((~g3317));
assign g25408 = (g22682&g9772);
assign g29764 = (g28219)|(g28226);
assign g31796 = ((~g29385));
assign II26693 = ((~g27930));
assign g32776 = ((~g31672));
assign g8059 = ((~g3171));
assign II32794 = ((~g34580));
assign II15144 = ((~g5659));
assign II31216 = (g30937&g31834&g32766&g32767);
assign g24111 = ((~g19890));
assign g31497 = (g20041&g29930);
assign g34870 = (g34820&g19882);
assign g7439 = ((~g6351));
assign g33949 = (g32446)|(g33459);
assign II22712 = ((~g21434))|((~II22710));
assign g34484 = (g34407&g18939);
assign g18262 = (g1259&g16000);
assign g11360 = ((~g3763)&(~g8669));
assign g14379 = ((~g5723))|((~g11907));
assign g18539 = (g2763&g15277);
assign g8255 = ((~g2028));
assign g8365 = ((~g2060));
assign g30011 = (g29183&g12930);
assign g19444 = ((~g17192)&(~g14295));
assign g23211 = ((~g21308));
assign g27330 = (g2541&g26744);
assign g12525 = ((~g7522))|((~g6668));
assign g19593 = (g17145)|(g14210);
assign g31808 = ((~g29385));
assign g27596 = (g26207)|(g24775);
assign g33570 = (g33420)|(g18405);
assign g28292 = (g23781&g27762);
assign g32330 = (g31320&g20631);
assign g18894 = ((~g16000));
assign g26690 = (g10776)|(g24433);
assign g13492 = (g9856&g11865);
assign g34839 = ((~II33053));
assign g15700 = (g3089&g13483);
assign g29511 = (g1736&g28783);
assign g19352 = ((~g15758));
assign g8587 = ((~g3689));
assign g17182 = (g8579&g13016);
assign g14321 = ((~g10874));
assign g20103 = ((~g17433));
assign g33799 = ((~g33299));
assign g13901 = ((~g11480));
assign g25099 = ((~g22369));
assign g25947 = ((~g1199)&(~g24591));
assign g6960 = ((~g1));
assign g18957 = ((~II19734));
assign II15295 = ((~g8515));
assign g26701 = ((~g25341));
assign g33035 = (g32019)|(g21872);
assign g28732 = (g27505)|(g16734);
assign g13771 = (g11441&g11355&g11302&II16111);
assign g22590 = (g19274&g19452);
assign II14259 = ((~g3133))|((~II14257));
assign g10355 = ((~g6816));
assign g34582 = (g7764&g34313);
assign g10029 = ((~II13548));
assign g28206 = ((~g12546))|((~g26105))|((~g27985));
assign g7684 = (g4072)|(g4176);
assign g27337 = ((~g8334)&(~g26616));
assign g7475 = ((~g896));
assign g31481 = (g29768&g23417);
assign g34280 = (g26833)|(g34213);
assign II32439 = ((~g34227))|((~g34220));
assign g28357 = (g27148)|(g15836);
assign g14930 = ((~g12609))|((~g12515));
assign g28488 = (g27969&g17713);
assign g24137 = ((~g20998));
assign II13779 = ((~g6868));
assign g18929 = ((~g16100));
assign g14871 = ((~g6653))|((~g12211))|((~g6661))|((~g12471));
assign g31913 = (g31485)|(g21999);
assign g24201 = (g22848)|(g18104);
assign g26935 = ((~II25677));
assign g28707 = (g27461)|(g16673);
assign g34145 = ((~II32096));
assign g24665 = ((~g23067));
assign II24067 = (g3731&g3736&g8553);
assign g8273 = ((~g2453));
assign g34330 = (g34069)|(g33717);
assign g32983 = (g31990)|(g18222);
assign g28747 = (g27521)|(g13942);
assign g8912 = ((~g4180));
assign g22531 = (g20773)|(g20922);
assign g9056 = ((~g3017));
assign g24466 = ((~II23671));
assign g13103 = ((~g10905));
assign g30314 = (g28268)|(g27266);
assign g9829 = ((~g2250));
assign g15011 = ((~g12716))|((~g12632));
assign g29692 = (g28197)|(g10873);
assign II14016 = ((~g9104));
assign g18157 = (g15057&g17433);
assign g34561 = (g34368&g17410);
assign g18634 = (g3813&g17096);
assign II31007 = (g32466&g32467&g32468&g32469);
assign g19533 = ((~g16261));
assign gbuf96 = (g3976);
assign g11381 = ((~g9660))|((~g3274));
assign g22664 = (g19139)|(g15694);
assign g32068 = (g31515&g10862);
assign g19880 = ((~g16201)&(~g13634));
assign g33361 = (g32257&g20911);
assign g33545 = (g33399)|(g18324);
assign g24303 = (g4369&g22228);
assign g11935 = ((~g9485)&(~g7267));
assign g25001 = ((~g23666));
assign g25748 = (g25078)|(g18799);
assign g16813 = ((~g3614))|((~g13799))|((~g3625))|((~g8542));
assign g31967 = (g31755&g22167);
assign g13528 = ((~g11294))|((~g7549))|((~g1008));
assign g9529 = ((~g6561));
assign g22936 = ((~g20283));
assign g32707 = ((~g31579));
assign g25160 = ((~g5390)&(~g23659));
assign g16212 = (g6167&g14321);
assign g27122 = (g22537)|(g25917);
assign g16283 = (g11547&g11592&g6789&II17606);
assign II19927 = ((~g17408));
assign g33386 = (g32258)|(g29951);
assign II22622 = ((~g21209));
assign gbuf12 = (g4809);
assign II22046 = ((~g19330));
assign g22005 = (g5759&g21562);
assign g6825 = ((~g979));
assign g29523 = (g28930&g22417);
assign g24408 = (g23989&g18946);
assign g12059 = ((~g9853)&(~g7004));
assign g33955 = (g33505)|(II31858)|(II31859);
assign g28144 = (g4608&g27020);
assign g24103 = ((~g21209));
assign g7887 = ((~II12278))|((~II12279));
assign g26923 = (g25923)|(g18290);
assign II14212 = ((~g9252))|((~II14211));
assign g20077 = (g16025)|(g13320);
assign g21127 = ((~g18065)&(~g12099));
assign g13892 = ((~g11653))|((~g11473));
assign g18116 = (g168&g17015);
assign g19540 = (g1124&g15904);
assign g9391 = ((~II13110))|((~II13111));
assign II17938 = ((~g3676));
assign g26672 = ((~g25275));
assign II18861 = ((~g14307));
assign g29751 = (g28297&g23216);
assign g23334 = ((~g20785));
assign g34765 = (g34692&g20057);
assign g12832 = (g10347)|(g10348);
assign g30614 = (g20154&g29814);
assign g34576 = ((~II32654));
assign g8889 = ((~g3684))|((~g4871));
assign g10351 = ((~g6802));
assign g13017 = ((~II15633));
assign g34816 = ((~II33030));
assign g21954 = (g5381&g21514);
assign g9607 = ((~g5046));
assign g18326 = (g1664&g17873);
assign g33310 = (g29631)|(g32165);
assign II30192 = (g29385)|(g31376)|(g30735)|(g30825);
assign g19930 = ((~g17200));
assign g24591 = ((~g22833))|((~g22642));
assign g23923 = ((~g18997));
assign g11405 = ((~g2741))|((~g2735))|((~g6856))|((~g2748));
assign g8009 = ((~g3106));
assign g29879 = (g28289)|(g26096);
assign g8235 = ((~II12463));
assign g22519 = ((~g19801));
assign g20130 = ((~g17328));
assign g32104 = (g31616&g29906);
assign g33580 = (g33330)|(g18442);
assign g27161 = (g26166&g8241&g1783);
assign g14613 = (g10602&g10585);
assign g18273 = (g1287&g16031);
assign g28157 = ((~II26670));
assign g21886 = (g4153&g19801);
assign g16744 = ((~II17964));
assign g21735 = (g3057&g20330);
assign II25692 = ((~g25689));
assign g11490 = ((~g8666))|((~g3639))|((~g3694));
assign g12907 = ((~g10415));
assign g15115 = (g2946&g14454);
assign g23308 = ((~g21024));
assign g34588 = (g26082&g34323);
assign g22329 = (g11940&g20329);
assign g12311 = ((~g6109)&(~g10136));
assign g19383 = (g16893&g13223);
assign g13555 = ((~g12692));
assign g34763 = (g34689&g19915);
assign g22647 = ((~II21959));
assign II15307 = ((~g10116))|((~II15306));
assign g33917 = ((~II31779));
assign g16203 = (g5821&g14297);
assign g24687 = (g5827&g23666);
assign g18903 = ((~g15758));
assign g20007 = ((~g11512))|((~g17794));
assign g26820 = ((~II25534));
assign g24966 = ((~g22763));
assign g24675 = (g17568&g22342);
assign g27854 = ((~g21228))|((~g25283))|((~g26424))|((~g26195));
assign g20598 = ((~g17929));
assign g25592 = (g24672)|(g21706);
assign g29536 = (g28969&g22432);
assign g30115 = (g28489)|(g11449);
assign g18668 = (g4322&g17367);
assign g9590 = ((~g1882));
assign g18518 = (g2657&g15509);
assign II22557 = ((~g20695));
assign g14570 = ((~g3933))|((~g11255))|((~g4023))|((~g8595));
assign II18560 = ((~g5969));
assign g30373 = (g30111)|(g18461);
assign g8808 = ((~g595));
assign g24211 = (g23572)|(g18138);
assign g10800 = (g7517)|(g952);
assign II26638 = ((~g27965));
assign g10921 = (g1548&g8685);
assign g10553 = ((~g8971));
assign g25241 = ((~g23651));
assign g24115 = ((~g20998));
assign g25870 = (g24840&g16182);
assign g25085 = (g4912&g22908);
assign g33353 = (g32240&g20732);
assign g25981 = (g2051&g25007);
assign g18185 = (g790&g17328);
assign g11966 = ((~II14800));
assign g15708 = ((~g7340))|((~g13083));
assign g25742 = (g25093)|(g22057);
assign g20577 = ((~g15483));
assign g32487 = ((~g30825));
assign g33460 = ((~II30998));
assign g28713 = ((~g27907));
assign g24729 = (g22719&g23018);
assign g9965 = ((~g127));
assign g32142 = (g31616&g29965);
assign II30400 = (g31021)|(g30937)|(g31327)|(g30614);
assign g34367 = (g7404&g34042);
assign g20219 = ((~II20495));
assign g14959 = ((~g12695))|((~g12798));
assign g9958 = ((~g6148));
assign g18278 = (g1345&g16136);
assign g29185 = ((~II27481));
assign g26253 = (g2327&g25435);
assign g33658 = ((~g33080));
assign g12074 = ((~II14932));
assign g18470 = (g2403&g15224);
assign g23720 = (g20165)|(g16801);
assign g28613 = (g27350)|(g26310);
assign g24548 = ((~g22942));
assign g8475 = ((~II12608));
assign g33434 = (g32239&g29702);
assign II12075 = ((~g996))|((~II12074));
assign II31031 = (g30614&g31801&g32499&g32500);
assign g14027 = ((~g8734)&(~g11363));
assign g28856 = ((~g27738))|((~g8093));
assign g19786 = ((~g17062));
assign g29263 = (g28239)|(g18617);
assign II15577 = ((~g10430));
assign II16875 = ((~g6675));
assign g29608 = (g28568&g11385);
assign g13041 = ((~II15667));
assign g34475 = (g27450&g34327);
assign g25542 = ((~g22763));
assign g33621 = (g33365)|(g18775);
assign g29368 = ((~II27730));
assign g17741 = ((~g12972));
assign II12287 = ((~g1484))|((~g1300));
assign g19890 = ((~g16987)&(~g8058));
assign g23381 = (g7239&g21413);
assign g13299 = (g437&g11048);
assign g26954 = (g26380)|(g24292);
assign g28271 = ((~g10533))|((~g27004))|((~g26990));
assign g34516 = (g34289&g19492);
assign g13300 = (g10656)|(g10676);
assign g18126 = (g15054&g16971);
assign g21924 = (g5057&g21468);
assign II22485 = ((~g21308));
assign g17501 = ((~II18434));
assign g27412 = (g26576&g17529);
assign g23388 = ((~g21070));
assign g15836 = (g3187&g14104);
assign II13182 = ((~g6500))|((~g6505));
assign g8721 = (g385&g376&g365);
assign g28214 = (g27731&g26625);
assign II14301 = ((~g8571));
assign g29595 = (g28475&g11833);
assign g20561 = ((~g17873));
assign II17446 = ((~g13336))|((~g956));
assign II17671 = ((~g13280));
assign g18135 = (g136&g17249);
assign g16811 = (g8690)|(g13914);
assign g26287 = (g2138&g25225);
assign g13822 = ((~g8160))|((~g11306));
assign II25612 = (g25567)|(g25568)|(g25569)|(g25570);
assign g8579 = ((~g2771));
assign g13010 = ((~II15620));
assign g28442 = (g27278&g20072);
assign g20028 = ((~g15371));
assign g23841 = ((~g19074));
assign II31162 = (g32689&g32690&g32691&g32692);
assign g21921 = (g5109&g21468);
assign g20268 = ((~g18008));
assign g23682 = (g16970&g20874);
assign g29859 = (g28388&g23307);
assign g32645 = ((~g30825));
assign g23427 = ((~II22542));
assign g12052 = ((~g7387))|((~g2465));
assign g17239 = ((~g11119)&(~g13518));
assign g24468 = (g10925)|(g22400);
assign g12152 = ((~g2485))|((~g8324));
assign g9554 = ((~g5105));
assign g32509 = ((~g31070));
assign II15208 = ((~g637));
assign g8442 = ((~g3476));
assign II12572 = ((~g51));
assign g13675 = ((~g10556));
assign g34342 = (g34103&g19998);
assign g31488 = (g1779&g30302);
assign g29914 = (g22531)|(g22585)|(II28147);
assign g11373 = ((~g7566));
assign g11866 = ((~g9883));
assign g28892 = ((~g27779))|((~g1772))|((~g7275));
assign g30021 = ((~g28994));
assign g17614 = ((~II18571));
assign II15918 = ((~g12381));
assign g29274 = (g28360)|(g18642);
assign II20830 = ((~g17657));
assign g18490 = (g2504&g15426);
assign g25528 = ((~g22594));
assign II24078 = ((~g22360));
assign g13312 = ((~g11048));
assign g29154 = ((~g27937))|((~g9835));
assign g34774 = (g34695&g20180);
assign g25047 = ((~g23733));
assign g32457 = ((~g30735));
assign g34873 = (g34830&g20046);
assign g33980 = (g33843)|(g18370);
assign g9564 = ((~g6120));
assign g18146 = (g595&g17533);
assign II31096 = (g31376&g31812&g32594&g32595);
assign g33469 = (g32519&II31041&II31042);
assign g30081 = (g28454)|(g11366);
assign g26778 = (g25501&g20923);
assign g27933 = ((~g21228))|((~g25356))|((~g26424))|((~g26236));
assign g33247 = (g32130&g19980);
assign g34667 = (g34471&g33424);
assign g25955 = (g24720&g19580);
assign g27264 = (g25941&g19714);
assign g16233 = (g6137&g14251);
assign g26179 = (g2504&g25155);
assign II22912 = (g21555)|(g21364)|(g21357);
assign g8785 = ((~II12767));
assign II14550 = ((~g10072));
assign g32269 = (g31253&g20443);
assign II21992 = ((~g7670))|((~g19638));
assign g20058 = ((~g16782));
assign g12914 = ((~g12235));
assign g16964 = ((~II18120));
assign g28385 = (g27201)|(g15857);
assign g33335 = ((~II30861));
assign g12221 = ((~II15079))|((~II15080));
assign g33496 = (g32714&II31176&II31177);
assign g12997 = ((~g11826));
assign g32754 = ((~g30825));
assign g30002 = (g28481&g23487);
assign g19961 = ((~g17328));
assign g21697 = ((~II21258));
assign g18875 = ((~g15171));
assign g30240 = ((~g7004)&(~g28982));
assign II12819 = ((~g4277));
assign g23030 = ((~g20453));
assign g20049 = ((~II20318));
assign II12538 = ((~g58));
assign g28107 = (g27970&g18874);
assign II18855 = ((~g13745));
assign g32595 = ((~g30825));
assign g25217 = (g12418&g23698);
assign g27040 = (g7812&g6565&g6573&g26226);
assign g11255 = ((~g8623)&(~g6928));
assign g12381 = ((~II15223));
assign g34264 = (g34081)|(g18701);
assign II32186 = ((~g33665))|((~II32185));
assign g18739 = (g5008&g16826);
assign g32648 = ((~g30614));
assign g8713 = ((~g4826));
assign II31625 = ((~g33197));
assign g32303 = (g27550&g31376);
assign g22107 = (g6411&g18833);
assign g28542 = (g27405&g20275);
assign g34807 = (g34764)|(g18596);
assign g15815 = (g3594&g14075);
assign g24843 = (g3010&g23211&II24015);
assign g30353 = (g30095)|(g18355);
assign II16575 = ((~g3298));
assign g18216 = (g967&g15979);
assign g15812 = (g3227&g13915);
assign g6954 = ((~g4138));
assign g32955 = ((~g30735));
assign g8417 = (g1056)|(g1116)|(II12583);
assign g33381 = (g11842&g32318);
assign g17199 = (g2236&g13034);
assign g25348 = ((~g22763));
assign g18097 = ((~II18897));
assign g19997 = ((~g16231)&(~g13739));
assign g12864 = ((~g10373));
assign g27129 = (g26026&g16584);
assign g33368 = (g32275&g21057);
assign g22306 = ((~g4584))|((~g4616))|((~g13202))|((~g19071));
assign II17615 = ((~g13251));
assign II15814 = ((~g11129));
assign g28239 = (g27135&g19659);
assign g30277 = (g28817&g23987);
assign g13622 = ((~g278)&(~g11166));
assign g14664 = ((~g5220))|((~g12059))|((~g5339))|((~g12497));
assign g19062 = (g446&g16180);
assign g25877 = (g25502)|(g23919);
assign g27234 = (g26055&g16814);
assign g30572 = ((~g29945));
assign g23314 = (g9104&g19200);
assign g28602 = (g27509&g20515);
assign g16313 = ((~g8005)&(~g13600));
assign g9478 = ((~II13152));
assign g32686 = ((~g31579));
assign g34349 = (g26019)|(g34104);
assign g24925 = ((~g20092))|((~g23154));
assign II15036 = ((~g799));
assign g31154 = (g19128&g29814);
assign g18623 = (g3484&g17062);
assign g10821 = ((~g7503)&(~g1384));
assign II18872 = ((~g13745));
assign g30186 = (g28641&g23839);
assign II25359 = ((~g24715));
assign g20323 = ((~g17873));
assign g23190 = ((~II22286));
assign g17192 = (g1677&g13022);
assign g14663 = ((~g5236))|((~g12002))|((~g5290))|((~g12239));
assign g29191 = ((~g7738)&(~g28010));
assign g31985 = (g4722&g30614);
assign g9772 = ((~II13352));
assign g34573 = ((~II32645));
assign g34052 = ((~g33635));
assign g10288 = ((~II13718));
assign g17059 = ((~II18151));
assign g12477 = ((~II15295));
assign g27493 = (g246&g26837);
assign g31246 = (g25965)|(g29518);
assign g29236 = (g28313)|(g18287);
assign g26377 = (g24700)|(g23007);
assign g14416 = ((~g12148)&(~g9541));
assign g25109 = ((~g23666));
assign g14565 = (g11934&g11952);
assign g21289 = ((~g14616))|((~g17493));
assign g34976 = (g34872)|(g34965);
assign II31859 = (g33501)|(g33502)|(g33503)|(g33504);
assign II12120 = ((~g632));
assign g34988 = ((~II33264));
assign g12939 = (g405&g11048);
assign g25187 = (g12296&g23629);
assign g33263 = (g32393&g25481);
assign g15743 = ((~g5893))|((~g14497))|((~g6005))|((~g9935));
assign g24347 = (g23754)|(g18790);
assign g20194 = ((~g16897));
assign g18946 = ((~g16100));
assign g33084 = ((~g31978)&(~g7655));
assign II17379 = ((~g13336))|((~g1129));
assign g29788 = (g28335&g23250);
assign gbuf7 = (g4408);
assign g29870 = (g2421&g29130);
assign g34878 = ((~II33106));
assign g13523 = (g7046&g12246);
assign g26689 = (g15754&g24431);
assign g18953 = ((~g16077));
assign g15783 = (g3215&g14098);
assign g30517 = (g30244)|(g22038);
assign g8584 = ((~g3639));
assign g13156 = (g10816&g10812&g10805);
assign g13378 = ((~g11374)&(~g11017));
assign g16866 = (g13492)|(g11044);
assign g22661 = ((~g20136))|((~g94));
assign g20977 = (g10123&g17301);
assign g34716 = ((~II32878));
assign g9822 = ((~g125));
assign g32735 = ((~g31021));
assign g27601 = (g26766&g26737);
assign g11149 = ((~g1564))|((~g7948));
assign g11678 = ((~II14563));
assign g28134 = (g27958)|(g27962);
assign g18833 = ((~II19661));
assign g10928 = ((~g8181))|((~g8137))|((~g417));
assign g8957 = (g2338)|(g2357);
assign g11929 = ((~II14745));
assign g20557 = ((~II20647));
assign g27650 = (g26519&g15479);
assign g30176 = (g23392)|(g28531);
assign g34183 = (g33695&g24385);
assign g14761 = ((~g12651))|((~g10281));
assign g16695 = ((~g14454));
assign g21988 = (g5583&g19074);
assign g22210 = ((~II21792));
assign g29491 = ((~II27777));
assign g13079 = ((~g1312))|((~g11336));
assign g6946 = ((~II11721));
assign g13322 = ((~g10918));
assign g26887 = (g26542)|(g24193);
assign g7891 = ((~g2994));
assign g34567 = (g34377&g17491);
assign g23503 = ((~g21468));
assign g30129 = ((~g28739)&(~g14537));
assign II18653 = ((~g5681));
assign g12014 = ((~g7197))|((~g703));
assign g25488 = (g6404&g23865&II24603);
assign g10033 = ((~g655));
assign g34613 = (g34515)|(g18567);
assign g7806 = ((~g4681));
assign g9253 = ((~g5037));
assign g20869 = ((~g15615));
assign g33728 = (g22626&g10851&g33187);
assign g27045 = (g10295&g3171&g3179&g26244);
assign g24819 = ((~II23998));
assign g23084 = ((~g19954));
assign g29007 = ((~g9269)&(~g28010));
assign g14170 = ((~g11715))|((~g11537));
assign gbuf41 = (g5976);
assign g20717 = ((~g5037)&(~g17217));
assign g8990 = ((~g146));
assign g25369 = ((~g22228));
assign II17125 = ((~g13809));
assign II24060 = ((~g22202));
assign g20146 = ((~g17533));
assign g24957 = ((~g21359))|((~g23462));
assign g8021 = ((~g3512));
assign g11037 = (g6128&g9184);
assign g23792 = ((~g19074));
assign II14797 = ((~g9636));
assign g13567 = (g10102&g11948);
assign g25886 = ((~g24537));
assign g20605 = ((~g17955));
assign g14065 = ((~g11048));
assign g27325 = (g12478&g26724);
assign g27541 = (g26278&g23334);
assign g32231 = (g30590)|(g29346);
assign g32834 = ((~g31672));
assign g8215 = ((~II12451));
assign g14422 = ((~g3187))|((~g11194))|((~g3298))|((~g8481));
assign g18763 = (g5481&g17929);
assign g14644 = (g10610&g10605);
assign g32480 = ((~g31070));
assign II14509 = ((~g370))|((~II14508));
assign g21282 = ((~II21019));
assign g9506 = ((~g5774));
assign g16300 = ((~II17626));
assign g34093 = (g20114&g33755&g9104);
assign g14848 = ((~g12651))|((~g12453));
assign g11217 = ((~g8531)&(~g6875));
assign g34639 = (g34486)|(g18722);
assign g17088 = ((~II18160));
assign g33047 = (g31944)|(g21927);
assign g18598 = (g3003&g16349);
assign g14586 = (g11953&g11970);
assign II16515 = ((~g12477));
assign g17771 = (g13288&g13190);
assign g15793 = (g3219&g13873);
assign g34555 = (g34349&g20512);
assign g27098 = (g25868&g22528);
assign g17399 = ((~g9626))|((~g9574))|((~g14535));
assign g16604 = ((~g3251))|((~g11194))|((~g3267))|((~g13877));
assign II16345 = ((~g881));
assign g19852 = ((~g17015));
assign g32195 = (g30734&g25451);
assign g21713 = (g298&g20283);
assign g30225 = (g28705&g23897);
assign g23189 = ((~g20060));
assign g19594 = (g11913&g17268);
assign gbuf19 = (g5283);
assign g34796 = (g34745)|(g18573);
assign g7195 = ((~g25));
assign g34322 = (g14188&g34174);
assign g23957 = (g4138&g19589);
assign g28690 = (g27436)|(g16641);
assign g32922 = ((~g31710));
assign g7041 = ((~g5644));
assign g7526 = ((~II12013));
assign g25008 = ((~g22432));
assign g22208 = (g19906&g20739);
assign g18562 = ((~II19384));
assign g14363 = ((~II16521));
assign g9381 = ((~g5527));
assign g7932 = (g4072)|(g4153);
assign g28814 = (g27545)|(g16841);
assign g17154 = ((~g14348));
assign g21403 = ((~g11652))|((~g17157));
assign g27648 = (g25882&g8974);
assign g16618 = (g6609&g15039);
assign g27551 = (g26091)|(g24675);
assign g31541 = (g22536&g29348);
assign g21788 = (g3401&g20391);
assign II15677 = ((~g5654));
assign g22215 = ((~g19277));
assign II32613 = ((~g34329));
assign g33069 = (g32009)|(g22113);
assign gbuf54 = (g6365);
assign g11269 = ((~g7516));
assign g10802 = (g7533)|(g1296);
assign g34179 = (g33686&g24372);
assign g26625 = ((~g23560)&(~g25144));
assign g29128 = ((~g27800));
assign II14935 = ((~g9902));
assign g14913 = (g1442&g10939);
assign g14497 = ((~g5990)&(~g12705));
assign g29894 = (g2070&g29169);
assign g33686 = ((~g33187));
assign II22958 = (g21603)|(g21386)|(g21365);
assign g18297 = (g1478&g16449);
assign g34045 = (g33766&g22942);
assign g19968 = ((~g17062)&(~g11223));
assign g28609 = (g27346)|(g16483);
assign g16239 = (g7892)|(g13432);
assign g9754 = ((~g2020));
assign g25972 = (g2217&g24993);
assign g20635 = ((~g18008));
assign g33370 = (g32279&g21139);
assign g29953 = ((~g28907));
assign g24416 = (g4939&g22870);
assign g30108 = (g28561&g20910);
assign g32681 = ((~g30735));
assign g11510 = ((~g7633));
assign g21808 = (g3570&g20924);
assign II22967 = ((~g21228))|((~II22965));
assign g8389 = ((~g3125));
assign g19950 = ((~g15885));
assign g23482 = ((~g18833));
assign g19147 = ((~II19786));
assign g9887 = ((~g5802));
assign g10589 = (g7223)|(g7201);
assign g34940 = ((~g34924));
assign g30040 = ((~g29025));
assign g28323 = (g27118)|(g15810);
assign II18385 = (g14413)|(g14391)|(g14360);
assign g15822 = (g3925&g13960);
assign g31140 = (g2102&g30037);
assign g28726 = ((~g27937));
assign g33719 = (g33141&g19433);
assign g20283 = ((~II20529));
assign g18302 = (g1514&g16489);
assign g21272 = ((~g11268))|((~g17157));
assign II12893 = ((~g4226));
assign g17287 = ((~g7262))|((~g14228));
assign g33628 = (g33071)|(g32450);
assign g23573 = ((~g20248));
assign g13583 = ((~II16028));
assign g21855 = (g3925&g21070);
assign g27384 = (g26400&g17496);
assign g17816 = ((~g6657))|((~g14602))|((~g6668))|((~g10061));
assign g14290 = ((~II16460));
assign g29985 = (g28127&g20532);
assign g31218 = (g30271&g23909);
assign g14432 = ((~g12311));
assign g18881 = ((~II19671));
assign g28733 = (g27507)|(g16735);
assign g11384 = ((~g8538)&(~g8540));
assign g29254 = (g28725)|(g18512);
assign g10500 = ((~II13875));
assign g29569 = (g29028&g22498);
assign g15134 = ((~g13638)&(~g12884));
assign g7046 = ((~g5791));
assign g19357 = ((~II19837));
assign g34054 = (g33778&g22942);
assign g31223 = (g20028&g29689);
assign g20765 = ((~g17748));
assign g34207 = (g33835)|(g33304);
assign II33131 = ((~g34906));
assign II22788 = ((~g18940));
assign g10002 = ((~g6195));
assign II18571 = ((~g13074));
assign g20374 = ((~g18065));
assign g23017 = ((~g20453));
assign g27036 = (g26329&g11038);
assign g27240 = (g25883)|(g24467);
assign g9537 = ((~g1748));
assign g7473 = ((~g6697));
assign g31269 = (g26024)|(g29569);
assign g19719 = ((~g16897));
assign g29869 = (g2331&g29129);
assign g10156 = ((~g2675));
assign g20624 = ((~g18065));
assign g18546 = (g2795&g15277);
assign g34120 = (g33930&g25158);
assign g33943 = (g33384&g21609);
assign g9746 = ((~II13326));
assign II25242 = ((~g490))|((~g24744));
assign g26090 = (g1624&g25081);
assign g17709 = ((~g14761));
assign g8177 = ((~g4966)&(~g4991)&(~g4983));
assign g8748 = ((~g776));
assign g32860 = ((~g30673));
assign g22159 = ((~II21744));
assign g32456 = ((~g31376));
assign g32706 = ((~g30673));
assign g10354 = ((~g6811));
assign g18604 = (g3125&g16987);
assign g21654 = ((~g17619));
assign II28591 = ((~g29371));
assign g28458 = (g27187&g12730&g20887&II26948);
assign g23266 = ((~g18918))|((~g2894));
assign g22530 = (g16751)|(g20171);
assign g21514 = ((~II21189));
assign g13543 = (g10543)|(g10565);
assign g27572 = (g26129)|(g24724);
assign g9653 = ((~g2441));
assign g13596 = ((~g10971));
assign g15829 = ((~g4112))|((~g13831));
assign g9014 = ((~g3004));
assign g16712 = ((~g13223));
assign g25498 = ((~g22498))|((~g2610))|((~g8418));
assign g19565 = ((~g16000));
assign g34188 = ((~g33875));
assign g21833 = (g15096&g20453);
assign g8833 = ((~g794));
assign g11932 = ((~g843)&(~g9166));
assign g20089 = ((~g17533));
assign g22017 = (g5763&g21562);
assign II31869 = (g33519)|(g33520)|(g33521)|(g33522);
assign g31601 = ((~II29207));
assign g33584 = (g33406)|(g18449);
assign g15125 = (g10363)|(g13605);
assign g24498 = (g14036&g23850);
assign g17179 = (g1041&g13211);
assign g10111 = ((~g1858));
assign g24095 = ((~g21209));
assign g20330 = ((~II20542));
assign II14497 = ((~g9020))|((~g8737));
assign g31929 = (g31540)|(g22093);
assign g25327 = ((~g22161));
assign g18551 = (g2811&g15277);
assign g31873 = (g31270)|(g21728);
assign II17094 = ((~g14331));
assign g24175 = ((~II23369));
assign g21329 = ((~g16577));
assign g22863 = (g9547&g20388);
assign g21380 = ((~g17955));
assign g32159 = (g31658&g30040);
assign II32234 = ((~g34126));
assign g14609 = ((~II16724));
assign g24271 = (g23451)|(g18628);
assign g25849 = ((~g24491));
assign g8922 = ((~II12907));
assign II13483 = ((~g6035));
assign g28819 = ((~II27271));
assign g13000 = ((~g7228))|((~g10598));
assign g23944 = ((~g19147));
assign g28765 = ((~g27800))|((~g7374))|((~g7280));
assign g25192 = (g20276&g23648);
assign II14225 = (g8457&g255&g8406&g262);
assign g24380 = ((~II23601))|((~II23602));
assign g23350 = ((~g20785));
assign g21011 = ((~g14504))|((~g17399))|((~g9629));
assign g18314 = (g1585&g16931);
assign g10775 = ((~g7960))|((~g7943))|((~g8470));
assign g20179 = ((~g17249));
assign g20080 = ((~g17328));
assign g28097 = (g27682)|(g22005);
assign g15699 = (g1437&g13861);
assign g24040 = ((~g19919));
assign g34598 = (g34541)|(g18136);
assign g22054 = (g6120&g21611);
assign g23286 = ((~g6875))|((~g20887));
assign g34271 = ((~g34160));
assign g27594 = (g26721&g26694);
assign II29337 = ((~g30286));
assign g15803 = (g12924)|(g10528);
assign g25156 = ((~g22498));
assign g18253 = (g1211&g16897);
assign g24327 = (g4549&g22228);
assign g32089 = (g27261&g31021);
assign g32631 = ((~g30825));
assign g14679 = ((~g12437)&(~g9911));
assign g34843 = (g33924)|(g34782);
assign g25396 = ((~g22384))|((~g2208))|((~g8259));
assign II32921 = ((~g34650));
assign g14773 = ((~g12711))|((~g12581));
assign g24114 = ((~g20720));
assign g9852 = ((~g3684))|((~g4871));
assign g13007 = ((~g11852));
assign g29719 = ((~g28406))|((~g13739));
assign g13509 = (g9951&g11889);
assign g33701 = (g33162&g16305);
assign II18903 = ((~g16872));
assign g32786 = ((~g31021));
assign g31284 = (g29575)|(g28290);
assign g28306 = (g27104)|(g15794);
assign g8291 = ((~II12503));
assign g21396 = ((~g17955));
assign g34162 = ((~g785))|((~g33823))|((~g11679));
assign g14166 = ((~g11048));
assign g17471 = ((~g14454));
assign g12972 = ((~g7209))|((~g10578));
assign g34287 = (g11370&g34124);
assign g34231 = (g33898)|(g33902);
assign g32285 = (g31222)|(g29740);
assign g32808 = ((~g30937));
assign g23285 = ((~g20887));
assign g27988 = (g26781&g23941);
assign g24278 = (g23201)|(g18648);
assign g32424 = ((~g8721)&(~g31294));
assign g23617 = ((~II22761))|((~II22762));
assign g22525 = (g13006&g19411);
assign g24659 = (g5134&g23590);
assign g34452 = (g34401)|(g18665);
assign g29880 = (g1936&g29149);
assign g9064 = ((~g4983));
assign g29331 = (g29143&g22169);
assign g26793 = (g24478)|(g7520);
assign g14252 = ((~II16438));
assign g25677 = (g24684)|(g21834);
assign g29993 = ((~g29018));
assign g19581 = (g15843&g1500&g10918);
assign II21784 = ((~g19638));
assign g10612 = ((~g10233));
assign II33246 = ((~g34970));
assign g20538 = ((~g15348));
assign g16595 = (g5921&g14697);
assign II16713 = ((~g5331));
assign g34235 = (g32585)|(g33953);
assign g15590 = (g3139&g13530);
assign g27027 = ((~g26398)&(~g26484));
assign g15673 = (g182&g13437);
assign g32964 = ((~g31672));
assign g34915 = ((~II33137));
assign II15663 = ((~g5308));
assign g24032 = ((~g21256));
assign g10856 = (g4269&g8967);
assign g19794 = ((~g16489));
assign g25093 = (g12831&g23493);
assign g29758 = (g28306&g23222);
assign g29891 = (g28420&g23356);
assign g13110 = ((~g7841)&(~g10741));
assign II18265 = ((~g13350));
assign g30192 = (g28649&g23847);
assign g27020 = (g4601&g25852);
assign g15024 = ((~g12780))|((~g10421));
assign g26605 = ((~g25293));
assign g27969 = ((~g7170)&(~g25821));
assign II13276 = ((~g5798));
assign g16588 = ((~g13929));
assign g32124 = (g24488)|(g30920);
assign g20442 = ((~g15171));
assign g29657 = ((~g28363))|((~g13634));
assign g22490 = (g21513)|(g12795);
assign g22881 = ((~II22096));
assign II21100 = ((~g16284));
assign g21785 = (g3431&g20391);
assign g26261 = (g24688&g10678&g8778&g8757);
assign g12859 = ((~g10366));
assign g14792 = ((~g10653)&(~g10623)&(~g10618)&(~g10611));
assign g8818 = ((~II12808));
assign II12106 = ((~g626));
assign g13856 = ((~II16160));
assign g34529 = (g34306&g19634);
assign g14905 = ((~g12785))|((~g7142));
assign g8358 = ((~II12541));
assign II26952 = ((~g27972));
assign g32816 = ((~g31327));
assign g17530 = ((~g14947));
assign g26548 = ((~g25255));
assign g28250 = ((~g27074));
assign g11610 = ((~g7980)&(~g3155));
assign g32848 = ((~g30825));
assign g29775 = (g25966)|(g28232);
assign II11826 = ((~g4601))|((~II11824));
assign II13715 = ((~g71));
assign g7541 = ((~g344));
assign g9721 = ((~g5097));
assign g29373 = (g13832)|(g28453);
assign g18577 = (g2988&g16349);
assign g19468 = ((~g15938));
assign g25578 = (g19402&g24146);
assign g23630 = ((~g20739))|((~g11123));
assign g31908 = (g31519)|(g21955);
assign g28557 = (g27772&g15647);
assign g18619 = (g3466&g17062);
assign g26291 = (g2681&g25439);
assign II18063 = ((~g14357));
assign g17819 = ((~II18825));
assign g27249 = (g25929&g19678);
assign II20999 = ((~g16709));
assign g22135 = (g6657&g19277);
assign g27225 = (g2975)|(g26364);
assign g23291 = ((~g21070));
assign g19450 = ((~g11471))|((~g17794));
assign g26906 = (g26423)|(g24223);
assign g32847 = ((~g30735));
assign g34731 = (g34662)|(g18272);
assign II15263 = ((~g10081))|((~II15262));
assign g24809 = ((~g19965))|((~g23132));
assign g14333 = ((~g12042))|((~g12014))|((~g11990))|((~g11892));
assign II15878 = ((~g11249));
assign g25141 = ((~g22228)&(~g10334));
assign g18099 = ((~II18903));
assign g8858 = ((~g671));
assign g23087 = (g19487)|(g15852);
assign II22719 = ((~g21434))|((~II22717));
assign g13394 = ((~II15915));
assign g23230 = ((~II22327));
assign g32130 = (g30921)|(g30925);
assign g9819 = ((~g92));
assign g15859 = (g3610&g13923);
assign II25369 = ((~g24891));
assign g34068 = ((~g33728));
assign g29770 = (g28320&g23238);
assign g14278 = ((~g562)&(~g12259)&(~g9217));
assign II14424 = ((~g4005));
assign g20905 = (g7216)|(g17264);
assign g17592 = ((~II18530))|((~II18531));
assign g23653 = ((~II22788));
assign g7824 = ((~g4169));
assign g10541 = ((~g9407));
assign g14271 = ((~g10002)&(~g10874));
assign II24414 = ((~g23751))|((~g14382));
assign g31710 = (g29814&g19128);
assign gbuf39 = (g6012);
assign g13247 = (g8964&g11316);
assign g17579 = ((~g14959));
assign g12182 = ((~II15030));
assign g15739 = ((~g13284));
assign g7086 = ((~g4826));
assign II33134 = ((~g34906));
assign g26789 = (g10776)|(g24471);
assign g14024 = ((~g7121))|((~g11763));
assign g34519 = (g34293&g19504);
assign g33405 = (g32354&g21398);
assign II12117 = ((~g586));
assign g19528 = ((~g16349));
assign g33708 = ((~II31555));
assign g18468 = (g2393&g15224);
assign g33407 = (g32357&g21406);
assign g24143 = (g17694&g21659);
assign g29808 = (g28361&g23273);
assign g24389 = ((~g22908));
assign II22542 = ((~g19773));
assign g31260 = (g25993)|(g29555);
assign II15089 = ((~g2393))|((~II15087));
assign g32400 = (g4743&g30989);
assign g34166 = (g33785)|(g19752);
assign g15056 = ((~g6809)&(~g13350));
assign g23461 = ((~g18833));
assign g30413 = (g30001)|(g21772);
assign g30465 = (g30164)|(g21936);
assign g32763 = ((~g31710));
assign g31183 = (g30249&g25174);
assign g32403 = (g31117&g15842);
assign g28046 = (g27667)|(g18157);
assign g11592 = ((~II14537));
assign g30276 = ((~g7074)&(~g29073));
assign g9816 = ((~g6167));
assign II21480 = ((~g18696));
assign g23544 = ((~g21562));
assign II16698 = ((~g12077));
assign g27959 = (g25948&g19374);
assign II22286 = ((~g19446));
assign g23360 = ((~II22461));
assign g32857 = ((~g30937));
assign g24789 = ((~g23309));
assign g32978 = (g32197)|(g18145);
assign g26724 = ((~g25341));
assign g14841 = ((~g12593))|((~g12443));
assign g16023 = (g3813&g13584);
assign II13730 = ((~g4534))|((~II13729));
assign g18395 = (g12849&g15373);
assign g29147 = ((~II27449));
assign g33606 = (g33369)|(g18522);
assign g21143 = ((~g15348)&(~g9517));
assign g26516 = (g24968&g8876);
assign g25815 = (g8155&g24603);
assign II11903 = ((~g4414));
assign g32676 = ((~g30614));
assign II11908 = ((~g4449));
assign g29849 = (g26049)|(g28273);
assign g7260 = ((~II11908));
assign g10022 = ((~g6474))|((~g6466));
assign g25711 = (g25105)|(g21962);
assign g29547 = (g1748&g28857);
assign g33837 = (g33251&g20233);
assign g30418 = (g29751)|(g21802);
assign g24526 = ((~g22942));
assign g10736 = (g4040&g8751);
assign g15109 = (g4269&g14454);
assign g29381 = (g28135&g19399);
assign g19752 = (g2771&g15864);
assign g25785 = ((~g25488)&(~g25462));
assign g19553 = ((~g16782));
assign g26972 = (g26780)|(g25229);
assign g19364 = ((~g15825));
assign g23721 = (g21401)|(g21385)|(II22852);
assign g33725 = (g22626&g10851&g33176);
assign g30433 = (g29899)|(g21817);
assign g27682 = (g25777&g23565);
assign g27102 = ((~g26750)&(~g26779));
assign g32463 = ((~g31566));
assign g15165 = ((~g12907)&(~g13835));
assign g31841 = ((~g29385));
assign g32971 = ((~g31672));
assign g14635 = ((~II16741));
assign g13302 = ((~g12321));
assign g19772 = ((~g17183));
assign II29149 = ((~g29384));
assign g11997 = ((~g2319))|((~g8316));
assign g23508 = ((~g21562));
assign g24865 = (g11323&g23253);
assign g25203 = ((~g6428)&(~g23756));
assign g32165 = (g31669&g27742);
assign II30766 = ((~g32363));
assign g32616 = ((~g30735));
assign g21138 = ((~g15634));
assign gbuf113 = (g4210);
assign g7063 = ((~g4831));
assign g18794 = (g6154&g15348);
assign g15102 = ((~g14591)&(~g6954));
assign g31785 = (g30071)|(g30082);
assign g10898 = (g3706&g9100);
assign II28588 = ((~g29368));
assign g13994 = ((~g4049)&(~g11363));
assign g25026 = (g22929&g10503);
assign g24501 = (g14000&g23182);
assign g20510 = ((~g17226));
assign g21290 = ((~II21029));
assign g29170 = ((~g27907));
assign g19523 = ((~g16100));
assign g18100 = ((~II18906));
assign g33595 = (g33368)|(g18489);
assign II17884 = ((~g13336))|((~II17883));
assign g34215 = (g33778&g22670);
assign g28772 = (g27534)|(g16802);
assign g9180 = ((~g3719));
assign g18639 = (g3831&g17096);
assign II22792 = ((~g11956))|((~g21434));
assign II17609 = ((~g13510));
assign g24508 = ((~g23577)&(~g23618));
assign g13436 = (g9721&g11811);
assign g12114 = ((~g8241))|((~g8146));
assign g7496 = ((~g5969));
assign g28986 = ((~g5517)&(~g28010));
assign II23919 = ((~g9333))|((~II23917));
assign II12204 = ((~g1094))|((~II12203));
assign g24751 = ((~g3034)&(~g23105));
assign g23420 = ((~g21514));
assign g12936 = ((~g12601));
assign g16122 = (g9491&g14291);
assign g29586 = (g1886&g28927);
assign g18351 = (g1760&g17955);
assign g27721 = ((~g9672)&(~g25805));
assign g32826 = ((~g30825));
assign g15656 = ((~II17198));
assign g26160 = (g2453&g25138);
assign II32684 = ((~g34430));
assign g22060 = (g6151&g21611);
assign g24437 = ((~g22654));
assign g23447 = ((~g21562));
assign g28347 = (g27138)|(g15822);
assign g25560 = ((~g22550));
assign II17590 = ((~g14591));
assign g29217 = ((~II27567));
assign g8450 = ((~g3821));
assign g16128 = (g14333&g14166);
assign g14391 = ((~g12112)&(~g9585));
assign g23777 = ((~II22918));
assign II18125 = ((~g13191));
assign g22844 = ((~g21163));
assign g34680 = ((~II32820));
assign g19680 = (g12028&g17013);
assign II31221 = (g31327&g31835&g32773&g32774);
assign g30054 = ((~g29134));
assign g21962 = (g5428&g21514);
assign g20629 = ((~g17955));
assign g22072 = (g6259&g19210);
assign g30487 = (g30187)|(g21983);
assign g9099 = ((~g3706));
assign g7223 = ((~II11878))|((~II11879));
assign g24931 = (g23153&g20178);
assign g26864 = (g2907&g24548);
assign g23401 = (g7262&g21460);
assign g24560 = ((~g22942));
assign g21816 = (g3602&g20924);
assign g28777 = (g27539)|(g16807);
assign g22189 = ((~II21769));
assign g30165 = (g28619&g23788);
assign g18150 = (g604&g17533);
assign g16025 = (g446&g14063);
assign g33867 = (g33277&g20529);
assign g32409 = (g4754&g30996);
assign gbuf104 = (g4277);
assign g28217 = (g27733&g23391);
assign g8561 = ((~g3782))|((~g3774));
assign II23318 = ((~g21689));
assign g22311 = ((~g18935));
assign g29862 = ((~g28406));
assign g20230 = ((~II20499));
assign g23581 = (g20183&g11900);
assign g25236 = ((~II24415))|((~II24416));
assign g22711 = ((~g19581))|((~g7888));
assign II12151 = ((~g604));
assign g27451 = (g26400&g17599);
assign g32565 = ((~g30735));
assign g33904 = (g33321&g21059);
assign g11974 = ((~g2185))|((~g8259));
assign g27151 = (g26026&g16626);
assign II31874 = (g33528)|(g33529)|(g33530)|(g33531);
assign g10664 = ((~g8928));
assign g18781 = (g5831&g18065);
assign II23348 = ((~g23384));
assign g11280 = ((~g8647)&(~g3408));
assign g24917 = ((~g19913))|((~g23172));
assign g29197 = (g27187)|(g27163);
assign g32324 = (g31315&g23537);
assign g24334 = (g23991)|(g18676);
assign g11153 = ((~II14205))|((~II14206));
assign g12019 = ((~g7322))|((~g1906));
assign g32203 = (g4249&g31327);
assign g26810 = ((~g25220));
assign g21862 = (g3953&g21070);
assign g24391 = ((~g22190)&(~g14645));
assign g27203 = (g26026&g16688);
assign II17496 = ((~g1448))|((~II17494));
assign g26233 = (g2279&g25309);
assign g21555 = ((~g17846))|((~g14946))|((~g17686))|((~g17650));
assign g8851 = ((~g590));
assign g34415 = (g34207&g21458);
assign g17735 = ((~g14807));
assign g31813 = ((~g29385));
assign II19857 = ((~g16640));
assign g15904 = ((~II17380))|((~II17381));
assign g14186 = ((~g11346));
assign g9662 = ((~g3983));
assign II22564 = ((~g20857));
assign g20982 = ((~g17929)&(~g12065));
assign g25903 = ((~II25005));
assign II24438 = ((~g23771))|((~g14411));
assign g27727 = (g22432&g25211&g26424&g26195);
assign g32119 = (g31609&g29939);
assign g18452 = (g2311&g15224);
assign g34070 = ((~g33725));
assign II32758 = ((~g25779))|((~II32756));
assign g34087 = (g33766&g9104&g18957);
assign g28649 = (g27390)|(g16597);
assign II12761 = ((~g4188));
assign g15850 = (g3606&g14151);
assign g21949 = (g5264&g18997);
assign II16596 = ((~g12640));
assign g17780 = (g6772&g11592&g11640&II18782);
assign g29803 = (g28414&g26836);
assign g28114 = (g25869&g27051);
assign g32353 = (g29853)|(g31283);
assign g25617 = (g25466)|(g18189);
assign g29933 = ((~g8808)&(~g28500)&(~g12259));
assign g9614 = ((~g5128));
assign g27837 = (g17401)|(g26725);
assign g16885 = (g6605&g14950);
assign g25381 = ((~g538))|((~g23088));
assign g33810 = (g33427&g12768);
assign g30349 = (g30051)|(g18333);
assign g10671 = ((~g1526)&(~g8466));
assign g12084 = ((~g2342))|((~g8211));
assign g24364 = ((~g22722));
assign g30391 = (g30080)|(g18557);
assign g29688 = (g2509&g28713);
assign II24690 = (g24043&g24044&g24045&g24046);
assign g12189 = ((~g1917)&(~g8302));
assign II31984 = ((~g33653))|((~II31983));
assign II17355 = ((~g14591));
assign g19911 = (g14707&g17748);
assign II24700 = (g24057&g24058&g24059&g24060);
assign II31276 = (g31376&g31844&g32854&g32855);
assign II17744 = ((~g14912));
assign g28653 = (g7544&g27014);
assign II25743 = ((~g25903));
assign g6903 = ((~g3502));
assign g11735 = ((~g8534));
assign g30536 = (g30234)|(g22082);
assign g14831 = (g1152&g10909);
assign g21363 = ((~g17708))|((~g14664))|((~g17640))|((~g14598));
assign g27373 = (g26488&g17477);
assign g27343 = ((~g8005)&(~g26616));
assign g33270 = (g32119)|(g29547);
assign g9516 = ((~g6116));
assign g30562 = (g30289)|(g22133);
assign g29737 = ((~g28421))|((~g13779));
assign g9968 = (g1339&g1500);
assign g31778 = (g21369&g29385);
assign g21344 = ((~g11428))|((~g17157));
assign g11479 = ((~g6875))|((~g3288))|((~g3347));
assign g21466 = ((~g15509));
assign g32224 = (g4300&g31327);
assign g14587 = (g10584&g10567);
assign g23303 = ((~g20785));
assign g22359 = ((~g19495));
assign g16222 = (g6513&g14348);
assign g18647 = (g4040&g17271);
assign g26334 = (g1171)|(g24591);
assign g19854 = ((~II20222))|((~II20223));
assign g25685 = (g24476)|(g21866);
assign g30335 = (g29746)|(g18174);
assign g9020 = ((~g4287));
assign g7649 = ((~g1345));
assign g33488 = (g32658&II31136&II31137);
assign g33294 = (g32152)|(g29604);
assign g18376 = (g1913&g15171);
assign g7109 = ((~g5011));
assign g24890 = ((~g13852))|((~g22929));
assign g24939 = (g23771&g21012);
assign g11493 = ((~g8964)&(~g8967));
assign g26801 = ((~II25511));
assign II33070 = ((~g34810));
assign II24576 = (g5390&g5396&g9792);
assign g33784 = (g33107&g20531);
assign g24075 = ((~g19935));
assign g18109 = (g437&g17015);
assign g34753 = (g34676&g19586);
assign g30496 = (g30231)|(g21992);
assign II31131 = (g31542&g31819&g32643&g32644);
assign g12646 = ((~g9234)&(~g9206));
assign g34018 = (g33887)|(g18505);
assign g24294 = (g4452&g22550);
assign g24718 = ((~g22182));
assign g33024 = (g32324)|(g21752);
assign g31858 = ((~g29385));
assign g34402 = (g34179)|(g25084);
assign g28179 = (g27494)|(g27474)|(g27445)|(g27421);
assign g11036 = (g9806&g5774);
assign g17762 = ((~g13000));
assign g31892 = (g31019)|(g21825);
assign g20217 = (g16221)|(g13523);
assign II31042 = (g32515&g32516&g32517&g32518);
assign g32038 = ((~g30934));
assign II14734 = ((~g9732))|((~II14733));
assign g13565 = ((~g11006));
assign II26439 = ((~g26549))|((~II26438));
assign g8829 = ((~g5011))|((~g4836));
assign g33590 = (g33358)|(g18470);
assign g34929 = ((~II33179));
assign g9334 = ((~g827))|((~g832));
assign g15064 = ((~g6820)&(~g13394));
assign g27664 = (g1024&g25911);
assign g25129 = (g17682&g23527);
assign g28475 = ((~g3863)&(~g27635));
assign II31146 = (g30735&g31821&g32666&g32667);
assign g32046 = (g10925&g30735);
assign g15715 = ((~g336))|((~g305))|((~g13385));
assign g32907 = ((~g30937));
assign g32230 = (g30589)|(g29345);
assign g32551 = ((~g30735));
assign g7563 = ((~g6322));
assign g28867 = ((~g27800))|((~g2227))|((~g2153));
assign g25579 = (g19422&g24147);
assign g32515 = ((~g30825));
assign g27088 = ((~g26694));
assign g25449 = (g6946&g22496);
assign g29202 = (g24088&II27508&II27509);
assign g23848 = ((~g19210));
assign g13706 = ((~g11280));
assign II24674 = (g19919&g24019&g24020&g24021);
assign g29625 = (g28514&g14226);
assign g17596 = ((~g8686))|((~g14367));
assign g32935 = ((~g31672));
assign g10142 = ((~II13637));
assign g11489 = ((~g9661))|((~g3618));
assign g10421 = ((~g6227)&(~g9518));
assign g21941 = (g5232&g18997);
assign g27131 = (g26055&g16588);
assign g31286 = (g30159&g27858);
assign g32580 = ((~g30825));
assign g11571 = ((~g10323)&(~g3512)&(~g3506));
assign g32517 = ((~g31194));
assign g9618 = ((~g5794));
assign II31659 = ((~g33219));
assign II22143 = ((~g20189));
assign g34622 = (g34520)|(g18584);
assign g25836 = (g25368)|(g23856);
assign g11941 = ((~II14761));
assign g11915 = (g1802&g7315);
assign g27351 = (g10218&g26804);
assign g27984 = ((~g26737));
assign g9779 = ((~g5156));
assign g33163 = ((~g32099)&(~g7809));
assign II22470 = ((~g21326));
assign g8181 = ((~g424));
assign g7611 = ((~g4057))|((~g4064));
assign g29223 = (g28341)|(g18131);
assign g26766 = (g10776)|(g24460);
assign g11780 = ((~g4899)&(~g8822));
assign g16539 = (g11547&g6782&g6789&II17741);
assign g32148 = (g31631&g29981);
assign g29637 = (g2533&g29134);
assign g14313 = ((~g12016)&(~g9250));
assign g9890 = ((~g6058));
assign g18682 = (g4646&g15885);
assign g24198 = (g351&g22722);
assign g34949 = ((~g34939));
assign II31810 = ((~g33164));
assign II24462 = ((~g23796))|((~II24461));
assign g21728 = (g3010&g20330);
assign II24455 = ((~g22541));
assign g34648 = ((~II32752));
assign g31213 = ((~II29013));
assign g11607 = ((~g8848)&(~g8993)&(~g376));
assign g30453 = (g29902)|(g21862);
assign g26026 = ((~II25105));
assign II11726 = ((~g4273));
assign g23492 = ((~g21562));
assign g18345 = (g1736&g17955);
assign g32822 = ((~g30937));
assign g23888 = ((~g18997));
assign g13058 = ((~g10544))|((~g1312));
assign g18182 = (g776&g17328);
assign II21226 = ((~g16540));
assign g32163 = (g3502&g31170);
assign II24278 = ((~g23440));
assign II30261 = (g29385)|(g31376)|(g30735)|(g30825);
assign g31672 = (g29814&g19050);
assign g31789 = (g30201&g24013);
assign g34003 = (g33866)|(g18452);
assign g15652 = (g174&g13437);
assign g32218 = (g31130)|(g29619);
assign g32729 = ((~g30937));
assign g28644 = (g27387)|(g16593);
assign II22945 = ((~g9492))|((~II22944));
assign g18776 = (g5813&g18065);
assign g19360 = ((~g16249));
assign g29842 = (g28372&g23284);
assign g10838 = (g7738&g5527&g5535);
assign g19266 = (g246&g16214);
assign II30718 = (g32348)|(g32356)|(g32097)|(g32020);
assign g26483 = ((~II25359));
assign g30529 = (g30212)|(g22075);
assign g9104 = ((~II12987));
assign g28668 = (g27411)|(g16617);
assign II14516 = ((~g10147))|((~g661));
assign g34846 = ((~II33064));
assign g29798 = (g28348&g23260);
assign g14000 = ((~g8766)&(~g12259));
assign g34226 = (g33914&g21467);
assign g7166 = ((~g4311));
assign g23008 = (g1570&g19783);
assign g8609 = ((~g1171))|((~g1157));
assign g29902 = (g28430&g23377);
assign gbuf122 = (g344);
assign g8594 = ((~g3849));
assign g22129 = (g6633&g19277);
assign g22681 = ((~II21993))|((~II21994));
assign g27136 = (g26026&g16605);
assign g18133 = (g15055&g17249);
assign g7845 = ((~g1146));
assign II31727 = ((~g33076));
assign gbuf129 = (g881);
assign g19644 = ((~g17953));
assign g24635 = (g19874&g22883);
assign II31770 = ((~g33197));
assign g25850 = (g3502&g24636);
assign g28286 = (g27090)|(g15757);
assign g26964 = (g26259)|(g24316);
assign g29747 = (g28286&g23196);
assign g12364 = ((~g10102)&(~g10224));
assign g22853 = ((~g20219))|((~g2922));
assign g13998 = (g6589&g12629);
assign II14923 = ((~g9558))|((~g5835));
assign g31757 = (g29992)|(g30010);
assign g32798 = ((~g31672));
assign g18626 = (g3498&g17062);
assign g25111 = ((~g23699));
assign II32449 = ((~g34127));
assign II17314 = ((~g14078));
assign g29505 = ((~g29186));
assign g14093 = ((~g8833)&(~g11083));
assign g34979 = (g34875)|(g34968);
assign g26226 = (g24688&g8812&g10658&g10627);
assign g24980 = ((~g22384));
assign g30212 = (g28687&g23879);
assign g23354 = ((~g20453));
assign g6820 = ((~g1070));
assign g8572 = ((~II12654));
assign g30138 = (g28595&g21182);
assign g20097 = ((~g17691));
assign II31071 = (g31170&g31808&g32557&g32558);
assign g30406 = (g29783)|(g21765);
assign g26842 = (g2894&g24522);
assign g33491 = (g32679&II31151&II31152);
assign g16349 = ((~II17661));
assign g20498 = ((~g15348));
assign g30171 = ((~g28880)&(~g7431));
assign g26897 = (g26611)|(g18176);
assign II30123 = (g29385)|(g31376)|(g30735)|(g30825);
assign g24422 = (g4771&g22896);
assign g32946 = ((~g31327));
assign g29385 = ((~g28180));
assign II17159 = ((~g13350));
assign g28958 = ((~g27833))|((~g8249));
assign II22755 = ((~g21434))|((~II22753));
assign g33015 = (g32343)|(g18507);
assign g32660 = ((~g30825));
assign g11206 = ((~II14276))|((~II14277));
assign g17688 = ((~II18667));
assign g32749 = ((~g31021));
assign g25016 = ((~g23666));
assign g7994 = ((~II12336));
assign g25779 = ((~g19694))|((~g24362));
assign g11988 = ((~II14836));
assign g21760 = (g3207&g20785);
assign g34655 = (g34573&g18885);
assign g15804 = (g3223&g13889);
assign II13382 = ((~g269))|((~g246));
assign g29134 = ((~g9762))|((~g27907));
assign g32449 = ((~II29977));
assign g34395 = (g34193&g21336);
assign g21421 = ((~g15171));
assign g25653 = (g24664)|(g18602);
assign g25459 = (g6058&g23844&II24582);
assign g12249 = ((~g5763)&(~g10096));
assign g18617 = (g3462&g17062);
assign g25258 = ((~II24439))|((~II24440));
assign g15669 = ((~g11945)&(~g14272));
assign g32740 = ((~g31672));
assign g14899 = ((~g12744))|((~g10421));
assign II14570 = ((~g7932));
assign g15153 = ((~g13745)&(~g12897));
assign g16291 = ((~g13551))|((~g13545));
assign g32156 = (g31639&g30018);
assign g12899 = ((~g10407));
assign g32732 = ((~g30825));
assign II20462 = ((~g14187))|((~II20460));
assign g28630 = (g27544&g20575);
assign g24299 = (g4456&g22550);
assign g24708 = (g16474&g22998);
assign g12025 = ((~g9705)&(~g7461));
assign II20954 = ((~g16228));
assign g22026 = (g5913&g19147);
assign II18633 = ((~g2504))|((~g14713));
assign g25989 = (g25258&g21012);
assign g8346 = ((~g3845));
assign g9217 = (g632&g626);
assign g29324 = (g29078&g18883);
assign g24028 = ((~g20841));
assign g29651 = (g2537&g29134);
assign g13510 = ((~II15981));
assign g31327 = (g19200&g29814);
assign g32504 = ((~g30673));
assign g30918 = (g8681&g29707);
assign II25586 = ((~g25537));
assign g17846 = ((~g6271))|((~g14575))|((~g6365))|((~g12672));
assign g22543 = ((~g19801));
assign II31820 = ((~g33323));
assign g28194 = (g22540)|(g27122);
assign g23575 = ((~II22711))|((~II22712));
assign g20514 = ((~g15348));
assign g25703 = (g25087)|(g21922);
assign g25569 = (II24684&II24685);
assign g12035 = ((~g10000))|((~g6144));
assign g21359 = ((~g11509))|((~g17157));
assign g26649 = ((~g9037)&(~g24732));
assign II17173 = ((~g13716));
assign g21348 = (g10121&g17625);
assign g22668 = ((~g20219))|((~g2912));
assign g34432 = ((~II32467));
assign g28124 = (g27368&g22842);
assign II30740 = (g31776)|(g32188)|(g32083)|(g32087);
assign g24994 = ((~g22432));
assign g24081 = ((~g21209));
assign g27992 = (g26800&g23964);
assign g19783 = ((~g16931));
assign g7980 = ((~g3161));
assign II28851 = ((~g29317));
assign g9745 = ((~g6537));
assign g28247 = (g27147&g19675);
assign II18135 = ((~g13144));
assign g26086 = (g9672&g25255);
assign g33147 = ((~g32090)&(~g7788));
assign g32624 = ((~g30825));
assign g18457 = (g2319&g15224);
assign g23025 = (g16021&g19798);
assign g27588 = (g26690&g26673);
assign g33820 = (g33075&g26830);
assign g14445 = ((~g12188)&(~g9693));
assign g33814 = (g33098&g28144);
assign g19689 = ((~g16795));
assign g16162 = ((~g13437));
assign II29233 = ((~g30295));
assign g29650 = (g28949&g22472);
assign g30566 = (g26247&g29507);
assign g31323 = (g30150&g27907);
assign g29040 = ((~g6209)&(~g26977));
assign g6928 = ((~II11716));
assign g30247 = (g28735&g23937);
assign II18681 = ((~g2638))|((~II18680));
assign g14681 = (g4392&g10476);
assign g25992 = (g2485&g25024);
assign g29015 = ((~g27742))|((~g9586));
assign g14515 = ((~g12225)&(~g9761));
assign g33113 = (g31964&g22339);
assign II12218 = ((~g1437))|((~II12217));
assign g34304 = ((~II32309));
assign g34495 = (g34274&g19365);
assign g20242 = ((~g16308));
assign g24585 = ((~g23063));
assign g34690 = ((~II32840));
assign g25962 = (g9258&g24971);
assign g23858 = ((~g18997));
assign g8286 = ((~g53));
assign II22589 = ((~g21340));
assign g11398 = ((~II14409));
assign g13479 = ((~g12686))|((~g12639))|((~g12590))|((~g12526));
assign g22537 = ((~g19720)&(~g1367));
assign g22926 = ((~g20391));
assign g12228 = ((~g10222)&(~g10206)&(~g10184)&(~g10335));
assign g25056 = (g12779&g23456);
assign g28637 = (g22399&g27011);
assign g27273 = ((~g10504))|((~g26131))|((~g26105));
assign g25700 = (g25040)|(g21919);
assign g31897 = (g31237)|(g24322);
assign g18752 = (g15146&g17926);
assign g34202 = ((~II32161));
assign g24086 = ((~g20998));
assign g22069 = (g6227&g19210);
assign g33892 = (g33312&g20701);
assign II22930 = ((~g12223))|((~II22929));
assign g11123 = (g5644&g7028&g5630&g9864);
assign II29263 = ((~g12046))|((~II29261));
assign g30095 = (g28545&g20768);
assign g11130 = ((~g1221))|((~g7918));
assign g33587 = (g33363)|(g18463);
assign g24326 = (g4552&g22228);
assign II12468 = ((~g405))|((~g392));
assign g8292 = ((~g218))|((~g215));
assign g24258 = (g22851)|(g18311);
assign g18590 = (g2917&g16349);
assign II31474 = ((~g33212));
assign g32578 = ((~g31376));
assign g20505 = ((~g15426));
assign II15128 = ((~g9914))|((~g2527));
assign g10812 = ((~II14050));
assign g19273 = ((~g16100));
assign g26187 = ((~II25190));
assign II13862 = (g7232&g7219&g7258);
assign II14790 = ((~g6167))|((~II14788));
assign g23864 = ((~g19210));
assign gbuf21 = (g5327);
assign g17774 = ((~g14902));
assign g23816 = ((~g21308));
assign g32589 = ((~g31070));
assign g26424 = ((~II25356));
assign g27434 = (g26549&g17584);
assign II31046 = (g29385&g32521&g32522&g32523);
assign g25765 = (g24989&g24973);
assign g29768 = (g22760)|(g28229);
assign g30551 = (g30235)|(g22122);
assign g22093 = (g6423&g18833);
assign g11011 = ((~g10274));
assign g17520 = ((~g5260))|((~g12002))|((~g5276))|((~g14631));
assign g31746 = (g30093&g23905);
assign g22984 = ((~g20114))|((~g2868));
assign g26147 = (g6513&g25133);
assign g20774 = ((~g18008));
assign g28577 = (g27326)|(g26272);
assign g17015 = ((~II18143));
assign II29981 = ((~g31591));
assign g33120 = ((~II30686));
assign g24290 = (g4430&g22550);
assign g22688 = ((~g20219))|((~g2936));
assign g24269 = (g23131)|(g18613);
assign g18535 = (g2741&g15277);
assign g29814 = ((~II28062));
assign g16842 = (g6279&g14861);
assign g16643 = ((~II17839));
assign II13581 = ((~g6727));
assign II24364 = ((~g23687))|((~II24363));
assign g19521 = (g513&g16739);
assign g22516 = (g21559)|(g12817);
assign g29967 = ((~g28946));
assign g24317 = (g4534&g22228);
assign g29989 = (g29006&g10489);
assign g13955 = ((~g11621))|((~g11527));
assign g14276 = ((~II16452));
assign g34800 = (g34752)|(g18586);
assign II27238 = ((~g27320));
assign g19984 = ((~g17096)&(~g8171));
assign g7888 = ((~g1536));
assign g18527 = ((~II19345));
assign g14720 = ((~g12593))|((~g10266));
assign g20154 = ((~II20412));
assign g14177 = ((~g11741))|((~g11721))|((~g753));
assign g21937 = (g5208&g18997);
assign g32264 = (g31187)|(g29711);
assign g18166 = (g655&g17433);
assign g28592 = (g27333)|(g26288);
assign g30549 = (g30215)|(g22120);
assign g24935 = (g22937)|(g19749);
assign II15569 = ((~g11965));
assign II24331 = ((~g22976));
assign g32373 = (g29894)|(g31321);
assign g13933 = ((~g11419));
assign g31834 = ((~g29385));
assign g10883 = (g3355&g9061);
assign g33964 = (g33817)|(g18146);
assign g17763 = ((~g15011));
assign g25698 = (g25104)|(g21917);
assign g10601 = ((~g896))|((~g7397));
assign g21301 = ((~g11371))|((~g17157));
assign g30067 = ((~g29060));
assign II27561 = ((~g28163));
assign g21975 = (g5523&g19074);
assign II22343 = ((~g19371));
assign II22180 = ((~g21366));
assign g11312 = ((~g8565))|((~g3794));
assign II22972 = ((~g9657))|((~g19638));
assign g30597 = (g13564)|(g29693);
assign g29486 = (g28537)|(g27595);
assign II17650 = ((~g13271));
assign g28317 = (g27114)|(g15805);
assign g11427 = (g5706&g7158);
assign g33640 = (g33387&g18831);
assign g34865 = (g16540&g34836);
assign g12461 = ((~g7536))|((~g6000));
assign g15728 = ((~g5200))|((~g14399))|((~g5313))|((~g9780));
assign g19865 = ((~g15885));
assign g19596 = (g1094&g16681);
assign g16178 = (g5845&g14297);
assign g24162 = ((~II23330));
assign g33314 = (g29663)|(g32174);
assign g8522 = ((~g298));
assign g18716 = (g4878&g15915);
assign g32050 = (g11003&g30825);
assign g11497 = (g6398&g7192);
assign g33760 = (g33143&g20328);
assign g15752 = ((~g5921))|((~g12129))|((~g5983))|((~g14701));
assign g22134 = (g6653&g19277);
assign g16246 = ((~g13551)&(~g11169));
assign g23232 = ((~II22331));
assign g22487 = (g21512)|(g12794);
assign g26335 = (g1526)|(g24609);
assign g12357 = ((~g7439))|((~g6329));
assign g33859 = (g33426&g10531);
assign g32296 = ((~g9044)&(~g31509)&(~g12259));
assign g32043 = (g31482&g16173);
assign g16299 = ((~g8160))|((~g8112))|((~g13706));
assign g31624 = ((~II29218));
assign g32679 = ((~g31579));
assign g18245 = (g1193&g16431);
assign g6867 = ((~II11685));
assign II26530 = (g26365&g24096&g24097&g24098);
assign g9229 = ((~g5052));
assign g32801 = ((~g30937));
assign g31945 = ((~g31189));
assign g7266 = ((~g35));
assign g22450 = ((~g19345)&(~g15724));
assign g28768 = (g21434&g26424&g25308&g27421);
assign g21802 = (g3562&g20924);
assign g31468 = (g29641)|(g29656);
assign g9880 = ((~g5787));
assign II13623 = ((~g4294));
assign g28133 = (g27367&g23108);
assign g24019 = ((~g19968));
assign g12119 = ((~g2351))|((~g8267));
assign g28332 = (g27130)|(g15815);
assign g19393 = (g691&g16325);
assign g10909 = ((~g7304))|((~g1116));
assign g13289 = (g10619)|(g10624);
assign g24667 = ((~g23112));
assign g33535 = (g33233)|(g21711);
assign g12042 = ((~g9086))|((~g703));
assign g6959 = ((~g4420));
assign g21401 = ((~g17755))|((~g14730))|((~g17712))|((~g14695));
assign g19556 = (g11932&g16809);
assign g16592 = (g5579&g14688);
assign g33455 = ((~II30983));
assign g34855 = ((~II33079));
assign g29889 = ((~g6905)&(~g28471));
assign g33197 = (g32342)|(II30745)|(II30746);
assign g31843 = ((~g29385));
assign g29519 = (g2295&g28840);
assign g33647 = (g33390&g18878);
assign g23258 = ((~g20924));
assign g7858 = ((~g947));
assign g12881 = ((~g10388));
assign g33712 = ((~II31561));
assign g25293 = ((~g21190))|((~g23726));
assign g31994 = (g31775&g22215);
assign II33232 = ((~g34957));
assign g27376 = (g26549&g17481);
assign g17010 = ((~II18138));
assign g12295 = ((~g7139));
assign g13919 = ((~g3347)&(~g11276));
assign g27501 = (g26400&g17673);
assign g13029 = (g8359&g11030);
assign gbuf32 = (g5673);
assign gbuf48 = (g6351);
assign g16476 = ((~g8119)&(~g13667));
assign II29199 = ((~g30237));
assign g14707 = ((~g10143)&(~g12259));
assign g23375 = ((~g20924));
assign g13823 = ((~g11313))|((~g3774));
assign g10623 = ((~g10181))|((~g9976));
assign g9730 = ((~g5436));
assign g18483 = (g2453&g15426);
assign g18088 = ((~g13267));
assign g11449 = (g6052&g7175);
assign II23375 = ((~g23403));
assign gbuf28 = (g5666);
assign II28925 = ((~g29987));
assign g22529 = ((~g19549));
assign g25926 = (g25005&g24839);
assign g33289 = (g32148)|(g29588);
assign g7343 = ((~g5290));
assign g10412 = ((~g7072));
assign g21757 = (g3187&g20785);
assign II22000 = ((~g20277));
assign II24759 = ((~g24229));
assign g34198 = (g33688&g24491);
assign gbuf87 = (g3668);
assign II15004 = ((~g1700))|((~II15002));
assign g15138 = ((~g13680)&(~g6993));
assign g21416 = ((~g17775))|((~g14781))|((~g17744))|((~g14706));
assign g15344 = ((~g14851));
assign g21893 = (g20094)|(g18655);
assign g15097 = ((~g12868)&(~g13191));
assign g22150 = ((~g21280));
assign g7917 = ((~g1157));
assign g28998 = (g17424&g25212&g26424&g27474);
assign g14216 = (g7631&g10608);
assign g28699 = (g27452)|(g16667);
assign g32018 = (g4146&g30937);
assign g31314 = (g30183&g27937);
assign g11846 = ((~g7635)&(~g7518)&(~g7548));
assign g23058 = ((~g20453));
assign g16522 = ((~g13889));
assign II23384 = ((~g23362));
assign g16053 = ((~II17442));
assign g12471 = ((~II15288))|((~II15289));
assign II20116 = ((~g15737));
assign g10573 = ((~g7992))|((~g8179));
assign g11252 = ((~g8620)&(~g3057));
assign g18307 = (g1559&g16931);
assign g33993 = (g33646)|(g18413);
assign g24504 = (g22226&g19410);
assign g33449 = ((~g10311)&(~g31950));
assign g33136 = ((~g32057));
assign g34058 = ((~g33660));
assign g26878 = (g25578)|(g25579);
assign II27749 = ((~g28917));
assign g24981 = ((~g22763));
assign g22227 = ((~g19801));
assign g32361 = (g29869)|(g31300);
assign gbuf154 = (g1116);
assign g29730 = (g28150)|(g28141);
assign II29939 = ((~g31667));
assign g30671 = (g29319&g22317);
assign g31857 = ((~g29385));
assign g27771 = ((~g9809)&(~g25839));
assign g25729 = (g25091)|(g22012);
assign g17419 = ((~g14965));
assign g23868 = ((~g19277));
assign g21829 = (g3770&g20453);
assign g7369 = ((~g1996));
assign g24036 = ((~g20982));
assign g32899 = ((~g31021));
assign g10178 = ((~g2126));
assign g27364 = ((~g8426)&(~g26616));
assign g33394 = ((~g10159))|((~g4474))|((~g32426));
assign g25173 = (g12234&g23589);
assign g34627 = (g34534)|(g18644);
assign g18721 = (g15138&g16077);
assign g25523 = ((~g22550));
assign g20452 = ((~g17200));
assign g16676 = ((~II17876));
assign g33440 = (g32250&g29719);
assign g28685 = (g27433)|(g16637);
assign g25761 = (g25152)|(g18812);
assign g32974 = ((~g30937));
assign g22761 = ((~g21024));
assign gbuf140 = (g1570);
assign g33850 = ((~II31701));
assign g13121 = ((~g11117))|((~g8411));
assign g29298 = (g28571)|(g18793);
assign g23248 = ((~g20924));
assign g14347 = ((~g9309)&(~g11123));
assign g14640 = ((~g12371)&(~g9824));
assign g13035 = (g8497&g11033);
assign g21781 = (g3408&g20391);
assign II11716 = ((~g4054));
assign gbuf59 = (g6697);
assign g28512 = ((~g10857))|((~g27155))|((~g27142));
assign g34500 = (g34276&g30568);
assign g15074 = ((~g12845)&(~g13416));
assign g24057 = ((~g20841));
assign g15678 = (g1094&g13846);
assign g12641 = (g10295&g3171&g3179);
assign g12821 = ((~g7132)&(~g10223)&(~g7149)&(~g10261));
assign g28232 = (g27732&g23586);
assign g19495 = ((~g15969))|((~g10841))|((~g7781));
assign g34437 = ((~II32482));
assign g8405 = ((~II12572));
assign g31639 = ((~II29225));
assign g21874 = (g4112&g19801);
assign g26347 = (g262&g24850);
assign g29884 = (g2555&g29153);
assign g34448 = (g34365)|(g18553);
assign II33027 = ((~g34767));
assign g14921 = ((~g12492))|((~g10266));
assign g31516 = (g29848&g23476);
assign g14546 = ((~g12125))|((~g9613));
assign g10388 = ((~g6983));
assign II21941 = ((~g18918));
assign g21670 = ((~g16540));
assign g33254 = (g32104)|(g29512);
assign g15588 = ((~II17166));
assign g34119 = (g20516&g9104&g33755);
assign g30198 = (g28662&g23860);
assign g18749 = (g5148&g17847);
assign g28079 = ((~II26578));
assign g34982 = ((~II33246));
assign II29579 = ((~g30565));
assign II24508 = (g9434&g9672&g5401);
assign g18930 = ((~g15789));
assign g6811 = ((~g714));
assign g26852 = (g24975&g24958);
assign g12976 = ((~II15587));
assign g17125 = ((~II18177));
assign g23678 = ((~g9809)&(~g21190));
assign g8770 = ((~g749));
assign g18238 = (g1152&g16326);
assign g26182 = (g9978&g25317);
assign g31069 = (g29793&g14150);
assign g28152 = (g26297&g27279);
assign g16599 = (g6601&g15030);
assign II14409 = ((~g8364));
assign g24757 = (g7004&g23563);
assign g19768 = (g2803&g15833);
assign g24773 = (g22832&g19872);
assign g31297 = (g30144&g27837);
assign g13907 = ((~g3941))|((~g11225))|((~g4023))|((~g11631));
assign g12543 = ((~g9417));
assign g18512 = (g2619&g15509);
assign g34266 = (g34076)|(g18719);
assign g23896 = ((~g19210));
assign g24574 = ((~g22709))|((~g22687));
assign g30144 = ((~g28789)&(~g7322));
assign g31520 = (g29879&g23507);
assign g19577 = ((~g16129));
assign g20040 = ((~g17271));
assign g11317 = ((~II14346));
assign g34429 = ((~II32458));
assign g33359 = (g32252&g20853);
assign g15081 = (g2689&g12983);
assign g17312 = ((~g7297))|((~g14248));
assign g8093 = ((~g1624));
assign g25714 = (g25056)|(g21965);
assign g8300 = ((~g1242));
assign g27796 = ((~g21228))|((~g25263))|((~g26424))|((~g26171));
assign g34957 = (g34948)|(g21662);
assign g18222 = (g1024&g16100);
assign g29474 = ((~II27758));
assign g6998 = ((~g4932));
assign g11888 = ((~g10160));
assign g21186 = ((~g14616))|((~g17363));
assign g29570 = (g2763&g28598);
assign g32249 = (g31169)|(g29687);
assign g21294 = ((~g11324))|((~g17157));
assign g7517 = ((~g962));
assign g26940 = (g25908)|(g21886);
assign II31106 = (g30825&g31814&g32608&g32609);
assign II18323 = ((~g13680));
assign g19493 = ((~g16349));
assign II31231 = (g31376&g31836&g32789&g32790);
assign II26095 = ((~g13539))|((~II26093));
assign g30297 = ((~g28758));
assign g15088 = ((~g13144)&(~g6874));
assign g19482 = ((~g16349));
assign II29441 = ((~g30917));
assign g23414 = ((~II22525));
assign g24491 = (g10727&g22332);
assign g23823 = ((~II22989));
assign g17576 = ((~g14953));
assign g11283 = ((~g7953)&(~g4991)&(~g9064));
assign g18815 = (g6523&g15483);
assign g25246 = ((~g23828));
assign g12778 = ((~g9856));
assign g30244 = (g28732&g23930);
assign g33928 = ((~II31800));
assign g25534 = ((~g22763));
assign g31241 = (g25959)|(g29510);
assign g17656 = ((~II18626))|((~II18627));
assign g26671 = (g316&g24429);
assign g11294 = ((~g7598));
assign g8792 = ((~II12790));
assign II31597 = ((~g33187));
assign g15103 = (g4180&g14454);
assign g17603 = ((~g14993));
assign g10796 = ((~g7537))|((~g7523));
assign g30101 = (g28551&g20780);
assign g24671 = (g5481&g23630);
assign g11920 = ((~II14730));
assign g18442 = (g2259&g18008);
assign g24964 = ((~II24128));
assign g25212 = ((~g22763));
assign g23477 = ((~g21468));
assign g33884 = (g33295&g20590);
assign g31149 = (g29508&g23021);
assign g13133 = ((~g11330));
assign g27391 = (g26549&g17505);
assign g25079 = (g21011&g23483);
assign g14590 = ((~g3546))|((~g11207))|((~g3680))|((~g8542));
assign g23273 = ((~g21070));
assign g22995 = ((~g20330));
assign g34984 = ((~II33252));
assign g29760 = (g28309&g23227);
assign g16959 = (g13542)|(g11142);
assign II15255 = ((~g1848))|((~II15253));
assign II15149 = ((~g5659))|((~II15147));
assign g19653 = ((~g16897));
assign g25631 = (g24554)|(g18275);
assign II12729 = ((~g4291))|((~II12728));
assign g11753 = ((~g8587));
assign g23237 = ((~g20924));
assign g12755 = ((~g6555)&(~g9407));
assign g21279 = ((~g15680));
assign g18212 = (g947&g15979);
assign g29056 = ((~g27800));
assign g33574 = (g33362)|(g18416);
assign g22130 = (g6637&g19277);
assign g13929 = ((~g11669))|((~g11763));
assign g17926 = ((~II18852));
assign g29187 = ((~g7704)&(~g27999));
assign g14780 = ((~g6275))|((~g12101))|((~g6329))|((~g12423));
assign g9280 = ((~II13054));
assign II20753 = ((~g16677));
assign g13260 = ((~g1116))|((~g10666));
assign g26249 = (g1858&g25300);
assign g19657 = ((~g16349));
assign g29576 = (g2177&g28903);
assign II16741 = ((~g5677));
assign g28522 = ((~g10857))|((~g26131))|((~g27142));
assign g14510 = ((~II16629));
assign g21990 = (g5591&g19074);
assign II29913 = ((~g30605));
assign g24748 = (g17656&g22457);
assign g31793 = (g28031)|(g30317);
assign g28227 = (g9397&g27583);
assign II13424 = ((~g5689));
assign g30289 = (g28884&g24000);
assign g29285 = (g28639)|(g18750);
assign g22172 = (g8064&g19857);
assign g23132 = ((~g8155))|((~g19932));
assign g18759 = (g5467&g17929);
assign g22049 = (g6082&g21611);
assign II31361 = ((~g33120));
assign II22425 = ((~g19379));
assign g18410 = (g2079&g15373);
assign g9024 = ((~g4358));
assign II29313 = ((~g29501))|((~g12154));
assign g29167 = ((~g9576)&(~g26994));
assign g30591 = ((~II28851));
assign g27599 = (g26337&g20033);
assign g27238 = (g25879)|(g24464);
assign g23239 = ((~g21308));
assign g8538 = ((~g3412));
assign g34285 = ((~II32284));
assign g26351 = (g239&g24869);
assign II15121 = ((~g9910))|((~g2102));
assign g25076 = (g12805&g23479);
assign g18420 = (g1996&g15373);
assign g19200 = ((~II19789));
assign g29343 = ((~g28174));
assign g12219 = (g1189&g7532);
assign g7133 = ((~II11825))|((~II11826));
assign g16430 = (g182)|(g13657);
assign g29708 = (g1955&g29082);
assign g22097 = (g6451&g18833);
assign II14567 = ((~g9708));
assign g9250 = ((~g1600));
assign g17490 = (g14364)|(g14337)|(g11958)|(II18421);
assign g23435 = ((~g18833));
assign g30135 = (g28592&g21180);
assign g23695 = ((~g17420)&(~g21140));
assign II14205 = ((~g8508))|((~II14204));
assign II13606 = ((~g74));
assign II31302 = (g32891&g32892&g32893&g32894);
assign g23946 = ((~g19210));
assign II19786 = ((~g17844));
assign g7870 = ((~g1193));
assign g25944 = ((~g7716)&(~g24591));
assign g32311 = (g31295&g20582);
assign g19374 = ((~g16047));
assign g23151 = (g18994&g7162);
assign g24660 = (g22648&g19737);
assign g22884 = ((~g20453));
assign g18678 = (g66&g15758);
assign g29307 = (g28706)|(g18814);
assign g10567 = ((~g1862))|((~g7405));
assign II25219 = ((~g482))|((~g24718));
assign II17976 = ((~g13638));
assign g29275 = (g28165)|(g21868);
assign g10116 = ((~g2413));
assign g23319 = (g19717)|(g16193);
assign g32607 = ((~g31542));
assign g16782 = ((~II18006));
assign g21336 = ((~g17367));
assign g19466 = ((~g11562))|((~g17794));
assign g23014 = ((~g20391));
assign g28063 = (g27541)|(g21773);
assign g32333 = (g31326&g23559);
assign g10654 = (g3085&g8434);
assign g17754 = ((~g14262));
assign g24555 = (g23184&g21024);
assign g10093 = ((~g5703));
assign II18434 = ((~g13782));
assign g27158 = (g26609&g16645);
assign II14727 = ((~g7753));
assign g26575 = ((~g25268));
assign g23938 = ((~g18997));
assign II12523 = ((~g3794));
assign g34522 = ((~g34271));
assign II29253 = ((~g29482))|((~g12017));
assign g10590 = (g7246&g7392&II13937);
assign g13833 = (g4546&g10613);
assign g11303 = ((~g8497)&(~g8500));
assign g9687 = ((~II13287));
assign g17746 = ((~g14825));
assign II17148 = ((~g14442));
assign g25574 = (II24709&II24710);
assign g22872 = (g19372)|(g19383);
assign g34729 = (g34666)|(g18270);
assign g22062 = (g6093&g21611);
assign g13099 = ((~II15732));
assign II20488 = ((~g16757))|((~II20486));
assign g25051 = ((~II24215));
assign g15566 = ((~II17143));
assign g8285 = ((~II12497));
assign g24152 = ((~II23300));
assign g34463 = (g34338)|(g18686);
assign II11825 = ((~g4593))|((~II11824));
assign g11003 = (g7880&g1300);
assign g25410 = ((~g22228));
assign g16320 = ((~g14454));
assign g21742 = (g3050&g20330);
assign II11801 = ((~g6395));
assign g6808 = ((~g554));
assign g30533 = (g30203)|(g22079);
assign II17166 = ((~g14536));
assign g31493 = (g29791&g23434);
assign II18089 = ((~g13144));
assign g31863 = ((~II29447));
assign g28585 = (g27063&g10530);
assign g18918 = ((~II19704));
assign g30339 = (g29629)|(g18244);
assign g29338 = (g29145&g22181);
assign g28572 = (g27829&g15669);
assign II13057 = ((~g112));
assign II32763 = ((~g34511));
assign g25420 = (g6058&g22220&II24555);
assign g18267 = (g1266&g16000);
assign g34459 = (g34415)|(g18673);
assign gbuf80 = (g3096);
assign g25882 = ((~g25026));
assign II24237 = ((~g23823));
assign g22113 = (g6561&g19277);
assign g34241 = ((~II32222));
assign g17690 = (g11547&g11592&g11640&II18671);
assign g8085 = ((~II12382));
assign g34703 = ((~g8899)&(~g34545)&(~g11083));
assign g21765 = (g3231&g20785);
assign II12884 = ((~g4213));
assign g7072 = ((~g6199));
assign g24892 = (g11559&g23264);
assign g22542 = ((~g19801));
assign g18651 = (g15102&g16249);
assign g23780 = ((~II22930))|((~II22931));
assign g19743 = ((~g17125));
assign g33238 = (g32048)|(g32051);
assign g32577 = ((~g31554));
assign g16227 = ((~g1554)&(~g13574));
assign g33803 = (g33231&g20071);
assign g11044 = (g5343&g10124);
assign g29068 = (g27628)|(g17119);
assign g14232 = ((~g11083));
assign g31922 = (g31525)|(g22047);
assign g19434 = ((~g16326));
assign g28672 = (g7577&g27017);
assign g18293 = (g1484&g16449);
assign g24071 = ((~g20841));
assign g33228 = ((~II30766));
assign g22991 = (g645&g20248);
assign g26382 = ((~g577))|((~g24953))|((~g12323));
assign g32185 = ((~II29717));
assign g21912 = (g5052&g21468);
assign g24534 = ((~g22670));
assign g12845 = ((~g10358));
assign g12001 = ((~II14854))|((~II14855));
assign g10198 = ((~II13672));
assign II26644 = (g27057)|(g27044)|(g27039)|(g27032);
assign g28031 = ((~g21209)&(~II26522)&(~II26523));
assign g30600 = (g30287&g18975);
assign g28752 = ((~II27232));
assign g23418 = ((~g21468));
assign g18205 = (g904&g15938);
assign g18381 = (g1882&g15171);
assign g18463 = (g2375&g15224);
assign g24643 = (g22636&g19696);
assign II12631 = ((~g1242));
assign g13239 = ((~g10632));
assign g27313 = (g1982&g26701);
assign g29621 = (g2449&g28994);
assign II15299 = ((~g10112))|((~II15298));
assign g14069 = ((~g11653))|((~g8864));
assign II13694 = ((~g117));
assign II18104 = ((~g13177));
assign g8038 = ((~II12360));
assign g25100 = ((~g22384));
assign II17456 = ((~g13680));
assign II15937 = ((~g11676));
assign g10336 = ((~II13750))|((~II13751));
assign II12418 = ((~g55));
assign II19802 = ((~g15727));
assign II14399 = ((~g8542))|((~II14398));
assign II15080 = ((~g1968))|((~II15078));
assign g25943 = (g24423)|(g22299);
assign II17964 = ((~g3661));
assign g30201 = (g23412)|(g28557);
assign II13705 = ((~g63));
assign g16487 = ((~II17695));
assign II29977 = ((~g31596));
assign g25622 = (g24546)|(g18217);
assign g7952 = ((~g3774));
assign g24000 = ((~g19277));
assign g9826 = ((~g1844));
assign g25273 = ((~g23978));
assign g24516 = ((~g22670));
assign g21228 = ((~g17531));
assign g33060 = (g31992)|(g22022);
assign g29645 = (g1714&g29018);
assign g20200 = ((~II20461))|((~II20462));
assign g23566 = ((~g21562));
assign g27179 = (g25816)|(g24409);
assign g23928 = ((~g21562));
assign g13414 = ((~g11048));
assign g14638 = ((~g9626))|((~g12361));
assign g8914 = ((~g4264));
assign g28427 = (g27258&g20008);
assign g30237 = ((~II28480));
assign II29262 = ((~g29485))|((~II29261));
assign g23820 = ((~g19147));
assign II31803 = ((~g33176));
assign g14361 = ((~g12079)&(~g9413));
assign g27406 = (g26488&g17521);
assign II32956 = ((~g34654));
assign g20107 = ((~g11404))|((~g17794));
assign g12945 = ((~g12467));
assign g31963 = (g30731&g18895);
assign g24046 = ((~g21256));
assign g12951 = ((~II15569));
assign II11734 = ((~g4473));
assign g29978 = ((~g28927));
assign g11323 = ((~II14351))|((~II14352));
assign g20584 = ((~g17873));
assign g34480 = ((~II32535));
assign g24250 = (g22633)|(g18295);
assign g11118 = ((~II14170))|((~II14171));
assign g25271 = ((~II24462))|((~II24463));
assign g20112 = (g13540&g16661);
assign g23747 = ((~II22865))|((~II22866));
assign g18772 = (g5689&g15615);
assign g16171 = ((~g13530));
assign g34387 = ((~g34188));
assign g25736 = (g25536)|(g18785);
assign g26399 = (g15572&g25566);
assign g32391 = (g31502)|(g29982);
assign g31238 = (g29583&g20053);
assign g14088 = ((~g3901))|((~g11255))|((~g4000))|((~g11631));
assign II23962 = ((~g23184))|((~II23961));
assign g29697 = ((~g28336));
assign g25724 = (g25043)|(g22007);
assign g25604 = (g24717)|(g18115);
assign g34034 = (g33719)|(g18713);
assign g29920 = ((~g28824));
assign g32071 = (g27236&g31070);
assign g34658 = (g34574&g18896);
assign g12521 = ((~g7471))|((~g5969));
assign g21606 = (g15959&g13763);
assign g21866 = (g4072&g19801);
assign g22898 = ((~g20283));
assign gbuf132 = (g365);
assign g33571 = (g33367)|(g18409);
assign g13594 = ((~g11012));
assign g13496 = ((~g1351))|((~g11336))|((~g11815));
assign g14696 = ((~g5567))|((~g12093))|((~g5685))|((~g12563));
assign g21997 = (g5619&g19074);
assign g20500 = ((~g17873));
assign g33029 = (g32332)|(g21798);
assign II29444 = ((~g30928));
assign g13143 = ((~g10695))|((~g7661))|((~g979))|((~g1061));
assign g29476 = (g28108)|(g28112);
assign gbuf149 = (g1227);
assign g33323 = (g31936)|(g32442);
assign g34926 = ((~II33170));
assign g23719 = ((~II22845))|((~II22846));
assign g16723 = ((~g3606))|((~g13730))|((~g3676))|((~g11576));
assign g18479 = (g2449&g15426);
assign g11747 = ((~g3530)&(~g8114));
assign g23260 = ((~g21070));
assign g25780 = (g25532&g25527);
assign g20545 = ((~g15373));
assign g18693 = (g4717&g16053);
assign g24228 = (g862&g22594);
assign II20388 = ((~g17724));
assign g27734 = ((~g9733)&(~g25821));
assign g28368 = (g27158)|(g27184);
assign g20073 = ((~g16540));
assign g12129 = ((~g9992)&(~g7051));
assign g8650 = ((~g4664));
assign g25120 = ((~g22432));
assign g7503 = ((~g1351));
assign g20661 = ((~g15171));
assign g34938 = ((~g34920));
assign g22084 = (g6291&g19210);
assign g27187 = ((~II25882));
assign g18890 = (g10158&g17625);
assign II13751 = ((~g4584))|((~II13749));
assign g34836 = ((~II33050));
assign gbuf58 = (g6144);
assign g13100 = ((~g6581))|((~g12137))|((~g6692))|((~g10061));
assign g6772 = ((~II11629));
assign g28823 = ((~g27738))|((~g14565));
assign g33601 = (g33422)|(g18508);
assign g31991 = (g4912&g30673);
assign g26653 = ((~g25337));
assign g32695 = ((~g30735));
assign g21252 = ((~g15656));
assign g30557 = (g30247)|(g22128);
assign g34786 = ((~II32988));
assign g25552 = ((~g22594));
assign g10966 = (g9226&g7948);
assign g7446 = ((~g1256));
assign g30381 = (g30126)|(g18497);
assign g23554 = (g20390&g13024);
assign g21061 = ((~II20929));
assign g21919 = (g15144&g21468);
assign g15860 = (g3889&g14160);
assign II15175 = ((~g9977))|((~II15174));
assign g9733 = ((~g5736));
assign II15238 = ((~g6351));
assign g9693 = ((~g1886));
assign g16667 = (g5268&g14659);
assign g13943 = ((~II16231));
assign g19690 = ((~g16826));
assign g18780 = (g5827&g18065);
assign g31302 = (g29590)|(g28302);
assign g12805 = ((~g9511));
assign g31596 = ((~II29204));
assign g11912 = ((~g8989));
assign g23906 = ((~g19074));
assign g32532 = ((~g31170));
assign g32341 = (g31472&g23610);
assign g24713 = (g5831&g23666);
assign g19632 = ((~g1413))|((~g1542))|((~g16047));
assign g7659 = ((~II12141));
assign g30153 = (g28610&g23768);
assign g11985 = ((~II14827));
assign g27486 = (g26519&g17645);
assign II15788 = ((~g10430));
assign II33143 = ((~g34903));
assign g22653 = (g18993)|(g15654);
assign g13188 = ((~g10909));
assign g10409 = ((~g7087));
assign g10404 = ((~g7026));
assign g18149 = (g608&g17533);
assign g28618 = (g27357)|(g16516);
assign g24836 = ((~II24008));
assign g16703 = (g5889&g15002);
assign g15704 = (g3440&g13504);
assign g17134 = (g5619&g14851);
assign g19906 = ((~g16209)&(~g13672));
assign g10398 = ((~g6999));
assign g31227 = ((~g29744));
assign g31591 = (g29358)|(g29353);
assign g24369 = ((~II23586))|((~II23587));
assign II31786 = ((~g33197));
assign II30468 = (g29385)|(g31376)|(g30735)|(g30825);
assign g9018 = ((~g4273));
assign g16896 = (g262&g13120);
assign g33473 = (g32549&II31061&II31062);
assign II32601 = ((~g34319));
assign g31501 = (g2047&g29310);
assign g13094 = ((~g7487)&(~g10762));
assign g32190 = (g142&g31233);
assign g25284 = ((~II24474));
assign g8136 = ((~g269));
assign g33744 = ((~II31604));
assign g13335 = ((~g7851)&(~g10741));
assign g28182 = (g8770&g27349);
assign g8933 = ((~g4709)&(~g4785));
assign g33074 = (g32387&g18830);
assign g26939 = (g25907)|(g21884);
assign g19443 = ((~g16449));
assign g20630 = ((~g17955));
assign g25222 = ((~II24400));
assign g24976 = ((~g671)&(~g23324));
assign g34043 = (g33903)|(g33905);
assign g25636 = (g24507)|(g18305);
assign g33538 = (g33252)|(g18144);
assign g32288 = (g31226)|(g31229);
assign g11903 = ((~g9099))|((~g3712));
assign II12411 = ((~g4809));
assign g27738 = ((~g21228))|((~g25243))|((~g26424))|((~g26148));
assign II14671 = ((~g7717));
assign II15148 = ((~g9864))|((~II15147));
assign g9954 = ((~g6128))|((~g6120));
assign g26051 = (g24896&g14169);
assign g34997 = ((~II33291));
assign g11164 = ((~g8085));
assign g26268 = ((~g283)&(~g24825));
assign g32919 = ((~g30735));
assign II31037 = (g32508&g32509&g32510&g32511);
assign g13655 = ((~g10573));
assign g27291 = (g11969&g26653);
assign g34631 = (g34562)|(g15118);
assign g30424 = (g29760)|(g21808);
assign g12009 = ((~II14862));
assign g13384 = (g4944&g11804);
assign g31779 = (g30050)|(g28673);
assign g22904 = ((~II22111));
assign g22190 = ((~g2827)&(~g18949));
assign g9976 = ((~g2537));
assign II20223 = ((~g11170))|((~II20221));
assign g23517 = ((~g21070));
assign II33276 = ((~g34985));
assign g31763 = (g30127&g23965);
assign g31306 = (g29595)|(g29610);
assign g17499 = ((~g14885));
assign g24065 = ((~g20982));
assign g26279 = (g4249&g25213);
assign g15910 = (g13025)|(g10654);
assign g27699 = (g26396&g20766);
assign g12749 = ((~g7074));
assign II22665 = ((~g21308));
assign g22156 = ((~g19147));
assign g29092 = ((~g27800));
assign g25506 = ((~g22228));
assign g18197 = (g854&g17821);
assign g26759 = (g24468)|(g7511);
assign II31091 = (g29385&g32586&g32587&g32588);
assign g33044 = (g32199)|(g24327);
assign g23298 = (g19693)|(g16179);
assign g21772 = (g3259&g20785);
assign g8506 = ((~g3782));
assign g9910 = ((~g2108));
assign g22331 = (g21405)|(g17809);
assign g10130 = ((~g5694));
assign g24345 = (g23606)|(g18788);
assign g17137 = ((~g13727))|((~g13511))|((~g13527));
assign g24375 = ((~g22722));
assign g12944 = ((~g12659));
assign g21739 = (g3080&g20330);
assign g33414 = (g32367&g21421);
assign g34337 = (g34095&g19881);
assign g26715 = ((~g23711)&(~g25203));
assign g33277 = (g32129)|(g29568);
assign g26830 = ((~g24411));
assign g10129 = ((~g5352));
assign g27426 = (g25967)|(g24588);
assign II29371 = ((~g30325));
assign II18301 = ((~g12976));
assign g17479 = ((~g14855));
assign g34424 = ((~II32440))|((~II32441));
assign g25230 = ((~g23314));
assign g13664 = ((~g11252));
assign g15967 = (g3913&g14058);
assign g14382 = ((~g9390)&(~g11139));
assign II31207 = (g32754&g32755&g32756&g32757);
assign g21790 = (g3454&g20391);
assign g26511 = (g19265&g24364);
assign g24924 = ((~g20007))|((~g23172));
assign g24907 = (g21558)|(g24015);
assign g11560 = ((~g7647));
assign g28293 = (g7424&g2495&g27474);
assign g19050 = ((~II19759));
assign g24401 = (g23811)|(g21298);
assign g24900 = (g3752&g23582&II24067);
assign g29304 = (g28588)|(g18810);
assign g18819 = (g6541&g15483);
assign g34538 = (g34330&g20054);
assign g8672 = ((~g4669));
assign g23802 = (g9104&g19050);
assign II17857 = ((~g3969));
assign g32415 = ((~g31591));
assign g34292 = (g26853)|(g34223);
assign g11861 = ((~g8070));
assign g30222 = (g28701&g23894);
assign II16639 = ((~g4000));
assign II12016 = ((~g772));
assign g27722 = ((~g7247)&(~g25805));
assign g7542 = ((~II12030));
assign II28480 = ((~g28652));
assign g28210 = (g9229&g27554);
assign g7618 = ((~II12092));
assign g24319 = (g4561&g22228);
assign g12590 = ((~g7097))|((~g7110))|((~g10229));
assign II31974 = ((~g33631))|((~II31972));
assign g34063 = (g33806&g23121);
assign g9543 = ((~g2217))|((~g2185));
assign g34513 = (g9003&g34346);
assign g14227 = ((~g9863)&(~g10838));
assign g34903 = (g34859)|(g21690);
assign g21690 = ((~g16540));
assign g33699 = (g32409)|(g33433);
assign g31860 = ((~II29438));
assign g23982 = ((~g19147));
assign g14123 = ((~g10685))|((~g10928));
assign g30068 = ((~g29157));
assign g21794 = (g15094&g20924);
assign g23139 = ((~g21163))|((~g10756));
assign II32976 = ((~g34699));
assign g13973 = (g11024)|(g11028);
assign g34358 = ((~II32364));
assign g33817 = (g33235&g20102);
assign g30037 = ((~g29121));
assign g33846 = (g33259&g20380);
assign g27180 = (g26026&g16654);
assign g20924 = ((~II20895));
assign g31904 = (g31780)|(g21923);
assign g6997 = ((~g4578));
assign g29314 = (g29005&g22144);
assign g33879 = (g33289&g20566);
assign II23303 = ((~g21669));
assign g24758 = (g6523&g23733);
assign II20467 = ((~g16663))|((~g16728));
assign g33617 = (g33263)|(g24326);
assign II18224 = ((~g13793));
assign g25803 = (g24798&g21024);
assign g26305 = (g24556)|(g24564);
assign g13986 = ((~g10323))|((~g11747));
assign g8870 = ((~II12837));
assign g23837 = (g21160&g10804);
assign g31273 = (g30143&g27779);
assign g20188 = (g5849&g17772);
assign g31194 = (g19128&g29814);
assign g30092 = (g28466)|(g16699);
assign g9657 = ((~g2763));
assign II30901 = ((~g32407));
assign g25590 = (g21694)|(g24160);
assign II27533 = (g21143&g24125&g24126&g24127);
assign g17145 = (g7469&g13249);
assign g14136 = ((~g11571))|((~g8906));
assign g32756 = ((~g31021));
assign g23026 = ((~g20391));
assign g34223 = (g33744&g22876);
assign g16758 = (g5220&g14758);
assign g28167 = ((~g925))|((~g27046));
assign g34277 = ((~II32274));
assign g26811 = ((~g25206));
assign g34724 = (g34702)|(g18152);
assign II23327 = ((~g22647));
assign g7245 = ((~II11896));
assign g21747 = (g3061&g20330);
assign g26631 = ((~g25467));
assign g31851 = ((~g29385));
assign g22990 = (g19555&g19760);
assign g30473 = (g30196)|(g21944);
assign g25584 = (g21670)|(g24154);
assign g29783 = (g28329&g23246);
assign g32248 = (g31616&g30299);
assign g18287 = (g1442&g16449);
assign g19575 = (g15693)|(g13042);
assign g9637 = ((~II13252));
assign g33105 = (g26298&g32138);
assign II31316 = (g29385&g32911&g32912&g32913);
assign g32865 = ((~g31327));
assign g29114 = (g27646)|(g26602);
assign II14713 = ((~g9671))|((~II14712));
assign g31290 = (g29734&g23335);
assign g12840 = ((~g10356));
assign g27336 = (g2675&g26777);
assign g10704 = (g2145&g10200&g2130);
assign g31258 = (g25991)|(g29550);
assign g34373 = (g26292)|(g34138);
assign g21753 = (g3179&g20785);
assign g23111 = ((~g20391));
assign g30304 = (g28255)|(g27259);
assign g34025 = (g33927)|(g18672);
assign g11025 = (g2980)|(g7831);
assign g24351 = (g23774)|(g18807);
assign g33948 = (g32442)|(g33458);
assign g33731 = (g33116&g19520);
assign g20541 = ((~g17821));
assign g32318 = ((~g31596));
assign II31226 = (g29385&g32781&g32782&g32783);
assign g17678 = ((~II18653));
assign g28240 = (g27356&g17239);
assign g24183 = ((~II23393));
assign g30429 = (g29844)|(g21813);
assign g13191 = ((~II15788));
assign g13107 = ((~g10476));
assign g26280 = (g13051&g25248);
assign g34100 = (g33690)|(g33697);
assign g18807 = (g6386&g15656);
assign g8919 = ((~II12896));
assign g33797 = ((~g33306));
endmodule
