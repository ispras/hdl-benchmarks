module s13207_bench(
  blif_clk_net,
  blif_reset_net,
  g43,
  g49,
  g633,
  g634,
  g635,
  g645,
  g647,
  g648,
  g690,
  g694,
  g698,
  g702,
  g722,
  g723,
  g751,
  g752,
  g753,
  g754,
  g755,
  g756,
  g757,
  g781,
  g941,
  g962,
  g1000,
  g1008,
  g1016,
  g1080,
  g1234,
  g1553,
  g1554,
  g206,
  g291,
  g372,
  g453,
  g534,
  g594,
  g785,
  g1006,
  g1015,
  g1017,
  g1246,
  g1724,
  g1783,
  g1798,
  g1804,
  g1810,
  g1817,
  g1824,
  g1829,
  g1870,
  g1871,
  g1894,
  g1911,
  g1944,
  g2662,
  g2844,
  g2888,
  g3077,
  g3096,
  g3130,
  g3159,
  g3191,
  g3829,
  g3859,
  g3860,
  g4267,
  g4316,
  g4370,
  g4371,
  g4372,
  g4373,
  g4655,
  g4657,
  g4660,
  g4661,
  g4663,
  g4664,
  g5143,
  g5164,
  g5571,
  g5669,
  g5678,
  g5682,
  g5684,
  g5687,
  g5729,
  g6207,
  g6212,
  g6223,
  g6236,
  g6269,
  g6425,
  g6648,
  g6653,
  g6675,
  g6849,
  g6850,
  g6895,
  g6909,
  g7048,
  g7063,
  g7103,
  g7283,
  g7284,
  g7285,
  g7286,
  g7287,
  g7288,
  g7289,
  g7290,
  g7291,
  g7292,
  g7293,
  g7294,
  g7295,
  g7298,
  g7423,
  g7424,
  g7425,
  g7474,
  g7504,
  g7505,
  g7506,
  g7507,
  g7508,
  g7514,
  g7729,
  g7730,
  g7731,
  g7732,
  g8216,
  g8217,
  g8218,
  g8219,
  g8234,
  g8661,
  g8663,
  g8872,
  g8958,
  g9128,
  g9132,
  g9204,
  g9280,
  g9297,
  g9299,
  g9305,
  g9308,
  g9310,
  g9312,
  g9314,
  g9378);
input blif_clk_net;
input blif_reset_net;
input g43;
input g49;
input g633;
input g634;
input g635;
input g645;
input g647;
input g648;
input g690;
input g694;
input g698;
input g702;
input g722;
input g723;
input g751;
input g752;
input g753;
input g754;
input g755;
input g756;
input g757;
input g781;
input g941;
input g962;
input g1000;
input g1008;
input g1016;
input g1080;
input g1234;
input g1553;
input g1554;
output g206;
output g291;
output g372;
output g453;
output g534;
output g594;
output g785;
output g1006;
output g1015;
output g1017;
output g1246;
output g1724;
output g1783;
output g1798;
output g1804;
output g1810;
output g1817;
output g1824;
output g1829;
output g1870;
output g1871;
output g1894;
output g1911;
output g1944;
output g2662;
output g2844;
output g2888;
output g3077;
output g3096;
output g3130;
output g3159;
output g3191;
output g3829;
output g3859;
output g3860;
output g4267;
output g4316;
output g4370;
output g4371;
output g4372;
output g4373;
output g4655;
output g4657;
output g4660;
output g4661;
output g4663;
output g4664;
output g5143;
output g5164;
output g5571;
output g5669;
output g5678;
output g5682;
output g5684;
output g5687;
output g5729;
output g6207;
output g6212;
output g6223;
output g6236;
output g6269;
output g6425;
output g6648;
output g6653;
output g6675;
output g6849;
output g6850;
output g6895;
output g6909;
output g7048;
output g7063;
output g7103;
output g7283;
output g7284;
output g7285;
output g7286;
output g7287;
output g7288;
output g7289;
output g7290;
output g7291;
output g7292;
output g7293;
output g7294;
output g7295;
output g7298;
output g7423;
output g7424;
output g7425;
output g7474;
output g7504;
output g7505;
output g7506;
output g7507;
output g7508;
output g7514;
output g7729;
output g7730;
output g7731;
output g7732;
output g8216;
output g8217;
output g8218;
output g8219;
output g8234;
output g8661;
output g8663;
output g8872;
output g8958;
output g9128;
output g9132;
output g9204;
output g9280;
output g9297;
output g9299;
output g9305;
output g9308;
output g9310;
output g9312;
output g9314;
output g9378;
reg g31;
reg g30;
reg g29;
reg g28;
reg g27;
reg g26;
reg g25;
reg g24;
reg g23;
reg g22;
reg g12;
reg g11;
reg g9;
reg g8;
reg g7;
reg g6;
reg g5;
reg g4;
reg g2;
reg g3;
reg g48;
reg g21;
reg g10;
reg g1;
reg g47;
reg g46;
reg g45;
reg g44;
reg g42;
reg g41;
reg g37;
reg g32;
reg g1207;
reg g1211;
reg g1214;
reg g1217;
reg g1220;
reg g1223;
reg g1224;
reg g1225;
reg g1226;
reg g1227;
reg g1228;
reg g1229;
reg g1230;
reg g1240;
reg g1236;
reg g1231;
reg g1244;
reg g1245;
reg g1243;
reg g1272;
reg g1276;
reg g1280;
reg g1284;
reg g1288;
reg g1292;
reg g1300;
reg g1296;
reg g1253;
reg g1308;
reg g1309;
reg g1310;
reg g1311;
reg g1312;
reg g1304;
reg g1307;
reg g1330;
reg g1333;
reg g1336;
reg g1339;
reg g1342;
reg g1345;
reg g1348;
reg g1351;
reg g1354;
reg g1357;
reg g1360;
reg g1190;
reg g1191;
reg g1192;
reg g1193;
reg g1194;
reg g1195;
reg g1196;
reg g1197;
reg g1198;
reg g1199;
reg g1200;
reg g1201;
reg g1202;
reg g1203;
reg g1204;
reg g1205;
reg g1206;
reg g1252;
reg g1250;
reg g1251;
reg g1247;
reg g1254;
reg g1266;
reg g1260;
reg g1257;
reg g1263;
reg g1267;
reg g1268;
reg g1269;
reg g1271;
reg g1270;
reg g172;
reg g1313;
reg g1317;
reg g1318;
reg g1319;
reg g1320;
reg g1321;
reg g1322;
reg g1323;
reg g1324;
reg g1325;
reg g1326;
reg g1327;
reg g1328;
reg g13;
reg g1329;
reg g20;
reg g1366;
reg g1364;
reg g1370;
reg g1368;
reg g1374;
reg g1372;
reg g1375;
reg g1365;
reg g1363;
reg g1369;
reg g1367;
reg g1373;
reg g1371;
reg g1389;
reg g1379;
reg g1377;
reg g1383;
reg g1381;
reg g1387;
reg g1385;
reg g1388;
reg g1378;
reg g1376;
reg g1382;
reg g1380;
reg g1386;
reg g1384;
reg g1390;
reg g1391;
reg g1392;
reg g1393;
reg g1395;
reg g1394;
reg g1396;
reg g1398;
reg g1397;
reg g1399;
reg g1401;
reg g1400;
reg g1402;
reg g1403;
reg g1404;
reg g16;
reg g1189;
reg g1412;
reg g1415;
reg g1409;
reg g1416;
reg g1421;
reg g1405;
reg g1408;
reg g1429;
reg g1428;
reg g1431;
reg g1430;
reg g1424;
reg g1524;
reg g1513;
reg g1486;
reg g1481;
reg g1489;
reg g1494;
reg g1499;
reg g1504;
reg g1509;
reg g1514;
reg g1519;
reg g1462;
reg g1467;
reg g1472;
reg g1477;
reg g727;
reg g1532;
reg g1528;
reg g1537;
reg g1541;
reg g1545;
reg g1549;
reg g1435;
reg g1439;
reg g1432;
reg g1443;
reg g33;
reg g38;
reg g1461;
reg g1444;
reg g1450;
reg g1454;
reg g1459;
reg g1460;
reg g979;
reg g966;
reg g969;
reg g963;
reg g970;
reg g971;
reg g972;
reg g973;
reg g976;
reg g984;
reg g985;
reg g990;
reg g995;
reg g1004;
reg g1005;
reg g998;
reg g999;
reg g1007;
reg g1012;
reg g1014;
reg g1013;
reg g1029;
reg g1018;
reg g1021;
reg g1025;
reg g1033;
reg g1034;
reg g1030;
reg g1081;
reg g1156;
reg g1157;
reg g1159;
reg g1158;
reg g1084;
reg g1146;
reg g1147;
reg g1148;
reg g1087;
reg g1098;
reg g1102;
reg g1106;
reg g1110;
reg g1114;
reg g1118;
reg g1122;
reg g1126;
reg g1142;
reg g1173;
reg g1170;
reg g1167;
reg g1166;
reg g1077;
reg g1153;
reg g1154;
reg g1155;
reg g1185;
reg g1097;
reg g1092;
reg g1130;
reg g1134;
reg g1138;
reg g1149;
reg g1037;
reg g1041;
reg g1045;
reg g1049;
reg g1053;
reg g1057;
reg g1061;
reg g1065;
reg g1069;
reg g1073;
reg g1163;
reg g1160;
reg g1182;
reg g1186;
reg g1179;
reg g1176;
reg g68;
reg g71;
reg g74;
reg g77;
reg g80;
reg g83;
reg g86;
reg g52;
reg g55;
reg g62;
reg g58;
reg g65;
reg g199;
reg g200;
reg g201;
reg g190;
reg g195;
reg g196;
reg g179;
reg g186;
reg g187;
reg g180;
reg g205;
reg g202;
reg g181;
reg g210;
reg g207;
reg g182;
reg g146;
reg g173;
reg g150;
reg g174;
reg g154;
reg g158;
reg g162;
reg g168;
reg g183;
reg g184;
reg g185;
reg g92;
reg g89;
reg g93;
reg g94;
reg g95;
reg g98;
reg g99;
reg g100;
reg g103;
reg g104;
reg g105;
reg g108;
reg g109;
reg g110;
reg g113;
reg g114;
reg g117;
reg g118;
reg g121;
reg g122;
reg g125;
reg g126;
reg g129;
reg g130;
reg g133;
reg g134;
reg g137;
reg g138;
reg g141;
reg g142;
reg g145;
reg g287;
reg g290;
reg g255;
reg g258;
reg g261;
reg g264;
reg g267;
reg g270;
reg g281;
reg g284;
reg g211;
reg g216;
reg g212;
reg g219;
reg g213;
reg g222;
reg g214;
reg g225;
reg g215;
reg g228;
reg g231;
reg g237;
reg g232;
reg g240;
reg g233;
reg g243;
reg g234;
reg g246;
reg g235;
reg g249;
reg g236;
reg g252;
reg g273;
reg g275;
reg g274;
reg g278;
reg g368;
reg g371;
reg g336;
reg g339;
reg g342;
reg g345;
reg g348;
reg g351;
reg g362;
reg g365;
reg g292;
reg g297;
reg g293;
reg g300;
reg g294;
reg g303;
reg g295;
reg g306;
reg g296;
reg g309;
reg g312;
reg g318;
reg g313;
reg g321;
reg g314;
reg g324;
reg g315;
reg g327;
reg g316;
reg g330;
reg g317;
reg g333;
reg g354;
reg g356;
reg g355;
reg g359;
reg g449;
reg g452;
reg g417;
reg g420;
reg g423;
reg g426;
reg g429;
reg g432;
reg g443;
reg g446;
reg g373;
reg g378;
reg g374;
reg g381;
reg g375;
reg g384;
reg g376;
reg g387;
reg g377;
reg g390;
reg g393;
reg g399;
reg g394;
reg g402;
reg g395;
reg g405;
reg g396;
reg g408;
reg g397;
reg g411;
reg g398;
reg g414;
reg g435;
reg g437;
reg g436;
reg g440;
reg g530;
reg g533;
reg g498;
reg g501;
reg g504;
reg g507;
reg g510;
reg g513;
reg g524;
reg g527;
reg g454;
reg g459;
reg g455;
reg g462;
reg g456;
reg g465;
reg g457;
reg g468;
reg g458;
reg g471;
reg g474;
reg g480;
reg g475;
reg g483;
reg g476;
reg g486;
reg g477;
reg g489;
reg g478;
reg g492;
reg g479;
reg g495;
reg g516;
reg g518;
reg g517;
reg g521;
reg g535;
reg g536;
reg g539;
reg g540;
reg g543;
reg g544;
reg g547;
reg g550;
reg g553;
reg g556;
reg g557;
reg g566;
reg g567;
reg g579;
reg g580;
reg g583;
reg g584;
reg g587;
reg g560;
reg g563;
reg g570;
reg g588;
reg g591;
reg g573;
reg g576;
reg g595;
reg g596;
reg g597;
reg g598;
reg g599;
reg g600;
reg g601;
reg g602;
reg g603;
reg g604;
reg g605;
reg g606;
reg g607;
reg g608;
reg g609;
reg g610;
reg g611;
reg g612;
reg g613;
reg g614;
reg g615;
reg g616;
reg g617;
reg g618;
reg g619;
reg g620;
reg g621;
reg g622;
reg g623;
reg g624;
reg g625;
reg g626;
reg g627;
reg g628;
reg g629;
reg g630;
reg g631;
reg g632;
reg g646;
reg g652;
reg g661;
reg g665;
reg g669;
reg g673;
reg g677;
reg g681;
reg g685;
reg g706;
reg g710;
reg g714;
reg g718;
reg g734;
reg g730;
reg g689;
reg g758;
reg g759;
reg g760;
reg g761;
reg g762;
reg g763;
reg g764;
reg g765;
reg g766;
reg g767;
reg g768;
reg g769;
reg g770;
reg g771;
reg g772;
reg g773;
reg g774;
reg g795;
reg g792;
reg g782;
reg g799;
reg g803;
reg g806;
reg g809;
reg g812;
reg g775;
reg g778;
reg g815;
reg g819;
reg g822;
reg g825;
reg g828;
reg g786;
reg g789;
reg g955;
reg g959;
reg g945;
reg g948;
reg g949;
reg g950;
reg g951;
reg g952;
reg g953;
reg g954;
reg g943;
reg g936;
reg g940;
reg g942;
reg g944;
reg g855;
reg g859;
reg g863;
reg g831;
reg g834;
reg g837;
reg g840;
reg g843;
reg g846;
reg g849;
reg g852;
reg g890;
reg g878;
reg g926;
reg g875;
reg g866;
reg g929;
reg g933;
reg g871;
reg g874;
reg g891;
reg g896;
reg g901;
reg g906;
reg g911;
reg g916;
reg g921;
reg g883;
reg g887;
reg g888;
reg g889;
reg g741;
reg g746;
wire g3491;
wire II11158;
wire g8902;
wire g6579;
wire II13463;
wire II10924;
wire II6524;
wire g7168;
wire g3892;
wire II15147;
wire II15405;
wire g3783;
wire g4111;
wire g3603;
wire g2887;
wire g6136;
wire II14712;
wire g7555;
wire g3885;
wire g6034;
wire g7658;
wire II14260;
wire II12226;
wire II16103;
wire g8278;
wire g6426;
wire g9023;
wire g8946;
wire g8932;
wire II8486;
wire II10315;
wire g9338;
wire g4960;
wire g6045;
wire g3221;
wire g7246;
wire g2039;
wire g3313;
wire g7100;
wire g5845;
wire g7440;
wire II5689;
wire g7600;
wire II15871;
wire g8801;
wire g7756;
wire g5119;
wire g5099;
wire g2282;
wire g5607;
wire II10039;
wire g4097;
wire g7252;
wire II10856;
wire g3864;
wire g7115;
wire g8862;
wire II8052;
wire g8904;
wire g8641;
wire II9929;
wire II13622;
wire g8938;
wire g8976;
wire g5589;
wire gbuf10;
wire g9034;
wire g4276;
wire g1794;
wire g2651;
wire g8941;
wire II12041;
wire g7521;
wire g6358;
wire II10250;
wire II10587;
wire II11069;
wire g9184;
wire II11440;
wire g2403;
wire II11150;
wire II16161;
wire g1736;
wire g8717;
wire g6890;
wire gbuf3;
wire II16040;
wire II15187;
wire II11894;
wire g3922;
wire II9804;
wire g1822;
wire g6847;
wire g6818;
wire g5491;
wire g8645;
wire g4883;
wire II7616;
wire g6015;
wire g7136;
wire g5726;
wire g4150;
wire g2177;
wire g3029;
wire g8885;
wire II11971;
wire g6827;
wire II12088;
wire g5673;
wire II15720;
wire II13509;
wire g6743;
wire g6101;
wire II5432;
wire g5302;
wire g6279;
wire II12250;
wire g6605;
wire II6615;
wire g9109;
wire II12678;
wire II15882;
wire g4919;
wire II14489;
wire g6594;
wire g8817;
wire II15519;
wire II6540;
wire g6155;
wire g1976;
wire II9597;
wire g8704;
wire II13544;
wire II15539;
wire II7053;
wire II11164;
wire II11773;
wire g2709;
wire g6333;
wire II13858;
wire g2703;
wire g9276;
wire g2315;
wire g6108;
wire g6389;
wire II15099;
wire g6142;
wire g4899;
wire II11171;
wire g7264;
wire II12406;
wire g5363;
wire g3848;
wire g6364;
wire II9250;
wire g1567;
wire g1784;
wire g3931;
wire g5185;
wire g3129;
wire g9347;
wire g8384;
wire g4413;
wire g4127;
wire g8804;
wire g1813;
wire g1958;
wire II11018;
wire g2780;
wire g7297;
wire II11758;
wire II8901;
wire g5258;
wire g2941;
wire II6009;
wire g3990;
wire g2727;
wire II12259;
wire II15711;
wire g8669;
wire g2340;
wire g3851;
wire g3936;
wire g4925;
wire g7132;
wire g3013;
wire II10001;
wire g9360;
wire g6822;
wire g2767;
wire g7238;
wire g2673;
wire II15803;
wire g9011;
wire g8678;
wire II13413;
wire g4699;
wire g5512;
wire g4028;
wire g4168;
wire g6488;
wire g4930;
wire g4720;
wire g7588;
wire g6150;
wire II14288;
wire II6643;
wire II15324;
wire g7537;
wire g6662;
wire g5489;
wire g3869;
wire II11028;
wire g2627;
wire II15211;
wire II8333;
wire g1698;
wire g2328;
wire g5305;
wire II13281;
wire II9341;
wire g9357;
wire II13962;
wire II13341;
wire g8461;
wire II11086;
wire g2157;
wire g2954;
wire g3973;
wire II7950;
wire II8460;
wire II8394;
wire II14996;
wire g5971;
wire g2014;
wire II12085;
wire g9271;
wire g4702;
wire g4031;
wire g3778;
wire g4120;
wire g8982;
wire II9630;
wire g6900;
wire II14148;
wire g5074;
wire g6147;
wire g8257;
wire g7681;
wire g5565;
wire g1675;
wire g1728;
wire II13882;
wire g6371;
wire g2246;
wire II16126;
wire g4777;
wire II9992;
wire g8227;
wire II5920;
wire g5525;
wire g6654;
wire g4249;
wire g3991;
wire g3465;
wire g9374;
wire g4637;
wire g9211;
wire g7364;
wire II8613;
wire g6174;
wire g2265;
wire II7487;
wire g1887;
wire g4285;
wire g7316;
wire II12319;
wire g2614;
wire II15042;
wire g6961;
wire g7339;
wire g5210;
wire II9422;
wire II13054;
wire g6225;
wire g3051;
wire g9207;
wire g5820;
wire g7747;
wire g1960;
wire II15702;
wire g1637;
wire g5142;
wire g5268;
wire g7713;
wire g6416;
wire g5038;
wire II8935;
wire II11714;
wire II8546;
wire II14315;
wire II10485;
wire II7655;
wire II9169;
wire II10801;
wire g4812;
wire g8293;
wire II14178;
wire g7449;
wire II7341;
wire II12193;
wire g7024;
wire II9639;
wire g6176;
wire g8668;
wire II10834;
wire g9200;
wire II16033;
wire g2683;
wire II5667;
wire g8915;
wire II16020;
wire g7787;
wire g3398;
wire II11034;
wire g3515;
wire g5244;
wire g7143;
wire II13261;
wire II12550;
wire II13653;
wire g6884;
wire II15962;
wire g6049;
wire g7147;
wire g1916;
wire II5997;
wire g7593;
wire g7676;
wire g4732;
wire g9111;
wire g5894;
wire II6112;
wire II15863;
wire g7105;
wire g2334;
wire II13695;
wire II13786;
wire g1949;
wire g7734;
wire g7495;
wire g2724;
wire II15292;
wire g7761;
wire g1752;
wire II11212;
wire g6252;
wire II13831;
wire g4435;
wire II10421;
wire g8891;
wire II5933;
wire g5766;
wire g4283;
wire g4824;
wire II8046;
wire II8558;
wire g7018;
wire II8186;
wire g7049;
wire g8640;
wire II5883;
wire g6569;
wire II11948;
wire g5624;
wire II7198;
wire g8844;
wire II7036;
wire II6872;
wire g8837;
wire g7137;
wire g8664;
wire g5160;
wire II6454;
wire g4219;
wire g4790;
wire g6977;
wire g3517;
wire II11149;
wire II15052;
wire II10265;
wire g7180;
wire II14427;
wire g7307;
wire g6804;
wire gbuf35;
wire g2253;
wire g3082;
wire g3874;
wire II9672;
wire II11832;
wire g6899;
wire II9938;
wire g6465;
wire II10292;
wire II11622;
wire II5696;
wire II8757;
wire g1583;
wire II7520;
wire g4678;
wire g7709;
wire g3631;
wire g5582;
wire II15334;
wire II8040;
wire II15085;
wire II12478;
wire II13484;
wire g3871;
wire II8904;
wire II14747;
wire II14094;
wire g2373;
wire g6064;
wire g2918;
wire g2959;
wire g9060;
wire g4873;
wire g7330;
wire g3945;
wire g4596;
wire g4613;
wire g6771;
wire g8131;
wire g7610;
wire g8781;
wire g3549;
wire g6553;
wire g4048;
wire II12989;
wire II7554;
wire g8854;
wire g6601;
wire g5460;
wire g5712;
wire g4840;
wire g2647;
wire II11431;
wire II9310;
wire II6416;
wire g8152;
wire g5138;
wire II9396;
wire g3721;
wire g5747;
wire II14974;
wire II11317;
wire g8335;
wire II5401;
wire g7268;
wire II6996;
wire g9366;
wire g6308;
wire II6075;
wire g3560;
wire g9158;
wire II12832;
wire g9048;
wire II8240;
wire II8998;
wire g3903;
wire g2354;
wire II10702;
wire g5829;
wire g8962;
wire II13018;
wire II15729;
wire II8823;
wire g7070;
wire II13004;
wire g3076;
wire g5395;
wire II13589;
wire II8436;
wire g5689;
wire II7172;
wire g8455;
wire g7191;
wire II8504;
wire g4957;
wire g7492;
wire II12968;
wire II12535;
wire g2832;
wire II13669;
wire g6402;
wire II13906;
wire II15030;
wire gbuf23;
wire g3189;
wire II13822;
wire g4054;
wire g2964;
wire II13296;
wire g1581;
wire gbuf76;
wire g8768;
wire II12141;
wire g7193;
wire g5984;
wire g7358;
wire g4044;
wire g7112;
wire g7695;
wire g6094;
wire II5512;
wire g4574;
wire II10460;
wire g9124;
wire II14807;
wire g6924;
wire g1842;
wire g6070;
wire gbuf72;
wire II11958;
wire II10919;
wire II10373;
wire II6940;
wire g7603;
wire g4094;
wire II14816;
wire II14695;
wire g7095;
wire g1820;
wire g1924;
wire II15340;
wire g6005;
wire II13106;
wire g6541;
wire g3611;
wire g6995;
wire g3950;
wire g8091;
wire II7797;
wire g5693;
wire g4611;
wire g2222;
wire g2891;
wire g4356;
wire g9095;
wire II6758;
wire g8620;
wire g6970;
wire g3160;
wire II5989;
wire II10430;
wire g4307;
wire g8883;
wire II11880;
wire g4343;
wire II7567;
wire II9001;
wire g8362;
wire II10491;
wire g3833;
wire g2926;
wire II9512;
wire II10223;
wire g5514;
wire g8069;
wire g7227;
wire II6500;
wire II8472;
wire II10457;
wire g2274;
wire II6178;
wire II9162;
wire g2548;
wire g5026;
wire II6936;
wire II10154;
wire g4395;
wire g8846;
wire g2213;
wire g4134;
wire g5547;
wire g5087;
wire II8449;
wire II8225;
wire g6356;
wire II9071;
wire II10207;
wire g6309;
wire II13193;
wire II11574;
wire II7087;
wire g9029;
wire g7791;
wire g6395;
wire II9382;
wire g3984;
wire II15818;
wire II15950;
wire g1833;
wire II9152;
wire II12659;
wire g4115;
wire II13213;
wire g7531;
wire g5477;
wire II11870;
wire g3095;
wire g5062;
wire g8788;
wire II7332;
wire g7185;
wire g5149;
wire g7538;
wire II9333;
wire g5540;
wire g3920;
wire g4650;
wire g3911;
wire g3760;
wire II11132;
wire g8681;
wire g2239;
wire g6186;
wire II8165;
wire g1772;
wire II13499;
wire g3767;
wire g8727;
wire II9987;
wire g7022;
wire g9214;
wire g4179;
wire g5197;
wire g5217;
wire II7374;
wire g6373;
wire II8034;
wire g6865;
wire II13588;
wire g4601;
wire II7460;
wire g7678;
wire II9624;
wire gbuf30;
wire g6952;
wire II10791;
wire II11323;
wire g9385;
wire g8682;
wire g1750;
wire g4669;
wire g9252;
wire II10519;
wire g3901;
wire g3429;
wire g6588;
wire g1848;
wire II12652;
wire g7810;
wire II14439;
wire g7056;
wire g6524;
wire g6196;
wire II6949;
wire II6894;
wire g6941;
wire II7179;
wire II10512;
wire g4409;
wire g5412;
wire II6234;
wire II9747;
wire g9052;
wire II7970;
wire II10973;
wire II8643;
wire g6685;
wire g9160;
wire g1827;
wire g2306;
wire II15533;
wire g8072;
wire g4527;
wire g4145;
wire g6392;
wire II15251;
wire g5231;
wire II6064;
wire II15275;
wire g2134;
wire g4309;
wire g2509;
wire II7365;
wire g5782;
wire g8985;
wire II6376;
wire g7157;
wire g1854;
wire g4237;
wire g7937;
wire g2392;
wire II10992;
wire g4667;
wire II5646;
wire II13147;
wire g8953;
wire II13173;
wire II6124;
wire g5069;
wire g8978;
wire g4226;
wire g8926;
wire gbuf55;
wire II6118;
wire g2043;
wire II12526;
wire g4411;
wire g6322;
wire II10439;
wire g3238;
wire g7702;
wire g5234;
wire g9233;
wire II12131;
wire II8847;
wire II13682;
wire g2554;
wire g8341;
wire g6698;
wire II12870;
wire g7752;
wire II15020;
wire g4196;
wire II11004;
wire II9126;
wire II11254;
wire g4457;
wire g9351;
wire II6849;
wire II11596;
wire g5574;
wire g7156;
wire II16049;
wire II10678;
wire g5202;
wire g2295;
wire II12508;
wire g6799;
wire g5835;
wire II8045;
wire g5526;
wire g6435;
wire g7487;
wire g7544;
wire II8400;
wire II14193;
wire II11633;
wire g8710;
wire g7129;
wire g8081;
wire II16058;
wire g1759;
wire II13869;
wire g3080;
wire II10190;
wire g5048;
wire g4513;
wire II9493;
wire g7726;
wire II13631;
wire g6858;
wire II5521;
wire g6302;
wire g4312;
wire g4388;
wire g6706;
wire g4075;
wire II8127;
wire gbuf15;
wire g6511;
wire g2625;
wire II7964;
wire g5178;
wire g5125;
wire II13060;
wire II8763;
wire g6754;
wire g7320;
wire g5228;
wire g6660;
wire g3579;
wire II14231;
wire II9606;
wire g6472;
wire II5368;
wire II9576;
wire g6764;
wire II11449;
wire II12466;
wire g8690;
wire g2379;
wire g5537;
wire g1664;
wire II6148;
wire II9663;
wire II7278;
wire gbuf63;
wire g6421;
wire g6314;
wire II8392;
wire II6522;
wire g6368;
wire II5562;
wire II6209;
wire II11841;
wire g5120;
wire g9092;
wire II7888;
wire g1769;
wire g4482;
wire g8238;
wire II8140;
wire g6458;
wire g4901;
wire II15073;
wire g7836;
wire g4559;
wire II15625;
wire II9582;
wire g8327;
wire g4067;
wire II7505;
wire II14124;
wire g9202;
wire g2992;
wire g8994;
wire g9298;
wire II11503;
wire II7629;
wire II7241;
wire g5436;
wire g4503;
wire II12463;
wire II7712;
wire g2969;
wire II11887;
wire II10525;
wire g3650;
wire II15283;
wire II5789;
wire II12649;
wire gbuf5;
wire g7066;
wire II6425;
wire g6841;
wire g6871;
wire g9100;
wire II11858;
wire II10384;
wire g4035;
wire II12124;
wire g6617;
wire g5787;
wire g7161;
wire g2999;
wire II15160;
wire g2936;
wire g6167;
wire g3985;
wire g4095;
wire g1683;
wire g6736;
wire g4181;
wire II10980;
wire g8288;
wire g7002;
wire II5868;
wire g1785;
wire II15660;
wire g2907;
wire g4662;
wire g9369;
wire g6255;
wire g9316;
wire g6792;
wire II14246;
wire g2290;
wire II8796;
wire II14952;
wire g5170;
wire g9087;
wire g6768;
wire g6217;
wire g5053;
wire g5847;
wire II6826;
wire II15759;
wire g9177;
wire g8065;
wire g2137;
wire g6227;
wire II5757;
wire g6838;
wire gbuf43;
wire II10198;
wire II8495;
wire II14330;
wire II13228;
wire g5209;
wire g9267;
wire II10940;
wire II12415;
wire g6162;
wire II16084;
wire g8638;
wire g1852;
wire II14759;
wire g4917;
wire II12888;
wire II7899;
wire g1235;
wire II11224;
wire g5763;
wire g5041;
wire g6780;
wire g8877;
wire g4804;
wire g8301;
wire II14772;
wire II13719;
wire g1574;
wire g4545;
wire II11425;
wire g6628;
wire g4564;
wire II8005;
wire g9135;
wire g7174;
wire g4056;
wire II9823;
wire g6739;
wire g5313;
wire g4328;
wire g4606;
wire II7938;
wire g3828;
wire g6112;
wire g4332;
wire g2982;
wire g3884;
wire g7107;
wire g6362;
wire g5051;
wire g8382;
wire II9531;
wire g5183;
wire II15880;
wire g7500;
wire g6140;
wire g3757;
wire II15974;
wire g8830;
wire g9355;
wire g9027;
wire g5987;
wire II9242;
wire g9274;
wire II13335;
wire II7186;
wire g7236;
wire g3562;
wire g6157;
wire II5380;
wire g6335;
wire g2671;
wire II7311;
wire II8966;
wire g8702;
wire g6294;
wire g4062;
wire g6250;
wire II9103;
wire g4129;
wire g8815;
wire g2551;
wire g3084;
wire g2052;
wire II5365;
wire II11368;
wire g8653;
wire g2051;
wire g4116;
wire g3805;
wire g2923;
wire g1556;
wire g6050;
wire g7326;
wire g6745;
wire II5621;
wire g9001;
wire g5151;
wire g2943;
wire g2375;
wire II8573;
wire g9307;
wire g3933;
wire g8018;
wire g3728;
wire g4786;
wire II13595;
wire g8944;
wire II7436;
wire II11533;
wire g8909;
wire g8698;
wire II14754;
wire g5028;
wire II14184;
wire g5443;
wire II11751;
wire II5801;
wire g7021;
wire II9954;
wire g6731;
wire II13267;
wire g6406;
wire g1831;
wire g5147;
wire g6298;
wire g5552;
wire II5718;
wire g3680;
wire g8676;
wire g2769;
wire II14980;
wire g8735;
wire II8014;
wire g2913;
wire II9099;
wire g7535;
wire II7082;
wire II8739;
wire II10073;
wire II13350;
wire g5105;
wire II7070;
wire II10475;
wire g5668;
wire g7528;
wire g8856;
wire II15062;
wire g8281;
wire g6593;
wire II6784;
wire g3915;
wire II15836;
wire g2230;
wire g1721;
wire II15669;
wire g6230;
wire g6975;
wire g6259;
wire II11551;
wire II7101;
wire II8745;
wire g7711;
wire g6340;
wire II11272;
wire II14801;
wire g4540;
wire g8603;
wire g2692;
wire II6217;
wire g5563;
wire II15230;
wire g2332;
wire g4608;
wire g9013;
wire g5632;
wire g7586;
wire g4560;
wire II10900;
wire g8709;
wire g6902;
wire g9311;
wire g6263;
wire II15833;
wire II7305;
wire g5706;
wire g8652;
wire g7777;
wire g4933;
wire II6160;
wire II9555;
wire g7576;
wire g8647;
wire II14828;
wire II10783;
wire II14413;
wire g2632;
wire g7549;
wire g6966;
wire g6351;
wire g9036;
wire II11293;
wire g7442;
wire g7754;
wire g8657;
wire g6074;
wire II8805;
wire g9054;
wire g7113;
wire g5519;
wire g3862;
wire g2366;
wire g2787;
wire g3841;
wire g7634;
wire II9041;
wire g6992;
wire g4871;
wire g8936;
wire g2989;
wire II15040;
wire II6305;
wire g5227;
wire II6800;
wire II8079;
wire g7552;
wire II8373;
wire g695;
wire II15738;
wire g6505;
wire g8643;
wire g4493;
wire II12996;
wire g6229;
wire II15889;
wire g5439;
wire II14039;
wire II15571;
wire g9309;
wire g6032;
wire g2106;
wire II8913;
wire II9654;
wire g7178;
wire g5609;
wire II13701;
wire g4549;
wire g5246;
wire g4524;
wire II11764;
wire g4274;
wire g5117;
wire II14403;
wire II15705;
wire g8753;
wire II10538;
wire II11689;
wire g5101;
wire II5528;
wire II13903;
wire g6013;
wire II12481;
wire g7000;
wire II14457;
wire g1918;
wire II11311;
wire II15019;
wire g8315;
wire g2653;
wire g8959;
wire g7616;
wire g2956;
wire g6796;
wire g4385;
wire g3867;
wire g3893;
wire II8895;
wire II9177;
wire g6276;
wire g1578;
wire g9174;
wire g6475;
wire g6118;
wire g6829;
wire II13897;
wire II5559;
wire g7163;
wire g5058;
wire g7428;
wire g6124;
wire g6382;
wire II15726;
wire II8665;
wire II15054;
wire g6379;
wire g4553;
wire II15784;
wire g2774;
wire g7244;
wire g5140;
wire g4700;
wire g6741;
wire g9186;
wire g2881;
wire g2533;
wire g6483;
wire g3633;
wire g6931;
wire II8114;
wire g9223;
wire II6291;
wire g2645;
wire g1838;
wire II12643;
wire II11178;
wire g3876;
wire g3498;
wire g1011;
wire g7745;
wire g8563;
wire g5256;
wire II9369;
wire g5165;
wire g6189;
wire II12295;
wire g8806;
wire II7495;
wire II12205;
wire g3735;
wire II9884;
wire g2971;
wire g2497;
wire g8720;
wire II6183;
wire g6704;
wire II13457;
wire g4914;
wire g5584;
wire g1803;
wire g8619;
wire II9484;
wire II12854;
wire g6133;
wire g1796;
wire II15915;
wire II8865;
wire g4598;
wire g4681;
wire g6439;
wire II15083;
wire g9345;
wire II13997;
wire g6213;
wire g7234;
wire g4819;
wire II5505;
wire g3341;
wire g2826;
wire II9528;
wire g3488;
wire II13912;
wire II7680;
wire II7064;
wire g6844;
wire g6893;
wire II12924;
wire II10835;
wire II14480;
wire g2934;
wire g5745;
wire II11978;
wire II9005;
wire g7254;
wire g3513;
wire g7305;
wire g2939;
wire g8967;
wire g7512;
wire g9038;
wire g8631;
wire II9347;
wire II15291;
wire g6057;
wire II11156;
wire g6571;
wire g1682;
wire g7654;
wire g2208;
wire g6447;
wire g8511;
wire II11043;
wire g1872;
wire g7110;
wire II7609;
wire g2916;
wire g6486;
wire II10347;
wire g9062;
wire II7788;
wire II9907;
wire g5076;
wire II7545;
wire g3644;
wire g3929;
wire II5954;
wire II15672;
wire g8310;
wire II12304;
wire g8795;
wire g3857;
wire g8960;
wire g8338;
wire g1569;
wire g3837;
wire II14245;
wire II11835;
wire g3905;
wire II7973;
wire g8333;
wire II12373;
wire g738;
wire g8623;
wire g2293;
wire g8276;
wire II15657;
wire g8295;
wire g4353;
wire g6824;
wire II7211;
wire II7752;
wire g6870;
wire II7611;
wire II6998;
wire II6323;
wire II7838;
wire g9199;
wire II11803;
wire II7618;
wire II5676;
wire g8581;
wire II6924;
wire II11143;
wire g4511;
wire II12268;
wire g7315;
wire II7443;
wire g9081;
wire g5112;
wire g2020;
wire g7497;
wire g7683;
wire g3971;
wire II11422;
wire II9549;
wire g7480;
wire g5813;
wire g7275;
wire II15856;
wire g8924;
wire g4265;
wire g9021;
wire g5670;
wire g4920;
wire II12337;
wire g5594;
wire g4287;
wire g2323;
wire g6172;
wire II11236;
wire g5603;
wire g8662;
wire g7140;
wire g4399;
wire g6650;
wire II13432;
wire g6621;
wire g3542;
wire II7268;
wire g5738;
wire g2834;
wire g8260;
wire g7344;
wire II11522;
wire g6243;
wire g4690;
wire II11842;
wire II6033;
wire g2995;
wire g6468;
wire g7141;
wire II10874;
wire g8997;
wire II7697;
wire g9376;
wire II13773;
wire g6673;
wire II13687;
wire II9021;
wire g8233;
wire g6968;
wire g7362;
wire II11961;
wire II14933;
wire g2845;
wire g7145;
wire II7098;
wire II7944;
wire II7575;
wire g2751;
wire g8930;
wire g4895;
wire g9008;
wire II7804;
wire g2721;
wire g2505;
wire g9320;
wire g7047;
wire II9209;
wire II15765;
wire II11129;
wire g9194;
wire g6886;
wire II10009;
wire g5434;
wire g4795;
wire II13035;
wire g2272;
wire g9327;
wire II6286;
wire II11096;
wire g2460;
wire g6345;
wire II15530;
wire g2229;
wire II8826;
wire g1677;
wire II8877;
wire g8282;
wire g1744;
wire g6659;
wire g5260;
wire II7485;
wire g2866;
wire g2484;
wire g6329;
wire g5628;
wire g7139;
wire g4501;
wire II8581;
wire II14172;
wire II7856;
wire II7814;
wire g6287;
wire g6859;
wire g3496;
wire g1896;
wire g7598;
wire g5822;
wire g4825;
wire g4622;
wire g4422;
wire g7591;
wire II7925;
wire II10758;
wire II13704;
wire g9259;
wire g6863;
wire II10561;
wire g4706;
wire II12881;
wire II14436;
wire II9360;
wire II5616;
wire II14106;
wire g3091;
wire g4584;
wire g3540;
wire g4065;
wire II13344;
wire II14657;
wire g4239;
wire g5757;
wire g5475;
wire g8041;
wire g3769;
wire g7079;
wire II12939;
wire g4630;
wire II13493;
wire g5545;
wire II8327;
wire g5956;
wire g5199;
wire g6623;
wire g6184;
wire II13628;
wire II7540;
wire g8765;
wire g5780;
wire g7456;
wire g2359;
wire II13140;
wire g4365;
wire g6681;
wire g5568;
wire g4228;
wire g6776;
wire II8205;
wire g4491;
wire II14831;
wire g3913;
wire g8296;
wire g6179;
wire g7522;
wire g8542;
wire II11386;
wire II5577;
wire g6692;
wire g5219;
wire g1923;
wire g6056;
wire g5344;
wire g2900;
wire g6687;
wire g9387;
wire II13365;
wire g8074;
wire g7769;
wire II12834;
wire g6380;
wire II10976;
wire g4354;
wire g8111;
wire g7159;
wire II14022;
wire II14397;
wire g7101;
wire gbuf50;
wire g8666;
wire II12561;
wire g5521;
wire g7038;
wire II6012;
wire g8983;
wire II15423;
wire g4379;
wire II6368;
wire g5488;
wire II7538;
wire g9069;
wire g4617;
wire g5734;
wire g6190;
wire g4123;
wire II12167;
wire g4797;
wire g4724;
wire II14822;
wire g2525;
wire g2242;
wire II15072;
wire g5714;
wire g5060;
wire g5824;
wire g8225;
wire II11920;
wire g4187;
wire g6657;
wire II8889;
wire II5377;
wire II13403;
wire g7351;
wire II14789;
wire II7389;
wire II16154;
wire g8313;
wire II6232;
wire g5744;
wire II11251;
wire g9148;
wire g6645;
wire g6984;
wire g4624;
wire g5576;
wire II12181;
wire g3187;
wire g6023;
wire II12592;
wire g4001;
wire g9264;
wire g8722;
wire g6400;
wire g4305;
wire g7418;
wire II7356;
wire g7081;
wire II5359;
wire II15007;
wire II7371;
wire II10608;
wire g3993;
wire g6316;
wire g7211;
wire g6635;
wire II10256;
wire II10888;
wire g6957;
wire II9561;
wire g7044;
wire g6555;
wire II12187;
wire II8537;
wire g9121;
wire g4838;
wire g4146;
wire g6926;
wire II6457;
wire g7097;
wire g6280;
wire II6437;
wire g5698;
wire g4420;
wire g3533;
wire II10469;
wire g6877;
wire II15897;
wire g3957;
wire g8742;
wire g7601;
wire gbuf74;
wire g9331;
wire g4543;
wire g2824;
wire II7640;
wire g7065;
wire g3287;
wire g9042;
wire g2385;
wire II12699;
wire II13131;
wire II13478;
wire II14780;
wire II9460;
wire g9318;
wire g4393;
wire g4433;
wire g8325;
wire g7983;
wire g2262;
wire II11110;
wire g5417;
wire II15510;
wire g6366;
wire g4132;
wire g4643;
wire g7625;
wire II12145;
wire II11461;
wire g6567;
wire g3613;
wire g7779;
wire II11929;
wire II8357;
wire II7931;
wire II11945;
wire g6076;
wire II5945;
wire g4959;
wire II7599;
wire g8996;
wire g4341;
wire II7290;
wire g8303;
wire II8412;
wire g7221;
wire II16180;
wire II14009;
wire II6956;
wire g8898;
wire g5768;
wire II9047;
wire g6562;
wire II8244;
wire II13397;
wire g7743;
wire II10933;
wire g5067;
wire II10770;
wire g3555;
wire g7313;
wire II12779;
wire II15010;
wire II14064;
wire II10062;
wire II14133;
wire g4310;
wire II12918;
wire g4740;
wire II13583;
wire g8067;
wire g5785;
wire II15285;
wire II8431;
wire g1704;
wire g6215;
wire II9837;
wire g2313;
wire II6752;
wire g2664;
wire g2901;
wire II11815;
wire g8443;
wire g5223;
wire g4334;
wire g5806;
wire g9107;
wire II8736;
wire g8875;
wire g6160;
wire g6914;
wire II6795;
wire g5621;
wire g3577;
wire II5565;
wire g8798;
wire g1934;
wire II15243;
wire g4579;
wire II14042;
wire g3659;
wire g3523;
wire II11851;
wire II15616;
wire g7119;
wire II9692;
wire II15110;
wire g4108;
wire gbuf33;
wire II14378;
wire II14076;
wire g7547;
wire II10684;
wire g5704;
wire g7632;
wire g7176;
wire g1782;
wire g5467;
wire g3970;
wire g1825;
wire g6910;
wire g9114;
wire g8778;
wire g6437;
wire g3771;
wire II6054;
wire II11556;
wire II6834;
wire g6809;
wire g4058;
wire g6716;
wire II10196;
wire II8811;
wire g8524;
wire gbuf17;
wire II8006;
wire g8820;
wire II15732;
wire g8784;
wire g1562;
wire II11874;
wire g4537;
wire g724;
wire II8856;
wire II8781;
wire g7082;
wire g5653;
wire g8803;
wire g4453;
wire g5287;
wire g8275;
wire g9133;
wire II9446;
wire g6457;
wire II12364;
wire g1576;
wire g3965;
wire g2790;
wire II15645;
wire g4802;
wire g4258;
wire II9964;
wire II9826;
wire g8712;
wire II15199;
wire II5842;
wire g7054;
wire g8758;
wire g2267;
wire g3093;
wire g3233;
wire II7864;
wire II13764;
wire g4489;
wire g5618;
wire g2539;
wire g2183;
wire g7826;
wire g3505;
wire II12597;
wire g9288;
wire g4639;
wire g2532;
wire g2921;
wire g8671;
wire II13879;
wire g2898;
wire g2962;
wire g6152;
wire II7174;
wire II14142;
wire g8613;
wire II8299;
wire II15507;
wire g3679;
wire II11233;
wire II8945;
wire g5206;
wire II10277;
wire g6708;
wire II8089;
wire g5200;
wire II9564;
wire II12214;
wire II12079;
wire g9235;
wire g2810;
wire II12138;
wire II12445;
wire g5084;
wire g7750;
wire II7149;
wire g3835;
wire II12451;
wire g4572;
wire g2345;
wire g658;
wire g4784;
wire g4685;
wire g7904;
wire II9502;
wire II6428;
wire g5232;
wire II10899;
wire II14276;
wire g6938;
wire g4072;
wire g8860;
wire g5192;
wire II8551;
wire g6789;
wire II12289;
wire g8176;
wire g8738;
wire II11347;
wire g5840;
wire g7724;
wire II10406;
wire II11218;
wire g4567;
wire II11821;
wire II15631;
wire II13656;
wire g7329;
wire g3002;
wire g8755;
wire g5127;
wire g1980;
wire II14169;
wire g6766;
wire g6490;
wire g4923;
wire II8932;
wire g6752;
wire II13326;
wire g4881;
wire II7216;
wire II10463;
wire II11242;
wire g8605;
wire g5441;
wire II12891;
wire g9073;
wire g1857;
wire g5158;
wire II9910;
wire g9212;
wire II14049;
wire II13807;
wire II14302;
wire g5078;
wire II9222;
wire II8502;
wire g3982;
wire II12397;
wire II7009;
wire II9979;
wire g2495;
wire g8719;
wire g5397;
wire g7208;
wire g3960;
wire g6797;
wire II10286;
wire g4466;
wire II8607;
wire g4295;
wire II15265;
wire II14959;
wire g5172;
wire g2562;
wire g6238;
wire g8629;
wire g3260;
wire g2477;
wire g6790;
wire g9090;
wire g3359;
wire II11470;
wire II8511;
wire g7783;
wire g4737;
wire II11967;
wire II14151;
wire II14127;
wire II14496;
wire g6713;
wire g9302;
wire g2206;
wire g7686;
wire g6807;
wire gbuf65;
wire g4021;
wire II15811;
wire g5672;
wire g3338;
wire g9348;
wire g9197;
wire g5605;
wire g8289;
wire g3085;
wire g8659;
wire II9271;
wire II8157;
wire II15429;
wire g6646;
wire II11392;
wire II12379;
wire II6045;
wire II10436;
wire g2479;
wire II10359;
wire g7470;
wire g7596;
wire II11122;
wire g5520;
wire g6888;
wire II12541;
wire II13834;
wire g3995;
wire g5071;
wire II13305;
wire II8243;
wire II14668;
wire g2215;
wire II14190;
wire g2256;
wire g7751;
wire g6695;
wire g7560;
wire g7772;
wire II13640;
wire gbuf26;
wire II11838;
wire g6461;
wire II5831;
wire II6021;
wire II11848;
wire g5033;
wire II15641;
wire II12190;
wire g8421;
wire g3999;
wire II5936;
wire II11704;
wire II14416;
wire II6431;
wire II14257;
wire g4304;
wire II7262;
wire g3097;
wire g8612;
wire g7543;
wire II15912;
wire g8290;
wire g6707;
wire g4793;
wire g2161;
wire g8636;
wire II9366;
wire II13876;
wire g4656;
wire g3643;
wire g7215;
wire II13454;
wire g2556;
wire g6469;
wire g5708;
wire g3895;
wire II15898;
wire g6639;
wire g2331;
wire g8655;
wire II13234;
wire II11014;
wire g5224;
wire g6775;
wire g6170;
wire g8859;
wire II13063;
wire g6116;
wire g6153;
wire II6974;
wire g8377;
wire II11506;
wire g5560;
wire II6419;
wire II12051;
wire g8774;
wire g5080;
wire g5723;
wire II8538;
wire g5031;
wire g7792;
wire g8737;
wire g5599;
wire g9300;
wire II10442;
wire g1671;
wire g4263;
wire II5923;
wire II7893;
wire II12552;
wire g8966;
wire g6324;
wire g4426;
wire g4912;
wire g2131;
wire g3882;
wire II8583;
wire g7540;
wire g7259;
wire g4081;
wire g6973;
wire g3907;
wire II11942;
wire II14311;
wire gbuf47;
wire II9235;
wire II15252;
wire g4538;
wire II11809;
wire II6248;
wire g4809;
wire II13527;
wire g5094;
wire g4788;
wire II10952;
wire g8583;
wire g7184;
wire II6233;
wire g5241;
wire g4514;
wire g2377;
wire II7995;
wire g5825;
wire g9192;
wire g1913;
wire II11172;
wire II5507;
wire II9195;
wire II12722;
wire g5139;
wire II8288;
wire II11936;
wire II9827;
wire II14460;
wire II12334;
wire g4592;
wire II5407;
wire g3812;
wire g7303;
wire g9115;
wire g9025;
wire g4250;
wire g8626;
wire g2644;
wire g6802;
wire g4521;
wire II11796;
wire g8173;
wire II12499;
wire II7326;
wire g1667;
wire g8336;
wire g8331;
wire g6038;
wire II10125;
wire g6288;
wire II5356;
wire g3545;
wire g7014;
wire g5017;
wire II14199;
wire II7558;
wire II13716;
wire II8134;
wire g655;
wire II7118;
wire II13258;
wire II12669;
wire g3753;
wire g6624;
wire g6315;
wire g5639;
wire g3949;
wire g3940;
wire g5014;
wire g5793;
wire g8236;
wire II12223;
wire II12582;
wire g5550;
wire g5482;
wire II15678;
wire g7438;
wire g3230;
wire II12951;
wire g5107;
wire g5569;
wire g7090;
wire II7811;
wire g7334;
wire g3942;
wire II15681;
wire II16006;
wire g3967;
wire g4038;
wire g6019;
wire II13277;
wire g8359;
wire g2825;
wire II10295;
wire g3520;
wire II6814;
wire II9081;
wire II5410;
wire g8852;
wire g6582;
wire g3978;
wire g4133;
wire g6432;
wire g4739;
wire g3918;
wire g6904;
wire g4878;
wire g5917;
wire g3822;
wire g4113;
wire II7204;
wire g8147;
wire g9127;
wire II5984;
wire g2634;
wire g6964;
wire g9031;
wire II15017;
wire II7919;
wire g3898;
wire g8439;
wire II10579;
wire g5116;
wire g2623;
wire II14531;
wire g5132;
wire II6451;
wire II14970;
wire g9188;
wire g1670;
wire II13215;
wire II11627;
wire II6805;
wire g3787;
wire II13416;
wire g2890;
wire II8024;
wire II6134;
wire g7239;
wire II14485;
wire g8089;
wire g4050;
wire II5605;
wire g3790;
wire g6875;
wire II9076;
wire g8514;
wire g3855;
wire II14121;
wire g8265;
wire II7085;
wire II9181;
wire II14766;
wire g7574;
wire g3955;
wire II10528;
wire g6341;
wire II15849;
wire g5299;
wire II15193;
wire II12244;
wire g9140;
wire II13017;
wire g9321;
wire g4893;
wire g2922;
wire II14091;
wire II11206;
wire II10247;
wire II5548;
wire g5677;
wire II8253;
wire g8284;
wire g6274;
wire g7232;
wire g9131;
wire g6728;
wire II7908;
wire g9171;
wire II15391;
wire g3889;
wire g5100;
wire g1975;
wire II6220;
wire g5182;
wire g7692;
wire g5731;
wire g6816;
wire II12017;
wire II11066;
wire g2487;
wire II9069;
wire II11686;
wire II11094;
wire g2746;
wire g8812;
wire g9065;
wire II11428;
wire g4934;
wire g5613;
wire g2344;
wire g8649;
wire II11800;
wire g2270;
wire g8729;
wire g4490;
wire g5841;
wire II13728;
wire g2677;
wire g5029;
wire II13435;
wire g7118;
wire II11666;
wire g2940;
wire g4686;
wire II9788;
wire g3865;
wire g8979;
wire g7411;
wire II7181;
wire g3849;
wire II13320;
wire g6832;
wire II7588;
wire g6498;
wire g7551;
wire g4272;
wire II14985;
wire g2362;
wire II12400;
wire II12032;
wire II5709;
wire g5772;
wire g2706;
wire II14709;
wire g7519;
wire II5682;
wire II15264;
wire II13854;
wire II12179;
wire II6087;
wire g5189;
wire g6476;
wire g9218;
wire II15190;
wire g8730;
wire g4041;
wire g3938;
wire g3802;
wire g5818;
wire II15648;
wire g1563;
wire II12062;
wire g5286;
wire g7780;
wire II5568;
wire g4820;
wire II11790;
wire g8878;
wire II12412;
wire II6676;
wire II9525;
wire II6229;
wire g8868;
wire II11410;
wire g1800;
wire II13918;
wire II12430;
wire g6296;
wire g1757;
wire II12409;
wire g7009;
wire II15178;
wire g9244;
wire II10479;
wire II6036;
wire g2784;
wire g3878;
wire g1694;
wire II9171;
wire g5719;
wire g6846;
wire II9965;
wire g8329;
wire g2945;
wire g6137;
wire g8708;
wire g6347;
wire g6003;
wire II5715;
wire g2311;
wire II11677;
wire II6839;
wire g6412;
wire g6385;
wire g3705;
wire g6414;
wire g8934;
wire g5314;
wire g6332;
wire II8237;
wire II6905;
wire g4887;
wire II15824;
wire g3844;
wire g7581;
wire II10011;
wire g8866;
wire g5155;
wire II7422;
wire g7532;
wire g4713;
wire g7443;
wire g2911;
wire g5145;
wire g4707;
wire II10018;
wire g5811;
wire g7510;
wire g7189;
wire g8908;
wire g4410;
wire g6145;
wire g7584;
wire g3935;
wire g7966;
wire II13676;
wire g4465;
wire g6122;
wire g8014;
wire g3723;
wire g3358;
wire II12577;
wire g8881;
wire II9947;
wire II7167;
wire g5163;
wire II10617;
wire II16107;
wire g5779;
wire g2324;
wire g8274;
wire g8267;
wire g8692;
wire II7438;
wire II11011;
wire g8297;
wire g7631;
wire II8150;
wire g2665;
wire g6733;
wire g6758;
wire g3011;
wire g7767;
wire II7953;
wire g2316;
wire II5392;
wire II10739;
wire g9015;
wire g6025;
wire g2006;
wire g8832;
wire II13749;
wire II6646;
wire g1868;
wire g8839;
wire g8697;
wire g8150;
wire g9057;
wire II15546;
wire g7256;
wire II16043;
wire g4245;
wire II8121;
wire II13410;
wire g7502;
wire II9840;
wire g8714;
wire g6306;
wire g2872;
wire II5948;
wire g6709;
wire g4015;
wire g2506;
wire g2350;
wire II15553;
wire g6580;
wire II8315;
wire II6629;
wire g4013;
wire II8078;
wire g9237;
wire g2209;
wire g7172;
wire II9845;
wire g7741;
wire II10400;
wire g7722;
wire g6474;
wire II16119;
wire g5578;
wire II5911;
wire g5064;
wire II14374;
wire g5174;
wire II9515;
wire g4905;
wire II7778;
wire g4906;
wire g6826;
wire II6578;
wire II12869;
wire g8895;
wire g6370;
wire g1802;
wire g3780;
wire II11389;
wire g6318;
wire g7832;
wire g7690;
wire g7697;
wire g6683;
wire g4463;
wire g6337;
wire II14643;
wire II5852;
wire g4101;
wire g4298;
wire II6877;
wire g8635;
wire g4541;
wire g8828;
wire g1793;
wire g6912;
wire g5121;
wire g6515;
wire II12894;
wire g7710;
wire g7050;
wire g2498;
wire g5839;
wire II8709;
wire II7498;
wire g4003;
wire g8180;
wire II7044;
wire g8379;
wire g5643;
wire II14015;
wire g3048;
wire II13635;
wire g6854;
wire II12340;
wire g8694;
wire g8272;
wire g4928;
wire g5238;
wire II15152;
wire g9055;
wire g6724;
wire II15385;
wire II15924;
wire g5592;
wire g3988;
wire II12111;
wire II11021;
wire g5832;
wire g4785;
wire II15501;
wire g1877;
wire g6927;
wire g2996;
wire g7121;
wire g5751;
wire g4632;
wire g7125;
wire g6787;
wire II8132;
wire II8547;
wire g8761;
wire g7033;
wire gbuf67;
wire g3677;
wire g4172;
wire II15041;
wire g8911;
wire g7150;
wire II11278;
wire g4746;
wire II15276;
wire II8853;
wire g2903;
wire g9088;
wire gbuf11;
wire g4486;
wire II11184;
wire g1565;
wire g5735;
wire g6407;
wire g2467;
wire g8060;
wire g7361;
wire g7177;
wire g1742;
wire II14118;
wire g6166;
wire g7265;
wire II11353;
wire II8011;
wire II8490;
wire II7568;
wire II9496;
wire II9636;
wire g2517;
wire g5118;
wire g4568;
wire II14046;
wire g6906;
wire g4270;
wire g4185;
wire g2877;
wire g2510;
wire g6783;
wire g8873;
wire g2238;
wire g4025;
wire g6188;
wire g6834;
wire II11221;
wire g3657;
wire II12826;
wire II10503;
wire gbuf31;
wire g5020;
wire g7353;
wire II13003;
wire g3511;
wire g2804;
wire g8794;
wire g7198;
wire g5205;
wire g4582;
wire g2291;
wire g6105;
wire g4577;
wire g5427;
wire II13039;
wire g6058;
wire II10743;
wire g9282;
wire g4086;
wire g8786;
wire g2234;
wire g4476;
wire g9105;
wire g1680;
wire II15308;
wire g7920;
wire II6422;
wire g1707;
wire II15985;
wire II6048;
wire II10424;
wire II15492;
wire g7346;
wire g2269;
wire g6448;
wire II8883;
wire II10387;
wire g2896;
wire g642;
wire II16176;
wire II11729;
wire II8733;
wire g7459;
wire g9083;
wire g5523;
wire II5649;
wire g8322;
wire II13930;
wire g8745;
wire II13924;
wire g5742;
wire g7036;
wire g5027;
wire g2557;
wire g4590;
wire g5716;
wire II5599;
wire g5705;
wire g5808;
wire g3850;
wire g5091;
wire g8810;
wire II8196;
wire g6573;
wire g3500;
wire g8809;
wire II13075;
wire II9505;
wire g5800;
wire II11269;
wire II12286;
wire II8784;
wire II14479;
wire g7719;
wire g6919;
wire II14031;
wire g1809;
wire g6430;
wire g1689;
wire II11230;
wire II6143;
wire g4255;
wire II12696;
wire II8817;
wire II5963;
wire g1789;
wire II6317;
wire II10172;
wire II15684;
wire II14798;
wire II15583;
wire g4627;
wire g2584;
wire II6274;
wire II6843;
wire g7599;
wire g8305;
wire g7607;
wire g5683;
wire g1815;
wire II11137;
wire II10597;
wire g6503;
wire g1585;
wire g6041;
wire g1580;
wire g2286;
wire II10393;
wire II6115;
wire II11725;
wire g8406;
wire g6793;
wire g7087;
wire g6949;
wire g1919;
wire g7120;
wire II11320;
wire g1760;
wire g3557;
wire g6637;
wire g4605;
wire II12912;
wire II8360;
wire II6930;
wire g4831;
wire g8740;
wire g4070;
wire II13428;
wire II11380;
wire II9935;
wire g6381;
wire g6282;
wire g3531;
wire g2957;
wire g7006;
wire II12325;
wire g4589;
wire II11998;
wire g4090;
wire g8092;
wire g7099;
wire g6641;
wire g2383;
wire II10236;
wire g2520;
wire g6920;
wire g6658;
wire g6051;
wire II8680;
wire g8827;
wire g5213;
wire II7368;
wire g6932;
wire II6170;
wire g7349;
wire g9075;
wire g5567;
wire II12247;
wire g8843;
wire II7511;
wire g6565;
wire II6741;
wire g8980;
wire II11864;
wire g4383;
wire g2365;
wire g8723;
wire II5619;
wire g9165;
wire g4718;
wire II9476;
wire g5458;
wire g5267;
wire g7276;
wire II7602;
wire II7157;
wire g7776;
wire g6264;
wire II13317;
wire II10377;
wire g5686;
wire g3285;
wire g7206;
wire g2979;
wire g2100;
wire g8763;
wire II13395;
wire II7592;
wire g4522;
wire g7337;
wire II8986;
wire g5558;
wire g6861;
wire g6204;
wire g4571;
wire g6971;
wire g6894;
wire g8318;
wire II13599;
wire g6868;
wire II10987;
wire g5221;
wire g6377;
wire g6939;
wire g8222;
wire g4614;
wire II15478;
wire II10143;
wire g8606;
wire II14181;
wire g9045;
wire g4654;
wire II5763;
wire g3527;
wire g8441;
wire g8544;
wire gbuf51;
wire g6177;
wire II5692;
wire II15696;
wire g4138;
wire g6688;
wire g6497;
wire II9600;
wire g9146;
wire II7377;
wire g6131;
wire g4555;
wire II12806;
wire II14837;
wire g6097;
wire g7527;
wire g4131;
wire II5975;
wire gbuf8;
wire II12511;
wire II11109;
wire II6163;
wire g4192;
wire II8351;
wire II15229;
wire g3124;
wire g4106;
wire g2543;
wire II9767;
wire II15101;
wire g4352;
wire II6258;
wire g5970;
wire II13009;
wire II15504;
wire II13134;
wire g7308;
wire g8857;
wire II14433;
wire g6193;
wire g5473;
wire g4391;
wire g6062;
wire g2970;
wire II7755;
wire II6065;
wire g3916;
wire g4646;
wire g1776;
wire g2641;
wire gbuf27;
wire g7310;
wire g4119;
wire g6955;
wire II7296;
wire g3071;
wire g6092;
wire g6945;
wire II5812;
wire g8974;
wire g6590;
wire g8989;
wire g3632;
wire II15172;
wire II11116;
wire g4005;
wire g3692;
wire gbuf20;
wire g5257;
wire g7217;
wire II14804;
wire II13801;
wire II15516;
wire g4455;
wire II10454;
wire II6499;
wire II10071;
wire g3083;
wire gbuf42;
wire II8636;
wire II12382;
wire g4692;
wire II12180;
wire g5150;
wire II12460;
wire II11778;
wire g8776;
wire g1970;
wire g5008;
wire g9139;
wire II14969;
wire II11718;
wire g6069;
wire II13743;
wire II9057;
wire g9370;
wire II5374;
wire II7734;
wire g6773;
wire II16145;
wire II16138;
wire g6908;
wire II15909;
wire g7301;
wire g2092;
wire g7829;
wire II15051;
wire II12958;
wire II10780;
wire g9063;
wire II11362;
wire g7993;
wire II10412;
wire II13813;
wire II8939;
wire II8063;
wire II14318;
wire g6525;
wire II15536;
wire g5005;
wire II9645;
wire II15762;
wire II13605;
wire g8759;
wire g7068;
wire g5082;
wire g6445;
wire II14904;
wire g4437;
wire g6936;
wire g3846;
wire g4688;
wire g6249;
wire II7532;
wire g6756;
wire g6996;
wire g1834;
wire g8029;
wire g6632;
wire g3648;
wire II7891;
wire II6018;
wire g2642;
wire g6169;
wire g5626;
wire g2349;
wire g3462;
wire II11787;
wire II10605;
wire g4741;
wire g5016;
wire II10649;
wire II14728;
wire g5243;
wire g6630;
wire II8898;
wire g6700;
wire g5403;
wire g6897;
wire II11497;
wire g7182;
wire g5438;
wire g9323;
wire II15262;
wire g5137;
wire g6237;
wire g4474;
wire II15181;
wire II10761;
wire II5422;
wire g5749;
wire II11047;
wire II11515;
wire II8868;
wire II7978;
wire II6203;
wire g3653;
wire g8791;
wire II10313;
wire g8271;
wire g3518;
wire g4036;
wire II10954;
wire II9443;
wire g8700;
wire II13425;
wire g2470;
wire g3853;
wire g5480;
wire g2649;
wire g8334;
wire g6603;
wire g6800;
wire g6087;
wire g6216;
wire II16168;
wire II7010;
wire g7332;
wire g5161;
wire g2985;
wire g5096;
wire II7800;
wire g8964;
wire II13332;
wire g4694;
wire g6036;
wire g5114;
wire g7092;
wire g4594;
wire II6072;
wire g3947;
wire II12813;
wire II10818;
wire g6917;
wire g2621;
wire II7551;
wire g9102;
wire g639;
wire g3547;
wire g3909;
wire g8585;
wire g6674;
wire II13787;
wire II14219;
wire g2264;
wire g8154;
wire g8971;
wire II5847;
wire II13559;
wire II15495;
wire g4424;
wire II11482;
wire II5861;
wire g1686;
wire II11078;
wire II10361;
wire g7436;
wire g1582;
wire g8819;
wire g6947;
wire g4868;
wire II6695;
wire II9009;
wire II10962;
wire II10000;
wire II12472;
wire g3605;
wire g2395;
wire g7688;
wire II10789;
wire g9304;
wire g2346;
wire g2210;
wire g8231;
wire g3567;
wire g5538;
wire g1603;
wire g9205;
wire g7594;
wire g8928;
wire II11124;
wire gbuf62;
wire g5362;
wire g4023;
wire II9534;
wire g8913;
wire II12544;
wire II11479;
wire II9025;
wire g9372;
wire II7069;
wire g2284;
wire g6143;
wire g3588;
wire g6303;
wire II8401;
wire II6151;
wire II8568;
wire II14157;
wire g1819;
wire II6326;
wire g6696;
wire g8906;
wire II15610;
wire II9609;
wire g6367;
wire g8299;
wire g6652;
wire g6291;
wire g5587;
wire g6008;
wire II10369;
wire II12307;
wire g4444;
wire II8245;
wire g3900;
wire g6760;
wire II16026;
wire II15842;
wire g3997;
wire II16132;
wire g5168;
wire g7770;
wire g7493;
wire II8180;
wire g6596;
wire g5843;
wire g5580;
wire g4580;
wire II10488;
wire II9850;
wire II15113;
wire g2821;
wire g7790;
wire g5648;
wire II13311;
wire II15595;
wire g8752;
wire II15817;
wire g1673;
wire g2880;
wire g6855;
wire g9067;
wire g4269;
wire g7130;
wire g1897;
wire II8841;
wire II10592;
wire II12424;
wire g6467;
wire g2862;
wire g6677;
wire g7476;
wire g6010;
wire g5597;
wire II14687;
wire g4389;
wire g4748;
wire g3641;
wire II14473;
wire g4302;
wire g4735;
wire g4078;
wire g4280;
wire II12632;
wire II10448;
wire II13666;
wire II6917;
wire II12256;
wire g1639;
wire g9003;
wire g6881;
wire g5615;
wire II12316;
wire II13164;
wire g7736;
wire g7479;
wire II12564;
wire g4909;
wire g5590;
wire g9005;
wire g8178;
wire II10614;
wire g5056;
wire g9190;
wire g4791;
wire g5827;
wire g6387;
wire II13752;
wire g4528;
wire II6471;
wire II11245;
wire II15298;
wire g7765;
wire g2326;
wire II7429;
wire II9963;
wire g6452;
wire g1805;
wire g8706;
wire g9178;
wire g6410;
wire g8732;
wire g6095;
wire g8016;
wire g7703;
wire II15589;
wire g6661;
wire g6267;
wire g7582;
wire g4408;
wire g4099;
wire g5284;
wire g4673;
wire II6538;
wire g2502;
wire II11747;
wire II14758;
wire g8691;
wire g4142;
wire g1770;
wire g5790;
wire g5180;
wire II8152;
wire II10946;
wire II5419;
wire g1864;
wire g4125;
wire II5386;
wire II13506;
wire g3808;
wire II5795;
wire g4885;
wire II12672;
wire g6722;
wire g9333;
wire g5187;
wire II8108;
wire II12993;
wire II9980;
wire g8864;
wire g5784;
wire g1739;
wire g1779;
wire g9358;
wire g8220;
wire g7530;
wire g5730;
wire g8386;
wire g4367;
wire II6680;
wire g6735;
wire g6353;
wire g6983;
wire g9017;
wire g1781;
wire g2782;
wire II12717;
wire II15021;
wire II11404;
wire II9095;
wire g7016;
wire II8057;
wire g7524;
wire g2947;
wire II8642;
wire g8155;
wire gbuf57;
wire II8588;
wire g9162;
wire II6006;
wire II15239;
wire g7187;
wire g6120;
wire gbuf1;
wire g8269;
wire II14282;
wire II7922;
wire g9258;
wire II8659;
wire II11615;
wire g4313;
wire g3587;
wire g7445;
wire g4963;
wire II10565;
wire g2952;
wire g5795;
wire g7034;
wire g1866;
wire II9166;
wire g9010;
wire II15717;
wire g9368;
wire g4705;
wire g5701;
wire II13725;
wire g5484;
wire g9019;
wire II6774;
wire II12575;
wire g3937;
wire II6663;
wire g4711;
wire II13255;
wire II14743;
wire g2628;
wire g8739;
wire II9145;
wire g8888;
wire g7273;
wire g2869;
wire II8020;
wire II10558;
wire II11549;
wire g4105;
wire II14055;
wire II10472;
wire g1879;
wire g3226;
wire II15776;
wire g7225;
wire II9573;
wire g3574;
wire II14381;
wire g4841;
wire g4154;
wire II10541;
wire II12496;
wire g2240;
wire II15044;
wire g4814;
wire g7545;
wire g6149;
wire II15498;
wire II12053;
wire g8311;
wire g7134;
wire g3316;
wire II8164;
wire II15753;
wire g7248;
wire II9277;
wire II7564;
wire II13837;
wire II11951;
wire g2636;
wire g7558;
wire g1646;
wire g7758;
wire II6733;
wire g8463;
wire g1715;
wire g6273;
wire g6814;
wire g2639;
wire g5739;
wire g8948;
wire II7635;
wire II9774;
wire II9148;
wire g1952;
wire g8675;
wire g691;
wire II9183;
wire g7557;
wire g3953;
wire g7280;
wire II6764;
wire g3746;
wire g7261;
wire g4296;
wire g4231;
wire II10046;
wire g2699;
wire g6339;
wire g1812;
wire II14298;
wire II10166;
wire II7875;
wire g3222;
wire II11419;
wire g8464;
wire g6278;
wire II8536;
wire g6103;
wire g4781;
wire g4696;
wire g5019;
wire g6343;
wire II9946;
wire II6443;
wire g2828;
wire g2963;
wire II7548;
wire g8263;
wire g9047;
wire g4167;
wire gbuf6;
wire g3888;
wire g3976;
wire g6054;
wire II13761;
wire g6607;
wire g4279;
wire g6001;
wire g7694;
wire II12980;
wire g9033;
wire II14474;
wire g8145;
wire g9126;
wire II11900;
wire g4937;
wire g3832;
wire g8939;
wire g6874;
wire g6254;
wire II6354;
wire II8261;
wire g2660;
wire II15254;
wire II11485;
wire g3924;
wire II10336;
wire II9746;
wire g2360;
wire g6726;
wire g2801;
wire g703;
wire g6570;
wire II7107;
wire II8962;
wire g7413;
wire g4083;
wire II8748;
wire II12753;
wire g2616;
wire g4876;
wire g6071;
wire II5478;
wire II8273;
wire g3863;
wire II10548;
wire g4497;
wire g5089;
wire g7715;
wire g5109;
wire II12760;
wire II14085;
wire g2353;
wire II7473;
wire g5104;
wire II12385;
wire g4807;
wire g7748;
wire g5425;
wire g7406;
wire g3485;
wire gbuf16;
wire g3655;
wire II14079;
wire g7165;
wire g5633;
wire g9103;
wire II6440;
wire II8678;
wire II15379;
wire g9226;
wire II8268;
wire g2965;
wire g2873;
wire g8871;
wire II14267;
wire g4318;
wire g6836;
wire g7448;
wire g4007;
wire g5335;
wire g6769;
wire II10321;
wire g7325;
wire II15791;
wire g1727;
wire II13909;
wire g5453;
wire g9216;
wire g2879;
wire g4376;
wire g3509;
wire II7792;
wire II12280;
wire g9159;
wire II9123;
wire g6164;
wire II10868;
wire II10626;
wire II15628;
wire II11867;
wire g9380;
wire g9208;
wire g6552;
wire g9079;
wire g3830;
wire g1910;
wire II12930;
wire II9325;
wire II10804;
wire g5573;
wire II14960;
wire II11586;
wire g8816;
wire II13126;
wire g1787;
wire g1807;
wire g9137;
wire g5022;
wire g6245;
wire II10415;
wire g4562;
wire g2894;
wire g8320;
wire g8743;
wire g7433;
wire g1687;
wire g6702;
wire g3961;
wire II12265;
wire g4911;
wire II9666;
wire II14130;
wire II12439;
wire g6934;
wire g4253;
wire II10826;
wire II11981;
wire g9070;
wire g5093;
wire g7578;
wire g4201;
wire II7617;
wire g3666;
wire g7258;
wire g4535;
wire g8825;
wire g5802;
wire II8072;
wire g7421;
wire g4665;
wire g2960;
wire g1571;
wire II13447;
wire II12532;
wire II6195;
wire g4088;
wire g8955;
wire II12961;
wire II9612;
wire II7844;
wire g7717;
wire II8218;
wire g9278;
wire g2655;
wire II12394;
wire g3839;
wire II10306;
wire g1666;
wire g9118;
wire II11102;
wire g2794;
wire g6256;
wire II13377;
wire g2236;
wire g5688;
wire II8594;
wire g7127;
wire g1587;
wire II7299;
wire g7123;
wire g4721;
wire g5645;
wire g3590;
wire g8893;
wire g7720;
wire II8989;
wire g5043;
wire g6409;
wire g8482;
wire g6718;
wire g2225;
wire g8258;
wire g4052;
wire g4073;
wire II11338;
wire g2180;
wire g6785;
wire II14109;
wire g4011;
wire g7788;
wire g6211;
wire g9239;
wire II8255;
wire g7738;
wire g5123;
wire g8079;
wire g1849;
wire g3492;
wire g5789;
wire g1856;
wire g6517;
wire II7467;
wire II13042;
wire II10896;
wire g6325;
wire g6046;
wire g8771;
wire g8008;
wire II8393;
wire g6423;
wire g9353;
wire g8633;
wire II9241;
wire g4092;
wire II7148;
wire g7705;
wire g7699;
wire II12274;
wire g4368;
wire g6383;
wire II14061;
wire II10535;
wire II9107;
wire g1795;
wire g4918;
wire g5126;
wire g6781;
wire II14783;
wire gbuf45;
wire gbuf69;
wire II13900;
wire g4891;
wire g9077;
wire gbuf13;
wire II8838;
wire g3602;
wire II12514;
wire II13707;
wire g1938;
wire g7340;
wire g5153;
wire II6750;
wire g5674;
wire g9247;
wire g7366;
wire g3675;
wire g7220;
wire g5679;
wire g6711;
wire g6470;
wire g7059;
wire II10350;
wire g5236;
wire g9059;
wire g7322;
wire g2232;
wire II13685;
wire g7564;
wire II8172;
wire II12022;
wire g7271;
wire g4926;
wire g7155;
wire II11284;
wire g5176;
wire g7727;
wire g5834;
wire II16052;
wire gbuf38;
wire II7454;
wire II5620;
wire II12008;
wire g7319;
wire g8608;
wire g7031;
wire g7152;
wire g4243;
wire g4618;
wire g3712;
wire II6093;
wire g8458;
wire g4198;
wire II15240;
wire g5658;
wire g3078;
wire II13843;
wire g4659;
wire g1909;
wire g8625;
wire II11693;
wire II7882;
wire g4903;
wire g5517;
wire g3764;
wire II13600;
wire II12454;
wire II7561;
wire II13659;
wire g7040;
wire gbuf40;
wire g5073;
wire II13028;
wire II10409;
wire II15887;
wire g2308;
wire g2837;
wire g4652;
wire II9111;
wire g8769;
wire g5753;
wire g6026;
wire g2928;
wire g4642;
wire II13144;
wire II9044;
wire g5549;
wire II13537;
wire g4648;
wire g3525;
wire g6235;
wire II14025;
wire II12232;
wire gbuf29;
wire g3819;
wire II7400;
wire II16183;
wire II11329;
wire g1649;
wire g4728;
wire g3614;
wire II12666;
wire g2480;
wire g5235;
wire g6060;
wire g6990;
wire g4027;
wire g7463;
wire II13888;
wire II8417;
wire g6612;
wire II7702;
wire gbuf22;
wire g4121;
wire g6762;
wire g5469;
wire g1748;
wire g8961;
wire g7267;
wire g4969;
wire II6251;
wire II12903;
wire g6502;
wire g8733;
wire II10907;
wire g4359;
wire g5761;
wire g5542;
wire II11090;
wire g4235;
wire g4350;
wire g6194;
wire II11371;
wire g7355;
wire g2910;
wire II9974;
wire II11824;
wire II15053;
wire II12176;
wire g6372;
wire II7956;
wire g5254;
wire g5760;
wire II11464;
wire g6369;
wire g8886;
wire II12953;
wire g7590;
wire II10403;
wire g5471;
wire g8987;
wire II15273;
wire g6950;
wire g5401;
wire g6978;
wire g3634;
wire g6393;
wire II14166;
wire II6564;
wire II14819;
wire II8871;
wire g6626;
wire g2841;
wire II14187;
wire g7827;
wire g5555;
wire II10328;
wire g2245;
wire II12885;
wire II15947;
wire II6371;
wire II8520;
wire II11177;
wire g9050;
wire g7025;
wire g6953;
wire II10675;
wire g6390;
wire g6586;
wire II11040;
wire II6460;
wire g7106;
wire g8039;
wire g8229;
wire II10687;
wire g6090;
wire II15864;
wire II10093;
wire g7605;
wire g6999;
wire II9372;
wire g7416;
wire g4361;
wire II5897;
wire II11933;
wire g2885;
wire g9195;
wire g7209;
wire g7350;
wire g2381;
wire g2458;
wire II15965;
wire g6220;
wire g4300;
wire g5718;
wire II6333;
wire II7129;
wire g8360;
wire g6428;
wire II12370;
wire g6509;
wire II5966;
wire II7188;
wire g6643;
wire g5470;
wire g7516;
wire g7760;
wire g4629;
wire g4587;
wire g9260;
wire II15003;
wire II7644;
wire g6922;
wire g5494;
wire g8725;
wire g5215;
wire g7028;
wire g6284;
wire II15568;
wire g6805;
wire II9064;
wire II7781;
wire g4033;
wire g1926;
wire II10516;
wire II7150;
wire g2522;
wire II15940;
wire g7774;
wire g8070;
wire II14224;
wire II6776;
wire g5756;
wire g2396;
wire g7061;
wire II5772;
wire g8404;
wire II12708;
wire g6320;
wire g9221;
wire g4620;
wire II9050;
wire g9097;
wire II11473;
wire g6404;
wire II8778;
wire g7196;
wire g8841;
wire g8848;
wire g7491;
wire g9144;
wire g2266;
wire g8684;
wire g8062;
wire II10745;
wire g3739;
wire g7278;
wire II8925;
wire g8991;
wire g4398;
wire g2074;
wire g7838;
wire g6929;
wire II15527;
wire g8457;
wire g6202;
wire gbuf70;
wire g4199;
wire II7380;
wire II6517;
wire II11308;
wire g4182;
wire II15959;
wire g7498;
wire g4069;
wire g2938;
wire II10848;
wire g6129;
wire g1844;
wire g6610;
wire g9335;
wire g4000;
wire g5194;
wire g8687;
wire II8718;
wire g6819;
wire g3062;
wire g8307;
wire II5751;
wire g6360;
wire g9389;
wire g5024;
wire g8968;
wire g7179;
wire II7691;
wire II14771;
wire g5367;
wire g3774;
wire g7089;
wire g3610;
wire II7683;
wire g4355;
wire g3951;
wire g7026;
wire II6959;
wire g4610;
wire g4396;
wire g2386;
wire II10773;
wire g6365;
wire II12128;
wire II8512;
wire II6501;
wire g8995;
wire II6051;
wire II15943;
wire g8090;
wire II8413;
wire II14227;
wire g6542;
wire g7763;
wire g4556;
wire II10849;
wire II15400;
wire g2368;
wire g4311;
wire g6293;
wire g5788;
wire g6577;
wire g5711;
wire II14163;
wire g6201;
wire g5748;
wire g5805;
wire II12771;
wire g5216;
wire g7352;
wire g5025;
wire g6629;
wire II11603;
wire g7314;
wire g5462;
wire II9301;
wire II10224;
wire II14941;
wire g4342;
wire g4623;
wire g5445;
wire II13214;
wire g3761;
wire g7367;
wire II7994;
wire g8361;
wire II12915;
wire g5680;
wire g4835;
wire g7030;
wire II5942;
wire g4197;
wire II16036;
wire II8166;
wire g6419;
wire II7344;
wire g7696;
wire II11305;
wire g8319;
wire g6022;
wire g8892;
wire g8728;
wire g7019;
wire g4009;
wire II14786;
wire g4236;
wire g8403;
wire II6208;
wire II14139;
wire g6222;
wire II13649;
wire II7132;
wire g6872;
wire g2298;
wire g5765;
wire II10690;
wire g3188;
wire gbuf75;
wire g1589;
wire g5874;
wire gbuf71;
wire g2680;
wire II7512;
wire II12355;
wire II6214;
wire g4956;
wire II8437;
wire II5957;
wire g6958;
wire g7604;
wire II8529;
wire g4454;
wire g8780;
wire g4830;
wire II12877;
wire g7192;
wire g6853;
wire g8749;
wire g1828;
wire II11994;
wire g7064;
wire g1925;
wire g4811;
wire g8779;
wire g4091;
wire II10790;
wire g8314;
wire II9769;
wire g5459;
wire g7194;
wire g3548;
wire g4421;
wire g6879;
wire II15205;
wire g6837;
wire g3716;
wire II6259;
wire g5743;
wire II8291;
wire II7651;
wire g8075;
wire II6254;
wire g7626;
wire II15990;
wire II7145;
wire II10694;
wire g6923;
wire II15274;
wire II7688;
wire g6994;
wire g7450;
wire II14291;
wire g3128;
wire II7905;
wire g8385;
wire g6587;
wire g7523;
wire g4649;
wire II15250;
wire II6941;
wire II6970;
wire II13515;
wire g1876;
wire II10993;
wire II10807;
wire g6523;
wire II16158;
wire II7279;
wire II12199;
wire g4068;
wire g4526;
wire g6391;
wire g2925;
wire g7158;
wire g8017;
wire g8757;
wire g4619;
wire II8787;
wire II15956;
wire II12576;
wire g4644;
wire II15475;
wire g9251;
wire g2307;
wire g4114;
wire g6556;
wire g1665;
wire II12900;
wire II14005;
wire g5758;
wire g4634;
wire II6096;
wire g5478;
wire g4839;
wire g6401;
wire g1922;
wire g6951;
wire II7353;
wire II11257;
wire II9381;
wire II14573;
wire II13562;
wire g2833;
wire II9363;
wire g1907;
wire II7584;
wire g6396;
wire g6866;
wire g2547;
wire II15033;
wire II8455;
wire II12238;
wire g6208;
wire g8787;
wire g7677;
wire II8612;
wire g5814;
wire II7086;
wire g8228;
wire g7045;
wire II11275;
wire II6463;
wire II9018;
wire g1853;
wire g3768;
wire g7023;
wire II9986;
wire g9053;
wire II10322;
wire g5141;
wire g1695;
wire g5541;
wire g5198;
wire g3912;
wire II10639;
wire g8680;
wire II13490;
wire II13231;
wire II14100;
wire g9384;
wire g4600;
wire g5269;
wire g6065;
wire g8766;
wire gbuf46;
wire g4030;
wire g9028;
wire g6055;
wire g4266;
wire II15411;
wire g8986;
wire g2915;
wire g7199;
wire g1751;
wire g1847;
wire g3958;
wire II13802;
wire II7423;
wire g4542;
wire g7539;
wire g9317;
wire g4603;
wire II16142;
wire II6509;
wire g6093;
wire g6185;
wire g6753;
wire g9215;
wire II15225;
wire g2876;
wire g1983;
wire II13369;
wire g6459;
wire II13469;
wire II14370;
wire gbuf60;
wire g5047;
wire II14964;
wire g4019;
wire g9072;
wire II9499;
wire II6574;
wire g5916;
wire II13524;
wire g1768;
wire II8190;
wire g7321;
wire g5159;
wire g2389;
wire g5396;
wire II9217;
wire gbuf64;
wire g4071;
wire g4803;
wire g3094;
wire II10329;
wire g8673;
wire g6239;
wire g4333;
wire II13287;
wire g8324;
wire g4294;
wire g9203;
wire g7784;
wire II6868;
wire g7222;
wire II15881;
wire g8750;
wire II6703;
wire g9361;
wire II12170;
wire g3651;
wire II8543;
wire II11165;
wire II13679;
wire II7626;
wire g8340;
wire g9093;
wire II15055;
wire II12871;
wire g2712;
wire g2561;
wire g3779;
wire II15433;
wire II13475;
wire g7680;
wire g4628;
wire g4566;
wire g4029;
wire II10866;
wire g4698;
wire g3834;
wire II8084;
wire II14305;
wire g6857;
wire g7725;
wire II15382;
wire g4880;
wire g6327;
wire g9122;
wire g9136;
wire g5548;
wire II14115;
wire II6275;
wire g2371;
wire II13137;
wire g6434;
wire g4002;
wire II5531;
wire II8983;
wire II8606;
wire II7215;
wire g4012;
wire g8876;
wire g7202;
wire g2393;
wire II12469;
wire II11239;
wire g8456;
wire g8064;
wire II8517;
wire g8741;
wire g9181;
wire g2781;
wire g2961;
wire II11332;
wire II7350;
wire g4387;
wire II9038;
wire g9084;
wire g7169;
wire g5054;
wire g3028;
wire g6301;
wire II15894;
wire g5191;
wire II10906;
wire g6197;
wire II12502;
wire g5203;
wire g4900;
wire g4259;
wire g7328;
wire g8302;
wire II14468;
wire g4076;
wire II6201;
wire g5177;
wire g7055;
wire g9319;
wire II12091;
wire g2930;
wire g3506;
wire II5466;
wire g5040;
wire g8716;
wire II11562;
wire g6226;
wire II11151;
wire g4382;
wire II11080;
wire g6767;
wire II8769;
wire II12927;
wire g4225;
wire g4565;
wire II12933;
wire g7173;
wire g2899;
wire g6420;
wire g7093;
wire II13639;
wire g5312;
wire g7828;
wire g2494;
wire II7937;
wire II6127;
wire g4607;
wire II10965;
wire g4595;
wire g6456;
wire g1575;
wire g3966;
wire II15756;
wire g8068;
wire g6214;
wire II13220;
wire g6444;
wire g6376;
wire g7207;
wire II12217;
wire g7069;
wire g6355;
wire g9261;
wire II8760;
wire II5781;
wire g5797;
wire g2091;
wire II10569;
wire II5978;
wire g6429;
wire g7162;
wire g5085;
wire g5515;
wire g3986;
wire g2343;
wire g4096;
wire g5617;
wire g5435;
wire II7112;
wire II7539;
wire g8823;
wire g8970;
wire II12343;
wire II13460;
wire g3684;
wire g1684;
wire g6937;
wire II11287;
wire II12262;
wire II10981;
wire II13323;
wire g7905;
wire II11263;
wire g5242;
wire g7003;
wire g4585;
wire g4180;
wire g1933;
wire II15666;
wire II9693;
wire g4502;
wire II12388;
wire II12025;
wire II13362;
wire g2816;
wire g6044;
wire II8029;
wire g3658;
wire g5846;
wire II6468;
wire II8264;
wire g6616;
wire g2906;
wire II15690;
wire II13241;
wire II13921;
wire II9182;
wire g5937;
wire g4916;
wire II9953;
wire g4954;
wire II6226;
wire g5492;
wire g6812;
wire g2626;
wire II5706;
wire g5310;
wire g6102;
wire II12687;
wire g4103;
wire g6828;
wire g1821;
wire II5383;
wire g3894;
wire g6848;
wire II8916;
wire g2104;
wire g3840;
wire g6817;
wire g4451;
wire II10028;
wire g2288;
wire g5009;
wire g3923;
wire II14472;
wire II10873;
wire II10092;
wire g8972;
wire g2184;
wire II12487;
wire g3902;
wire II10923;
wire II11203;
wire g5294;
wire II8844;
wire g2631;
wire g3972;
wire g6111;
wire II8177;
wire II12986;
wire g7160;
wire g8646;
wire II7605;
wire II9243;
wire g9354;
wire g4494;
wire II7444;
wire g3743;
wire II13740;
wire g6135;
wire g6543;
wire g3754;
wire g7562;
wire II15522;
wire II11669;
wire g7417;
wire g1711;
wire g7114;
wire g4155;
wire g7243;
wire g3886;
wire g8703;
wire g4961;
wire g7556;
wire II8886;
wire g9035;
wire g9337;
wire II7430;
wire II13672;
wire g8651;
wire g7606;
wire g6427;
wire II7317;
wire g6697;
wire gbuf4;
wire II7452;
wire g4931;
wire II14410;
wire g2663;
wire g3220;
wire II11170;
wire II7302;
wire g3314;
wire g8981;
wire g6896;
wire II8053;
wire g5608;
wire II14739;
wire II8105;
wire g8261;
wire g6350;
wire g8287;
wire g2314;
wire g6614;
wire g8642;
wire g7757;
wire g8975;
wire g7282;
wire g8462;
wire g7251;
wire II11179;
wire g5049;
wire g649;
wire g9363;
wire II5939;
wire II14270;
wire g8863;
wire g1886;
wire g4057;
wire g4898;
wire II6673;
wire g7149;
wire g8940;
wire II11701;
wire II15420;
wire g7589;
wire g6268;
wire II6900;
wire g6663;
wire II10555;
wire II13373;
wire II14349;
wire g4160;
wire g4932;
wire II13737;
wire g6770;
wire g7228;
wire g2595;
wire g8239;
wire g5006;
wire g6125;
wire II14285;
wire II10390;
wire II6571;
wire g5106;
wire g2015;
wire g5610;
wire g9330;
wire g4374;
wire II8742;
wire g8172;
wire II15074;
wire g4703;
wire g7513;
wire II8461;
wire g7536;
wire II14448;
wire g2329;
wire g6738;
wire g8884;
wire II11037;
wire g4778;
wire II10128;
wire II13850;
wire II10243;
wire g6334;
wire g1977;
wire g7108;
wire g3963;
wire g6755;
wire g8383;
wire g3883;
wire II15098;
wire g1555;
wire g6744;
wire g7657;
wire II14825;
wire g8087;
wire g6363;
wire g3649;
wire g1568;
wire g9275;
wire II8772;
wire g9240;
wire II8907;
wire g7135;
wire g6035;
wire II6860;
wire g3891;
wire II10646;
wire II9648;
wire g7595;
wire g2672;
wire II11855;
wire II7648;
wire g5186;
wire g4884;
wire g4126;
wire g6493;
wire g1690;
wire II13713;
wire g8807;
wire g7131;
wire g1959;
wire g8679;
wire g4924;
wire g5253;
wire II10908;
wire II15315;
wire g6310;
wire II12629;
wire II6358;
wire g4414;
wire II15586;
wire g3930;
wire g1797;
wire g7237;
wire II14052;
wire g8736;
wire g6507;
wire II8952;
wire g6156;
wire g6141;
wire II10882;
wire g7230;
wire II7445;
wire II5404;
wire g4597;
wire II7270;
wire g5709;
wire g7615;
wire g2882;
wire g7592;
wire II6166;
wire II13638;
wire II7041;
wire g4047;
wire g9125;
wire g2372;
wire g4733;
wire g6219;
wire g2202;
wire II11964;
wire g4821;
wire II5636;
wire II14492;
wire II6652;
wire g6417;
wire II15550;
wire II7785;
wire II12558;
wire g7148;
wire g8630;
wire g8905;
wire II11740;
wire g6144;
wire II12567;
wire g2953;
wire II11197;
wire g7017;
wire II13794;
wire II6003;
wire g3921;
wire g3568;
wire g9193;
wire g6464;
wire II8326;
wire g6572;
wire g9009;
wire g1655;
wire g8277;
wire g6048;
wire g2223;
wire g4670;
wire g7144;
wire g8294;
wire II15426;
wire II7928;
wire g6883;
wire g1676;
wire II11974;
wire II9233;
wire g8890;
wire II11296;
wire g5035;
wire g6803;
wire II6918;
wire II6104;
wire g5524;
wire g7441;
wire II12301;
wire II5515;
wire II9548;
wire g7714;
wire g8198;
wire g7701;
wire II15111;
wire II9139;
wire II13776;
wire g8925;
wire II8115;
wire II10445;
wire g6962;
wire g7682;
wire g6655;
wire g6710;
wire g3858;
wire g8363;
wire g8834;
wire g8845;
wire II13225;
wire g7008;
wire II9558;
wire g6117;
wire g5166;
wire II12229;
wire II9543;
wire II9136;
wire II13419;
wire g9375;
wire g4636;
wire II7417;
wire g7274;
wire II11525;
wire g7733;
wire II8706;
wire g2734;
wire II10854;
wire g8667;
wire g6175;
wire g1948;
wire g5821;
wire II11781;
wire g6930;
wire g5211;
wire II10274;
wire g3052;
wire II15557;
wire II6911;
wire g9230;
wire II12313;
wire g3192;
wire II5926;
wire II9993;
wire II13487;
wire II7338;
wire II7807;
wire g7317;
wire g9210;
wire II7576;
wire II11383;
wire II7526;
wire II12457;
wire II15862;
wire g5196;
wire g6720;
wire II7466;
wire g8916;
wire g4805;
wire g9157;
wire II11652;
wire g2273;
wire II9344;
wire g8767;
wire g6130;
wire g6554;
wire g5245;
wire II13314;
wire g9382;
wire g2917;
wire II13376;
wire g2038;
wire g7167;
wire g5218;
wire g6915;
wire g6028;
wire II7269;
wire II12220;
wire g3639;
wire g7432;
wire g7331;
wire II12376;
wire II8339;
wire g3946;
wire II8721;
wire g5075;
wire g2933;
wire g6173;
wire g7111;
wire g7357;
wire g4093;
wire g7188;
wire II11912;
wire gbuf2;
wire II13553;
wire g9119;
wire g3229;
wire II11614;
wire g6701;
wire g2407;
wire g9068;
wire II10752;
wire g6600;
wire g4798;
wire II11060;
wire g4800;
wire g8622;
wire g9049;
wire g4789;
wire g2646;
wire g7306;
wire II6963;
wire g8151;
wire g2174;
wire II6997;
wire II12833;
wire g3499;
wire g7342;
wire g1746;
wire g4436;
wire g7269;
wire g5623;
wire II13209;
wire g3845;
wire II15169;
wire g5562;
wire g3992;
wire g7746;
wire II12442;
wire II13570;
wire II14244;
wire II14058;
wire II14196;
wire g4403;
wire II10815;
wire II13550;
wire g4443;
wire II16061;
wire g6976;
wire g3315;
wire II15857;
wire g3629;
wire g8256;
wire II6716;
wire II8161;
wire II8754;
wire g1941;
wire g6604;
wire g8814;
wire II13785;
wire g5725;
wire II12052;
wire II6078;
wire g3873;
wire II5609;
wire g6622;
wire II12080;
wire g7094;
wire g6109;
wire g1573;
wire II11926;
wire g4472;
wire II12490;
wire g6319;
wire II7459;
wire II15086;
wire g9206;
wire II7523;
wire g5433;
wire II14932;
wire II9681;
wire g7455;
wire g3514;
wire g3854;
wire g7483;
wire g5595;
wire II7239;
wire g8782;
wire g5583;
wire II14725;
wire II7195;
wire g9344;
wire g3516;
wire II11991;
wire g1584;
wire II14035;
wire g4053;
wire II7287;
wire II6309;
wire g8921;
wire g6940;
wire II9918;
wire II13359;
wire II8033;
wire g4712;
wire II7293;
wire g3583;
wire g6568;
wire g6063;
wire g9147;
wire g8695;
wire g3529;
wire II8277;
wire g4363;
wire g8077;
wire II8775;
wire g8998;
wire II9591;
wire g8850;
wire II9678;
wire gbuf44;
wire g7781;
wire g8954;
wire g4412;
wire g7768;
wire g5068;
wire g5752;
wire g6431;
wire g8226;
wire II16135;
wire g6300;
wire II9440;
wire g4658;
wire II13577;
wire II7232;
wire II13012;
wire II13066;
wire II15071;
wire g4238;
wire II8724;
wire g8977;
wire g8882;
wire g4417;
wire g1743;
wire II11827;
wire II12196;
wire g5696;
wire g9151;
wire g1774;
wire II8751;
wire g3075;
wire g5823;
wire gbuf36;
wire g6864;
wire g9386;
wire g6398;
wire II15031;
wire g4066;
wire g5230;
wire g4583;
wire g6589;
wire II9383;
wire II5908;
wire g4631;
wire II9785;
wire g3541;
wire g3019;
wire g4796;
wire g7078;
wire II6853;
wire II9336;
wire g8789;
wire II13196;
wire g2453;
wire g7043;
wire g5476;
wire g4246;
wire g7146;
wire II8510;
wire g6779;
wire g4366;
wire g7096;
wire II14777;
wire II6099;
wire g3286;
wire II6267;
wire g6969;
wire g9061;
wire g2016;
wire g7679;
wire II11326;
wire g7347;
wire g6374;
wire g1611;
wire II12154;
wire II8524;
wire g6183;
wire II14273;
wire II15855;
wire g8541;
wire II13587;
wire II7959;
wire g7010;
wire g8689;
wire g4109;
wire II11135;
wire gbuf56;
wire g4394;
wire II7164;
wire g5681;
wire II9567;
wire II6337;
wire g6684;
wire g6006;
wire II6561;
wire g5713;
wire gbuf9;
wire g1826;
wire II11144;
wire g3928;
wire g7312;
wire g3612;
wire g4135;
wire g8061;
wire g1929;
wire g7609;
wire II8224;
wire g7778;
wire II11055;
wire g8621;
wire g3578;
wire g6878;
wire g5546;
wire g7486;
wire g5309;
wire II9053;
wire II8814;
wire g7365;
wire g5513;
wire II13293;
wire II6608;
wire g5733;
wire g5767;
wire g7744;
wire II9463;
wire g4378;
wire II11200;
wire g8899;
wire II15100;
wire g9074;
wire g6281;
wire g5418;
wire g7138;
wire g8309;
wire II9466;
wire II8922;
wire II12776;
wire g2351;
wire II8446;
wire gbuf73;
wire II5413;
wire II10836;
wire g5343;
wire II8456;
wire II7392;
wire g9168;
wire II9684;
wire g3532;
wire g4186;
wire II5901;
wire g4314;
wire g3983;
wire g2798;
wire g5750;
wire g4100;
wire II14603;
wire II8064;
wire g4958;
wire g7212;
wire g4625;
wire g4837;
wire II6273;
wire g9129;
wire g6021;
wire II10982;
wire II16151;
wire g1773;
wire g4832;
wire II15329;
wire g7359;
wire g5452;
wire II11890;
wire g4004;
wire II13828;
wire II8715;
wire II13663;
wire g8874;
wire g7602;
wire II6939;
wire g2384;
wire II6728;
wire II13045;
wire g2752;
wire g3340;
wire g7080;
wire g7190;
wire g6815;
wire g3777;
wire g6198;
wire g3969;
wire g9339;
wire g7062;
wire g3190;
wire g6830;
wire g8777;
wire II15723;
wire g1679;
wire g4380;
wire g8747;
wire g4546;
wire g9086;
wire g5045;
wire II16165;
wire g6839;
wire g6228;
wire g5649;
wire II7255;
wire g3232;
wire II15018;
wire g9113;
wire g8821;
wire g8826;
wire g4220;
wire g5070;
wire II10197;
wire g8802;
wire g8523;
wire II14202;
wire II8133;
wire g7197;
wire II11873;
wire II14795;
wire II14012;
wire II13979;
wire II15601;
wire g4456;
wire II11722;
wire II9158;
wire g7426;
wire II11194;
wire g5741;
wire II10969;
wire II5425;
wire II8859;
wire g1663;
wire II6198;
wire II7981;
wire II15638;
wire g1577;
wire g7164;
wire g8670;
wire g8718;
wire II13846;
wire II7104;
wire g7825;
wire g6913;
wire g2268;
wire g4257;
wire II12598;
wire II14400;
wire g3504;
wire II13816;
wire g2474;
wire II12639;
wire II14088;
wire g4227;
wire g4327;
wire II11025;
wire II11736;
wire g4701;
wire II13122;
wire g4536;
wire II15622;
wire II10875;
wire II7126;
wire g5128;
wire II16173;
wire II15619;
wire II14211;
wire g1967;
wire g4335;
wire g6618;
wire g5061;
wire g9091;
wire II11939;
wire g8945;
wire g4195;
wire II14338;
wire g2929;
wire II5362;
wire g8764;
wire g2275;
wire g7566;
wire II15242;
wire g6729;
wire g7354;
wire g8562;
wire g6504;
wire g2818;
wire g5786;
wire g5807;
wire g6321;
wire II8338;
wire II13112;
wire g5222;
wire g5233;
wire II11136;
wire g6206;
wire II13861;
wire II11186;
wire II15284;
wire g4349;
wire g7546;
wire g1935;
wire II13092;
wire g3522;
wire II13099;
wire II14662;
wire II7662;
wire g7001;
wire g5001;
wire g5171;
wire II14951;
wire II13894;
wire g9108;
wire g3989;
wire g7633;
wire g2908;
wire II12829;
wire g3842;
wire g6765;
wire g8797;
wire II15388;
wire g7067;
wire II14646;
wire II14420;
wire g8639;
wire g5468;
wire g4006;
wire g8066;
wire g5208;
wire g5642;
wire g2892;
wire g4017;
wire g9098;
wire g2096;
wire II8552;
wire II7314;
wire II15708;
wire g2743;
wire II14848;
wire II11001;
wire g4430;
wire II13185;
wire g8783;
wire g8984;
wire II8977;
wire g2073;
wire g7628;
wire g6313;
wire g1889;
wire g8711;
wire II10283;
wire g5836;
wire II14070;
wire II6887;
wire II11645;
wire II6553;
wire gbuf49;
wire g9213;
wire g4500;
wire g8628;
wire II7383;
wire g8762;
wire g9183;
wire g6956;
wire g7224;
wire g7753;
wire g5077;
wire II12976;
wire g1586;
wire II15845;
wire g6751;
wire g7835;
wire g5529;
wire g6693;
wire g8918;
wire II12003;
wire II6820;
wire g4609;
wire II13329;
wire g3815;
wire II12684;
wire gbuf18;
wire g2555;
wire g6842;
wire II7233;
wire g8602;
wire II8000;
wire II14925;
wire II9978;
wire g4561;
wire II12161;
wire g6514;
wire g5201;
wire g6151;
wire g4558;
wire g6361;
wire g3502;
wire g1733;
wire g9142;
wire II10901;
wire g6644;
wire g9120;
wire g7071;
wire g6168;
wire g5059;
wire II13347;
wire II12135;
wire II12782;
wire gbuf66;
wire II11344;
wire g2897;
wire g2924;
wire g9234;
wire g8342;
wire II12655;
wire g6705;
wire g5193;
wire g8790;
wire g6436;
wire g4783;
wire II13338;
wire II7277;
wire g2777;
wire g5575;
wire II11452;
wire II12866;
wire g4492;
wire II12517;
wire II7347;
wire g6014;
wire II14019;
wire g4306;
wire II15735;
wire II13388;
wire g7723;
wire g4575;
wire g7327;
wire II14145;
wire II13613;
wire g7039;
wire g4889;
wire g4512;
wire II10719;
wire g8175;
wire g5129;
wire g7205;
wire g6715;
wire g5052;
wire g4010;
wire II7492;
wire g8510;
wire g5612;
wire g4922;
wire g5444;
wire II15417;
wire g2768;
wire II11750;
wire g5148;
wire g7587;
wire g7520;
wire II12571;
wire g3259;
wire g7855;
wire II13755;
wire g6299;
wire g5179;
wire g8800;
wire II12403;
wire g8677;
wire II5471;
wire II8015;
wire II15228;
wire II10072;
wire g6258;
wire II12646;
wire g8901;
wire II9034;
wire II12484;
wire g5737;
wire g5812;
wire g1557;
wire II7987;
wire g6262;
wire g4882;
wire g3681;
wire II7486;
wire g6231;
wire g3914;
wire g2330;
wire II15231;
wire g6123;
wire II11443;
wire g6592;
wire g6336;
wire II9425;
wire g6171;
wire g7529;
wire g7534;
wire II12011;
wire g3678;
wire g7263;
wire g9185;
wire g6798;
wire II16046;
wire g5207;
wire II12253;
wire g8965;
wire g9367;
wire II11215;
wire g6489;
wire g6901;
wire g2728;
wire g2057;
wire g4826;
wire g5050;
wire II13512;
wire g5184;
wire g5794;
wire g3861;
wire II11488;
wire g7296;
wire g4128;
wire g1869;
wire g3939;
wire g8699;
wire II13541;
wire II12909;
wire II14732;
wire II9985;
wire II15927;
wire g6107;
wire g8381;
wire g4117;
wire II10925;
wire g9022;
wire II13734;
wire g7235;
wire g8861;
wire g6158;
wire II15830;
wire II10271;
wire g6330;
wire g4714;
wire g6295;
wire g2650;
wire g4677;
wire II11281;
wire II5545;
wire g6974;
wire g5152;
wire g9273;
wire g3932;
wire II8820;
wire g4169;
wire II12391;
wire II8071;
wire II12078;
wire g6312;
wire g2618;
wire g8280;
wire II8617;
wire II13915;
wire g4059;
wire g8937;
wire g2695;
wire II15580;
wire g4548;
wire g8012;
wire g6357;
wire g8756;
wire g3630;
wire II8574;
wire g3852;
wire g5988;
wire II12068;
wire gbuf53;
wire II10180;
wire g1832;
wire g7170;
wire II11559;
wire g8903;
wire g8316;
wire g6892;
wire g3770;
wire g2624;
wire II15850;
wire g5265;
wire g2686;
wire g9000;
wire II9419;
wire II10889;
wire II10397;
wire II16100;
wire g7338;
wire g5018;
wire g2659;
wire II5552;
wire II13873;
wire g2870;
wire g4599;
wire g2496;
wire g3512;
wire g9285;
wire II8892;
wire g7241;
wire g7229;
wire II14763;
wire g9012;
wire g7494;
wire g5551;
wire g4684;
wire g6012;
wire II12675;
wire g3539;
wire II13746;
wire g4386;
wire g6115;
wire g7577;
wire II6363;
wire II7504;
wire g4477;
wire g2333;
wire g8831;
wire g9191;
wire g4552;
wire g5939;
wire II10169;
wire g7427;
wire g2955;
wire g5724;
wire g4736;
wire g5057;
wire g6795;
wire g6277;
wire g1718;
wire II11050;
wire II5855;
wire II12757;
wire g6148;
wire II6523;
wire II8471;
wire II11494;
wire g8460;
wire g2367;
wire g2944;
wire g3847;
wire II15714;
wire g2312;
wire g6033;
wire II9633;
wire II11157;
wire II10582;
wire g5872;
wire g9037;
wire g5969;
wire g6810;
wire II11163;
wire II8712;
wire g5518;
wire II11683;
wire II11550;
wire II15043;
wire g2105;
wire g4110;
wire g5622;
wire g6110;
wire II15651;
wire II11476;
wire g6993;
wire g6352;
wire II10930;
wire g3556;
wire g2689;
wire II7706;
wire g2633;
wire g1814;
wire II12712;
wire g3390;
wire II12763;
wire g8644;
wire g1758;
wire g7253;
wire II11359;
wire II7832;
wire g8943;
wire II11341;
wire g3014;
wire g7553;
wire g6506;
wire g7554;
wire g7175;
wire g7712;
wire g9134;
wire g7834;
wire II11696;
wire II11759;
wire g6699;
wire II13247;
wire g8931;
wire g4158;
wire II15543;
wire II7079;
wire II9999;
wire II5520;
wire II9258;
wire II10708;
wire g8855;
wire g4080;
wire II10914;
wire g2271;
wire g9272;
wire g6181;
wire II13271;
wire g7304;
wire g4308;
wire II10151;
wire II10366;
wire II10494;
wire g1643;
wire g5638;
wire g3750;
wire g7186;
wire II14674;
wire g4434;
wire g6925;
wire g3926;
wire g6446;
wire II8955;
wire g4445;
wire g2207;
wire g9328;
wire g5604;
wire g8332;
wire g6075;
wire II7323;
wire g2867;
wire II6856;
wire II10280;
wire g2294;
wire II7728;
wire g6730;
wire g3081;
wire g6307;
wire g8796;
wire II13646;
wire g3497;
wire g6253;
wire g3904;
wire II11299;
wire II11142;
wire II6923;
wire g7653;
wire g1888;
wire II14264;
wire g8304;
wire g3836;
wire g5108;
wire g1678;
wire II12331;
wire II8483;
wire g4915;
wire II7610;
wire g8658;
wire g7511;
wire II6925;
wire II11227;
wire g2931;
wire II13698;
wire g2889;
wire g3561;
wire II11576;
wire g2827;
wire II8862;
wire g6821;
wire g4679;
wire g8564;
wire g3881;
wire II6474;
wire g8648;
wire II12475;
wire g3994;
wire II7947;
wire II13533;
wire g1943;
wire g3784;
wire II13302;
wire II12921;
wire II5371;
wire II11413;
wire g6876;
wire g6742;
wire g4364;
wire g5345;
wire g5364;
wire g4427;
wire II12298;
wire II15084;
wire II11290;
wire g6898;
wire g6441;
wire II9520;
wire g2972;
wire g6481;
wire II12725;
wire g5585;
wire g5662;
wire g6703;
wire g6599;
wire II12853;
wire II14467;
wire II10268;
wire II10545;
wire II14753;
wire II10298;
wire II10259;
wire II6242;
wire g3732;
wire g3656;
wire II7569;
wire g3944;
wire g1638;
wire II9579;
wire II14097;
wire g7454;
wire g8951;
wire II7870;
wire g7951;
wire g5259;
wire g9332;
wire II9642;
wire g4264;
wire g9043;
wire g9112;
wire II13710;
wire g7233;
wire g3647;
wire g4779;
wire g9306;
wire II6299;
wire g4507;
wire II12346;
wire g2214;
wire g1917;
wire g1799;
wire II13084;
wire g7518;
wire g8654;
wire g6885;
wire g4020;
wire g5066;
wire g9201;
wire g5746;
wire g6405;
wire g2884;
wire II11314;
wire g2402;
wire II13810;
wire II7574;
wire g6634;
wire II15933;
wire II10451;
wire g7142;
wire g5487;
wire II14683;
wire g2221;
wire g9007;
wire II11350;
wire g3237;
wire g9123;
wire g5157;
wire II7581;
wire g6415;
wire g2044;
wire II11793;
wire g1737;
wire II12948;
wire gbuf24;
wire II13565;
wire II14342;
wire g1662;
wire g6083;
wire g6346;
wire II11659;
wire g8665;
wire g4616;
wire II8480;
wire II13797;
wire g9039;
wire II8254;
wire g6651;
wire g2241;
wire g7102;
wire II5670;
wire II8328;
wire g5627;
wire II7749;
wire g3896;
wire g8923;
wire g7766;
wire g7488;
wire g6286;
wire II13152;
wire II8582;
wire II9196;
wire II10334;
wire g5030;
wire II13103;
wire g5261;
wire g8897;
wire g7755;
wire g6656;
wire g9279;
wire g8380;
wire II8829;
wire g8836;
wire g4282;
wire II10160;
wire g4510;
wire II10506;
wire g4194;
wire g4823;
wire II8793;
wire g2485;
wire II5395;
wire g7363;
wire II9618;
wire II15773;
wire II5353;
wire II11398;
wire g8582;
wire II6103;
wire g3092;
wire II15598;
wire g2145;
wire g6224;
wire g3466;
wire g6980;
wire II8835;
wire g4284;
wire II5981;
wire g7460;
wire g5819;
wire g1745;
wire g6462;
wire g9080;
wire II10716;
wire g8059;
wire g9379;
wire g7439;
wire II8802;
wire g8660;
wire g7467;
wire g3875;
wire g7345;
wire II15481;
wire II8215;
wire g6672;
wire g1600;
wire g1961;
wire g1616;
wire g6089;
wire g6967;
wire g9030;
wire g6777;
wire II14810;
wire g8232;
wire g5037;
wire g4744;
wire II11843;
wire II10353;
wire II9547;
wire II14175;
wire g8224;
wire II7335;
wire II14851;
wire g9377;
wire g7708;
wire II10842;
wire g6960;
wire g4738;
wire g8611;
wire II9029;
wire g3706;
wire II6791;
wire II12737;
wire g2842;
wire g9343;
wire g2374;
wire g7475;
wire II14028;
wire II9892;
wire g7020;
wire II12586;
wire g5831;
wire g8063;
wire II13779;
wire g9277;
wire g7509;
wire g5570;
wire g8273;
wire g6712;
wire II5657;
wire g8912;
wire II6757;
wire g9056;
wire g2185;
wire g6004;
wire II10019;
wire g6686;
wire II11710;
wire g6471;
wire II13438;
wire g8223;
wire II7461;
wire g4929;
wire g4397;
wire II11434;
wire II13686;
wire gbuf68;
wire g2920;
wire II6770;
wire g9096;
wire g7360;
wire II12352;
wire II9070;
wire g9078;
wire g9219;
wire g4018;
wire g7614;
wire g8849;
wire g3047;
wire g1987;
wire g4743;
wire g3676;
wire g7277;
wire g8610;
wire II15604;
wire g2289;
wire gbuf12;
wire g7037;
wire g4633;
wire g6825;
wire g7226;
wire II9819;
wire g9089;
wire g9076;
wire II5535;
wire II7453;
wire g9154;
wire II10418;
wire g6788;
wire g2237;
wire g1564;
wire g7887;
wire II7173;
wire II7480;
wire II9129;
wire g8634;
wire II5428;
wire g5593;
wire g4904;
wire g6305;
wire II16072;
wire g4051;
wire g3980;
wire g5173;
wire g7698;
wire g4104;
wire g5736;
wire g9227;
wire II12505;
wire g6869;
wire g7728;
wire g8889;
wire II11248;
wire g8869;
wire II8605;
wire g4202;
wire g5239;
wire g6516;
wire g4147;
wire g8009;
wire g7721;
wire g8235;
wire II8727;
wire g4907;
wire g4464;
wire g1708;
wire g6477;
wire g4229;
wire II10466;
wire g3008;
wire II14279;
wire g9236;
wire II6878;
wire II11008;
wire g6221;
wire g6424;
wire g6680;
wire II7867;
wire g6386;
wire g3049;
wire II5633;
wire g5644;
wire g8724;
wire g5264;
wire II12031;
wire II12164;
wire g9352;
wire II8296;
wire II6751;
wire II5389;
wire g6242;
wire g5122;
wire II8340;
wire II5960;
wire II9669;
wire g1942;
wire II11266;
wire g6068;
wire g6449;
wire II13770;
wire g5762;
wire II9603;
wire g8156;
wire g6440;
wire g8808;
wire II9955;
wire g3503;
wire g5873;
wire II13250;
wire g2233;
wire g6933;
wire g7270;
wire g8824;
wire g7341;
wire g3956;
wire g4254;
wire g1570;
wire II10627;
wire g2793;
wire II12529;
wire g6187;
wire II15196;
wire g7718;
wire II7847;
wire II15635;
wire g3962;
wire g7151;
wire g5661;
wire g8607;
wire g1749;
wire g5432;
wire g5801;
wire g6574;
wire II10061;
wire g4299;
wire g1837;
wire II12731;
wire II14082;
wire g8952;
wire II11875;
wire g3665;
wire g1788;
wire g6040;
wire II14136;
wire II5732;
wire g6311;
wire g4517;
wire II13383;
wire g2973;
wire II15577;
wire g4532;
wire g8323;
wire II7765;
wire g3838;
wire g7833;
wire II10305;
wire g4666;
wire g4877;
wire II6590;
wire II15241;
wire g4808;
wire g7419;
wire g6408;
wire II12748;
wire g5044;
wire II7885;
wire g9106;
wire II12158;
wire II6081;
wire g5220;
wire II14623;
wire II6192;
wire g8721;
wire II8202;
wire II8491;
wire g4085;
wire II9202;
wire g5511;
wire II11185;
wire II11818;
wire g6438;
wire g6664;
wire II12101;
wire g7126;
wire g3654;
wire II8363;
wire g699;
wire g1801;
wire g2546;
wire g7742;
wire g8793;
wire g6210;
wire II6189;
wire II9393;
wire g7324;
wire g2511;
wire g8438;
wire g4719;
wire g2878;
wire II5598;
wire g7420;
wire g6342;
wire II7386;
wire g5090;
wire II15208;
wire g6784;
wire g8442;
wire II11884;
wire g2932;
wire II7939;
wire g2909;
wire II6446;
wire II10532;
wire g2490;
wire g1725;
wire g7098;
wire II15918;
wire II14234;
wire II7731;
wire g1681;
wire g5428;
wire g6165;
wire g6911;
wire II12520;
wire g7583;
wire g7210;
wire g6265;
wire II13598;
wire g5715;
wire II6171;
wire g7083;
wire g8174;
wire II12108;
wire g8969;
wire II12983;
wire g5466;
wire II9660;
wire g5654;
wire II8428;
wire g6359;
wire II11861;
wire II8432;
wire g5722;
wire g4588;
wire g7336;
wire II7158;
wire II8308;
wire g7348;
wire g8785;
wire II6102;
wire II13396;
wire II6130;
wire II6434;
wire II15414;
wire g4570;
wire g1579;
wire II12538;
wire g9044;
wire g3981;
wire g6972;
wire g6598;
wire g8775;
wire g6625;
wire g8604;
wire II16055;
wire g8713;
wire g4303;
wire II6723;
wire g1588;
wire g8760;
wire II10060;
wire II12965;
wire g5759;
wire g5740;
wire g8999;
wire g2843;
wire g6840;
wire g6954;
wire g6862;
wire g6566;
wire g8688;
wire II9687;
wire II15814;
wire g5095;
wire g8306;
wire g2902;
wire g2226;
wire II7911;
wire g2958;
wire g8407;
wire g3906;
wire g2364;
wire II6842;
wire g2382;
wire II8477;
wire g3589;
wire II10360;
wire g6636;
wire g6283;
wire II10829;
wire g9058;
wire II12120;
wire g4216;
wire g7565;
wire II7902;
wire g6640;
wire II15592;
wire g3530;
wire g8772;
wire g5516;
wire II8470;
wire g4573;
wire II11607;
wire gbuf7;
wire g6794;
wire II7479;
wire g8584;
wire g6052;
wire g8082;
wire II10433;
wire g8896;
wire II10744;
wire g3811;
wire g5697;
wire g7060;
wire g8957;
wire g5577;
wire g4525;
wire g2883;
wire g6384;
wire g4107;
wire g5065;
wire g8378;
wire g4638;
wire II15408;
wire g4118;
wire g3074;
wire g6946;
wire g5799;
wire II12148;
wire II11115;
wire II15693;
wire II7011;
wire g8071;
wire II9330;
wire II12277;
wire g8842;
wire g7992;
wire gbuf34;
wire g3693;
wire g6991;
wire g6091;
wire g3158;
wire gbuf41;
wire II12852;
wire g8990;
wire g4640;
wire g3642;
wire II8496;
wire g5442;
wire g8685;
wire II12547;
wire g6205;
wire II12098;
wire g2454;
wire g6774;
wire g2459;
wire g1661;
wire II11458;
wire II8193;
wire g6778;
wire g8013;
wire g6289;
wire g7171;
wire II13885;
wire II6066;
wire II11467;
wire g4232;
wire II6686;
wire g6591;
wire g6182;
wire II15953;
wire gbuf19;
wire g4022;
wire II8730;
wire II12044;
wire g7195;
wire g8317;
wire II8850;
wire II13109;
wire g8040;
wire g7356;
wire g1701;
wire g7608;
wire g7526;
wire II10681;
wire g7041;
wire II13290;
wire g6059;
wire g9349;
wire II14103;
wire g9381;
wire II12635;
wire II11491;
wire g4362;
wire II8523;
wire g6232;
wire g5559;
wire II15109;
wire g3258;
wire II7428;
wire gbuf54;
wire g6763;
wire II8956;
wire II6090;
wire g4604;
wire g7042;
wire g6132;
wire II9627;
wire g5474;
wire g4578;
wire g4008;
wire g3917;
wire g5754;
wire g3927;
wire II8354;
wire II10135;
wire II7716;
wire II9760;
wire g6397;
wire II13203;
wire g6689;
wire II13758;
wire g5440;
wire II8418;
wire g4034;
wire g7775;
wire g5463;
wire g4377;
wire g8094;
wire g8076;
wire g6178;
wire g4645;
wire g4193;
wire g5212;
wire g5690;
wire II15102;
wire II8679;
wire II12283;
wire g7309;
wire g8543;
wire II13299;
wire II7240;
wire g4653;
wire II6029;
wire g1597;
wire II8041;
wire g7737;
wire g5034;
wire g3996;
wire II10482;
wire g3519;
wire g2652;
wire g4879;
wire g6154;
wire g4794;
wire g8637;
wire II10144;
wire g2128;
wire g1860;
wire g5079;
wire g4191;
wire g7046;
wire II5747;
wire II9828;
wire II16122;
wire g7091;
wire II7180;
wire II10953;
wire II15565;
wire g9046;
wire II9539;
wire II13118;
wire II13051;
wire II13161;
wire II9615;
wire g8674;
wire II9116;
wire II14677;
wire II9768;
wire g8701;
wire II16090;
wire II7672;
wire g9032;
wire g2216;
wire g6348;
wire g6203;
wire g6482;
wire g1672;
wire g6965;
wire g5598;
wire g6611;
wire II12328;
wire g7499;
wire g4691;
wire g3691;
wire g8177;
wire g8748;
wire g8656;
wire II10820;
wire g5591;
wire g9371;
wire g5700;
wire II8282;
wire II15297;
wire g8754;
wire II15082;
wire II14112;
wire II8874;
wire II12436;
wire II8618;
wire g5830;
wire g7466;
wire g2007;
wire g5081;
wire g9014;
wire g1590;
wire gbuf61;
wire g6880;
wire g5032;
wire g6463;
wire g1867;
wire g2807;
wire g8833;
wire g5561;
wire g6088;
wire g4504;
wire II12310;
wire g5437;
wire g5671;
wire g9006;
wire g8627;
wire g9301;
wire II14838;
wire g7687;
wire g8963;
wire g5481;
wire II10183;
wire g3086;
wire II6711;
wire g8929;
wire II5519;
wire II6952;
wire g4687;
wire g7627;
wire II7214;
wire g1912;
wire g6073;
wire g8922;
wire II12292;
wire g5606;
wire g3707;
wire g8493;
wire g6460;
wire g7013;
wire g6647;
wire II7187;
wire II5664;
wire g7183;
wire g2376;
wire g1658;
wire g5072;
wire g3877;
wire g5566;
wire g5169;
wire g6009;
wire g6694;
wire g4286;
wire g2946;
wire g5039;
wire g1816;
wire g7782;
wire g2629;
wire g7029;
wire g2205;
wire g7773;
wire gbuf25;
wire II6669;
wire II16017;
wire g8291;
wire II7850;
wire g1964;
wire II13199;
wire g7335;
wire II9276;
wire g4079;
wire g7231;
wire g3521;
wire II12427;
wire g6039;
wire II13481;
wire II11757;
wire g9064;
wire g8330;
wire II14208;
wire II8832;
wire g6801;
wire g4872;
wire g5285;
wire II13444;
wire g5162;
wire g9322;
wire II8635;
wire g2914;
wire II14857;
wire II11955;
wire g2986;
wire g3528;
wire II15663;
wire g1558;
wire g5817;
wire g3868;
wire II15202;
wire II12702;
wire g8339;
wire g4801;
wire g6251;
wire g9270;
wire g3941;
wire g6487;
wire g9198;
wire II6815;
wire II9089;
wire g5796;
wire II7478;
wire g2259;
wire g9187;
wire II10862;
wire g6732;
wire g8818;
wire II13422;
wire g3968;
wire g3943;
wire g6843;
wire II6186;
wire II7878;
wire g2347;
wire g9116;
wire g4082;
wire II10262;
wire g7541;
wire g7548;
wire g3870;
wire g4425;
wire II15513;
wire II8090;
wire II12551;
wire g3231;
wire g9340;
wire II15263;
wire g5826;
wire g3582;
wire g8858;
wire g2285;
wire II10643;
wire II14722;
wire II15253;
wire g6323;
wire II13610;
wire II14424;
wire II14325;
wire g8935;
wire g3635;
wire II8560;
wire g6134;
wire II7061;
wire gbuf39;
wire II7531;
wire g7561;
wire g9329;
wire II7859;
wire g7086;
wire g2643;
wire g4913;
wire g4539;
wire II12117;
wire g4593;
wire g5732;
wire g5479;
wire II11512;
wire g4351;
wire g1775;
wire II6946;
wire g5402;
wire g4256;
wire II13617;
wire II9477;
wire g4163;
wire g7302;
wire g7007;
wire g8512;
wire g7691;
wire g4935;
wire g9141;
wire g2486;
wire g6275;
wire II9170;
wire g2617;
wire g4315;
wire g3934;
wire g7242;
wire g2363;
wire g3887;
wire g6106;
wire II5775;
wire g4734;
wire g5842;
wire g6326;
wire g1732;
wire g8128;
wire g3038;
wire g4936;
wire II11903;
wire g7104;
wire II11908;
wire g4251;
wire g7260;
wire II9194;
wire II11897;
wire II6767;
wire II9142;
wire II8119;
wire g8264;
wire g4780;
wire g4727;
wire g3977;
wire g5046;
wire g8015;
wire g6727;
wire II5865;
wire II15607;
wire g2325;
wire g6613;
wire g7255;
wire g4275;
wire g4547;
wire g6018;
wire g7412;
wire II12033;
wire II15921;
wire g3225;
wire II7775;
wire g6011;
wire g8283;
wire g8949;
wire g7437;
wire II10890;
wire g6139;
wire II13353;
wire g3604;
wire II14451;
wire g9180;
wire II6739;
wire II6135;
wire g6433;
wire II11377;
wire g6559;
wire g3897;
wire g1756;
wire II14160;
wire II7308;
wire g5115;
wire II7139;
wire g7496;
wire g1895;
wire II7892;
wire II5972;
wire g8483;
wire g2698;
wire II9588;
wire g2404;
wire g4159;
wire g6266;
wire g9294;
wire g2622;
wire II10186;
wire g3825;
wire g5298;
wire g8088;
wire II9132;
wire g3954;
wire II8808;
wire g3880;
wire II12839;
wire g7575;
wire g8917;
wire g9281;
wire II14366;
wire g4400;
wire g4569;
wire g4921;
wire g1904;
wire II12999;
wire g2635;
wire g1878;
wire II8001;
wire g4475;
wire g7764;
wire II12235;
wire g7247;
wire g3310;
wire g9099;
wire g2276;
wire g7223;
wire II11984;
wire g5586;
wire g2170;
wire g5918;
wire g4230;
wire II11500;
wire g8513;
wire g2895;
wire g4742;
wire II8233;
wire II15218;
wire II15290;
wire g1808;
wire II15232;
wire g3722;
wire II8452;
wire g8693;
wire g9313;
wire g7444;
wire II11101;
wire g4894;
wire II12151;
wire II6904;
wire II8101;
wire g7240;
wire II6539;
wire g5291;
wire g5810;
wire II9948;
wire g8851;
wire g5278;
wire g4695;
wire g7585;
wire g8298;
wire II9794;
wire II11365;
wire II11095;
wire g5002;
wire g1780;
wire II15839;
wire g3563;
wire g6121;
wire II12173;
wire II11638;
wire g7501;
wire g7117;
wire g4244;
wire g6823;
wire g8867;
wire g8880;
wire II13767;
wire g4122;
wire g4704;
wire g5146;
wire II8971;
wire g6903;
wire g2235;
wire g6024;
wire g2919;
wire II8589;
wire g4175;
wire g4962;
wire g2011;
wire g6740;
wire g9026;
wire g5614;
wire g2868;
wire g6338;
wire g8900;
wire g6714;
wire g5611;
wire g5334;
wire II15222;
wire g2310;
wire II5542;
wire g4870;
wire g9020;
wire g9222;
wire II6636;
wire II13692;
wire g6759;
wire II9151;
wire g6297;
wire g7109;
wire g6159;
wire g8707;
wire g3495;
wire g8879;
wire II6864;
wire g5156;
wire II15394;
wire g4888;
wire II14442;
wire g8328;
wire g8813;
wire g8266;
wire II6202;
wire II6532;
wire g6413;
wire g5631;
wire II6121;
wire II14484;
wire II16023;
wire g1830;
wire g8829;
wire II11591;
wire g9334;
wire II9621;
wire II12065;
wire g4910;
wire g1955;
wire II8565;
wire g6723;
wire II12367;
wire g7563;
wire II8790;
wire II13800;
wire II10786;
wire g2640;
wire g8744;
wire II11744;
wire g6257;
wire g6921;
wire g4563;
wire g4252;
wire g8840;
wire g6806;
wire g4483;
wire II12038;
wire g3501;
wire II8880;
wire II12690;
wire g1688;
wire II8940;
wire II8569;
wire g6510;
wire II10574;
wire g4813;
wire g1786;
wire II11401;
wire g5600;
wire g8181;
wire g7611;
wire g7434;
wire g4591;
wire g1572;
wire II10193;
wire g7579;
wire II10766;
wire g6496;
wire g2795;
wire g1908;
wire II12810;
wire II13072;
wire g7422;
wire II7623;
wire g4087;
wire g5092;
wire g8312;
wire g4200;
wire g2966;
wire g6851;
wire g2817;
wire II14388;
wire g9130;
wire II15982;
wire g8822;
wire II10010;
wire II13378;
wire II9058;
wire g8308;
wire g4130;
wire II12211;
wire g6508;
wire II8980;
wire g2424;
wire g9117;
wire g2654;
wire II13865;
wire g8321;
wire g5652;
wire g6317;
wire g6615;
wire g4271;
wire g7749;
wire g4806;
wire g5657;
wire II11616;
wire g6907;
wire g9388;
wire g6163;
wire g9209;
wire g9104;
wire g3617;
wire II11575;
wire II7320;
wire II10343;
wire g2904;
wire g7166;
wire g8609;
wire II7632;
wire g2352;
wire g9071;
wire g4026;
wire II5600;
wire II14073;
wire II8766;
wire g5426;
wire g2905;
wire g7032;
wire g1726;
wire g5769;
wire II10522;
wire g8146;
wire g2514;
wire II13189;
wire g4319;
wire g4452;
wire g6734;
wire II10625;
wire g5214;
wire g6737;
wire g6782;
wire II7517;
wire II6270;
wire II12358;
wire g2231;
wire II14334;
wire g6820;
wire g7311;
wire g4375;
wire g5204;
wire g5311;
wire II13580;
wire g4829;
wire g8042;
wire g4297;
wire II9889;
wire g9362;
wire II10157;
wire g4032;
wire g5572;
wire II10867;
wire g5042;
wire II6057;
wire II5697;
wire g5021;
wire II13048;
wire g9094;
wire g7035;
wire g3831;
wire g5579;
wire g8179;
wire II6740;
wire g5237;
wire II9585;
wire II10300;
wire g7058;
wire g3573;
wire II15484;
wire g3890;
wire II12681;
wire g7689;
wire g5522;
wire II12936;
wire g5897;
wire II13472;
wire g4190;
wire g3674;
wire g9217;
wire g6244;
wire g636;
wire II10380;
wire g4357;
wire g7279;
wire g8799;
wire g1901;
wire II10040;
wire II12609;
wire II8019;
wire II15261;
wire g7281;
wire g7323;
wire II8928;
wire g7318;
wire g2292;
wire g8847;
wire g5781;
wire II11656;
wire II13518;
wire gbuf14;
wire g5833;
wire II11732;
wire g6786;
wire g8993;
wire g4776;
wire II11191;
wire II9570;
wire II8593;
wire II5817;
wire g8910;
wire II9834;
wire g7124;
wire II8143;
wire g6928;
wire II7140;
wire g8632;
wire g9138;
wire II14792;
wire g4626;
wire II14637;
wire II11641;
wire g5086;
wire g7704;
wire g8715;
wire g8286;
wire g5190;
wire g2327;
wire II6876;
wire g2501;
wire II10509;
wire g7447;
wire g8459;
wire II7510;
wire g8259;
wire II11335;
wire g9238;
wire g4016;
wire g6835;
wire g7789;
wire II8503;
wire g2871;
wire g9350;
wire g8292;
wire II5416;
wire g6717;
wire g6473;
wire II10497;
wire g6020;
wire g4014;
wire II13002;
wire g4102;
wire gbuf21;
wire g6047;
wire II5969;
wire II15899;
wire II8919;
wire g8080;
wire II12945;
wire g3987;
wire g6682;
wire g4745;
wire II10998;
wire g9082;
wire II7667;
wire g4074;
wire g2764;
wire II10500;
wire g4676;
wire g8078;
wire g4369;
wire g5124;
wire II7468;
wire g2893;
wire II8799;
wire II11455;
wire g8887;
wire II7738;
wire II6657;
wire II14001;
wire g2528;
wire g5710;
wire g5871;
wire g6597;
wire II13956;
wire g9051;
wire g6944;
wire g6290;
wire II13088;
wire g8073;
wire g1855;
wire g8973;
wire g4523;
wire g6422;
wire II10320;
wire g5448;
wire g5556;
wire g5764;
wire II10307;
wire II13574;
wire g4384;
wire g8992;
wire II6257;
wire g7700;
wire g4320;
wire II6294;
wire II6788;
wire II11923;
wire II6015;
wire g6585;
wire g5175;
wire g4902;
wire g4668;
wire II15699;
wire g6520;
wire g7057;
wire g2573;
wire g6098;
wire g2840;
wire II16148;
wire g6979;
wire g4281;
wire g9143;
wire g4360;
wire g5685;
wire II10796;
wire II10299;
wire g3964;
wire g6538;
wire II15978;
wire II9791;
wire g9303;
wire II10094;
wire g4055;
wire II8528;
wire g2452;
wire II15272;
wire g6867;
wire II11648;
wire g5557;
wire II10991;
wire II12973;
wire g3818;
wire II14680;
wire g4651;
wire g7266;
wire g8230;
wire g3959;
wire g3591;
wire g8221;
wire g9383;
wire II7362;
wire g6027;
wire g4641;
wire g6378;
wire II9691;
wire g2942;
wire g3524;
wire g2949;
wire g6959;
wire g3510;
wire g7128;
wire g6042;
wire g4554;
wire gbuf52;
wire II14430;
wire g6218;
wire g2927;
wire g6916;
wire II14813;
wire g4729;
wire g8440;
wire g5013;
wire II6109;
wire g8683;
wire g4544;
wire g9315;
wire II10079;
wire gbuf32;
wire g4647;
wire g6791;
wire g4576;
wire gbuf48;
wire g9255;
wire II11752;
wire g1747;
wire g6180;
wire g7739;
wire g6394;
wire g4968;
wire gbuf28;
wire g2521;
wire g8545;
wire g4390;
wire g2309;
wire g9248;
wire g7343;
wire g6478;
wire g6761;
wire g5255;
wire g8734;
wire II12742;
wire g5755;
wire II13308;
wire g8835;
wire g2263;
wire II9657;
wire g2287;
wire II7156;
wire II14294;
wire g5266;
wire g9220;
wire g5461;
wire g6399;
wire g3700;
wire II14990;
wire g2378;
wire II5872;
wire II5754;
wire II9782;
wire II12952;
wire g3079;
wire II9475;
wire g5229;
wire g3264;
wire II9675;
wire g7216;
wire g6403;
wire II6172;
wire g3461;
wire g5007;
wire g1843;
wire g6860;
wire II9994;
wire II10327;
wire g8773;
wire II13825;
wire g5023;
wire g2478;
wire II13407;
wire II13496;
wire g9336;
wire g8326;
wire g4098;
wire g2471;
wire II6759;
wire g5144;
wire g6002;
wire g4615;
wire g7088;
wire g2937;
wire g8686;
wire g6627;
wire II10847;
wire II12271;
wire g3061;
wire g5195;
wire II6844;
wire II12241;
wire gbuf59;
wire g4955;
wire II7359;
wire g5063;
wire g6887;
wire g4301;
wire II12942;
wire g8405;
wire g7415;
wire II7115;
wire g2457;
wire g8950;
wire g7405;
wire g2380;
wire g1823;
wire II15888;
wire II10032;
wire II7138;
wire II6060;
wire g7740;
wire II6831;
wire II6154;
wire g2148;
wire g6948;
wire II12596;
wire g8894;
wire g6285;
wire g6638;
wire g2886;
wire g6811;
wire II13441;
wire II10937;
wire II10080;
wire g7116;
wire g4836;
wire g2348;
wire g8770;
wire II7595;
wire g1945;
wire g6195;
wire g4586;
wire g2397;
wire II15112;
wire II7758;
wire g6642;
wire g8726;
wire g6501;
wire g8093;
wire g8300;
wire II11260;
wire g5717;
wire II6239;
wire II9752;
wire g6998;
wire II9594;
wire g4621;
wire g5493;
wire g5699;
wire g4344;
wire g7517;
wire g4139;
wire g7077;
wire g2224;
wire II14214;
wire II13466;
wire II11806;
wire II11917;
wire g7580;
wire g4037;
wire II13356;
wire II6024;
wire II11374;
wire g8337;
wire g9101;
wire g5581;
wire II12361;
wire gbuf37;
wire g8270;
wire g7333;
wire g3546;
wire II16116;
wire g8792;
wire g6161;
wire g7837;
wire g2912;
wire g6061;
wire II14454;
wire II10314;
wire g3652;
wire g8237;
wire II13238;
wire g1685;
wire II13023;
wire II16009;
wire g6037;
wire II11356;
wire g4077;
wire g7300;
wire g2935;
wire II9014;
wire g2648;
wire g3948;
wire II11987;
wire g8853;
wire g3526;
wire g3640;
wire g6852;
wire g5113;
wire g4462;
wire g6466;
wire II15747;
wire g2401;
wire II10427;
wire II12059;
wire II11395;
wire II11407;
wire II13274;
wire II8094;
wire g6578;
wire g3908;
wire g1652;
wire g6918;
wire g8153;
wire II16129;
wire II6084;
wire g4084;
wire II12768;
wire II15741;
wire g5625;
wire II13782;
wire g2394;
wire g3872;
wire g8199;
wire g4423;
wire g9024;
wire II15068;
wire g9196;
wire g3430;
wire g7429;
wire g9179;
wire g6935;
wire g6633;
wire g8805;
wire g7133;
wire g1566;
wire II15687;
wire g9145;
wire II5679;
wire II12493;
wire II12448;
wire II14718;
wire g5083;
wire II14205;
wire II5766;
wire g6889;
wire II9745;
wire II13819;
wire g7870;
wire II6245;
wire II9234;
wire II8637;
wire g9324;
wire g5240;
wire II11680;
wire II7723;
wire g3131;
wire g4635;
wire g6631;
wire II9278;
wire II6597;
wire g1898;
wire II10705;
wire g1811;
wire g7515;
wire g4392;
wire II15337;
wire II15562;
wire g2283;
wire g4089;
wire II12523;
wire g1777;
wire g9066;
wire g4473;
wire II7503;
wire II12208;
wire g3879;
wire II14463;
wire g1674;
wire g5036;
wire g8751;
wire II8660;
wire g8285;
wire II11108;
wire g6891;
wire g6808;
wire g2481;
wire II15930;
wire II6916;
wire g2615;
wire II9059;
wire g4176;
wire II13057;
wire g2761;
wire g2536;
wire g5844;
wire II14844;
wire g4268;
wire g6856;
wire g4747;
wire II10204;
wire II8910;
wire g6246;
wire g7015;
wire g9002;
wire g5472;
wire II7658;
wire g9004;
wire II11437;
wire g4890;
wire g4792;
wire g4581;
wire g4448;
wire g5055;
wire II10142;
wire g6676;
wire g6418;
wire II11416;
wire g2668;
wire g4407;
wire II12322;
wire g6831;
wire g6096;
wire II8559;
wire g2863;
wire g4693;
wire g4317;
wire II9084;
wire II12202;
wire g8988;
wire g7735;
wire II13031;
wire g6595;
wire g8038;
wire II15937;
wire II12418;
wire g7652;
wire g6963;
wire g5483;
wire II14495;
wire g5167;
wire g4024;
wire g4787;
wire II15165;
wire g4602;
wire II14238;
wire g7027;
wire II6813;
wire g3974;
wire g4810;
wire II11031;
wire II7746;
wire II8938;
wire II11117;
wire II5839;
wire II14154;
wire g1612;
wire g7435;
wire g7793;
wire g8914;
wire g6649;
wire g6209;
wire g8279;
wire g9373;
wire g6304;
wire II8658;
wire II9535;
wire g3050;
wire g7811;
wire II7095;
wire g9110;
wire II7068;
wire g4697;
wire II13157;
wire g5539;
wire g6007;
wire g4689;
wire II11079;
wire II13502;
wire g7471;
wire II6000;
wire II11123;
wire II13451;
wire g7762;
wire g5015;
wire g4288;
wire g3339;
wire II12421;
wire g5384;
wire II12897;
wire g5868;
wire II9350;
wire g8942;
wire g6292;
wire g4469;
wire II5914;
wire g6602;
wire II14251;
wire g4358;
wire g7771;
wire II15613;
wire g5588;
wire II10776;
wire II5654;
wire g8927;
wire g4799;
wire g8865;
wire g5809;
wire g3018;
wire g9161;
wire g7525;
wire II5398;
wire g6873;
wire g5783;
wire g7559;
wire II8957;
wire g7272;
wire II10078;
wire II10356;
wire g8650;
wire g7503;
wire g4892;
wire II15574;
wire g6146;
wire II13891;
wire II7437;
wire gbuf58;
wire g6772;
wire II10289;
wire g8811;
wire g4869;
wire g3694;
wire g7446;
wire II8974;
wire g7550;
wire II11103;
wire II13264;
wire II10017;
wire g9359;
wire II7421;
wire II15175;
wire II15675;
wire g5490;
wire g2674;
wire II10177;
wire g6882;
wire g9182;
wire II12433;
wire II7676;
wire g3798;
wire g5616;
wire II7329;
wire II8028;
wire II6775;
wire g4153;
wire g1753;
wire g4242;
wire g9356;
wire g1974;
wire g1778;
wire II13940;
wire g5000;
wire g8624;
wire g3843;
wire g9018;
wire g3866;
wire g3899;
wire g9291;
wire II10949;
wire g4822;
wire II6587;
wire g4867;
wire g9085;
wire g8838;
wire g8268;
wire g4908;
wire g8933;
wire II6341;
wire II11707;
wire II15065;
wire II6302;
wire g6833;
wire g8705;
wire g6349;
wire g8746;
wire g8731;
wire g2976;
wire g2149;
wire II15770;
wire II8949;
wire II11446;
wire II6348;
wire II15029;
wire g5596;
wire g9016;
wire g5564;
wire g4529;
wire g1771;
wire II10038;
wire g1806;
wire II6906;
wire g6411;
wire g8696;
wire II6039;
wire g2540;
wire II14406;
wire g3012;
wire g3801;
wire g3910;
wire g9346;
wire II13547;
wire g4224;
wire II5506;
wire g6138;
wire g6721;
wire g6813;
wire II8151;
wire g3856;
wire II8058;
wire II15032;
wire g4927;
wire g6905;
wire g3219;
wire g6671;
wire g2948;
wire g1863;
wire II8109;
wire g6344;
wire II11672;
wire g5798;
wire II14394;
wire II9153;
wire II7967;
wire II9651;
wire g3998;
wire g5188;
wire g4886;
wire II13731;
wire g5154;
wire II12349;
wire II13016;
wire g2700;
wire II14839;
wire g4124;
wire II8097;
wire II10819;
wire g6331;
wire g3975;
wire g1738;
wire g6104;
wire g4710;
wire II12015;
wire II5555;
wire g6328;
wire II11209;
wire g6053;
wire g6606;
wire II15184;
wire g7299;
wire g6043;
wire g5665;
wire g8907;
wire g4612;
wire g7262;
wire II6157;
wire g7693;
wire g6725;
wire II10855;
wire II5879;
wire II5889;
wire g9189;
wire g8956;
wire g5181;
wire g5317;
wire g8672;
wire II13244;
wire g4938;
wire II13722;
wire II7762;
wire g2361;
wire II12016;
wire g2162;
wire g8262;
wire g6354;
wire g7542;
wire g6072;
wire g2637;
wire II5475;
wire II7029;
wire g2829;
wire II5894;
wire II7533;
wire g6757;
wire g2770;
wire g4049;
wire II10335;
wire g4782;
wire II14834;
wire g4273;
wire II10253;
wire g5707;
wire II10552;
wire II11662;
wire g7597;
wire II9407;
wire g4166;
wire g5938;
wire II11569;
wire g7257;
wire g5088;
wire g7414;
wire g6270;
wire g5828;
wire g1865;
wire II5435;
wire II15971;
wire g4438;
wire II8209;
wire II8120;
wire II6042;
wire II12906;
wire II9416;
wire II15819;
wire g3925;
wire g2605;
wire g6997;
wire g7122;
wire II7769;
wire II14614;
wire g9241;
wire II14445;
wire g8870;
wire g6388;
wire g8920;
wire II15848;
wire g7716;
wire g1818;
wire g6581;
wire II14067;
wire g3919;
wire II6133;
wire g4557;
wire g6719;
wire g3952;
wire g7245;
wire g2661;
wire II15654;
wire g6375;
wire g4381;
wire g1792;
wire g7533;
wire II13284;
wire II10810;
wire II11302;
wire II14942;
wire g6845;
wire g2630;
wire g4112;
wire g8481;
wire II14767;
wire II5695;
wire II6223;
wire g6119;
wire g1714;
wire g3979;
wire g7181;
wire II8994;
wire g2783;
wire g2638;
wire g7759;
wire g4680;
wire II10225;
wire II15075;
wire II13927;
wire II9457;
wire g8947;
wire II15014;
wire II9261;
wire g8919;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g31 <= 0;
  else
    g31 <= g6302;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g30 <= 0;
  else
    g30 <= g6301;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g29 <= 0;
  else
    g29 <= g6300;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g28 <= 0;
  else
    g28 <= g6298;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g27 <= 0;
  else
    g27 <= g6297;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g26 <= 0;
  else
    g26 <= g6296;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g25 <= 0;
  else
    g25 <= g6295;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g24 <= 0;
  else
    g24 <= g6294;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g23 <= 0;
  else
    g23 <= g6293;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g22 <= 0;
  else
    g22 <= g6292;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g12 <= 0;
  else
    g12 <= g8662;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g11 <= 0;
  else
    g11 <= g6290;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g9 <= 0;
  else
    g9 <= g6288;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g8 <= 0;
  else
    g8 <= g9376;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g7 <= 0;
  else
    g7 <= g9375;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g6 <= 0;
  else
    g6 <= g9374;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g5 <= 0;
  else
    g5 <= g9373;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g4 <= 0;
  else
    g4 <= g9372;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g2 <= 0;
  else
    g2 <= g9361;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g3 <= 0;
  else
    g3 <= g9360;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g48 <= 0;
  else
    g48 <= g9362;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g21 <= 0;
  else
    g21 <= g6299;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g10 <= 0;
  else
    g10 <= g6291;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1 <= 0;
  else
    g1 <= g6289;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g47 <= 0;
  else
    g47 <= g9389;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g46 <= 0;
  else
    g46 <= g8955;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g45 <= 0;
  else
    g45 <= g6308;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g44 <= 0;
  else
    g44 <= g6307;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g42 <= 0;
  else
    g42 <= g6306;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g41 <= 0;
  else
    g41 <= g6305;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g37 <= 0;
  else
    g37 <= g6304;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g32 <= 0;
  else
    g32 <= g6303;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1207 <= 0;
  else
    g1207 <= g5173;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1211 <= 0;
  else
    g1211 <= g5174;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1214 <= 0;
  else
    g1214 <= g5736;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1217 <= 0;
  else
    g1217 <= g6377;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1220 <= 0;
  else
    g1220 <= g6378;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1223 <= 0;
  else
    g1223 <= g6379;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1224 <= 0;
  else
    g1224 <= g6857;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1225 <= 0;
  else
    g1225 <= g6858;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1226 <= 0;
  else
    g1226 <= g6859;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1227 <= 0;
  else
    g1227 <= g7108;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1228 <= 0;
  else
    g1228 <= g7109;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1229 <= 0;
  else
    g1229 <= g7110;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1230 <= 0;
  else
    g1230 <= g7300;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1240 <= 0;
  else
    g1240 <= g1235;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1236 <= 0;
  else
    g1236 <= gbuf1;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1231 <= 0;
  else
    g1231 <= gbuf2;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1244 <= 0;
  else
    g1244 <= g2659;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1245 <= 0;
  else
    g1245 <= gbuf3;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1243 <= 0;
  else
    g1243 <= g2660;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1272 <= 0;
  else
    g1272 <= g6383;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1276 <= 0;
  else
    g1276 <= g6384;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1280 <= 0;
  else
    g1280 <= g7112;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1284 <= 0;
  else
    g1284 <= g7301;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1288 <= 0;
  else
    g1288 <= g7527;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1292 <= 0;
  else
    g1292 <= g7302;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1300 <= 0;
  else
    g1300 <= g7303;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1296 <= 0;
  else
    g1296 <= g7304;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1253 <= 0;
  else
    g1253 <= g5741;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1308 <= 0;
  else
    g1308 <= g6385;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1309 <= 0;
  else
    g1309 <= gbuf4;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1310 <= 0;
  else
    g1310 <= gbuf5;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1311 <= 0;
  else
    g1311 <= gbuf6;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1312 <= 0;
  else
    g1312 <= gbuf7;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1304 <= 0;
  else
    g1304 <= gbuf8;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1307 <= 0;
  else
    g1307 <= g3858;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1330 <= 0;
  else
    g1330 <= g6862;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1333 <= 0;
  else
    g1333 <= g6863;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1336 <= 0;
  else
    g1336 <= g6864;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1339 <= 0;
  else
    g1339 <= g6865;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1342 <= 0;
  else
    g1342 <= g7119;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1345 <= 0;
  else
    g1345 <= g7528;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1348 <= 0;
  else
    g1348 <= g7529;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1351 <= 0;
  else
    g1351 <= g7530;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1354 <= 0;
  else
    g1354 <= g7768;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1357 <= 0;
  else
    g1357 <= g8675;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1360 <= 0;
  else
    g1360 <= g8676;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1190 <= 0;
  else
    g1190 <= g8677;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1191 <= 0;
  else
    g1191 <= g6373;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1192 <= 0;
  else
    g1192 <= gbuf9;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1193 <= 0;
  else
    g1193 <= gbuf10;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1194 <= 0;
  else
    g1194 <= gbuf11;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1195 <= 0;
  else
    g1195 <= g6374;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1196 <= 0;
  else
    g1196 <= gbuf12;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1197 <= 0;
  else
    g1197 <= gbuf13;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1198 <= 0;
  else
    g1198 <= gbuf14;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1199 <= 0;
  else
    g1199 <= g6375;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1200 <= 0;
  else
    g1200 <= gbuf15;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1201 <= 0;
  else
    g1201 <= gbuf16;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1202 <= 0;
  else
    g1202 <= gbuf17;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1203 <= 0;
  else
    g1203 <= g6376;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1204 <= 0;
  else
    g1204 <= gbuf18;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1205 <= 0;
  else
    g1205 <= gbuf19;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1206 <= 0;
  else
    g1206 <= gbuf20;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1252 <= 0;
  else
    g1252 <= g2661;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1250 <= 0;
  else
    g1250 <= g7111;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1251 <= 0;
  else
    g1251 <= g6860;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1247 <= 0;
  else
    g1247 <= g6380;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1254 <= 0;
  else
    g1254 <= g6381;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1266 <= 0;
  else
    g1266 <= g5739;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1260 <= 0;
  else
    g1260 <= g6382;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1257 <= 0;
  else
    g1257 <= g5738;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1263 <= 0;
  else
    g1263 <= g5737;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1267 <= 0;
  else
    g1267 <= g4656;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1268 <= 0;
  else
    g1268 <= g5175;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1269 <= 0;
  else
    g1269 <= g5740;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1271 <= 0;
  else
    g1271 <= g5176;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1270 <= 0;
  else
    g1270 <= gbuf21;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g172 <= 0;
  else
    g172 <= gbuf22;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1313 <= 0;
  else
    g1313 <= g5742;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1317 <= 0;
  else
    g1317 <= g5743;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1318 <= 0;
  else
    g1318 <= g6861;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1319 <= 0;
  else
    g1319 <= g7113;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1320 <= 0;
  else
    g1320 <= g7114;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1321 <= 0;
  else
    g1321 <= g7115;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1322 <= 0;
  else
    g1322 <= g7116;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1323 <= 0;
  else
    g1323 <= g7117;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1324 <= 0;
  else
    g1324 <= g7118;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1325 <= 0;
  else
    g1325 <= g7305;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1326 <= 0;
  else
    g1326 <= g7306;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1327 <= 0;
  else
    g1327 <= g7307;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1328 <= 0;
  else
    g1328 <= g7309;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g13 <= 0;
  else
    g13 <= g7308;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1329 <= 0;
  else
    g1329 <= g2663;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g20 <= 0;
  else
    g20 <= g6386;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1366 <= 0;
  else
    g1366 <= g6866;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1364 <= 0;
  else
    g1364 <= g6878;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1370 <= 0;
  else
    g1370 <= g6876;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1368 <= 0;
  else
    g1368 <= g6874;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1374 <= 0;
  else
    g1374 <= g6872;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1372 <= 0;
  else
    g1372 <= g6870;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1375 <= 0;
  else
    g1375 <= g6869;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1365 <= 0;
  else
    g1365 <= g6867;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1363 <= 0;
  else
    g1363 <= g6877;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1369 <= 0;
  else
    g1369 <= g6875;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1367 <= 0;
  else
    g1367 <= g6873;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1373 <= 0;
  else
    g1373 <= g6871;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1371 <= 0;
  else
    g1371 <= g6868;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1389 <= 0;
  else
    g1389 <= g4658;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1379 <= 0;
  else
    g1379 <= g6879;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1377 <= 0;
  else
    g1377 <= g6891;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1383 <= 0;
  else
    g1383 <= g6889;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1381 <= 0;
  else
    g1381 <= g6887;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1387 <= 0;
  else
    g1387 <= g6885;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1385 <= 0;
  else
    g1385 <= g6883;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1388 <= 0;
  else
    g1388 <= g6882;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1378 <= 0;
  else
    g1378 <= g6880;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1376 <= 0;
  else
    g1376 <= g6890;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1382 <= 0;
  else
    g1382 <= g6888;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1380 <= 0;
  else
    g1380 <= g6886;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1386 <= 0;
  else
    g1386 <= g6884;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1384 <= 0;
  else
    g1384 <= g6881;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1390 <= 0;
  else
    g1390 <= g4659;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1391 <= 0;
  else
    g1391 <= gbuf23;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1392 <= 0;
  else
    g1392 <= g6387;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1393 <= 0;
  else
    g1393 <= g2664;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1395 <= 0;
  else
    g1395 <= gbuf24;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1394 <= 0;
  else
    g1394 <= g6388;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1396 <= 0;
  else
    g1396 <= g4662;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1398 <= 0;
  else
    g1398 <= gbuf25;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1397 <= 0;
  else
    g1397 <= g6389;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1399 <= 0;
  else
    g1399 <= g3861;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1401 <= 0;
  else
    g1401 <= gbuf26;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1400 <= 0;
  else
    g1400 <= g6390;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1402 <= 0;
  else
    g1402 <= g6391;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1403 <= 0;
  else
    g1403 <= gbuf27;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1404 <= 0;
  else
    g1404 <= gbuf28;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g16 <= 0;
  else
    g16 <= gbuf29;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1189 <= 0;
  else
    g1189 <= g6392;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1412 <= 0;
  else
    g1412 <= g5745;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1415 <= 0;
  else
    g1415 <= g5180;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1409 <= 0;
  else
    g1409 <= g5178;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1416 <= 0;
  else
    g1416 <= g4665;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1421 <= 0;
  else
    g1421 <= g5179;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1405 <= 0;
  else
    g1405 <= g5744;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1408 <= 0;
  else
    g1408 <= g5177;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1429 <= 0;
  else
    g1429 <= g2671;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1428 <= 0;
  else
    g1428 <= g2672;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1431 <= 0;
  else
    g1431 <= g2673;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1430 <= 0;
  else
    g1430 <= g4666;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1424 <= 0;
  else
    g1424 <= g3862;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1524 <= 0;
  else
    g1524 <= g6393;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1513 <= 0;
  else
    g1513 <= gbuf30;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1486 <= 0;
  else
    g1486 <= g8226;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1481 <= 0;
  else
    g1481 <= g7769;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1489 <= 0;
  else
    g1489 <= g7770;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1494 <= 0;
  else
    g1494 <= g7771;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1499 <= 0;
  else
    g1499 <= g7772;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1504 <= 0;
  else
    g1504 <= g7773;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1509 <= 0;
  else
    g1509 <= g7774;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1514 <= 0;
  else
    g1514 <= g7775;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1519 <= 0;
  else
    g1519 <= g8227;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1462 <= 0;
  else
    g1462 <= g8678;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1467 <= 0;
  else
    g1467 <= g8875;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1472 <= 0;
  else
    g1472 <= g8960;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1477 <= 0;
  else
    g1477 <= g9036;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g727 <= 0;
  else
    g727 <= g8228;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1532 <= 0;
  else
    g1532 <= g7781;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1528 <= 0;
  else
    g1528 <= g7776;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1537 <= 0;
  else
    g1537 <= g7777;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1541 <= 0;
  else
    g1541 <= g7778;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1545 <= 0;
  else
    g1545 <= g7779;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1549 <= 0;
  else
    g1549 <= g7780;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1435 <= 0;
  else
    g1435 <= g5181;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1439 <= 0;
  else
    g1439 <= g5182;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1432 <= 0;
  else
    g1432 <= g5183;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1443 <= 0;
  else
    g1443 <= g4667;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g33 <= 0;
  else
    g33 <= g5184;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g38 <= 0;
  else
    g38 <= g5746;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1461 <= 0;
  else
    g1461 <= g4669;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1444 <= 0;
  else
    g1444 <= g5185;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1450 <= 0;
  else
    g1450 <= g5186;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1454 <= 0;
  else
    g1454 <= g5187;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1459 <= 0;
  else
    g1459 <= g3863;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1460 <= 0;
  else
    g1460 <= g4668;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g979 <= 0;
  else
    g979 <= g7104;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g966 <= 0;
  else
    g966 <= g8223;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g969 <= 0;
  else
    g969 <= gbuf31;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g963 <= 0;
  else
    g963 <= g7764;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g970 <= 0;
  else
    g970 <= gbuf32;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g971 <= 0;
  else
    g971 <= g5171;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g972 <= 0;
  else
    g972 <= g2653;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g973 <= 0;
  else
    g973 <= g8672;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g976 <= 0;
  else
    g976 <= g8864;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g984 <= 0;
  else
    g984 <= g9133;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g985 <= 0;
  else
    g985 <= g7515;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g990 <= 0;
  else
    g990 <= g7516;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g995 <= 0;
  else
    g995 <= g7517;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1004 <= 0;
  else
    g1004 <= g7105;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1005 <= 0;
  else
    g1005 <= gbuf33;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g998 <= 0;
  else
    g998 <= gbuf34;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g999 <= 0;
  else
    g999 <= g8865;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1007 <= 0;
  else
    g1007 <= g8867;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1012 <= 0;
  else
    g1012 <= g6851;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1014 <= 0;
  else
    g1014 <= gbuf35;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1013 <= 0;
  else
    g1013 <= gbuf36;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1029 <= 0;
  else
    g1029 <= g2654;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1018 <= 0;
  else
    g1018 <= g8869;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1021 <= 0;
  else
    g1021 <= g8870;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1025 <= 0;
  else
    g1025 <= g8871;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1033 <= 0;
  else
    g1033 <= g9034;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1034 <= 0;
  else
    g1034 <= g8957;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1030 <= 0;
  else
    g1030 <= g7518;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1081 <= 0;
  else
    g1081 <= g6852;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1156 <= 0;
  else
    g1156 <= gbuf37;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1157 <= 0;
  else
    g1157 <= gbuf38;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1159 <= 0;
  else
    g1159 <= gbuf39;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1158 <= 0;
  else
    g1158 <= gbuf40;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1084 <= 0;
  else
    g1084 <= g7106;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1146 <= 0;
  else
    g1146 <= g1612;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1147 <= 0;
  else
    g1147 <= gbuf41;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1148 <= 0;
  else
    g1148 <= gbuf42;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1087 <= 0;
  else
    g1087 <= g6853;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1098 <= 0;
  else
    g1098 <= g6854;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1102 <= 0;
  else
    g1102 <= g6855;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1106 <= 0;
  else
    g1106 <= g7107;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1110 <= 0;
  else
    g1110 <= g7299;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1114 <= 0;
  else
    g1114 <= g7521;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1118 <= 0;
  else
    g1118 <= g7766;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1122 <= 0;
  else
    g1122 <= g8225;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1126 <= 0;
  else
    g1126 <= g8674;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1142 <= 0;
  else
    g1142 <= g8874;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1173 <= 0;
  else
    g1173 <= g7526;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1170 <= 0;
  else
    g1170 <= gbuf43;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1167 <= 0;
  else
    g1167 <= gbuf44;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1166 <= 0;
  else
    g1166 <= gbuf45;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1077 <= 0;
  else
    g1077 <= g7767;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1153 <= 0;
  else
    g1153 <= g6856;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1154 <= 0;
  else
    g1154 <= gbuf46;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1155 <= 0;
  else
    g1155 <= gbuf47;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1185 <= 0;
  else
    g1185 <= gbuf48;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1097 <= 0;
  else
    g1097 <= gbuf49;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1092 <= 0;
  else
    g1092 <= g7520;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1130 <= 0;
  else
    g1130 <= g7522;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1134 <= 0;
  else
    g1134 <= g7523;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1138 <= 0;
  else
    g1138 <= g7524;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1149 <= 0;
  else
    g1149 <= g7525;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1037 <= 0;
  else
    g1037 <= g7519;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1041 <= 0;
  else
    g1041 <= g7765;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1045 <= 0;
  else
    g1045 <= g8224;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1049 <= 0;
  else
    g1049 <= g8673;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1053 <= 0;
  else
    g1053 <= g8873;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1057 <= 0;
  else
    g1057 <= g8959;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1061 <= 0;
  else
    g1061 <= g9035;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1065 <= 0;
  else
    g1065 <= g9117;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1069 <= 0;
  else
    g1069 <= g9134;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1073 <= 0;
  else
    g1073 <= g9145;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1163 <= 0;
  else
    g1163 <= g2655;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1160 <= 0;
  else
    g1160 <= gbuf50;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1182 <= 0;
  else
    g1182 <= gbuf51;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1186 <= 0;
  else
    g1186 <= gbuf52;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1179 <= 0;
  else
    g1179 <= gbuf53;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g1176 <= 0;
  else
    g1176 <= g5172;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g68 <= 0;
  else
    g68 <= g6774;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g71 <= 0;
  else
    g71 <= g6775;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g74 <= 0;
  else
    g74 <= g6776;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g77 <= 0;
  else
    g77 <= g6777;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g80 <= 0;
  else
    g80 <= g6778;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g83 <= 0;
  else
    g83 <= g6779;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g86 <= 0;
  else
    g86 <= g6780;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g52 <= 0;
  else
    g52 <= g6781;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g55 <= 0;
  else
    g55 <= g7733;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g62 <= 0;
  else
    g62 <= g7509;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g58 <= 0;
  else
    g58 <= g7734;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g65 <= 0;
  else
    g65 <= g4598;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g199 <= 0;
  else
    g199 <= g3832;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g200 <= 0;
  else
    g200 <= gbuf54;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g201 <= 0;
  else
    g201 <= gbuf55;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g190 <= 0;
  else
    g190 <= gbuf56;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g195 <= 0;
  else
    g195 <= g3831;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g196 <= 0;
  else
    g196 <= g5731;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g179 <= 0;
  else
    g179 <= g5159;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g186 <= 0;
  else
    g186 <= g3830;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g187 <= 0;
  else
    g187 <= g5730;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g180 <= 0;
  else
    g180 <= g5158;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g205 <= 0;
  else
    g205 <= g3835;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g202 <= 0;
  else
    g202 <= g5732;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g181 <= 0;
  else
    g181 <= g5160;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g210 <= 0;
  else
    g210 <= g3834;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g207 <= 0;
  else
    g207 <= g5733;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g182 <= 0;
  else
    g182 <= g5161;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g146 <= 0;
  else
    g146 <= g7735;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g173 <= 0;
  else
    g173 <= g7736;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g150 <= 0;
  else
    g150 <= g7738;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g174 <= 0;
  else
    g174 <= g7737;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g154 <= 0;
  else
    g154 <= g7739;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g158 <= 0;
  else
    g158 <= g7740;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g162 <= 0;
  else
    g162 <= g7741;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g168 <= 0;
  else
    g168 <= g7742;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g183 <= 0;
  else
    g183 <= g6309;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g184 <= 0;
  else
    g184 <= g6310;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g185 <= 0;
  else
    g185 <= g4599;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g92 <= 0;
  else
    g92 <= g6794;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g89 <= 0;
  else
    g89 <= gbuf57;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g93 <= 0;
  else
    g93 <= g5145;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g94 <= 0;
  else
    g94 <= g6782;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g95 <= 0;
  else
    g95 <= gbuf58;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g98 <= 0;
  else
    g98 <= g5146;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g99 <= 0;
  else
    g99 <= g6783;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g100 <= 0;
  else
    g100 <= gbuf59;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g103 <= 0;
  else
    g103 <= g5157;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g104 <= 0;
  else
    g104 <= g6784;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g105 <= 0;
  else
    g105 <= gbuf60;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g108 <= 0;
  else
    g108 <= g5147;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g109 <= 0;
  else
    g109 <= g6785;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g110 <= 0;
  else
    g110 <= gbuf61;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g113 <= 0;
  else
    g113 <= g5148;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g114 <= 0;
  else
    g114 <= g6786;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g117 <= 0;
  else
    g117 <= g5153;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g118 <= 0;
  else
    g118 <= g6787;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g121 <= 0;
  else
    g121 <= g5154;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g122 <= 0;
  else
    g122 <= g6788;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g125 <= 0;
  else
    g125 <= g5155;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g126 <= 0;
  else
    g126 <= g6789;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g129 <= 0;
  else
    g129 <= g5156;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g130 <= 0;
  else
    g130 <= g6790;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g133 <= 0;
  else
    g133 <= g5149;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g134 <= 0;
  else
    g134 <= g6791;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g137 <= 0;
  else
    g137 <= g5150;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g138 <= 0;
  else
    g138 <= g6792;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g141 <= 0;
  else
    g141 <= g5151;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g142 <= 0;
  else
    g142 <= g6793;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g145 <= 0;
  else
    g145 <= g5152;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g287 <= 0;
  else
    g287 <= g3836;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g290 <= 0;
  else
    g290 <= gbuf62;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g255 <= 0;
  else
    g255 <= g9087;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g258 <= 0;
  else
    g258 <= g9088;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g261 <= 0;
  else
    g261 <= g9089;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g264 <= 0;
  else
    g264 <= g9090;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g267 <= 0;
  else
    g267 <= g9091;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g270 <= 0;
  else
    g270 <= g9092;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g281 <= 0;
  else
    g281 <= g9085;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g284 <= 0;
  else
    g284 <= g9086;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g211 <= 0;
  else
    g211 <= g4600;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g216 <= 0;
  else
    g216 <= g6311;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g212 <= 0;
  else
    g212 <= g4601;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g219 <= 0;
  else
    g219 <= g6312;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g213 <= 0;
  else
    g213 <= g4602;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g222 <= 0;
  else
    g222 <= g6313;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g214 <= 0;
  else
    g214 <= g4603;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g225 <= 0;
  else
    g225 <= g6314;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g215 <= 0;
  else
    g215 <= g4604;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g228 <= 0;
  else
    g228 <= g6315;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g231 <= 0;
  else
    g231 <= g4605;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g237 <= 0;
  else
    g237 <= g6316;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g232 <= 0;
  else
    g232 <= g4606;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g240 <= 0;
  else
    g240 <= g6317;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g233 <= 0;
  else
    g233 <= g4607;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g243 <= 0;
  else
    g243 <= g6318;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g234 <= 0;
  else
    g234 <= g4608;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g246 <= 0;
  else
    g246 <= g6319;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g235 <= 0;
  else
    g235 <= g4609;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g249 <= 0;
  else
    g249 <= g6320;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g236 <= 0;
  else
    g236 <= g4610;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g252 <= 0;
  else
    g252 <= g6321;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g273 <= 0;
  else
    g273 <= g4611;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g275 <= 0;
  else
    g275 <= g6322;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g274 <= 0;
  else
    g274 <= g4612;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g278 <= 0;
  else
    g278 <= g6323;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g368 <= 0;
  else
    g368 <= g3838;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g371 <= 0;
  else
    g371 <= gbuf63;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g336 <= 0;
  else
    g336 <= g9095;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g339 <= 0;
  else
    g339 <= g9096;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g342 <= 0;
  else
    g342 <= g9097;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g345 <= 0;
  else
    g345 <= g9098;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g348 <= 0;
  else
    g348 <= g9099;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g351 <= 0;
  else
    g351 <= g9100;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g362 <= 0;
  else
    g362 <= g9093;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g365 <= 0;
  else
    g365 <= g9094;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g292 <= 0;
  else
    g292 <= g4613;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g297 <= 0;
  else
    g297 <= g6324;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g293 <= 0;
  else
    g293 <= g4614;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g300 <= 0;
  else
    g300 <= g6325;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g294 <= 0;
  else
    g294 <= g4615;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g303 <= 0;
  else
    g303 <= g6326;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g295 <= 0;
  else
    g295 <= g4616;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g306 <= 0;
  else
    g306 <= g6327;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g296 <= 0;
  else
    g296 <= g4617;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g309 <= 0;
  else
    g309 <= g6328;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g312 <= 0;
  else
    g312 <= g4618;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g318 <= 0;
  else
    g318 <= g6329;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g313 <= 0;
  else
    g313 <= g4619;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g321 <= 0;
  else
    g321 <= g6330;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g314 <= 0;
  else
    g314 <= g4620;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g324 <= 0;
  else
    g324 <= g6331;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g315 <= 0;
  else
    g315 <= g4621;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g327 <= 0;
  else
    g327 <= g6332;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g316 <= 0;
  else
    g316 <= g4622;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g330 <= 0;
  else
    g330 <= g6333;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g317 <= 0;
  else
    g317 <= g4623;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g333 <= 0;
  else
    g333 <= g6334;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g354 <= 0;
  else
    g354 <= g4624;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g356 <= 0;
  else
    g356 <= g6335;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g355 <= 0;
  else
    g355 <= g4625;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g359 <= 0;
  else
    g359 <= g6336;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g449 <= 0;
  else
    g449 <= g3840;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g452 <= 0;
  else
    g452 <= gbuf64;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g417 <= 0;
  else
    g417 <= g9103;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g420 <= 0;
  else
    g420 <= g9104;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g423 <= 0;
  else
    g423 <= g9105;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g426 <= 0;
  else
    g426 <= g9106;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g429 <= 0;
  else
    g429 <= g9107;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g432 <= 0;
  else
    g432 <= g9108;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g443 <= 0;
  else
    g443 <= g9101;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g446 <= 0;
  else
    g446 <= g9102;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g373 <= 0;
  else
    g373 <= g4626;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g378 <= 0;
  else
    g378 <= g6337;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g374 <= 0;
  else
    g374 <= g4627;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g381 <= 0;
  else
    g381 <= g6338;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g375 <= 0;
  else
    g375 <= g4628;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g384 <= 0;
  else
    g384 <= g6339;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g376 <= 0;
  else
    g376 <= g4629;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g387 <= 0;
  else
    g387 <= g6340;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g377 <= 0;
  else
    g377 <= g4630;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g390 <= 0;
  else
    g390 <= g6341;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g393 <= 0;
  else
    g393 <= g4631;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g399 <= 0;
  else
    g399 <= g6342;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g394 <= 0;
  else
    g394 <= g4632;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g402 <= 0;
  else
    g402 <= g6343;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g395 <= 0;
  else
    g395 <= g4633;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g405 <= 0;
  else
    g405 <= g6344;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g396 <= 0;
  else
    g396 <= g4634;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g408 <= 0;
  else
    g408 <= g6345;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g397 <= 0;
  else
    g397 <= g4635;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g411 <= 0;
  else
    g411 <= g6346;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g398 <= 0;
  else
    g398 <= g4636;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g414 <= 0;
  else
    g414 <= g6347;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g435 <= 0;
  else
    g435 <= g4637;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g437 <= 0;
  else
    g437 <= g6348;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g436 <= 0;
  else
    g436 <= g4638;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g440 <= 0;
  else
    g440 <= g6349;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g530 <= 0;
  else
    g530 <= g3842;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g533 <= 0;
  else
    g533 <= gbuf65;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g498 <= 0;
  else
    g498 <= g9111;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g501 <= 0;
  else
    g501 <= g9112;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g504 <= 0;
  else
    g504 <= g9113;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g507 <= 0;
  else
    g507 <= g9114;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g510 <= 0;
  else
    g510 <= g9115;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g513 <= 0;
  else
    g513 <= g9116;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g524 <= 0;
  else
    g524 <= g9109;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g527 <= 0;
  else
    g527 <= g9110;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g454 <= 0;
  else
    g454 <= g4639;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g459 <= 0;
  else
    g459 <= g6350;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g455 <= 0;
  else
    g455 <= g4640;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g462 <= 0;
  else
    g462 <= g6351;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g456 <= 0;
  else
    g456 <= g4641;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g465 <= 0;
  else
    g465 <= g6352;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g457 <= 0;
  else
    g457 <= g4642;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g468 <= 0;
  else
    g468 <= g6353;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g458 <= 0;
  else
    g458 <= g4643;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g471 <= 0;
  else
    g471 <= g6354;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g474 <= 0;
  else
    g474 <= g4644;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g480 <= 0;
  else
    g480 <= g6355;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g475 <= 0;
  else
    g475 <= g4645;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g483 <= 0;
  else
    g483 <= g6356;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g476 <= 0;
  else
    g476 <= g4646;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g486 <= 0;
  else
    g486 <= g6357;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g477 <= 0;
  else
    g477 <= g4647;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g489 <= 0;
  else
    g489 <= g6358;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g478 <= 0;
  else
    g478 <= g4648;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g492 <= 0;
  else
    g492 <= g6359;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g479 <= 0;
  else
    g479 <= g4649;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g495 <= 0;
  else
    g495 <= g6360;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g516 <= 0;
  else
    g516 <= g4650;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g518 <= 0;
  else
    g518 <= g6361;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g517 <= 0;
  else
    g517 <= g4651;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g521 <= 0;
  else
    g521 <= g6362;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g535 <= 0;
  else
    g535 <= g3844;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g536 <= 0;
  else
    g536 <= g6363;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g539 <= 0;
  else
    g539 <= g3845;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g540 <= 0;
  else
    g540 <= g6364;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g543 <= 0;
  else
    g543 <= g3846;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g544 <= 0;
  else
    g544 <= g6365;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g547 <= 0;
  else
    g547 <= g9026;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g550 <= 0;
  else
    g550 <= g9027;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g553 <= 0;
  else
    g553 <= g9028;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g556 <= 0;
  else
    g556 <= g3847;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g557 <= 0;
  else
    g557 <= g6366;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g566 <= 0;
  else
    g566 <= g3848;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g567 <= 0;
  else
    g567 <= g6367;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g579 <= 0;
  else
    g579 <= g3850;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g580 <= 0;
  else
    g580 <= g6368;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g583 <= 0;
  else
    g583 <= g3851;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g584 <= 0;
  else
    g584 <= g6369;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g587 <= 0;
  else
    g587 <= g3852;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g560 <= 0;
  else
    g560 <= g6370;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g563 <= 0;
  else
    g563 <= g9029;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g570 <= 0;
  else
    g570 <= g9030;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g588 <= 0;
  else
    g588 <= g9031;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g591 <= 0;
  else
    g591 <= g9032;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g573 <= 0;
  else
    g573 <= g9033;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g576 <= 0;
  else
    g576 <= g3849;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g595 <= 0;
  else
    g595 <= gbuf66;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g596 <= 0;
  else
    g596 <= g6795;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g597 <= 0;
  else
    g597 <= g6796;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g598 <= 0;
  else
    g598 <= g6797;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g599 <= 0;
  else
    g599 <= g6798;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g600 <= 0;
  else
    g600 <= g6807;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g601 <= 0;
  else
    g601 <= g6799;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g602 <= 0;
  else
    g602 <= g6800;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g603 <= 0;
  else
    g603 <= g6801;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g604 <= 0;
  else
    g604 <= g6802;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g605 <= 0;
  else
    g605 <= g6803;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g606 <= 0;
  else
    g606 <= g6804;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g607 <= 0;
  else
    g607 <= g6805;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g608 <= 0;
  else
    g608 <= g6806;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g609 <= 0;
  else
    g609 <= g6808;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g610 <= 0;
  else
    g610 <= g6809;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g611 <= 0;
  else
    g611 <= g6810;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g612 <= 0;
  else
    g612 <= g6811;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g613 <= 0;
  else
    g613 <= g6820;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g614 <= 0;
  else
    g614 <= g6812;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g615 <= 0;
  else
    g615 <= g6813;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g616 <= 0;
  else
    g616 <= g6814;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g617 <= 0;
  else
    g617 <= g6815;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g618 <= 0;
  else
    g618 <= g6816;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g619 <= 0;
  else
    g619 <= g6817;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g620 <= 0;
  else
    g620 <= g6818;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g621 <= 0;
  else
    g621 <= g6819;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g622 <= 0;
  else
    g622 <= g6821;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g623 <= 0;
  else
    g623 <= g6822;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g624 <= 0;
  else
    g624 <= g6831;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g625 <= 0;
  else
    g625 <= g6823;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g626 <= 0;
  else
    g626 <= g6824;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g627 <= 0;
  else
    g627 <= g6825;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g628 <= 0;
  else
    g628 <= g6826;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g629 <= 0;
  else
    g629 <= g6827;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g630 <= 0;
  else
    g630 <= g6828;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g631 <= 0;
  else
    g631 <= g6829;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g632 <= 0;
  else
    g632 <= g6830;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g646 <= 0;
  else
    g646 <= g4652;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g652 <= 0;
  else
    g652 <= gbuf67;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g661 <= 0;
  else
    g661 <= g7743;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g665 <= 0;
  else
    g665 <= g7744;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g669 <= 0;
  else
    g669 <= g7745;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g673 <= 0;
  else
    g673 <= g7746;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g677 <= 0;
  else
    g677 <= g7747;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g681 <= 0;
  else
    g681 <= g7748;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g685 <= 0;
  else
    g685 <= g7749;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g706 <= 0;
  else
    g706 <= g7750;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g710 <= 0;
  else
    g710 <= g7751;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g714 <= 0;
  else
    g714 <= g7752;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g718 <= 0;
  else
    g718 <= g7753;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g734 <= 0;
  else
    g734 <= g7755;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g730 <= 0;
  else
    g730 <= g7754;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g689 <= 0;
  else
    g689 <= g6371;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g758 <= 0;
  else
    g758 <= g6840;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g759 <= 0;
  else
    g759 <= g6832;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g760 <= 0;
  else
    g760 <= g6833;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g761 <= 0;
  else
    g761 <= g6834;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g762 <= 0;
  else
    g762 <= g6835;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g763 <= 0;
  else
    g763 <= g6836;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g764 <= 0;
  else
    g764 <= g6837;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g765 <= 0;
  else
    g765 <= g6838;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g766 <= 0;
  else
    g766 <= g6839;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g767 <= 0;
  else
    g767 <= g6841;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g768 <= 0;
  else
    g768 <= g6842;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g769 <= 0;
  else
    g769 <= g6843;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g770 <= 0;
  else
    g770 <= g6844;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g771 <= 0;
  else
    g771 <= g6845;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g772 <= 0;
  else
    g772 <= g6846;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g773 <= 0;
  else
    g773 <= g6847;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g774 <= 0;
  else
    g774 <= g6848;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g795 <= 0;
  else
    g795 <= g3854;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g792 <= 0;
  else
    g792 <= g5162;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g782 <= 0;
  else
    g782 <= g5734;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g799 <= 0;
  else
    g799 <= g7756;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g803 <= 0;
  else
    g803 <= g7757;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g806 <= 0;
  else
    g806 <= g7510;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g809 <= 0;
  else
    g809 <= g7511;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g812 <= 0;
  else
    g812 <= g7758;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g775 <= 0;
  else
    g775 <= g7759;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g778 <= 0;
  else
    g778 <= g7296;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g815 <= 0;
  else
    g815 <= g7760;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g819 <= 0;
  else
    g819 <= g7761;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g822 <= 0;
  else
    g822 <= g7512;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g825 <= 0;
  else
    g825 <= g7513;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g828 <= 0;
  else
    g828 <= g7762;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g786 <= 0;
  else
    g786 <= g7763;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g789 <= 0;
  else
    g789 <= g7297;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g955 <= 0;
  else
    g955 <= g3857;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g959 <= 0;
  else
    g959 <= g5169;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g945 <= 0;
  else
    g945 <= g5170;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g948 <= 0;
  else
    g948 <= g8664;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g949 <= 0;
  else
    g949 <= g8665;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g950 <= 0;
  else
    g950 <= g8666;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g951 <= 0;
  else
    g951 <= g8667;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g952 <= 0;
  else
    g952 <= g8668;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g953 <= 0;
  else
    g953 <= g8669;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g954 <= 0;
  else
    g954 <= g8670;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g943 <= 0;
  else
    g943 <= g8671;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g936 <= 0;
  else
    g936 <= g5168;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g940 <= 0;
  else
    g940 <= g5735;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g942 <= 0;
  else
    g942 <= g2652;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g944 <= 0;
  else
    g944 <= g6372;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g855 <= 0;
  else
    g855 <= g8220;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g859 <= 0;
  else
    g859 <= g8221;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g863 <= 0;
  else
    g863 <= g8222;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g831 <= 0;
  else
    g831 <= g2651;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g834 <= 0;
  else
    g834 <= g2650;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g837 <= 0;
  else
    g837 <= g2649;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g840 <= 0;
  else
    g840 <= g2648;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g843 <= 0;
  else
    g843 <= g2647;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g846 <= 0;
  else
    g846 <= g2646;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g849 <= 0;
  else
    g849 <= g2645;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g852 <= 0;
  else
    g852 <= g2644;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g890 <= 0;
  else
    g890 <= g7102;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g878 <= 0;
  else
    g878 <= gbuf68;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g926 <= 0;
  else
    g926 <= gbuf69;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g875 <= 0;
  else
    g875 <= g5165;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g866 <= 0;
  else
    g866 <= g5163;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g929 <= 0;
  else
    g929 <= g3856;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g933 <= 0;
  else
    g933 <= g5166;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g871 <= 0;
  else
    g871 <= g5167;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g874 <= 0;
  else
    g874 <= g4654;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g891 <= 0;
  else
    g891 <= g3855;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g896 <= 0;
  else
    g896 <= gbuf70;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g901 <= 0;
  else
    g901 <= gbuf71;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g906 <= 0;
  else
    g906 <= gbuf72;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g911 <= 0;
  else
    g911 <= gbuf73;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g916 <= 0;
  else
    g916 <= gbuf74;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g921 <= 0;
  else
    g921 <= gbuf75;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g883 <= 0;
  else
    g883 <= gbuf76;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g887 <= 0;
  else
    g887 <= g7099;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g888 <= 0;
  else
    g888 <= g7100;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g889 <= 0;
  else
    g889 <= g7101;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g741 <= 0;
  else
    g741 <= g9386;
always @(posedge blif_clk_net or posedge blif_reset_net)
  if(blif_reset_net == 1)
    g746 <= 0;
  else
    g746 <= g8956;
assign g3491 = ((~g1800));
assign g3610 = ((~g2424));
assign II7683 = ((~g2573));
assign g4355 = (g390&g3160);
assign II11158 = ((~g3052))|((~II11156));
assign g7026 = (g4186)|(g6554);
assign g3951 = ((~II7648));
assign g8902 = (g8844)|(g8654);
assign g6579 = (g6098)|(g1975);
assign II13463 = ((~g7264));
assign II10924 = ((~g5525))|((~II10923));
assign II6524 = ((~g1102))|((~II6522));
assign II6959 = ((~g1558));
assign g4610 = ((~II8745));
assign g7168 = ((~II13072));
assign g3892 = ((~g3131));
assign g4396 = (g459&g3192);
assign g2386 = (g1130&g1092);
assign II10773 = ((~g5708));
assign g6365 = ((~II11422));
assign II12128 = ((~g5897));
assign II8512 = ((~g2807))|((~II8510));
assign II15147 = (g8483)|(g8464)|(g8514);
assign II15405 = ((~g8902));
assign g3783 = ((~II7255));
assign g4111 = ((~II7944));
assign g3603 = ((~g2092));
assign g2887 = ((~g2241));
assign g6136 = ((~II10773));
assign II6501 = ((~g1537))|((~II6499));
assign g8995 = (g8935)|(g8837);
assign II14712 = ((~g8059));
assign II6051 = ((~g440));
assign g7555 = ((~II13843));
assign g3885 = ((~g3310)&(~g3466));
assign II15943 = ((~g9214));
assign g6034 = ((~II10639));
assign g8090 = (g843&g7658);
assign g7658 = (g7367&g4150);
assign II8413 = (g3316&g3287&g3264&g1987);
assign II14260 = ((~g7717));
assign II12226 = ((~g6636));
assign II14227 = ((~g7552));
assign II16103 = ((~g9339));
assign g6542 = ((~II11718));
assign g8278 = (g4589&g7993);
assign g6426 = ((~II11559));
assign g7763 = ((~II14160));
assign g9023 = (g8888&g5317);
assign g8946 = (g4556&g8786);
assign g4556 = ((~g2895));
assign II10849 = ((~g2595))|((~II10847));
assign g8932 = (g3868&g8762);
assign II8486 = ((~g2824));
assign g5729 = ((~g5144));
assign II10315 = ((~g1041))|((~II10313));
assign II15400 = (g8736)|(g8748)|(g8740);
assign g2368 = (II6208)|(II6209);
assign g4311 = ((~II8282));
assign g7506 = ((~II13698));
assign g9338 = (g9258)|(g9334);
assign g4960 = ((~g4259));
assign g6045 = (g1472&g5591);
assign g3221 = ((~II6877))|((~II6878));
assign g7246 = ((~II13196));
assign g5788 = ((~II10409));
assign g2039 = ((~g1228));
assign g6293 = ((~II11206));
assign g3313 = (g2334&g2316&g2298);
assign g6577 = (g6142&g4160);
assign g5711 = (g4959)|(g4352);
assign II14163 = ((~g7533));
assign g7100 = ((~II12888));
assign g6201 = ((~II10946));
assign g5845 = ((~II10548));
assign g5748 = ((~II10306))|((~II10307));
assign g7440 = ((~II13577));
assign II5689 = ((~g906));
assign II12771 = ((~g6735));
assign g5805 = ((~II10448));
assign g5216 = (g5062)|(g4391);
assign g7352 = ((~II13472));
assign g2662 = ((~II6457));
assign g7600 = (g7460&g3466);
assign g6629 = (g6023&g4841);
assign g5025 = ((~II9363));
assign II15871 = ((~g9184));
assign II11603 = (g6193)|(g6197)|(g6175);
assign g8801 = ((~g8635)&(~g3790));
assign g7314 = ((~g7180)&(~g6972));
assign g7756 = ((~II14139));
assign g5119 = (g543&g4027);
assign g5462 = ((~g4886));
assign g5099 = ((~g4477));
assign g2282 = ((~g1400));
assign g5607 = ((~g4938));
assign II10224 = ((~g2522))|((~II10223));
assign II9301 = ((~g4295));
assign II14941 = (g8275)|(g8323)|(g8459)|(g8380);
assign II10039 = ((~g4893))|((~II10038));
assign g4097 = (g2624&g2614);
assign g4342 = (g228&g3097);
assign g7252 = (g3591&g6977);
assign g4623 = ((~II8784));
assign II10856 = ((~g2584))|((~II10854));
assign g5445 = ((~g5059));
assign g3864 = ((~g2943));
assign g7115 = ((~II12933));
assign II13214 = ((~g7065))|((~II13213));
assign g8862 = ((~g8493)&(~g8239)&(~II15172));
assign II8052 = (g2162&g2149&g2137&g2106);
assign g8904 = (g8090)|(g8080)|(g8706);
assign g8361 = (g426&g7920);
assign II7994 = (g3430&g3398&g3359&g3341);
assign g8641 = ((~g6559)&(~g162)&(~g7784)&(~g3591));
assign g7367 = ((~II13515));
assign II9929 = ((~g5052));
assign g3761 = ((~g1772));
assign II13622 = ((~g7279));
assign II12915 = ((~g7000));
assign g5680 = ((~g5101));
assign g4835 = ((~II9195))|((~II9196));
assign g8938 = (g3878&g8771);
assign g7030 = (g6705&g5723);
assign g8976 = (g8903&g6588);
assign II5942 = ((~g300));
assign g5589 = ((~II10061))|((~II10062));
assign II16036 = ((~g9282));
assign g4197 = ((~g3591));
assign gbuf10 = (g1192);
assign II8166 = ((~g3231))|((~II8164));
assign g9034 = ((~II15516));
assign g4276 = (g2216&g2618);
assign g1794 = ((~II5646));
assign g6419 = (g162&g6032);
assign g2651 = ((~II6437));
assign g7696 = (g7367&g4469);
assign II7344 = ((~g2964));
assign g8319 = (g255&g7838);
assign II11305 = ((~g5807));
assign g8941 = (g3882&g8776);
assign II12041 = ((~g5897));
assign g7521 = ((~II13743));
assign g6358 = ((~II11401));
assign g6022 = (g5595&g2424);
assign II10250 = ((~g5268));
assign g291 = ((~II5356));
assign g8892 = (g8681&g4969);
assign g8728 = (g3815&g8464);
assign g7019 = ((~II12771));
assign II10587 = ((~g5439));
assign II11069 = ((~g5671));
assign g4009 = ((~II7758));
assign II14786 = ((~g8606));
assign g9184 = ((~II15830));
assign II11440 = ((~g6009));
assign g4236 = (g3260&g3221);
assign g8403 = (g639&g7793);
assign II6208 = (g891)|(g896)|(g901)|(g906);
assign II14139 = ((~g7548));
assign g6222 = ((~g5654));
assign II13649 = ((~g7281));
assign II7132 = ((~g2554));
assign g6872 = ((~II12487));
assign g2403 = ((~g1176));
assign g2298 = ((~II6072));
assign g5765 = (g1695&g5428);
assign II11150 = ((~g5473))|((~II11149));
assign II10690 = ((~g5538));
assign g3188 = (g2298&g2316);
assign II16161 = ((~g9363));
assign g1736 = ((~II5577));
assign g8717 = (g2764&g8421);
assign g5874 = ((~II10565));
assign g1589 = ((~g746));
assign gbuf75 = (g916);
assign gbuf71 = (g896);
assign g6890 = ((~II12541));
assign g2680 = ((~g1665));
assign gbuf3 = (g1244);
assign II7512 = ((~g1711))|((~II7510));
assign II12355 = ((~g6756));
assign g4956 = (g295&g3892);
assign II6214 = ((~g7));
assign II8437 = (g3316&g3287&g3264&g1987);
assign g6958 = ((~II12675));
assign II5957 = ((~g110));
assign II16040 = ((~g9285));
assign II15187 = ((~g8682));
assign II11894 = ((~g5956));
assign g7604 = (g7456&g3466);
assign II8529 = (g3316&g2057&g3264&g3238);
assign g3922 = ((~II7561));
assign II9804 = ((~g5113));
assign g4454 = (g544&g2845);
assign g1822 = ((~g761));
assign g6847 = ((~II12412));
assign g6818 = ((~II12325));
assign g5491 = ((~g4918));
assign g8645 = (g550&g8094);
assign g4883 = (g3746&g3723&g4288);
assign g8780 = ((~g8524));
assign g4830 = (g4288&g3723);
assign II7616 = ((~g3008))|((~g1721));
assign g6015 = ((~II10617));
assign II12877 = ((~g6700));
assign g7136 = (g4057&g6953);
assign g7192 = (g7026&g3526);
assign g8749 = (g2989&g8493);
assign g5726 = ((~II10243));
assign g6853 = ((~II12430));
assign g4150 = (II8019&II8020);
assign g2177 = ((~g1322));
assign g1828 = ((~g769));
assign II11994 = ((~g6195));
assign g7064 = ((~II12829));
assign g3029 = ((~g1929));
assign g8885 = (g8723)|(g8806)|(II15243);
assign II11971 = ((~g6179));
assign g1925 = ((~g825));
assign g6827 = ((~II12352));
assign II12088 = ((~g5874));
assign g5673 = (g4823)|(g4872);
assign g4811 = ((~II9158));
assign II15720 = ((~g9053));
assign g8779 = (g8634&g7037);
assign g4091 = (g129&g3639);
assign II10790 = ((~g5512))|((~II10789));
assign II13509 = ((~g7137));
assign g6743 = (g730&g5916);
assign g6101 = ((~g5317));
assign g8314 = (g443&g7920);
assign II9769 = ((~g1114))|((~II9767));
assign II5432 = ((~g1176));
assign g5459 = ((~g4882));
assign g7194 = ((~II13118));
assign g5302 = ((~g5028));
assign g1829 = ((~II5715));
assign II12250 = ((~g6651));
assign g6279 = ((~II11132));
assign g6605 = ((~II11821));
assign g3548 = ((~g2185));
assign II6615 = ((~g1983));
assign g9109 = ((~II15717));
assign II12678 = ((~g6516));
assign II15882 = ((~g9179))|((~II15880));
assign g4421 = (g333&g3131);
assign g4919 = ((~g4104));
assign g6879 = ((~II12508));
assign II15205 = ((~g8809));
assign II14489 = ((~g7829));
assign g6594 = ((~II11796));
assign g6837 = ((~II12382));
assign g8817 = (g4545&g8482);
assign II15519 = ((~g9019));
assign g3716 = ((~g2522));
assign II6259 = ((~g901))|((~II6257));
assign II8291 = ((~g878));
assign g5743 = ((~II10286));
assign II6540 = ((~g2557))|((~II6538));
assign II7651 = ((~g2573));
assign g8075 = (g7460&g7634);
assign g6155 = ((~II10826));
assign II6254 = ((~g536));
assign g1976 = ((~g1269));
assign g7626 = (g7463&g3466);
assign II9597 = ((~g4738));
assign g8704 = (g2829&g8386);
assign II15990 = ((~g9239));
assign II13544 = ((~g1167));
assign II7145 = ((~g2501));
assign II15539 = ((~g9005));
assign II10694 = ((~g5445));
assign g6923 = (g6570&g5612);
assign II7053 = ((~g2452));
assign II11164 = ((~g5469))|((~II11163));
assign II11773 = ((~g6262));
assign II15274 = (g8306)|(g8361)|(g8299)|(g8687);
assign g2709 = ((~g1747));
assign g6333 = ((~II11326));
assign II13858 = ((~g7329));
assign g2703 = ((~g1809));
assign g9276 = (g9244&g5649);
assign g2315 = ((~II6103))|((~II6104));
assign g6108 = ((~g5345));
assign g6389 = ((~II11494));
assign II15099 = (g7855)|(g7838)|(g7905)|(g7870);
assign g6142 = ((~II10790))|((~II10791));
assign II7688 = ((~g3650));
assign g6994 = (g3658&g6538);
assign g4899 = ((~g4080));
assign g7450 = (g6090)|(g7195);
assign II11171 = ((~g5477))|((~II11170));
assign g7264 = ((~II13234));
assign II12406 = ((~g6773));
assign g5363 = ((~II9827))|((~II9828));
assign II14291 = ((~g7680));
assign g3128 = ((~II6839));
assign g3848 = ((~II7347));
assign II7905 = ((~g2863));
assign g6364 = ((~II11419));
assign II9250 = ((~g4134));
assign g1567 = ((~g655));
assign g8219 = ((~II14436));
assign g8385 = (g695&g7811);
assign g6587 = ((~II11781));
assign g1784 = ((~II5636));
assign g3931 = ((~II7592));
assign g5185 = ((~II9681));
assign g4649 = ((~II8862));
assign g7523 = ((~II13749));
assign II15250 = (g8238)|(g8265)|(g8272)|(g8292);
assign II6941 = ((~g2051))|((~II6939));
assign g3129 = ((~II6843))|((~II6844));
assign II6970 = ((~g1872));
assign II13515 = ((~g7152));
assign II10993 = ((~g2389))|((~II10991));
assign g9347 = (g9332&g6226);
assign g1876 = ((~g77));
assign g6523 = ((~II11707));
assign II10807 = ((~g5294));
assign g8384 = (g636&g7793);
assign II16158 = ((~g9363));
assign II7279 = ((~g1898))|((~II7277));
assign g4413 = (g2371)|(g3285);
assign g4127 = (g2628&g2618);
assign g4068 = (g121&g3540);
assign II12199 = ((~g6475));
assign g4526 = (g2642&g741);
assign g8804 = (g6060)|(g8609);
assign g2925 = ((~g2324));
assign g6391 = ((~II11500));
assign g7158 = ((~II13048));
assign g1813 = ((~g620));
assign g8017 = ((~g7692));
assign g8757 = ((~g8585));
assign g1958 = ((~g786));
assign II11018 = ((~g5626));
assign g3130 = ((~II6849));
assign g2780 = ((~II6517));
assign g7297 = ((~II13323));
assign II11758 = ((~g1758))|((~II11757));
assign II8901 = ((~g4122));
assign g4619 = ((~II8772));
assign g5258 = ((~II9774));
assign II15956 = ((~g9216));
assign II8787 = ((~g4012));
assign II12576 = ((~g6574))|((~II12575));
assign g2941 = ((~g2349));
assign g4644 = ((~II8847));
assign II6009 = ((~g359));
assign II15475 = ((~g8901));
assign g3990 = ((~g3160));
assign g2727 = ((~g2424));
assign II15711 = ((~g9075));
assign II12259 = ((~g6652));
assign g8669 = ((~II14801));
assign g9251 = (g4748&g9230);
assign g2340 = ((~g1327));
assign g3851 = ((~II7356));
assign g2307 = ((~II6078));
assign g6556 = ((~II11732));
assign g4114 = ((~II7953));
assign g3936 = ((~II7605));
assign g4925 = ((~g4114));
assign g7132 = ((~II12980));
assign g3013 = ((~II6764));
assign g1665 = ((~g1467));
assign II12900 = ((~g6947));
assign II14005 = ((~g7434));
assign g5758 = ((~II10347));
assign g4634 = ((~II8817));
assign II10001 = ((~g1929))|((~II9999));
assign II6096 = ((~g521));
assign g5478 = ((~g5025));
assign g4839 = ((~g1879))|((~g4269));
assign g9360 = ((~II16116));
assign g6822 = ((~II12337));
assign g2767 = ((~II6509));
assign g6401 = (g5971&g5367);
assign g7238 = (g6707&g7098);
assign g2673 = ((~II6474));
assign g6951 = (g5511&g6595);
assign g1922 = ((~g1251));
assign II7353 = ((~g2833));
assign II11257 = ((~g5805));
assign II9381 = ((~g4062))|((~g1908));
assign II14573 = ((~g8179));
assign II15803 = ((~g9148));
assign g9011 = (g6046)|(g8892);
assign g8678 = ((~II14828));
assign II13413 = ((~g7127));
assign II13562 = ((~g7179));
assign II9363 = ((~g4258));
assign g2833 = ((~II6561));
assign g4699 = (g1557&g4276);
assign g1907 = ((~g52));
assign II7584 = ((~g3062));
assign g5512 = ((~g1879))|((~g4877));
assign g6396 = (g661&g6008);
assign g4028 = ((~II7797));
assign g6866 = ((~II12469));
assign g4168 = (g1106&g3500);
assign g6488 = ((~II11652));
assign g4930 = ((~g4121));
assign g2547 = ((~II6371));
assign II15033 = (II15029)|(II15030)|(II15031)|(II15032);
assign II8455 = (g3430&g3398&g3359&g3341);
assign g4720 = (g190&g4055);
assign g7588 = ((~II13909));
assign g6150 = ((~g5287));
assign g7514 = ((~II13722));
assign II14288 = ((~g7705));
assign II12238 = ((~g6637));
assign g8787 = ((~g8564));
assign g6208 = ((~II10965));
assign II6643 = ((~g1970));
assign II8612 = (g3430&g3398&g3359&g3341);
assign II15324 = ((~g8779));
assign g7677 = (g7503&g5073);
assign g7537 = (g7363&g7411);
assign g5814 = ((~II10475));
assign g6662 = ((~II11964));
assign g5489 = (g4912&g5053);
assign g6269 = ((~II11090));
assign g3869 = ((~II7400));
assign II7086 = ((~g1753))|((~II7085));
assign g8228 = ((~II14463));
assign II11028 = ((~g5642));
assign g2627 = ((~g1572));
assign g7045 = ((~g6490));
assign II15211 = ((~g8808));
assign II8333 = ((~g3721));
assign II11275 = ((~g5768));
assign II6463 = ((~g1769));
assign g1698 = ((~II5542));
assign g2328 = ((~II6127));
assign II9018 = ((~g3872));
assign g5305 = ((~g5009))|((~g4335))|((~g4328));
assign II13281 = ((~g7155));
assign g3768 = ((~g2253));
assign g1853 = ((~g766));
assign g7023 = ((~II12779));
assign II9341 = ((~g4251));
assign II9986 = ((~g4836))|((~II9985));
assign g9357 = (g9278)|(g9347);
assign g9053 = ((~II15557));
assign II13962 = ((~g7413));
assign II13341 = ((~g7207));
assign II10322 = ((~g2573))|((~II10320));
assign g8461 = (g658&g7793);
assign g5141 = ((~II9548))|((~II9549));
assign II11086 = ((~g5397));
assign g2157 = ((~II5897));
assign g1695 = ((~g778));
assign g2954 = ((~g2374));
assign g5541 = ((~g4814));
assign g5198 = ((~g4969));
assign II10639 = ((~g5224));
assign g3912 = ((~g3192));
assign g3973 = ((~g3097));
assign g8680 = ((~g8493)&(~g8239)&(~II14834));
assign II7950 = ((~g2774));
assign II13490 = ((~g7130));
assign II13231 = ((~g6897));
assign II14100 = ((~g7580));
assign g785 = ((~II5407));
assign g9384 = (g9383&g6245);
assign II8460 = (g3430&g3398&g3359&g2106);
assign g5269 = ((~II9791));
assign g4600 = ((~II8715));
assign g8766 = ((~g8545));
assign g6065 = ((~II10684));
assign II8394 = ((~g1925))|((~II8392));
assign II14996 = ((~g8510));
assign g5971 = ((~II10587));
assign g4030 = ((~g3160));
assign gbuf46 = (g1153);
assign g2014 = ((~g1421)&(~g1416));
assign g9028 = ((~II15498));
assign II12085 = ((~g5971));
assign g9271 = (g4748&g9244);
assign g6055 = (g5239&g4202);
assign g4702 = (g4243&g1690);
assign g4266 = ((~II8202));
assign g4031 = ((~II7804));
assign g3778 = ((~g2145));
assign II15411 = ((~g8897));
assign g8986 = (g8926)|(g8825);
assign g4120 = ((~II7967));
assign g2915 = ((~II6643));
assign g7199 = (g1467&g7003);
assign g8982 = (g8922)|(g8820);
assign II9630 = ((~g4867));
assign g1847 = ((~g765));
assign g1751 = ((~g452));
assign II13802 = ((~g1061))|((~II13800));
assign g3958 = ((~g3097));
assign II7423 = ((~g2703))|((~II7421));
assign g6900 = ((~II12571));
assign g4542 = ((~g2884));
assign II14148 = ((~g7543));
assign g7539 = ((~II13797));
assign g9317 = ((~g9306));
assign g5074 = ((~II9440));
assign g6147 = ((~II10804));
assign II16142 = ((~g9366));
assign g6093 = ((~g5345));
assign II6509 = ((~g1684));
assign g4603 = ((~II8724));
assign g6185 = ((~g5305)&(~g1590));
assign g8257 = (g146&g8042);
assign g6753 = (g5939&g5384);
assign g7681 = (g7444&g5099);
assign g9215 = ((~II15921));
assign II15225 = ((~g8689));
assign g2876 = ((~g2231));
assign g1983 = ((~II5839));
assign g5565 = ((~g2044))|((~g4933));
assign II13369 = ((~g7268));
assign g1675 = ((~g1519));
assign g6459 = (g6259)|(g6185)|(II11603);
assign g1728 = (g1432&g1439);
assign II13469 = ((~g7123));
assign II13882 = ((~g7350));
assign g6371 = ((~II11440));
assign II14370 = ((~g7603));
assign g2246 = ((~II5989));
assign gbuf60 = (g104);
assign g5047 = (g373&g3964);
assign II16126 = ((~g9354));
assign II14964 = ((~g8406));
assign g4777 = ((~II9084));
assign II9992 = ((~g2145))|((~g4871));
assign g4019 = ((~II7778));
assign g9072 = ((~II15610));
assign g8227 = ((~II14460));
assign II5920 = ((~g219));
assign g5525 = ((~g4934));
assign II9499 = ((~g4382));
assign g6654 = ((~II11942));
assign g4249 = (g3617)|(g1639);
assign g3991 = ((~g3160));
assign g3465 = ((~II6963));
assign g9374 = ((~II16148));
assign g7283 = ((~II13281));
assign g4637 = ((~II8826));
assign g9211 = ((~II15909));
assign g7364 = ((~II13506));
assign g5916 = ((~g5384));
assign II6574 = ((~g576));
assign g6174 = ((~g1855)&(~g5305));
assign II8613 = (g2074&g3287&g3264&g1987);
assign II13524 = ((~g7151));
assign g2265 = ((~II6000));
assign II7487 = ((~g1708))|((~II7485));
assign g1887 = ((~g83));
assign g1768 = ((~g605));
assign g4285 = ((~II8233));
assign g7316 = ((~II13377))|((~II13378));
assign II12319 = ((~g6741));
assign II8190 = ((~g3545));
assign g2614 = ((~g1562));
assign II15042 = (g7951)|(g7920)|(g7983)|(g8181);
assign g6961 = ((~II12684));
assign g7339 = ((~II13435));
assign g7321 = ((~g7187)&(~g6990));
assign g5210 = (g5045)|(g4385);
assign II9422 = ((~g4360));
assign g5159 = ((~II9603));
assign II13054 = ((~g6960));
assign g2389 = ((~g1230));
assign g6225 = ((~II11014));
assign g3051 = ((~II6791));
assign g5396 = ((~g4692));
assign g9207 = ((~g9197));
assign g5820 = ((~II10485));
assign g7747 = ((~II14112));
assign II9217 = ((~g4443));
assign gbuf64 = (g449);
assign g1960 = ((~g1268));
assign II15702 = ((~g9064));
assign g4071 = ((~II7850));
assign g1637 = ((~g1087));
assign g5142 = (g1677&g4202);
assign g5268 = ((~II9788));
assign g4803 = ((~II9132));
assign g6416 = (g710&g6026);
assign g7713 = (g4403&g7367);
assign g5038 = ((~g4457));
assign II8935 = ((~g4005));
assign II10329 = ((~g2562))|((~II10327));
assign g3094 = (g945&g1898);
assign II11714 = ((~g5772));
assign g6239 = (g1514&g5314);
assign II8546 = (g3430&g3398&g3359&g3341);
assign g8673 = ((~II14813));
assign g4333 = (g1087&g2782);
assign II14315 = ((~g7676));
assign II10485 = ((~g5229));
assign II13287 = ((~g7157));
assign II7655 = ((~g2734));
assign II9169 = ((~g1935))|((~g4244));
assign II10801 = ((~g5463));
assign g4812 = (g2490)|(g4237);
assign g8293 = (g4510&g7855);
assign g8324 = ((~II14573));
assign II14178 = ((~g7562));
assign g7449 = (g7272&g6901);
assign II7341 = ((~g2931));
assign II12193 = ((~g6468));
assign g7024 = ((~II12782));
assign II9639 = ((~g4685));
assign g4294 = ((~II8244))|((~II8245));
assign g6176 = (g1149&g5198);
assign g8668 = ((~II14798));
assign II10834 = ((~g5514))|((~g2584));
assign g9203 = ((~II15888))|((~II15889));
assign g9200 = ((~g9189));
assign g6909 = ((~II12592));
assign g7784 = (g7406)|(g6664)|(g3492)|(II14219);
assign II16033 = ((~g9282));
assign g3077 = ((~II6805));
assign g7222 = (g6049)|(g6971);
assign II6868 = ((~g530));
assign g2683 = ((~g1666));
assign II5667 = ((~g916));
assign II15881 = ((~g9190))|((~II15880));
assign g8750 = ((~g8524));
assign II6703 = ((~g1983));
assign II12170 = ((~g5956));
assign g9361 = ((~II16119));
assign g8915 = (g8794&g8239);
assign II16020 = ((~g9264));
assign g7787 = (g4791)|(g7602);
assign g3398 = ((~II6952));
assign g4267 = ((~II8205));
assign II11034 = ((~g5644));
assign g3651 = ((~II7129));
assign II8543 = ((~g2810));
assign g3515 = ((~g1388)&(~g2262)&(~g2230)&(~g2214));
assign II11165 = ((~g3029))|((~II11163));
assign g5244 = (g5107)|(g4436);
assign II13679 = ((~g7259));
assign g7143 = ((~g6996));
assign II7626 = ((~g3632));
assign g8340 = (g423&g7920);
assign II13261 = ((~g7041));
assign II12550 = ((~g6689))|((~g1462));
assign g9093 = ((~II15669));
assign II13653 = ((~g7246));
assign II12871 = ((~g6618))|((~II12869));
assign II15055 = (II15051)|(II15052)|(II15053)|(II15054);
assign g6884 = ((~II12523));
assign II15962 = ((~g9218));
assign g2712 = ((~g2039));
assign g2561 = ((~g1555));
assign g3779 = ((~g2511));
assign II15433 = ((~g8911));
assign g7680 = (g7367&g4166);
assign II13475 = ((~g7125));
assign g4628 = ((~II8799));
assign g6049 = (g1045&g5597);
assign g7147 = ((~g6904));
assign g4566 = ((~g2902));
assign g1916 = ((~g775));
assign g4029 = ((~II7800));
assign II10866 = ((~g5480))|((~g2605));
assign II5997 = ((~g114));
assign g4698 = ((~II8989));
assign g7593 = ((~II13924));
assign II8084 = ((~g3706));
assign g3834 = ((~II7305));
assign II14305 = ((~g7537));
assign g7676 = (g7367&g4216);
assign g4732 = ((~II9034));
assign g9111 = ((~II15723));
assign g7725 = ((~II14046));
assign g6857 = ((~II12442));
assign II15382 = ((~g8883));
assign g4880 = ((~g4287))|((~g1879));
assign g6327 = ((~II11308));
assign g9122 = (g8953)|(g9084);
assign g5894 = (g1118&g5552);
assign g9136 = (g8952)|(g9131);
assign g5548 = (g1549&g4826);
assign II6112 = ((~g4));
assign II14115 = ((~g7563));
assign II15863 = ((~g9174))|((~II15862));
assign g7105 = ((~II12903));
assign II6275 = ((~g906))|((~II6273));
assign g2334 = ((~II6143));
assign II13695 = ((~g7345));
assign g2371 = ((~g944));
assign II13137 = ((~g7027));
assign II13786 = ((~g7427))|((~II13785));
assign g6434 = (g855&g6048);
assign g4002 = ((~g3192));
assign II8983 = ((~g4536));
assign g1949 = ((~g1292));
assign II5531 = ((~g866));
assign II8606 = ((~g2487))|((~II8605));
assign g4661 = ((~II8898));
assign g7734 = ((~II14073));
assign II7215 = ((~g815))|((~II7214));
assign g7495 = ((~II13663));
assign g2724 = ((~g1814));
assign II15292 = (g8704)|(g8710)|(g8805);
assign g4012 = ((~II7765));
assign g8876 = (g8769&g6102);
assign g7202 = (g6028)|(g7071);
assign g2393 = ((~II6267));
assign II12469 = ((~g6586));
assign g7761 = ((~II14154));
assign g8456 = (g703&g7811);
assign II11239 = ((~g6173));
assign II11212 = ((~g6146));
assign g1752 = ((~g603));
assign g6252 = ((~g5418));
assign g4435 = (g414&g3160);
assign II13831 = ((~g7322));
assign II10421 = ((~g5208));
assign g8891 = (g8705)|(g8811)|(II15297)|(II15298);
assign g8064 = (g7483&g7634);
assign II5933 = ((~g1158));
assign g5766 = ((~II10373));
assign II8517 = ((~g3014));
assign g4283 = (g3587)|(g2665);
assign g8741 = (g3787&g8464);
assign g4824 = ((~II9182))|((~II9183));
assign g9181 = ((~g9177));
assign II8046 = (g2074&g2057&g3264&g1987);
assign II8558 = ((~g2502))|((~g2790));
assign g2781 = (g1600&g976);
assign g7018 = ((~II12768));
assign g2961 = ((~II6711));
assign II8186 = (g3778&g3549&g3568&g3583);
assign g7049 = ((~II12813));
assign II11332 = ((~g5832));
assign g8640 = ((~II14728));
assign II5883 = ((~g80));
assign g6569 = ((~II11747));
assign II11948 = ((~g5897));
assign g4387 = (g378&g3160);
assign g5624 = (g5140&g2794);
assign II7350 = ((~g2971));
assign II7198 = ((~g2509));
assign g8844 = (g4056&g8602);
assign II9038 = (g4507)|(g4497)|(g4486);
assign II7036 = ((~g2454));
assign II6872 = ((~g2185));
assign g9084 = (g8964&g5345);
assign g7169 = ((~II13075));
assign g5054 = ((~g4457));
assign g3028 = ((~II6775))|((~II6776));
assign II15894 = ((~g9195));
assign g6301 = ((~II11230));
assign g5191 = ((~g4969));
assign II10906 = ((~g5492))|((~g2605));
assign g6197 = ((~g875)&(~g866)&(~g1590)&(~g5291));
assign g8837 = (g426&g8564);
assign g7137 = ((~II12993));
assign g8664 = ((~II14786));
assign II12502 = ((~g6604));
assign g5160 = ((~II9606));
assign g5203 = (g5032)|(g4378);
assign II6454 = ((~g1868));
assign g4900 = ((~II9258));
assign g4219 = ((~II8120))|((~II8121));
assign g4790 = (g4185)|(g4131)|(g4129)|(II9107);
assign g6977 = ((~g6664));
assign g3517 = ((~g2283));
assign g7328 = ((~g7196)&(~g7001));
assign g4259 = ((~II8196));
assign g8302 = (g4521&g7855);
assign II14468 = (g7937)|(g7887)|(g8029)|(g8018);
assign II11149 = ((~g5473))|((~g3038));
assign II15052 = (g7855)|(g7838)|(g7905)|(g7870);
assign II10265 = ((~g5468));
assign g4076 = ((~II7859));
assign g7180 = ((~II13092));
assign g7424 = ((~II13547));
assign II14427 = ((~g7835));
assign II6201 = ((~g831))|((~g891));
assign g5177 = ((~II9657));
assign g7307 = ((~II13353));
assign g7055 = ((~g6517));
assign g9319 = ((~g9309));
assign II12091 = ((~g5988));
assign g6804 = ((~II12283));
assign gbuf35 = (g1012);
assign g2253 = ((~g1323));
assign g2930 = ((~g2328));
assign g3506 = ((~g1781));
assign g3082 = ((~g1680));
assign II5466 = ((~g926));
assign g5040 = (g3900)|(g3895)|(g3890)|(g4363);
assign g8716 = (g3506&g8443);
assign g3874 = ((~g2957));
assign II11562 = ((~g5939));
assign g6226 = ((~g5658));
assign II9672 = ((~g4803));
assign II11832 = ((~g6274));
assign II11151 = ((~g3038))|((~II11149));
assign g6899 = ((~g6525));
assign II9938 = ((~g4878));
assign g4382 = ((~II8373));
assign II11080 = ((~g2511))|((~II11078));
assign g6767 = ((~II12170));
assign II8769 = ((~g3999));
assign g6465 = ((~g5403)&(~g5802)&(~g5769)&(~g5790));
assign g4225 = (g2686&g2689&g2692&g2695);
assign II12927 = ((~g7014));
assign II10292 = ((~g5577));
assign g4565 = ((~g2901));
assign II12933 = ((~g7018));
assign II11622 = ((~g5847));
assign II5696 = ((~g1513))|((~II5695));
assign g7173 = ((~g6980));
assign II8757 = ((~g3921));
assign g2899 = ((~g2272));
assign g1583 = ((~g718));
assign g6420 = (g5918&g5367);
assign g7093 = ((~II12870))|((~II12871));
assign g7474 = ((~II13628));
assign II7520 = ((~g2734));
assign II13639 = ((~g7257))|((~II13638));
assign g4678 = ((~II8935));
assign g5312 = ((~g5009))|((~g5002))|((~g4963));
assign g7828 = ((~II14245))|((~II14246));
assign g7709 = (g7367&g4529);
assign g3631 = ((~II7098));
assign g2494 = ((~g9));
assign g5687 = ((~II10190));
assign g5582 = ((~g4969));
assign II15334 = ((~g8800));
assign II8040 = (g3430&g3398&g3359&g3341);
assign II7937 = ((~g3614))|((~g1138));
assign II15085 = (g8363)|(g8342)|(g8407)|(g8386);
assign II6127 = ((~g471));
assign g3829 = ((~II7290));
assign II10965 = ((~g5719));
assign g4607 = ((~II8736));
assign II12478 = ((~g6603));
assign II13484 = ((~g7128));
assign g4595 = ((~g2942));
assign II8904 = ((~g4126));
assign g3871 = ((~g2953));
assign II14747 = ((~g8175));
assign g9305 = ((~II16033));
assign g6456 = (g6116&g2407);
assign II14094 = ((~g7593));
assign g1575 = ((~g685));
assign II15756 = ((~g9081));
assign g3966 = ((~g3160));
assign g2373 = ((~II6217));
assign g6064 = ((~II10681));
assign g1870 = ((~II5751));
assign g8068 = (g7687&g5610);
assign g2918 = ((~g2310));
assign g6214 = ((~g878)&(~g5284));
assign g2959 = ((~g1926));
assign II13220 = (g58)|(g6258)|(g5418);
assign g9060 = ((~II15574));
assign g4873 = ((~II9217));
assign g6444 = (g1676&g6125);
assign g7330 = ((~II13410));
assign g3945 = ((~g3097));
assign g6376 = ((~II11455));
assign g7207 = ((~II13137));
assign II12217 = ((~g6631));
assign g7069 = ((~g5435))|((~g6680));
assign g9261 = (g9238)|(g6227);
assign g6355 = ((~II11392));
assign II8760 = ((~g3931));
assign g4596 = ((~g3466));
assign II5781 = ((~g979));
assign g4613 = ((~II8754));
assign g6771 = (g146&g6004);
assign g5797 = ((~II10430));
assign g8131 = ((~II14378));
assign g2091 = ((~g819));
assign g7610 = ((~g7450));
assign II10569 = ((~g5417));
assign II5978 = ((~g414));
assign g6429 = (g168&g6035);
assign g7162 = ((~II13060));
assign g8781 = ((~g8585));
assign g5085 = ((~II9457));
assign g5515 = ((~g4923));
assign g3549 = ((~g2404));
assign g6553 = ((~II11725));
assign g3986 = (g202)|(g3129);
assign g2343 = ((~g1392));
assign g4048 = (g1288&g3513);
assign g4096 = ((~II7911));
assign II12989 = ((~g6932));
assign g5617 = ((~g4969));
assign II7554 = ((~g2573));
assign g8854 = (g443&g8564);
assign g5435 = ((~g5121));
assign II7112 = ((~g2546));
assign II7539 = ((~g2996))|((~II7538));
assign g8823 = (g4561&g8512);
assign g8970 = ((~II15414));
assign g6601 = ((~g6083));
assign g5460 = ((~g4684));
assign g5712 = ((~II10224))|((~II10225));
assign g4840 = (g4235&g1980);
assign II12343 = ((~g6731));
assign g2647 = ((~II6425));
assign II13460 = ((~g7263));
assign II11431 = ((~g5782));
assign g3684 = ((~g2180));
assign II9310 = ((~g4268));
assign II6416 = ((~g1794));
assign g1684 = ((~g1));
assign g8152 = ((~II14388));
assign g6937 = ((~II12632));
assign II11287 = ((~g5806));
assign II10981 = ((~g5625))|((~II10980));
assign II12262 = ((~g6656));
assign g5138 = (g4108)|(g3049);
assign II13323 = ((~g7145));
assign II9396 = ((~g3908));
assign g7905 = ((~II14279));
assign g7003 = (g1462&g6689);
assign II11263 = ((~g5784));
assign g5242 = (g5105)|(g4434);
assign g4585 = ((~g2925));
assign g3721 = ((~II7211));
assign g5747 = ((~II10299))|((~II10300));
assign g4180 = (g1114&g3511);
assign II14974 = ((~g8442));
assign II11317 = ((~g5787));
assign g1933 = ((~g1247));
assign II9693 = ((~g1037))|((~II9691));
assign g8335 = (g342&g7870);
assign II15666 = ((~g9070));
assign II5401 = ((~g723));
assign g7268 = ((~II13244));
assign g4502 = ((~II8559))|((~II8560));
assign II6996 = ((~g2275))|((~g2242));
assign II12388 = ((~g6403));
assign g9366 = ((~II16126));
assign II12025 = ((~g5918));
assign g6308 = ((~II11251));
assign II13362 = ((~g7265));
assign II6075 = ((~g2));
assign g3560 = ((~g2361));
assign g9158 = (g9137&g6070);
assign g2816 = ((~g1685));
assign II12832 = ((~g6722))|((~g6709));
assign g9048 = ((~II15546));
assign g6044 = (g1467&g5584);
assign II8240 = (g2298&g2316&g2334&g2354);
assign II8029 = (g2074&g2057&g3264&g1987);
assign II8998 = ((~g4576));
assign g3658 = ((~II7149))|((~II7150));
assign g5846 = ((~g5367));
assign g3903 = ((~II7498));
assign II8264 = ((~g3653));
assign II6468 = ((~g1917));
assign g2354 = ((~II6178));
assign g3859 = ((~II7380));
assign g6616 = ((~II11848));
assign II10702 = ((~g5529));
assign g5829 = ((~II10512));
assign g2906 = ((~g2288));
assign g8962 = (g8890&g5317);
assign II15690 = ((~g9074));
assign II13018 = ((~g1142))|((~II13016));
assign II15729 = ((~g9073));
assign II8823 = ((~g3965));
assign g7070 = ((~g6562));
assign II13004 = ((~g1053))|((~II13002));
assign g3076 = ((~g1831));
assign II13241 = ((~g7030));
assign g5395 = ((~II9840));
assign II13589 = ((~g7234))|((~II13587));
assign II13921 = ((~g7362));
assign II9182 = ((~g4231))|((~II9181));
assign II8436 = (g3430&g3398&g3359&g2106);
assign g5689 = ((~II10197))|((~II10198));
assign g5937 = (g5562&g2407);
assign g4916 = ((~g4202));
assign II7172 = ((~g1739))|((~g2006));
assign g8455 = (g652&g7793);
assign g7191 = (g7071)|(g6980);
assign II9953 = ((~g2131))|((~g4831));
assign g4954 = ((~g4319))|((~g2460));
assign II8504 = ((~g2038))|((~II8502));
assign g4957 = (g2746&g2728&g4320);
assign II6226 = ((~g408));
assign g5492 = ((~g4919));
assign g7492 = ((~II13656));
assign g6812 = ((~II12307));
assign g2626 = ((~g1571));
assign II12968 = ((~g6925));
assign II5706 = ((~g901));
assign II12535 = ((~g6599));
assign g5310 = ((~g5009))|((~g4335))|((~g4963));
assign g2832 = ((~g2184));
assign g6102 = ((~g5345));
assign II12687 = ((~g6745));
assign g4103 = ((~II7922));
assign II13669 = ((~g7240));
assign g6402 = (g665&g6012);
assign II13906 = ((~g7358));
assign II15030 = (g7855)|(g7838)|(g7905)|(g7870);
assign gbuf23 = (g1390);
assign g6828 = ((~II12355));
assign g3189 = ((~II6864));
assign II13822 = ((~g7459));
assign g4054 = (g3767&g2424);
assign g2964 = ((~II6716));
assign II13296 = ((~g7161));
assign g1821 = ((~g631));
assign II5383 = ((~g647));
assign g3894 = ((~II7460))|((~II7461));
assign g6848 = ((~II12415));
assign g1581 = ((~g710));
assign II8916 = ((~g4195));
assign g2104 = ((~II5879));
assign gbuf76 = (g921);
assign g8768 = ((~g8585));
assign II12141 = ((~g5897));
assign g3840 = ((~II7323));
assign g6817 = ((~II12322));
assign g7193 = (g6911&g1616);
assign g5984 = (g1041&g5484);
assign g7358 = ((~II13490));
assign g4044 = ((~g2595));
assign g7112 = ((~II12924));
assign g7695 = (g7367&g4466);
assign g4451 = (g359&g3131);
assign g6094 = ((~II10716));
assign II5512 = ((~g557));
assign II10028 = ((~g4825));
assign g4574 = ((~g3466));
assign g5009 = ((~g4344));
assign g2288 = ((~II6048));
assign II10460 = ((~g5219));
assign g3923 = ((~II7564));
assign g9124 = (g8876)|(g9038);
assign II14472 = ((~g8147))|((~g1069));
assign II10873 = ((~g5516))|((~g2595));
assign II10092 = ((~g4881))|((~g2177));
assign II14807 = ((~g8603));
assign g8972 = ((~II15420));
assign g6924 = (g6400)|(g6405);
assign g2184 = ((~II5911));
assign g1842 = ((~g764));
assign g6070 = ((~g5317));
assign gbuf72 = (g901);
assign II12487 = ((~g6623));
assign g3902 = ((~II7495));
assign II10923 = ((~g5525))|((~g2752));
assign II11958 = ((~g5874));
assign II11203 = ((~g6129));
assign g5294 = ((~g5087));
assign II10919 = ((~g5479));
assign II8844 = ((~g3992));
assign II10373 = ((~g5722));
assign g2631 = ((~g1586));
assign II6940 = ((~g2161))|((~II6939));
assign g7603 = ((~II13940));
assign g3972 = ((~II7691));
assign g4094 = ((~II7905));
assign II14816 = ((~g8642));
assign g6111 = ((~g5453));
assign II8177 = ((~g2810));
assign II12986 = ((~g6931));
assign g7160 = ((~II13054));
assign II14695 = ((~g8016));
assign g7095 = ((~II12877));
assign g1820 = ((~g621));
assign g8646 = (g553&g8094);
assign II7605 = ((~g2752));
assign g1924 = ((~g174));
assign II9243 = ((~g4305))|((~II9241));
assign II15340 = ((~g8856));
assign g9354 = (g9275)|(g9344);
assign g4494 = (II8546&II8547);
assign g6005 = (g5557&g2407);
assign II7444 = ((~g2973))|((~II7443));
assign II13106 = ((~g7056));
assign g3743 = ((~g1776));
assign II13740 = ((~g7364));
assign g6541 = (g6144&g3510);
assign g3611 = ((~II7079));
assign g6543 = (g6125)|(g1553);
assign g6135 = ((~II10770));
assign g7562 = ((~II13858));
assign g3754 = ((~g2543));
assign g7417 = (g7144&g1616);
assign g6995 = (g6435&g1616);
assign II15522 = ((~g9018));
assign II11669 = ((~g5918));
assign g1711 = ((~II5555));
assign g3950 = ((~g3131));
assign g8091 = (g7215)|(g6452)|(II14366);
assign II7797 = ((~g3019));
assign g5693 = ((~II10204));
assign g7114 = ((~II12930));
assign g4611 = ((~II8748));
assign g4155 = (II8028&II8029);
assign g7243 = ((~II13189));
assign g2222 = ((~II5939));
assign g3886 = ((~II7422))|((~II7423));
assign g8703 = (g3574&g8407);
assign g2891 = ((~g2265));
assign g4961 = (g377&g3904);
assign g7556 = ((~II13846));
assign II8886 = ((~g4308));
assign g9035 = ((~II15519));
assign g4356 = (g468&g3192);
assign g9337 = (g9240)|(g9327);
assign g9095 = ((~II15675));
assign II7430 = ((~g1541))|((~II7428));
assign II6758 = ((~g186))|((~II6757));
assign g8620 = (g751&g8199);
assign g8651 = ((~II14747));
assign II13672 = ((~g7242));
assign g7606 = (g7471&g3466);
assign g6970 = (g5035&g6490);
assign g6427 = ((~II11562));
assign g3160 = (g1751)|(g449);
assign II5989 = ((~g1460));
assign II10430 = ((~g5211));
assign g4307 = ((~g3700));
assign g8883 = ((~II15225));
assign g4343 = (g306&g3131);
assign II11880 = ((~g5748));
assign II7317 = ((~g2893));
assign g6697 = ((~II12025));
assign II7567 = ((~g2481))|((~g3780));
assign II9001 = ((~g4577));
assign gbuf4 = (g1308);
assign g8362 = (g504&g7966);
assign II7452 = ((~g3226))|((~g1106));
assign II10491 = ((~g5231));
assign g3833 = ((~II7302));
assign g4931 = ((~II9301));
assign II14410 = ((~g7697));
assign g2926 = ((~g2325));
assign g7508 = ((~II13704));
assign g4657 = ((~II8886));
assign g2663 = ((~II6460));
assign II9512 = ((~g3985));
assign II10223 = ((~g2522))|((~g4895));
assign g5514 = ((~g4922));
assign g8069 = (g7456&g7634);
assign g7227 = (g6992)|(g3128);
assign g3220 = ((~g1889));
assign II11170 = ((~g5477))|((~g3038));
assign II6500 = ((~g1913))|((~II6499));
assign II7302 = ((~g2825));
assign g3314 = ((~II6917))|((~II6918));
assign g8981 = (g8921)|(g8816);
assign II8472 = ((~g2821))|((~II8470));
assign II10457 = ((~g5218));
assign g2274 = ((~g782));
assign g6896 = ((~II12561));
assign II8053 = (g3316&g3287&g3264&g3238);
assign II6178 = ((~g1220));
assign II9162 = ((~g4272));
assign II14739 = ((~g8173));
assign g5608 = ((~g4969));
assign II8105 = ((~g3339));
assign g2548 = ((~g1351));
assign g5026 = ((~II9366));
assign II6936 = ((~g1878));
assign g5682 = ((~II10177));
assign g8261 = (g174&g8042);
assign g8287 = (g4500&g7855);
assign II10154 = ((~g5109));
assign g6350 = ((~II11377));
assign g4395 = (g405&g3160);
assign g2844 = ((~II6574));
assign g2213 = (g1367)|(g1368)|(g1369)|(g1370);
assign g8846 = (g510&g8585);
assign g4134 = ((~g3676));
assign g2314 = ((~II6099));
assign g5547 = (g4814&g1819);
assign g8642 = ((~II14732));
assign g6614 = ((~II11838));
assign g8975 = ((~II15429));
assign g534 = ((~II5365));
assign g7757 = ((~II14142));
assign g5087 = ((~II9463));
assign g7282 = (g5830&g6939);
assign II8449 = ((~g3630));
assign II8225 = (g3062)|(g2712)|(g2734)|(g2752);
assign g8462 = (g49&g8199);
assign g7251 = ((~II13203));
assign g6356 = ((~II11395));
assign II9071 = ((~g1149))|((~II9069));
assign II10207 = ((~g5075));
assign g6309 = ((~II11254));
assign II13193 = ((~g7007));
assign II11179 = ((~g3019))|((~II11177));
assign g5049 = (g474&g3969);
assign II11574 = ((~g5894))|((~g1122));
assign II7087 = ((~g1918))|((~II7085));
assign g9363 = (g9359)|(g6210);
assign g649 = ((~II5380));
assign g9029 = ((~II15501));
assign g7791 = (g4796)|(g7606);
assign II5939 = ((~g275));
assign g8863 = ((~g8493)&(~g8239)&(~II15175));
assign g6395 = (g2157&g6007);
assign II14270 = ((~g7703));
assign II9382 = ((~g4062))|((~II9381));
assign g3984 = (g2403&g3085);
assign g1886 = ((~II5766));
assign II15818 = ((~g9151))|((~II15817));
assign II15950 = ((~g9222));
assign g4057 = ((~II7832));
assign g1833 = ((~g770));
assign II9152 = ((~g3883))|((~II9151));
assign II12659 = ((~g6459));
assign g4115 = ((~II7956));
assign II13213 = ((~g7065))|((~g7082));
assign g7531 = ((~II13773));
assign g4898 = ((~g4079));
assign g7505 = ((~II13695));
assign g5477 = ((~g4908));
assign II6673 = ((~g2246));
assign g8940 = (g4543&g8775);
assign g7149 = ((~II13031));
assign II11870 = ((~g5752));
assign g3095 = ((~II6831));
assign II11701 = ((~g5772));
assign g5062 = (g235&g3973);
assign II15420 = ((~g8881));
assign g8788 = (g8620)|(g8658)|(II14990);
assign II7332 = ((~g2947));
assign g7589 = ((~II13912));
assign g6268 = (g1092&g5309);
assign II6900 = ((~g1866));
assign g6663 = ((~II11967));
assign II14349 = ((~g7588));
assign II13373 = ((~g7270));
assign g7185 = ((~II13099));
assign II10555 = ((~g5529));
assign g5149 = ((~II9573));
assign g7538 = ((~II13794));
assign g4160 = ((~g1231)&(~g2834));
assign II9333 = ((~g4245));
assign g5540 = ((~II9954))|((~II9955));
assign g3920 = ((~g3097));
assign g4650 = ((~II8865));
assign g3911 = ((~II7526));
assign g3760 = (II7232)|(II7233);
assign II11132 = ((~g5624));
assign g4932 = ((~g4202));
assign g8681 = ((~II14838))|((~II14839));
assign II13737 = ((~g7446));
assign g6770 = ((~II12180))|((~II12181));
assign g2239 = ((~II5978));
assign g7228 = (g6688&g7090);
assign g6186 = ((~II10919));
assign g2595 = ((~g1643));
assign II8165 = ((~g1943))|((~II8164));
assign g1772 = ((~g607));
assign II13499 = ((~g7134));
assign g7289 = ((~II13299));
assign g8239 = ((~g8073))|((~g8092));
assign g3767 = ((~II7240))|((~II7241));
assign g8727 = (g2724&g8421);
assign II14285 = ((~g7625));
assign g6125 = (g5548&g4202);
assign g5006 = ((~II9333));
assign II9987 = ((~g2096))|((~II9985));
assign II10390 = ((~g5195));
assign g7022 = ((~II12776));
assign g9214 = ((~II15918));
assign II6571 = ((~g1711));
assign g4179 = (g207)|(g3083);
assign g5197 = ((~g4938));
assign g5217 = (g5063)|(g4392);
assign II7374 = ((~g3084));
assign g6373 = ((~II11446));
assign II8034 = (g2074&g2057&g3264&g3238);
assign g5106 = (g398&g4015);
assign g2015 = ((~g33));
assign g9330 = ((~g9319));
assign g5610 = ((~g4938));
assign g6865 = ((~II12466));
assign II13588 = ((~g2556))|((~II13587));
assign g4374 = (g1182)|(g1186)|(g1179)|(II8363);
assign g4601 = ((~II8718));
assign g8172 = ((~II14397));
assign II8742 = ((~g3919));
assign II7460 = ((~g2506))|((~II7459));
assign II15074 = (g8363)|(g8342)|(g8407)|(g8386);
assign g4703 = ((~II8998));
assign g7678 = (g7367&g4158);
assign II9624 = ((~g4746));
assign gbuf30 = (g1524);
assign II8461 = (g3316&g3287&g2020&g3238);
assign g6952 = (g6633)|(g6204);
assign g7513 = ((~II13719));
assign g7290 = ((~II13302));
assign II10791 = ((~g2170))|((~II10789));
assign g9297 = ((~II16017));
assign g7536 = (g4414&g7367);
assign II11323 = ((~g5808));
assign II14448 = ((~g7792));
assign g9385 = ((~II16173));
assign g6738 = (g5847&g5367);
assign g2329 = ((~II6130));
assign g8884 = (g8735)|(g8818)|(II15232);
assign g8682 = ((~II14844));
assign II11037 = ((~g5299));
assign II10128 = ((~g4688));
assign g4778 = (g4169&g1760);
assign II13850 = ((~g7328));
assign g4669 = ((~II8922));
assign g1750 = ((~g602));
assign II10243 = ((~g5026));
assign g9252 = ((~II15982));
assign II10519 = ((~g5242));
assign g3901 = ((~II7492));
assign g1977 = ((~g1357));
assign g6334 = ((~II11329));
assign g3429 = (g1454&g1838&g1444);
assign g7108 = ((~II12912));
assign g6588 = ((~g5836));
assign g3963 = ((~II7672));
assign g1848 = ((~g772));
assign g6755 = ((~II12138));
assign II12652 = ((~g6664));
assign g7810 = (g4799)|(g7609);
assign g8383 = (g730&g7937);
assign g3883 = ((~g2276))|((~g3188));
assign II14439 = ((~g8063));
assign g7056 = ((~g6520));
assign II15098 = (g8131)|(g8111)|(g8042)|(g8156);
assign g6524 = ((~II11710));
assign g6196 = (g4927&g5615);
assign II6949 = ((~g2148));
assign g6744 = ((~II12124));
assign II6894 = ((~g1863));
assign g1555 = ((~II5428));
assign g7657 = (g7367&g4201);
assign g6941 = (g1126&g6582);
assign II7179 = ((~g2351))|((~g795));
assign II14825 = ((~g8651));
assign II10512 = ((~g5238));
assign g8087 = (g7471&g7634);
assign g4409 = (g384&g3160);
assign g5412 = ((~II9850));
assign II9747 = ((~g1549))|((~II9745));
assign II6234 = ((~g896))|((~II6232));
assign g594 = ((~II5368));
assign g9052 = (g8728)|(g8733)|(g9014)|(g8679);
assign II7970 = ((~g3557));
assign g6363 = ((~II11416));
assign II10973 = ((~g5726));
assign II8643 = (g2074&g3287&g3264&g1987);
assign g3649 = ((~g2424));
assign g9275 = (g9241&g5645);
assign g1568 = ((~g658));
assign g6685 = (g4067)|(g5969);
assign g9240 = (g9223&g5261);
assign g9160 = (g9139&g6092);
assign II8772 = ((~g4011));
assign g1827 = ((~g762));
assign II8907 = ((~g4095));
assign g2306 = ((~II6075));
assign II15533 = ((~g9002));
assign g8072 = ((~II14349));
assign g7135 = ((~II12989));
assign g4527 = ((~g3466));
assign g4145 = (g2639&g2635);
assign g6035 = ((~g5494));
assign g3891 = ((~g3097));
assign II6860 = ((~g2185));
assign g6392 = ((~II11503));
assign II10646 = ((~g5364));
assign II15251 = (g8302)|(g8288)|(g8311)|(g8296);
assign g7595 = ((~II13930));
assign g5231 = (g5081)|(g4411);
assign II9648 = ((~g4795));
assign II6064 = ((~g852))|((~g883));
assign II15275 = (g8693)|(g8703)|(g8712)|(g8717);
assign II11855 = ((~g5751));
assign g7298 = ((~II13326));
assign g2672 = ((~II6471));
assign II7648 = ((~g2712));
assign g2134 = ((~g1317));
assign g5186 = ((~II9684));
assign g4309 = ((~g3002))|((~g3124))|((~g3659));
assign g2509 = ((~g37));
assign II7365 = ((~g3061));
assign g5782 = ((~II10393));
assign g4884 = ((~g4492)&(~g4476)&(~g4456)&(~g4294));
assign g6493 = ((~II11659));
assign g4126 = ((~II7981));
assign g1690 = (g1021)|(g1025)|(g1018);
assign II13713 = ((~g7341));
assign g8985 = (g8925)|(g8824);
assign II6376 = ((~g38));
assign g7729 = ((~II14058));
assign g7157 = ((~II13045));
assign g1854 = ((~g773));
assign g8807 = ((~g8443)&(~g8421)&(~II15055));
assign g7131 = ((~g6976));
assign g8679 = ((~g8493)&(~g8239)&(~II14831));
assign g4237 = ((~II8151))|((~II8152));
assign g1959 = ((~g1252));
assign g7937 = ((~II14285));
assign g2392 = ((~g11));
assign g4924 = ((~g4113));
assign II10992 = ((~g5632))|((~II10991));
assign g5253 = (g5116)|(g4451);
assign g4667 = ((~II8916));
assign II10908 = ((~g2605))|((~II10906));
assign II15315 = ((~g8738));
assign II5646 = ((~g883));
assign g6310 = ((~II11257));
assign II13147 = ((~g7024));
assign II12629 = ((~g6523));
assign g4414 = (II8412&II8413);
assign II6358 = ((~g13));
assign II15586 = ((~g8987));
assign g3930 = ((~g3097));
assign g1797 = ((~g627));
assign g7237 = ((~g7050))|((~g3739));
assign g8953 = (g8758&g6093);
assign II13173 = ((~g7089));
assign II6124 = ((~g399));
assign II14052 = ((~g7494));
assign g8736 = (g3771&g8464);
assign g5069 = (g566&g3983);
assign g6507 = ((~II11683));
assign g8978 = (g8909&g5587);
assign II8952 = ((~g4197));
assign g4226 = ((~g3591));
assign g8926 = (g4593&g8755);
assign gbuf55 = (g200);
assign II6118 = ((~g243));
assign g6156 = ((~II10829));
assign g6141 = ((~II10786));
assign II10882 = ((~g5600));
assign g2043 = (g1263)|(g1257);
assign g7230 = (g4190)|(g6995);
assign II7445 = ((~g1701))|((~II7443));
assign II12526 = ((~g6626));
assign g4411 = (g462&g3192);
assign g6236 = ((~II11037));
assign II5404 = ((~g722));
assign g6322 = ((~II11293));
assign g6207 = ((~II10962));
assign g4597 = ((~II8706));
assign II7270 = ((~g955))|((~II7268));
assign II10439 = ((~g5214));
assign g7615 = (g7488&g3466);
assign g5709 = ((~g4841));
assign g8663 = ((~II14783));
assign g7592 = ((~II13921));
assign g2882 = ((~g2236));
assign II6166 = ((~g480));
assign II13638 = ((~g7257))|((~g7069));
assign II7041 = ((~g2401));
assign g4047 = (g1272&g3503);
assign g9125 = ((~II15753));
assign g3238 = ((~II6894));
assign g2372 = ((~II6214));
assign g6219 = ((~II10998));
assign g4733 = ((~g4202));
assign g7702 = ((~II13997));
assign II11964 = ((~g5971));
assign g2202 = ((~g1321));
assign g5234 = (g5090)|(g4421);
assign g9233 = ((~II15953));
assign g4821 = ((~g4220))|((~g3605));
assign II5636 = ((~g891));
assign II14492 = ((~g7829));
assign II12131 = ((~g5918));
assign II8847 = ((~g4025));
assign II13682 = ((~g7251));
assign g6417 = (g718&g6027);
assign II6652 = ((~g2016));
assign g2554 = ((~II6376));
assign g8341 = (g501&g7966);
assign g6698 = (g4073)|(g6001);
assign II12870 = ((~g2536))|((~II12869));
assign II15550 = ((~g9008));
assign II7785 = ((~g3029));
assign g7752 = ((~II14127));
assign II12558 = ((~g6449));
assign II15020 = (g8363)|(g8342)|(g8407)|(g8386);
assign g4196 = ((~II8097));
assign g8905 = (g8089)|(g8087)|(g8694);
assign g8630 = ((~g6110)&(~g7784)&(~g3591)&(~g1864));
assign g7148 = ((~II13028));
assign II11740 = ((~g6136));
assign II11004 = ((~g5613));
assign II9126 = ((~g3870));
assign II11254 = ((~g5793));
assign g4457 = ((~II8477));
assign g6144 = (g4175)|(g5458);
assign g9351 = ((~II16103));
assign II6849 = ((~g368));
assign II12567 = ((~g6721));
assign II11596 = ((~g6228));
assign g5574 = ((~g4969));
assign g2953 = ((~g2373));
assign g7156 = ((~II13042));
assign II11197 = ((~g6122));
assign II16049 = ((~g9288));
assign II10678 = ((~g5566));
assign II13794 = ((~g7346));
assign g7017 = (g3390&g6706);
assign g5202 = (g5031)|(g4377);
assign II6003 = ((~g228));
assign g2295 = ((~g995));
assign II12508 = ((~g6593));
assign g3921 = ((~II7558));
assign g6799 = ((~II12268));
assign g5835 = ((~II10528));
assign II8045 = (g3430&g3398&g3359&g2106);
assign g9193 = ((~g9181));
assign g5526 = ((~g5086));
assign g3568 = ((~g1935));
assign g6435 = ((~II11575))|((~II11576));
assign g7487 = ((~II13649));
assign g7544 = ((~II13816));
assign II8400 = (g3430&g3398&g3359&g3341);
assign II14193 = ((~g7532));
assign g6464 = (g6177&g2424);
assign II11633 = ((~g5897));
assign g8710 = (g2790&g8421);
assign II8326 = ((~g2011))|((~g2721));
assign g7129 = ((~II12973));
assign g6572 = ((~II11764));
assign g9009 = (g8949)|(g8858);
assign g8081 = (g834&g7658);
assign g1655 = ((~g1231));
assign g8277 = (g162&g8042);
assign II16058 = ((~g9294));
assign g1759 = ((~II5599))|((~II5600));
assign II13869 = ((~g7338));
assign II10190 = ((~g4670));
assign g3080 = ((~g1679));
assign g5048 = (g394&g3966);
assign g6048 = ((~g5246));
assign g4513 = ((~II8582))|((~II8583));
assign g7144 = ((~II13017))|((~II13018));
assign g4670 = ((~II8925));
assign g2223 = ((~II5942));
assign g8294 = (g281&g7838);
assign II15426 = ((~g8895));
assign II9493 = ((~g4426));
assign II7928 = ((~g2873));
assign g7726 = ((~II14049));
assign II13631 = ((~g7248));
assign g6883 = ((~II12520));
assign g6858 = ((~II12445));
assign g1676 = ((~g727));
assign II5521 = ((~g1098))|((~II5519));
assign II11974 = ((~g5956));
assign g6302 = ((~II11233));
assign II9233 = ((~g4310))|((~g2180));
assign g8890 = (II15290)|(II15291)|(II15292);
assign g4388 = (g402&g3160);
assign g4312 = (g3666&g3684&g3694&g3707);
assign g6706 = (g4077)|(g6002);
assign g5035 = ((~II9382))|((~II9383));
assign II11296 = ((~g5831));
assign g4075 = ((~II7856));
assign g4660 = ((~II8895));
assign g6803 = ((~II12280));
assign II6918 = ((~g1732))|((~II6916));
assign II6104 = ((~g921))|((~II6102));
assign II8127 = (g2699&g2674&g2677);
assign gbuf15 = (g1199);
assign g7441 = ((~II13580));
assign g5524 = ((~II9938));
assign II12301 = ((~g6703));
assign g6511 = ((~II11693));
assign II5515 = ((~g567));
assign II9548 = ((~g1952))|((~II9547));
assign g2625 = ((~g1570));
assign g8198 = ((~g7721));
assign g7714 = ((~II14019));
assign g7701 = (g7367&g4497);
assign II15111 = (g7951)|(g7920)|(g7983)|(g8181);
assign II9139 = ((~g4364));
assign II7964 = ((~g3488));
assign II13776 = ((~g7497));
assign g8925 = (g4592&g8754);
assign II8115 = (g2074&g3287&g3264&g1987);
assign g5178 = ((~II9660));
assign II10445 = ((~g5418));
assign g5125 = (g517&g4036);
assign g6962 = ((~II12687));
assign g7682 = (g6044)|(g7412);
assign g6655 = ((~II11945));
assign g6710 = (g55)|(g6264);
assign g8363 = ((~g7992));
assign g3858 = ((~II7377));
assign g8845 = (g432&g8564);
assign g8834 = (g7096)|(g8229);
assign II13060 = ((~g6959));
assign II8763 = ((~g3947));
assign II13225 = ((~g7095));
assign g6754 = ((~II12135));
assign g7320 = ((~II13388));
assign g7008 = (g6615&g5083);
assign II9558 = ((~g4597));
assign g6117 = ((~II10739));
assign g5166 = ((~II9624));
assign II12229 = ((~g6659));
assign g5228 = (g5078)|(g4408);
assign II9543 = ((~g4279));
assign g6660 = ((~II11958));
assign g3579 = ((~g1929));
assign II13419 = ((~g7277));
assign II9136 = ((~g4280));
assign II14231 = ((~g7566));
assign II7417 = ((~g3659));
assign g9375 = ((~II16151));
assign g4636 = ((~II8823));
assign II9606 = ((~g4687));
assign g7274 = ((~II13258));
assign II11525 = ((~g5874));
assign g7733 = ((~II14070));
assign II8706 = ((~g3828));
assign g2734 = ((~g2170));
assign II10854 = ((~g5521))|((~g2584));
assign g6472 = ((~g5971))|((~g5269));
assign II5368 = ((~g3853));
assign II9576 = ((~g4706));
assign g8667 = ((~II14795));
assign g6175 = (g4332&g5614);
assign II12466 = ((~g6687));
assign g6764 = ((~II12161));
assign II11449 = ((~g6068));
assign g8690 = (g3485&g8363);
assign g2379 = ((~II6239));
assign g5537 = (g3617)|(g4835);
assign g1664 = ((~g1462));
assign g1948 = ((~g1250));
assign II6148 = ((~g5));
assign II9663 = ((~g4809));
assign II7278 = ((~g2497))|((~II7277));
assign gbuf63 = (g368);
assign g5821 = ((~II10488));
assign g6421 = (g5847&g5384);
assign II11781 = ((~g6284));
assign g6930 = (g6414)|(g6420);
assign g5143 = ((~II9555));
assign g5211 = (g5046)|(g4386);
assign g6314 = ((~II11269));
assign II15557 = ((~g9010));
assign II10274 = ((~g5524));
assign g3052 = ((~g2096));
assign II6911 = ((~g1869));
assign II8392 = ((~g2949))|((~g1925));
assign II6522 = ((~g1919))|((~g1102));
assign g6368 = ((~II11431));
assign II5562 = ((~g1300));
assign II6209 = (g911)|(g916)|(g921)|(g883);
assign g9230 = ((~II15950));
assign II11841 = ((~g2548))|((~g6158));
assign g5120 = ((~II9512));
assign II12313 = ((~g6730));
assign g3192 = (g1756)|(g530);
assign g9092 = ((~II15666));
assign II5926 = ((~g297));
assign II7888 = ((~g3505));
assign g1769 = ((~II5609));
assign g4482 = ((~II8520));
assign g8238 = (g100&g8131);
assign II9993 = ((~g2145))|((~II9992));
assign II8140 = ((~g3429));
assign II13487 = ((~g7129));
assign g6458 = (g6184)|(g6259)|(g6174)|(g6214);
assign g4901 = (g3723&g4288&II9261);
assign g9210 = ((~g9200));
assign g7317 = ((~II13383));
assign II7807 = ((~g2595));
assign II7338 = ((~g2923));
assign II15073 = (g7951)|(g7920)|(g7983)|(g8181);
assign g7836 = ((~II14260));
assign II7576 = ((~g1718))|((~II7574));
assign g4559 = ((~g2898));
assign II11383 = ((~g5827));
assign II7526 = ((~g2752));
assign II15625 = ((~g9000));
assign II12457 = ((~g6671));
assign II9582 = ((~g4694));
assign II15862 = ((~g9174))|((~g9171));
assign g8327 = (g336&g7870);
assign g4067 = (g133&g3539);
assign g5196 = (g5020)|(g4369);
assign II7505 = ((~g3802))|((~II7503));
assign II14124 = ((~g7591));
assign g9202 = ((~II15881))|((~II15882));
assign g6720 = ((~g6254));
assign g2992 = ((~g1833));
assign g8994 = (g8934)|(g8836);
assign II7466 = ((~g2982))|((~g1704));
assign g8916 = ((~II15334));
assign g9298 = ((~II16020));
assign II11503 = ((~g6220));
assign g9157 = ((~g9141));
assign g4805 = ((~II9136));
assign II7629 = ((~g3633));
assign II7241 = ((~g2134))|((~II7239));
assign g5436 = (g1541&g4926);
assign II11652 = ((~g5939));
assign II9344 = ((~g4341));
assign g2273 = ((~II6024));
assign g8767 = ((~g8564));
assign g6130 = ((~II10761));
assign g4503 = ((~II8565));
assign g6554 = (g5762&g1616);
assign II12463 = ((~g6682));
assign II7712 = ((~g3657));
assign g2969 = ((~g2393));
assign II11887 = ((~g5918));
assign g5245 = (g5108)|(g4437);
assign II13314 = ((~g7160));
assign II10525 = ((~g5244));
assign g9382 = ((~II16168));
assign g3650 = ((~II7126));
assign g2917 = ((~g2309));
assign II15283 = (g8291)|(g8276)|(g8325)|(g8330);
assign II5789 = ((~g1524));
assign II12649 = ((~g6457));
assign gbuf5 = (g1309);
assign g7066 = ((~II12839));
assign II6425 = ((~g1811));
assign g6841 = ((~II12394));
assign II13376 = ((~g7199))|((~g1472));
assign g2038 = ((~g809));
assign g7167 = (g6438)|(g6915);
assign g5218 = (g5064)|(g4393);
assign g6871 = ((~II12484));
assign g9100 = ((~II15690));
assign g6915 = (g6493&g5246);
assign II11858 = ((~g6165));
assign g6028 = ((~g5529));
assign II10384 = ((~g5193));
assign g4035 = ((~II7814));
assign II12124 = ((~g5847));
assign II7269 = ((~g2486))|((~II7268));
assign g6617 = ((~II11851));
assign II12220 = ((~g6645));
assign g5787 = ((~II10406));
assign g3639 = ((~g2424));
assign g7432 = ((~II13559));
assign g7161 = ((~II13057));
assign g7331 = ((~II13413));
assign II12376 = ((~g6766));
assign g2999 = ((~g1823));
assign II15160 = ((~g8631));
assign II8339 = ((~g2966))|((~II8338));
assign g3946 = ((~g3097));
assign g2936 = ((~II6680));
assign II8721 = ((~g3918));
assign g6167 = ((~II10862));
assign g5075 = ((~II9443));
assign g3985 = ((~II7712));
assign g2933 = ((~II6673));
assign g4095 = ((~II7908));
assign g6173 = ((~II10882));
assign g7357 = ((~II13487));
assign g7111 = ((~II12921));
assign g1683 = ((~g795));
assign g7188 = ((~II13106));
assign g4093 = ((~II7902));
assign g6736 = ((~II12108));
assign II11912 = ((~g5897));
assign g4181 = (g1142&g3512);
assign gbuf2 = (g1236);
assign II10980 = ((~g5625))|((~g2210));
assign II13553 = (g1166)|(g1167)|(g1170);
assign g9119 = (g9049&g5345);
assign g8288 = (g270&g7838);
assign g7002 = (g6770&g5054);
assign g3229 = (g1728&g2015);
assign II5868 = ((~g74));
assign II15660 = ((~g9062));
assign g1785 = ((~g615));
assign II11614 = ((~g6239))|((~g1519));
assign g6701 = ((~II12032))|((~II12033));
assign g2407 = ((~II6286));
assign g2907 = ((~g2289));
assign g4662 = ((~II8901));
assign g9369 = ((~II16135));
assign g6255 = ((~II11066));
assign g9316 = ((~g9302));
assign g9068 = ((~II15598));
assign g6792 = ((~II12247));
assign g6600 = (g5443)|(g6055);
assign II10752 = ((~g5618));
assign II14246 = ((~g1065))|((~II14244));
assign g2290 = ((~II6054));
assign g4798 = (g4216&g1760);
assign II8796 = ((~g3934));
assign II14952 = (g8456)|(g8513)|(g8458)|(g8236);
assign g5170 = ((~II9636));
assign II11060 = ((~g5453));
assign g4800 = ((~II9123));
assign g8622 = (g738&g7811);
assign g9049 = (g8732)|(g8737)|(g9015)|(g8861);
assign g9087 = ((~II15651));
assign g6768 = ((~II12173));
assign g4789 = (g2751&g4202);
assign g6217 = ((~g5649));
assign g2646 = ((~II6422));
assign g8151 = (g849&g7658);
assign g5053 = ((~g4438));
assign II6963 = ((~g1558));
assign g7306 = ((~II13350));
assign g2174 = ((~g1319));
assign g5847 = ((~II10552));
assign II6826 = ((~g2185));
assign II6997 = ((~g2275))|((~II6996));
assign II15759 = ((~g9082));
assign II12833 = ((~g6722))|((~II12832));
assign g9177 = ((~II15811));
assign g7342 = ((~II13444));
assign g3499 = ((~g2185));
assign g4436 = (g492&g3192);
assign g7269 = ((~II13247));
assign g1746 = ((~g290));
assign g5623 = ((~g4969));
assign g8065 = ((~II14338));
assign II13209 = ((~g6912));
assign g3845 = ((~II7338));
assign II15169 = (g8483)|(g8464)|(g8514);
assign g2137 = ((~II5889));
assign g6227 = ((~II11018));
assign II5757 = (g969)|(g970)|(g966)|(g963);
assign g6838 = ((~II12385));
assign g5562 = ((~II10010))|((~II10011));
assign gbuf43 = (g1173);
assign g3992 = ((~II7723));
assign II12442 = ((~g6542));
assign g7746 = ((~II14109));
assign II13570 = ((~g7198));
assign II14244 = ((~g7683))|((~g1065));
assign II10198 = ((~g1958))|((~II10196));
assign g4403 = (II8400&II8401);
assign II14196 = ((~g7534));
assign II14058 = ((~g7544));
assign II8495 = (g3430&g3398&g3359&g2106);
assign II14330 = ((~g7538));
assign II13228 = ((~g6892));
assign II10815 = ((~g5418));
assign II13550 = ((~g1173));
assign g5209 = (g5044)|(g4384);
assign g4443 = ((~II8449));
assign II16061 = ((~g9294));
assign g6976 = (g4399&g6508);
assign g9267 = (g9251)|(g6225);
assign g3315 = ((~II6924))|((~II6925));
assign II10940 = ((~g5489));
assign II12415 = ((~g6410));
assign II15857 = ((~g9165))|((~II15855));
assign g8256 = (g95&g8131);
assign g3629 = ((~g2424));
assign g6162 = (g1134&g5724);
assign II8161 = ((~g3517));
assign II6716 = ((~g1721));
assign II16084 = ((~g9324));
assign g8638 = ((~II14722));
assign g1852 = ((~g887));
assign II14759 = (g7937)|(g7887)|(g8029)|(g8018);
assign g4917 = ((~g4102));
assign II8754 = ((~g3911));
assign g1941 = ((~II5812));
assign g6604 = ((~II11818));
assign II12888 = ((~g6948));
assign II7899 = ((~g3743));
assign g8814 = (g3880&g8463);
assign g1235 = ((~II5422));
assign II13785 = ((~g7427))|((~g1477));
assign II11224 = ((~g6255));
assign g5725 = ((~g4841));
assign g5763 = ((~II10366));
assign II12052 = ((~g5956))|((~II12051));
assign g5041 = ((~II9393));
assign II6078 = ((~g95));
assign g3873 = ((~g2956));
assign g6780 = ((~II12211));
assign g8877 = (g8773&g6104);
assign g4804 = (g952&g3876);
assign g8301 = (g182&g8156);
assign II5609 = ((~g16));
assign II14772 = (g7937)|(g7887)|(g8029)|(g8018);
assign II13719 = ((~g7334));
assign g6622 = ((~II11858));
assign g1574 = ((~g681));
assign II12080 = ((~g5971))|((~II12078));
assign g4545 = ((~g2887));
assign g7094 = ((~g6525));
assign g6109 = (g5453&g5335);
assign II11425 = ((~g5872));
assign g1573 = ((~g677));
assign II11926 = ((~g6190));
assign g4472 = (g440&g3160);
assign II12490 = ((~g6625));
assign g6628 = ((~II11880));
assign g6319 = ((~II11284));
assign g4564 = ((~II8665));
assign II7459 = ((~g2506))|((~g3815));
assign II8005 = (g3430&g3398&g3359&g2106);
assign II15086 = (II15082)|(II15083)|(II15084)|(II15085);
assign g9135 = (g8951)|(g9130);
assign g7174 = ((~g7097));
assign g4056 = ((~g3082));
assign II9823 = ((~g5138));
assign g9206 = ((~g9196));
assign II7523 = ((~g2562));
assign g6739 = (g4099)|(g6021);
assign g5433 = ((~g5024));
assign g5313 = (g4820&g2407);
assign g4328 = ((~g3086));
assign g7423 = ((~II13544));
assign II14932 = (g8278)|(g8329)|(g8461)|(g8382);
assign g4606 = ((~II8733));
assign g7455 = ((~II13613));
assign II9681 = ((~g4811));
assign g3514 = ((~g2424));
assign g3854 = ((~II7365));
assign II7938 = ((~g3614))|((~II7937));
assign g3828 = ((~II7287));
assign g7483 = ((~g7226));
assign g5595 = ((~II10079))|((~II10080));
assign II7239 = ((~g1658))|((~g2134));
assign g6112 = (g5673&g4841&g5541);
assign g8782 = (g8624)|(g8659)|(II14980);
assign g5583 = (g1775&g4969);
assign II14725 = ((~g8145));
assign II7195 = ((~g1795));
assign g9344 = (g9329&g6211);
assign II11991 = ((~g5939));
assign g3516 = ((~g2282)&(~g1401));
assign II14035 = ((~g7310));
assign g1584 = ((~g738));
assign g4053 = (g1292&g3523);
assign II7287 = ((~g2561));
assign II6309 = ((~g1336));
assign g4332 = ((~g3681))|((~g2368));
assign g8921 = (g4579&g8747);
assign g2982 = ((~g1848));
assign g3884 = ((~II7417));
assign g6940 = ((~II12639));
assign g7107 = ((~II12909));
assign II9918 = ((~g4968));
assign II13359 = ((~g7255));
assign g6362 = ((~II11413));
assign g5051 = ((~II9407));
assign g8382 = (g685&g7887);
assign II8033 = (g3430&g3398&g3359&g2106);
assign II9531 = ((~g4463));
assign g4712 = (g1179&g4276);
assign g5183 = ((~II9675));
assign II15880 = ((~g9190))|((~g9179));
assign g7500 = ((~II13676));
assign g6140 = ((~II10783));
assign g3757 = ((~g1977));
assign II15974 = ((~g9234));
assign g8830 = (g345&g8545);
assign II7293 = ((~g2955));
assign g9355 = (g9276)|(g9345);
assign g3583 = ((~g2128));
assign g6568 = ((~II11744));
assign g6063 = ((~II10678));
assign g9027 = ((~II15495));
assign g9147 = (g9136&g6103);
assign g8695 = (g2709&g8363);
assign g5987 = ((~g5294));
assign II9242 = ((~g2540))|((~II9241));
assign g9274 = (g4748&g9255);
assign II13335 = ((~g7206));
assign II7186 = ((~g2353))|((~g1834));
assign g7236 = ((~g6944));
assign g7295 = ((~II13317));
assign g3529 = ((~g2323));
assign g3562 = ((~II7044));
assign II8277 = ((~g3504));
assign g4363 = ((~II8339))|((~II8340));
assign g8077 = (g859&g7616);
assign g6157 = (g1130&g5717);
assign g6335 = ((~II11332));
assign II5380 = ((~g645));
assign II8775 = ((~g4019));
assign g8998 = (g8938)|(g8842);
assign g2671 = ((~II6468));
assign II7311 = ((~g2879));
assign II8966 = ((~g4444));
assign g8702 = (g2837&g8386);
assign g6294 = ((~II11209));
assign g4062 = (g809&g2986);
assign g6250 = ((~g5679));
assign II9591 = ((~g4710));
assign II9103 = ((~g4374));
assign g8850 = ((~g8493)&(~g8239)&(~II15152));
assign g4129 = (g2629&g2621);
assign g8815 = (g258&g8524);
assign g2551 = ((~g1360));
assign II9678 = ((~g4808));
assign g2052 = ((~II5865));
assign g3084 = ((~II6820));
assign gbuf44 = (g1170);
assign II5365 = ((~g3843));
assign II11368 = ((~g5833));
assign g8653 = (g573&g8094);
assign g4664 = ((~II8907));
assign g7781 = ((~II14214));
assign g2051 = ((~g1444))|((~g1450));
assign g8954 = (g8763&g6097);
assign g4412 = (g486&g3192);
assign g4116 = ((~II7959));
assign g3805 = ((~g1752));
assign g7768 = ((~II14175));
assign g2923 = ((~II6657));
assign g5068 = (g475&g3982);
assign g1556 = ((~g65));
assign g6431 = (g5847&g5494);
assign g5752 = ((~II10328))|((~II10329));
assign g6849 = ((~II12418));
assign g8226 = ((~II14457));
assign II16135 = ((~g9357));
assign g6050 = ((~g5246));
assign II9440 = ((~g4285));
assign g6300 = ((~II11227));
assign g7326 = ((~g7194)&(~g6999));
assign g6745 = (g1872&g6198);
assign g4658 = ((~II8889));
assign II13577 = ((~g7186));
assign II5621 = ((~g1130))|((~II5619));
assign II7232 = (g2367)|(g2352)|(g2378)|(g2330);
assign g9001 = (g8941)|(g8846);
assign II13012 = ((~g7071));
assign II13066 = ((~g6957));
assign g5151 = ((~II9579));
assign g2943 = ((~g2362));
assign II15071 = (g8131)|(g8111)|(g8042)|(g8156);
assign g3159 = ((~II6856));
assign g2375 = ((~II6223));
assign II8573 = (g3430&g3398&g3359&g2106);
assign g9307 = ((~g9300));
assign g3933 = ((~g3131));
assign g8018 = ((~II14315));
assign g3728 = ((~g2202));
assign g4786 = (g4107)|(g4097)|(g4124)|(II9099);
assign g4238 = (g2695&g2698&II8157);
assign II13595 = ((~g7216));
assign g8944 = (g4539&g8783);
assign II7436 = ((~g2517))|((~g3822));
assign g8977 = ((~II15433));
assign II8724 = ((~g3927));
assign g206 = ((~II5353));
assign g8882 = ((~II15222));
assign g4417 = (II8417&II8418);
assign II11533 = ((~g5847));
assign g1743 = ((~g598));
assign g8909 = (g6043)|(g8764);
assign II11827 = ((~g6231));
assign II12196 = ((~g6471));
assign g5696 = ((~II10207));
assign g8698 = (g3774&g8342);
assign II14754 = (g7937)|(g7887)|(g8029)|(g8018);
assign g5028 = ((~II9372));
assign g9151 = (g9144)|(g8961);
assign II14184 = ((~g7726));
assign g1774 = ((~II5616));
assign g5443 = (g1549&g4935);
assign II11751 = ((~g6112))|((~II11750));
assign II5801 = ((~g1424));
assign II8751 = ((~g4009));
assign g7021 = (g3390&g6673);
assign g3075 = ((~g2216));
assign g5823 = ((~II10494));
assign II9954 = ((~g2131))|((~II9953));
assign g6731 = ((~II12101));
assign II13267 = ((~g6913));
assign g6406 = (g154&g6018);
assign g1831 = ((~g689));
assign gbuf36 = (g1014);
assign g5147 = ((~II9567));
assign g6298 = ((~II11221));
assign g6864 = ((~II12463));
assign g9386 = ((~II16176));
assign g5552 = (g1114&g4832);
assign II5718 = ((~g896));
assign g6398 = ((~II11515));
assign g3680 = ((~II7187))|((~II7188));
assign II15031 = (g7951)|(g7920)|(g7983)|(g8181);
assign g8676 = ((~II14822));
assign g2769 = ((~g2424));
assign II14980 = (g8362)|(g8403)|(g8610);
assign g4066 = (g1280&g3532);
assign g8735 = (g2807&g8443);
assign II8014 = (g3430&g3398&g3359&g3341);
assign g5230 = (g5080)|(g4410);
assign g2913 = ((~g2307));
assign g4583 = ((~g2924));
assign II9099 = (g4127)|(g4123)|(g4117);
assign g7535 = ((~II13786))|((~II13787));
assign g6589 = ((~g6083));
assign II7082 = ((~g2470));
assign II9383 = ((~g1908))|((~II9381));
assign II8739 = ((~g3910));
assign II10073 = ((~g2253))|((~II10071));
assign II13350 = ((~g7223));
assign g5105 = (g354&g4013);
assign II5908 = ((~g196));
assign II7070 = ((~g1643))|((~II7068));
assign g4631 = ((~II8808));
assign II10475 = ((~g5529));
assign II9785 = ((~g4747));
assign g3541 = (g1663)|(g1421);
assign g5668 = ((~II10151));
assign g3019 = ((~g2007));
assign g7528 = ((~II13764));
assign g4796 = (g950&g4584);
assign g7078 = ((~g6683));
assign g8856 = ((~II15160));
assign II15062 = ((~g8632));
assign II6853 = ((~g2185));
assign g8281 = (g168&g8042);
assign II9336 = ((~g4493));
assign g8789 = ((~g8564));
assign II13196 = ((~g7008));
assign g6593 = ((~II11793));
assign g2453 = ((~II6291));
assign II6784 = ((~g2052));
assign g3915 = ((~II7539))|((~II7540));
assign g2230 = (g1380)|(g1381)|(g1382)|(g1383);
assign II15836 = ((~g9165));
assign g7043 = ((~g6543));
assign g1721 = ((~II5565));
assign II15669 = ((~g9045));
assign g4246 = (g1106&g3226);
assign g5476 = ((~g4907));
assign g6230 = ((~II11025));
assign g6975 = ((~II12712));
assign g6259 = ((~g3002)&(~g5312));
assign II11551 = ((~g1045))|((~II11549));
assign g7146 = ((~g6998));
assign II7101 = ((~g2478));
assign II8745 = ((~g3929));
assign II8510 = ((~g2517))|((~g2807));
assign g7711 = ((~II14012));
assign g6340 = ((~II11347));
assign g6779 = ((~II12208));
assign g4366 = (g216&g3097);
assign II11272 = ((~g5758));
assign II14801 = ((~g8608));
assign g7096 = (g6677&g5101);
assign g4540 = ((~g2882));
assign II14777 = ((~g8511));
assign II6099 = ((~g584));
assign g3286 = ((~II6905))|((~II6906));
assign g8603 = ((~II14674));
assign II6217 = ((~g105));
assign g2692 = ((~g1671));
assign g9061 = ((~II15577));
assign g6969 = ((~II12702));
assign II6267 = ((~g100));
assign g7679 = (g7447&g5084);
assign g2016 = ((~II5852));
assign g5563 = (g3390&g5070);
assign g7347 = ((~II13457));
assign II11326 = ((~g5819));
assign II15230 = (g8274)|(g8321)|(g8298)|(g8696);
assign g2332 = ((~g926));
assign g6374 = ((~II11449));
assign g4608 = ((~II8739));
assign g9013 = (g8907&g8239);
assign g5632 = ((~g2276))|((~g4901));
assign II12154 = ((~g5874));
assign g1611 = ((~g1073));
assign II8524 = (g3316&g2057&g3264&g1987);
assign g7586 = ((~II13903));
assign g4560 = ((~g2899));
assign g6183 = ((~II10914));
assign II14273 = ((~g7631));
assign II15855 = ((~g9168))|((~g9165));
assign II10900 = ((~g5520))|((~II10899));
assign g8541 = ((~g8094));
assign g8709 = (g2818&g8386);
assign II13587 = ((~g2556))|((~g7234));
assign g6902 = ((~II12576))|((~II12577));
assign g9311 = ((~II16049));
assign II7959 = ((~g2793));
assign g7010 = (g1049&g6574);
assign g6263 = ((~g5688));
assign g8689 = ((~II14857));
assign II15833 = ((~g9162));
assign II7305 = ((~g3048));
assign g4109 = (g990&g3790);
assign g5706 = (g4955)|(g4342);
assign II11135 = ((~g5476))|((~g3052));
assign g4394 = (g381&g3160);
assign gbuf56 = (g201);
assign g8652 = (g563&g8094);
assign g5681 = ((~g5132))|((~g2043));
assign g7777 = ((~II14202));
assign II7164 = ((~g2157));
assign g4933 = (g2746&g2728&g4320&g2770);
assign II9555 = ((~g4892));
assign II6160 = ((~g324));
assign g7576 = ((~II13873));
assign g8647 = ((~II14739));
assign g6684 = ((~II11998));
assign II9567 = ((~g4693));
assign II6337 = ((~g1348));
assign g6006 = (g5575&g2424);
assign II6561 = ((~g1715));
assign II14828 = ((~g8639));
assign g5713 = ((~g4841));
assign II10783 = ((~g5542));
assign gbuf9 = (g1191);
assign II14413 = ((~g7723));
assign g1826 = ((~g632));
assign II11144 = ((~g3062))|((~II11142));
assign g3928 = ((~g3097));
assign g2632 = ((~g1576));
assign g7549 = ((~II13831));
assign g6966 = (g6580&g5580);
assign g7312 = ((~g7178)&(~g6970));
assign g6351 = ((~II11380));
assign g9036 = ((~II15522));
assign g3612 = ((~II7082));
assign II11293 = ((~g5824));
assign g4135 = (II7994&II7995);
assign g8061 = ((~II14330));
assign g7442 = ((~II13583));
assign g1929 = ((~g1224));
assign g7609 = (g7467&g3466);
assign g7754 = ((~II14133));
assign II8224 = (g3019)|(g3029)|(g3038)|(g3052);
assign g8657 = ((~II14763));
assign g6074 = ((~g5317));
assign II8805 = ((~g3976));
assign g9054 = (g8724)|(g8729)|(g9013)|(g8680);
assign g7113 = ((~II12927));
assign g5519 = ((~II9929));
assign g7778 = ((~II14205));
assign II11055 = ((~g5696));
assign g8621 = (g734&g7937);
assign g3862 = ((~II7389));
assign g3578 = ((~II7053));
assign g2366 = ((~II6198));
assign g5546 = ((~II9964))|((~II9965));
assign g6878 = ((~II12505));
assign g7486 = ((~II13646));
assign g5309 = ((~g4969));
assign II9053 = ((~g4327));
assign g3841 = ((~II7326));
assign g2787 = ((~g1807));
assign g7634 = (g7367&g4549);
assign II8814 = ((~g4028));
assign g7365 = ((~II13509));
assign II9041 = (g4483)|(g4466)|(g4445);
assign g6992 = (g6610&g3519);
assign g4871 = ((~g3635))|((~g3605))|((~g4220))|((~g3644));
assign g8936 = (g3875&g8768);
assign g2989 = ((~g1843));
assign II15040 = (g8131)|(g8111)|(g8042)|(g8156);
assign g5513 = (g4889&g5071);
assign II13293 = ((~g7159));
assign II6305 = ((~g1333));
assign II6608 = ((~g1612));
assign g5227 = (g5077)|(g4407);
assign g5733 = ((~II10256));
assign II6800 = ((~g2016));
assign II8079 = (g3316&g3287&g2020&g1987);
assign g7552 = (g7319&g5749);
assign II8373 = ((~g3783));
assign g695 = ((~II5392));
assign II15738 = ((~g9079));
assign g6505 = ((~II11677));
assign g5767 = (g5344&g3079);
assign II9463 = ((~g3942));
assign g7744 = ((~II14103));
assign g8643 = (g547&g8094);
assign g4378 = (g321&g3131);
assign II11200 = ((~g6251));
assign g8899 = (g8839)|(g8652);
assign II15100 = (g7951)|(g7920)|(g7983)|(g8181);
assign g4493 = ((~II8543));
assign g9074 = ((~II15616));
assign g6281 = ((~II11143))|((~II11144));
assign II12996 = ((~g6934));
assign g6229 = ((~g5665));
assign II15889 = ((~g9191))|((~II15887));
assign g5439 = ((~g5058));
assign II14039 = ((~g7449));
assign g7138 = ((~II12996));
assign g5418 = ((~g5100));
assign II15571 = ((~g8982));
assign g8309 = (g550&g8181);
assign II9466 = ((~g3943));
assign g9309 = ((~II16043));
assign II12776 = ((~g6739));
assign g6032 = ((~g5494));
assign II8922 = ((~g4229));
assign g2106 = ((~II5883));
assign g2351 = ((~g792));
assign II8913 = ((~g4306));
assign II9654 = ((~g4792));
assign g7178 = ((~II13088));
assign II8446 = ((~g3014));
assign g5609 = ((~g4748));
assign II13701 = ((~g7349));
assign gbuf73 = (g906);
assign II5413 = ((~g1016));
assign II10836 = ((~g2584))|((~II10834));
assign g5343 = (g4690)|(g2862);
assign g4549 = (II8642&II8643);
assign II8456 = (g3316&g3287&g2020&g1987);
assign g5246 = ((~II9760));
assign II7392 = ((~g3230));
assign g9168 = (g9160)|(g9025);
assign II9684 = ((~g4813));
assign g4524 = ((~g2869));
assign II11764 = ((~g6056));
assign g3532 = ((~g2407));
assign g4186 = (g1118&g3520);
assign g4274 = ((~II8218));
assign g5117 = (g435&g4024);
assign II5901 = ((~g52));
assign g4314 = (g3694&g3684&g3666);
assign II14403 = ((~g7679));
assign g3983 = ((~g2845));
assign g5750 = ((~II10314))|((~II10315));
assign II15705 = ((~g9068));
assign g2798 = ((~g1787));
assign g8753 = ((~II14925));
assign II10538 = ((~g5255));
assign II11689 = ((~g5956));
assign g5101 = ((~g4259));
assign g4100 = (g113&g3648);
assign II5528 = ((~g43));
assign g6013 = (g5589&g2424);
assign II13903 = ((~g7357));
assign II14603 = ((~g7827));
assign II12481 = ((~g6616));
assign II8064 = (g3316&g3287&g3264&g1987);
assign II14457 = ((~g8093));
assign g7000 = ((~II12742));
assign g7212 = (g1053&g7010);
assign g4958 = (g296&g3897);
assign g4625 = ((~II8790));
assign g1918 = ((~g822));
assign II11311 = ((~g5760));
assign g4837 = (g2573&g2562&II9202);
assign II6273 = ((~g840))|((~g906));
assign II15019 = (g7951)|(g7920)|(g7983)|(g8181);
assign g8315 = (g4544&g7993);
assign g2653 = ((~II6443));
assign g9129 = ((~II15765));
assign g6021 = (g5594&g2424);
assign II10982 = ((~g2210))|((~II10980));
assign g8959 = ((~II15391));
assign II16151 = ((~g9369));
assign g1773 = ((~g610));
assign g7616 = (g7367&g4517);
assign g4832 = (g1110&g4246);
assign II15329 = ((~g8793));
assign g6796 = ((~II12259));
assign g2956 = ((~g2375));
assign g4385 = (g300&g3131);
assign g7359 = ((~II13493));
assign g3867 = ((~g2946));
assign g3893 = ((~II7453))|((~II7454));
assign II8895 = ((~g4130));
assign II9177 = ((~g4299));
assign g5452 = (g4876&g3499);
assign II11890 = ((~g6135));
assign g6276 = ((~II11116))|((~II11117));
assign g1578 = ((~g699));
assign g4372 = ((~II8357));
assign g4004 = ((~g2845));
assign II13828 = ((~g7321));
assign g9174 = (g9147)|(g8963);
assign g6475 = ((~II11633));
assign g6118 = ((~g5549));
assign II8715 = ((~g3903));
assign II13663 = ((~g7235));
assign g6829 = ((~II12358));
assign II13897 = ((~g7354));
assign g8874 = ((~II15208));
assign g7602 = (g7476&g3466);
assign II5559 = ((~g1292));
assign II6939 = ((~g2161))|((~g2051));
assign g7163 = ((~II13063));
assign g5058 = ((~II9416));
assign g2384 = ((~II6254));
assign g7428 = (g6040)|(g7175);
assign g6124 = (g5432)|(g4789);
assign II15726 = ((~g9069));
assign g6382 = ((~II11473));
assign II6728 = ((~g1959));
assign II13045 = ((~g6955));
assign II8665 = ((~g3051));
assign II15054 = (g8363)|(g8342)|(g8407)|(g8386);
assign g6379 = ((~II11464));
assign g2752 = ((~g2389));
assign g3340 = ((~g2474));
assign g7080 = (g4086)|(g6462);
assign g4553 = ((~g2891));
assign g7190 = ((~II13112));
assign II15784 = ((~g9125));
assign g6198 = ((~g5335));
assign g6815 = ((~II12316));
assign g2774 = ((~g1813));
assign g3777 = ((~g2170));
assign g3969 = ((~g3192));
assign g9339 = (g9259)|(g9335);
assign g7244 = ((~g7050))|((~g3757))|((~g3739));
assign g5140 = (g4333)|(g3509);
assign g4700 = ((~g2460))|((~g4271));
assign g7062 = (g4048)|(g6456);
assign g6741 = ((~II12117));
assign g3190 = (g1658&g2424);
assign g9186 = ((~II15836));
assign g6830 = ((~II12361));
assign g8777 = (II14969)|(II14970);
assign II15723 = ((~g9065));
assign g1679 = ((~II5512));
assign g2881 = ((~g2235));
assign g2533 = ((~g1336));
assign g4380 = (g584&g2845);
assign g8747 = ((~g8545));
assign g6483 = ((~II11645));
assign g4546 = (g2643&g746);
assign g5045 = (g293&g3961);
assign g9086 = ((~II15648));
assign g3633 = ((~II7104));
assign g6931 = (g6416)|(g6421);
assign II16165 = ((~g9377));
assign g6839 = ((~II12388));
assign g6228 = ((~II11021));
assign II8114 = (g2162&g2149&g2137&g2106);
assign g5649 = ((~g4748));
assign II7255 = ((~g1955));
assign g3232 = ((~g2298))|((~g2276));
assign II15018 = (g7855)|(g7838)|(g7905)|(g7870);
assign g9113 = ((~II15729));
assign g9223 = ((~II15943));
assign g8821 = (g339&g8545);
assign g8826 = (g420&g8564);
assign g4220 = (g3533&g3549&g3568&g3583);
assign g2645 = ((~II6419));
assign II6291 = ((~g46));
assign II10197 = ((~g4724))|((~II10196));
assign g5070 = (g4052)|(g4058);
assign g1838 = ((~g1450));
assign g8523 = ((~g7658)&(~g7616)&(~g8082)&(~g7634));
assign g8802 = ((~II15014));
assign II14202 = ((~g7708));
assign II12643 = ((~g6501));
assign II11178 = ((~g5466))|((~II11177));
assign II8133 = ((~g3232))|((~II8132));
assign g7197 = (g7093&g5055);
assign g3876 = ((~g3466));
assign g1011 = ((~II5413));
assign g3498 = ((~g1616));
assign II11873 = ((~g2543))|((~g6187));
assign II14795 = ((~g8604));
assign II14012 = ((~g7438));
assign g7745 = ((~II14106));
assign g8563 = ((~II14662));
assign g5256 = (g5119)|(g4454);
assign II13979 = ((~g7415));
assign II9369 = ((~g3901));
assign II15601 = ((~g8992));
assign g5165 = ((~II9621));
assign g6189 = ((~II10930));
assign g4456 = ((~II8471))|((~II8472));
assign II11722 = ((~g5772));
assign II12295 = ((~g6693));
assign II9158 = ((~g4256));
assign g8806 = ((~g8443)&(~g8421)&(~II15044));
assign II7495 = ((~g3562));
assign II12205 = ((~g6488));
assign g7426 = (g1173)|(g7217)|(II13553);
assign g3735 = ((~g1961));
assign II9884 = ((~g4868));
assign g2497 = ((~g945));
assign g2971 = ((~II6723));
assign g8720 = (g3825&g8421);
assign II11194 = ((~g6243));
assign II10969 = ((~g5606));
assign g5741 = ((~II10280));
assign II5425 = ((~g1245));
assign II8859 = ((~g3968));
assign II6183 = ((~g6));
assign g1663 = ((~g1416));
assign g6704 = ((~II12044));
assign II13457 = ((~g7120));
assign g4914 = ((~g4093));
assign II15638 = ((~g8978));
assign II7981 = ((~g3555));
assign II6198 = ((~g483));
assign g5584 = ((~g4841));
assign g3191 = ((~II6868));
assign g1803 = ((~g758));
assign g1577 = ((~g695));
assign g8619 = ((~II14695));
assign g7164 = ((~II13066));
assign II9484 = ((~g3957));
assign g8670 = ((~II14804));
assign g8718 = (g2774&g8386);
assign II12854 = ((~g6695))|((~II12852));
assign II13846 = ((~g7487));
assign g6133 = ((~II10766));
assign II7104 = ((~g2479));
assign g7825 = (g4801)|(g7615);
assign g6913 = (g6733)|(g6738);
assign g1796 = ((~g617));
assign g2268 = ((~II6009));
assign II12598 = ((~g1126))|((~II12596));
assign g4257 = ((~II8190));
assign II15915 = ((~g9194));
assign II14400 = ((~g7677));
assign II8865 = ((~g4032));
assign g4598 = ((~II8709));
assign g4681 = (g4255&g3533);
assign g3504 = ((~g1375)&(~g2229)&(~g2213)&(~g2206));
assign g6439 = (g789&g6150);
assign II15083 = (g7855)|(g7838)|(g7905)|(g7870);
assign g9345 = (g9330&g6217);
assign II13816 = ((~g7455));
assign g9310 = ((~II16046));
assign II13997 = ((~g7432));
assign g6213 = ((~II10976));
assign g2474 = ((~g1405))|((~g1412));
assign II12639 = ((~g6506));
assign g4371 = ((~II8354));
assign g7234 = ((~g3757))|((~g3739))|((~g7050))|((~g3770));
assign II14088 = ((~g7585));
assign g4227 = ((~II8133))|((~II8134));
assign II11736 = ((~g6076));
assign II11025 = ((~g5638));
assign g4819 = (g2573&g2562&II9166);
assign g4327 = (g2959&g1867);
assign II5505 = ((~g1532))|((~g1528));
assign g4701 = ((~II8994));
assign II13122 = ((~g7070));
assign g4536 = ((~g2877));
assign g3341 = ((~II6936));
assign II15622 = ((~g8999));
assign g2826 = ((~g2183));
assign II9528 = ((~g4006));
assign g3488 = ((~g1727));
assign II13912 = ((~g7359));
assign II7680 = ((~g2712));
assign II7064 = ((~g2458));
assign II10875 = ((~g2595))|((~II10873));
assign g6844 = ((~II12403));
assign g6893 = ((~II12551))|((~II12552));
assign II12924 = ((~g6983));
assign II10835 = ((~g5514))|((~II10834));
assign g5128 = ((~II9528));
assign II7126 = ((~g2494));
assign II16173 = ((~g9382));
assign II14480 = (g7937)|(g7887)|(g8029)|(g8018);
assign II15619 = ((~g8998));
assign II14211 = ((~g7712));
assign g2934 = ((~II6676));
assign g1967 = ((~g1432));
assign g6618 = ((~g6003));
assign g4335 = ((~g3659));
assign g5745 = ((~II10292));
assign g5061 = ((~II9425));
assign g9091 = ((~II15663));
assign II11939 = ((~g6015));
assign g8945 = (g4541&g8784);
assign II11978 = ((~g6186));
assign II14338 = ((~g7581));
assign g4195 = ((~II8094));
assign II9005 = ((~g4585));
assign g2929 = ((~g2327));
assign g7254 = (g6923)|(g5298);
assign g3513 = ((~g2407));
assign g7305 = ((~II13347));
assign II5362 = ((~g3841));
assign g8764 = (g8231&g4969);
assign g2939 = ((~g2348));
assign g8967 = ((~II15405));
assign g7512 = ((~II13716));
assign g2275 = ((~g990));
assign g9038 = (g8966&g5345);
assign g8631 = ((~II14709));
assign g7566 = ((~g7421)&(~g1597));
assign II9347 = ((~g3896));
assign II15242 = (g8697)|(g8714)|(g8718)|(g8719);
assign II15291 = (g8331)|(g8336)|(g8338)|(g8688);
assign g6057 = (g1061&g5617);
assign g6729 = ((~g6263));
assign g8562 = ((~g8094));
assign g7354 = ((~II13478));
assign II11156 = ((~g5482))|((~g3052));
assign g6504 = ((~g5269))|((~g5874));
assign g6571 = ((~II11758))|((~II11759));
assign g1682 = ((~II5520))|((~II5521));
assign g7654 = (g7367&g4142);
assign g5786 = ((~II10403));
assign g2208 = ((~II5923));
assign g2818 = ((~g1792));
assign g6447 = (g734&g6073);
assign g5807 = ((~II10454));
assign g8511 = ((~II14646));
assign g6321 = ((~II11290));
assign II11043 = ((~g5648));
assign II8338 = ((~g2966))|((~g1698));
assign g7110 = ((~II12918));
assign g1872 = (g971)|(g962)|(g972)|(II5757);
assign II13112 = ((~g7021));
assign g5233 = (g5089)|(g4420);
assign g5222 = (g5068)|(g4397);
assign II7609 = ((~g2471))|((~g3771));
assign g2916 = ((~II6646));
assign II11136 = ((~g5476))|((~II11135));
assign g6486 = ((~II11648));
assign II10347 = ((~g5706));
assign g9062 = ((~II15580));
assign II13861 = ((~g7330));
assign g6206 = ((~g5639));
assign II7788 = ((~g2595));
assign II9907 = ((~g4837));
assign g5076 = ((~II9446));
assign II11186 = ((~g3029))|((~II11184));
assign II15284 = (g8335)|(g8340)|(g8290)|(g8691);
assign g4349 = ((~g2496)&(~g3310));
assign g7546 = ((~II13822));
assign II7545 = ((~g3589));
assign g3644 = ((~g2131));
assign g1935 = ((~g1280));
assign II13092 = ((~g7047));
assign II13099 = ((~g7054));
assign g3522 = ((~g2407));
assign g3929 = ((~II7588));
assign II14662 = ((~g7783));
assign II5954 = ((~g89));
assign II15672 = ((~g9047));
assign g8310 = (g573&g8181);
assign II7662 = ((~g3642));
assign II12304 = ((~g6711));
assign g7001 = (g3722&g6562);
assign g8795 = (g8151)|(g8077)|(g8075)|(g8279);
assign g5001 = (g458&g3912);
assign g3857 = ((~II7374));
assign g5171 = ((~II9639));
assign g8960 = ((~II15394));
assign g8338 = (g570&g8181);
assign g3837 = ((~II7314));
assign g1569 = ((~g661));
assign II14951 = (g8328)|(g8316)|(g8455)|(g8378);
assign II14245 = ((~g7683))|((~II14244));
assign II13894 = ((~g7353));
assign II11835 = ((~g6181));
assign g3905 = ((~g3192));
assign II7973 = ((~g3071));
assign g3989 = ((~g3131));
assign g9108 = ((~II15714));
assign g7633 = ((~II13962));
assign g8333 = (g563&g8181);
assign II12373 = ((~g6763));
assign g738 = ((~II5404));
assign g2908 = ((~g2290));
assign g8623 = (g755&g8199);
assign II12829 = ((~g6441));
assign g2293 = ((~g888));
assign g8276 = (g150&g8042);
assign II15657 = ((~g9059));
assign g6765 = ((~II12164));
assign g3842 = ((~II7329));
assign g8295 = (g4512&g7905);
assign g4353 = ((~g3665));
assign g6824 = ((~II12343));
assign II7211 = ((~g1742));
assign g8797 = ((~II15003));
assign II15388 = ((~g8898));
assign g7067 = ((~g6658));
assign II14646 = ((~g7790));
assign II7752 = ((~g3591));
assign g6870 = ((~II12481));
assign II7611 = ((~g3771))|((~II7609));
assign II6998 = ((~g2242))|((~II6996));
assign g8639 = ((~II14725));
assign II14420 = ((~g7554));
assign II6323 = ((~g1342));
assign g5468 = ((~II9884));
assign g8066 = (g7488&g7634);
assign II7838 = ((~g2781));
assign g4006 = ((~II7749));
assign g9199 = ((~g9188));
assign II11803 = ((~g6280));
assign II7618 = ((~g1721))|((~II7616));
assign II5676 = ((~g911));
assign g8581 = ((~g8094));
assign g5208 = (g5043)|(g4383);
assign II11143 = ((~g5493))|((~II11142));
assign II6924 = ((~g1728))|((~II6923));
assign g5642 = ((~II10125));
assign II12268 = ((~g6661));
assign g4511 = ((~g2841));
assign g2892 = ((~g2266));
assign g7315 = ((~II13373));
assign g7285 = ((~II13287));
assign II7443 = ((~g2973))|((~g1701));
assign g9081 = ((~II15635));
assign g5112 = ((~II9496));
assign g2020 = ((~II5855));
assign g7497 = ((~II13669));
assign g4017 = ((~g2845));
assign g7683 = (g1061&g7429);
assign II8552 = (g3316&g2057&g3264&g1987);
assign II11422 = ((~g5842));
assign g3971 = ((~II7688));
assign g9098 = ((~II15684));
assign g2096 = ((~g1226));
assign II9549 = ((~g4307))|((~II9547));
assign II7314 = ((~g2916));
assign g7480 = ((~II13639))|((~II13640));
assign g5813 = ((~II10472));
assign II15708 = ((~g9072));
assign g2743 = ((~g1808));
assign g7275 = ((~II13261));
assign II14848 = ((~g8625));
assign II15856 = ((~g9168))|((~II15855));
assign g8924 = (g4588&g8752);
assign g4430 = (II8436&II8437);
assign II11001 = ((~g5698));
assign g4265 = ((~g3591));
assign g9021 = (g8886&g5317);
assign g8783 = ((~g8524));
assign II13185 = ((~g7020));
assign g7732 = ((~II14067));
assign g5670 = ((~II10157));
assign g4920 = ((~g4105));
assign g8984 = (g8924)|(g8822);
assign II8977 = ((~g3877));
assign g7628 = (g7367&g4532);
assign II12337 = ((~g6724));
assign g2073 = ((~g1254));
assign g5594 = ((~II10072))|((~II10073));
assign g4287 = (g3563&g2334&g3579&II8237);
assign g6313 = ((~II11266));
assign g1889 = ((~g1018));
assign g8711 = (g3542&g8407);
assign II10283 = ((~g5643));
assign g5836 = ((~g5529));
assign II14070 = ((~g7714));
assign II6887 = ((~g2528));
assign II11645 = ((~g5874));
assign II6553 = ((~g2246));
assign gbuf49 = (g1185);
assign g9378 = ((~II16158));
assign g2323 = ((~II6112));
assign g6172 = (g1514&g5192);
assign g9213 = ((~II15915));
assign II11236 = ((~g6148));
assign g8628 = (g753&g8199);
assign g4500 = ((~g2832));
assign g8762 = ((~g8585));
assign II7383 = ((~g3465));
assign g9183 = ((~g9161));
assign g5603 = ((~g4938));
assign g8662 = ((~II14780));
assign g7140 = ((~II13003))|((~II13004));
assign g6956 = ((~II12669));
assign g4399 = ((~II8393))|((~II8394));
assign g7224 = ((~II13164));
assign g6650 = ((~g6213));
assign II13432 = ((~g7280));
assign g5077 = (g236&g3988);
assign g6621 = ((~II11855));
assign g7753 = ((~II14130));
assign g3542 = ((~g1777));
assign II7268 = ((~g2486))|((~g955));
assign g5738 = ((~II10271));
assign II12976 = ((~g6928));
assign g2834 = ((~II6564));
assign g8260 = (g138&g8111);
assign g7344 = ((~g7150));
assign II11522 = ((~g5847));
assign g1586 = ((~g730));
assign II15845 = ((~g9174));
assign g6243 = ((~II11050));
assign g4690 = (g4081&g3078);
assign g6751 = ((~II12128));
assign g7835 = ((~II14257));
assign II11842 = ((~g2548))|((~II11841));
assign g5529 = ((~g4689));
assign II6033 = ((~g3));
assign g2995 = ((~II6740))|((~II6741));
assign g6693 = ((~II12011));
assign g6468 = ((~II11622));
assign g8918 = ((~II15340));
assign g7141 = ((~II13009));
assign II12003 = ((~g6202));
assign II10874 = ((~g5516))|((~II10873));
assign g8997 = (g8937)|(g8841);
assign II7697 = ((~g3052));
assign g9376 = ((~II16154));
assign II6820 = ((~g1707));
assign g4609 = ((~II8742));
assign II13329 = ((~g7247));
assign II12684 = ((~g6472));
assign g3815 = ((~g1822));
assign II13773 = ((~g7496));
assign g6673 = (g4053)|(g5937);
assign II13687 = ((~g7237))|((~II13685));
assign gbuf18 = (g1203);
assign II9021 = ((~g4489));
assign g2555 = ((~g936));
assign II7233 = (g2315)|(g2385)|(g2294)|(g2395);
assign g6842 = ((~II12397));
assign g8602 = ((~g8094));
assign g8233 = ((~g8199)&(~II14484)&(~II14485));
assign II8000 = (g3430&g3398&g3359&g3341);
assign g6968 = ((~II12699));
assign g7362 = ((~II13502));
assign II11961 = ((~g5988));
assign II14925 = ((~g8381));
assign II14933 = (g8385)|(g8404)|(g8441)|(g8462);
assign g2845 = (g1877)|(g576);
assign g7145 = ((~II13023));
assign II7098 = ((~g2477));
assign II9978 = ((~g4880))|((~g2092));
assign II12161 = ((~g5971));
assign g4561 = ((~g2900));
assign g6514 = ((~II11696));
assign g5201 = (g5030)|(g4376);
assign g6151 = (g1494&g5709);
assign II7944 = ((~g3774));
assign II7575 = ((~g2999))|((~II7574));
assign g4558 = ((~g2897));
assign g2751 = ((~II6500))|((~II6501));
assign g8930 = (g3866&g8760);
assign g4895 = ((~g4078));
assign g6361 = ((~II11410));
assign g9008 = (g8948)|(g8857);
assign g372 = ((~II5359));
assign II7804 = ((~g3029));
assign g2505 = ((~g28));
assign g2721 = ((~g1803));
assign g3502 = ((~g1616));
assign g9320 = ((~g9307));
assign g7047 = ((~g6498));
assign II9209 = ((~g4349));
assign g1733 = (g1489&g1481);
assign II15765 = ((~g9039));
assign II11129 = ((~g5418));
assign g9142 = (g9124&g6059);
assign II10901 = ((~g2752))|((~II10899));
assign g9194 = ((~g9182));
assign g6644 = ((~g6208));
assign g6886 = ((~II12529));
assign g9120 = (g9052&g5345);
assign g7071 = (g6639&g1872);
assign g6168 = (g1138&g5191);
assign II10009 = ((~g1949))|((~g4821));
assign g5059 = ((~II9419));
assign II13347 = ((~g7224));
assign II12135 = ((~g5988));
assign II12782 = ((~g6463));
assign gbuf66 = (g576);
assign II11344 = ((~g5820));
assign g2897 = ((~g2270));
assign g9234 = ((~II15956));
assign g2924 = ((~g2314));
assign g5434 = ((~g5112));
assign g4795 = ((~II9116));
assign II13035 = ((~g6964));
assign g8342 = ((~g8008));
assign II12655 = ((~g6458));
assign g2272 = ((~II6021));
assign g9327 = (g9316&g5757);
assign g6705 = (g6157)|(g5583);
assign II6286 = ((~g1307));
assign g5193 = (g5017)|(g4366);
assign g8790 = ((~g8585));
assign g6436 = (g6266)|(g5699);
assign g4783 = (g948&g4527);
assign II13338 = ((~g7190));
assign II7277 = ((~g2497))|((~g1898));
assign g2777 = ((~g1797));
assign II11096 = ((~g2734))|((~II11094));
assign g5575 = ((~II10039))|((~II10040));
assign g6345 = ((~II11362));
assign g2460 = ((~II6302));
assign g2229 = (g1371)|(g1372)|(g1373)|(g1374);
assign II15530 = ((~g8972));
assign II11452 = ((~g6071));
assign II8826 = ((~g4023));
assign g1677 = ((~g1532));
assign II12866 = ((~g6483));
assign g4492 = ((~II8537))|((~II8538));
assign II12517 = ((~g6613));
assign II8877 = ((~g4274));
assign g4663 = ((~II8904));
assign g8282 = (g179&g8156);
assign g6014 = ((~II10614));
assign g1744 = ((~g600));
assign II7347 = ((~g2985));
assign g6659 = ((~II11955));
assign g5260 = (g5123)|(g4473);
assign II7485 = ((~g2989))|((~g1708));
assign II14019 = ((~g7480));
assign g4306 = ((~II8273));
assign g2866 = ((~g2221));
assign II15735 = ((~g9078));
assign II13388 = ((~g7149));
assign g2484 = ((~g45));
assign g7723 = ((~II14042));
assign g6329 = ((~II11314));
assign g5628 = ((~g4748));
assign g4575 = ((~II8679))|((~II8680));
assign g7327 = ((~II13403));
assign g7139 = ((~II12999));
assign g4501 = ((~g2801));
assign II14145 = ((~g7542));
assign II13613 = ((~g7273));
assign II8581 = ((~g2498))|((~g2777));
assign II14172 = ((~g7545));
assign g7039 = ((~g6543));
assign g4889 = ((~II9242))|((~II9243));
assign II7856 = ((~g3805));
assign II7814 = ((~g2605));
assign g4512 = ((~g2842));
assign g8175 = ((~II14406));
assign II10719 = ((~g5559));
assign g6287 = ((~II11185))|((~II11186));
assign g6859 = ((~II12448));
assign g3496 = ((~II6974));
assign g1896 = ((~g86));
assign g5129 = ((~II9531));
assign g7598 = (g7483&g3466);
assign g5822 = ((~II10491));
assign g4825 = (g4228&g1964);
assign g6715 = (g677&g5843);
assign g7205 = ((~II13131));
assign g4622 = ((~II8781));
assign g4422 = (g411&g3160);
assign g5052 = (g4049)|(g4054);
assign g7591 = ((~II13918));
assign II7925 = ((~g2761));
assign II10758 = ((~g5662));
assign g4010 = ((~g3097));
assign II13704 = ((~g7352));
assign II7492 = ((~g3561));
assign g9259 = (g9230&g5639);
assign g8510 = ((~II14643));
assign g5612 = ((~g4814));
assign g6863 = ((~II12460));
assign II15417 = ((~g8893));
assign II10561 = ((~g5265));
assign g5444 = ((~g5074));
assign g4922 = ((~g4111));
assign g4706 = ((~II9005));
assign g2768 = (g1597&g973);
assign II14436 = ((~g7904));
assign II12881 = ((~g6478));
assign II11750 = ((~g6112))|((~g1486));
assign II9360 = ((~g4257));
assign g5148 = ((~II9570));
assign g7587 = ((~II13906));
assign II5616 = ((~g979));
assign g7520 = ((~II13740));
assign II14106 = ((~g7586));
assign II12571 = ((~g6729));
assign g3091 = ((~g1603));
assign g4584 = ((~g3466));
assign g3259 = (g1976&g1960);
assign g7855 = ((~II14267));
assign g3540 = ((~g2424));
assign II13755 = ((~g7317));
assign II13344 = ((~g7210));
assign g4065 = ((~II7838));
assign II14657 = ((~g7782));
assign g5179 = ((~II9663));
assign g6299 = ((~II11224));
assign g8800 = ((~II15010));
assign g4239 = (g1541&g3222);
assign II12403 = ((~g6769));
assign g5757 = ((~g5261));
assign g5475 = (g3801&g5022);
assign g8677 = ((~II14825));
assign II8015 = (g2074&g2057&g3264&g3238);
assign II5471 = ((~g1029));
assign II15228 = (g8270)|(g8258)|(g8281)|(g8273);
assign g8041 = ((~g7701));
assign II10072 = ((~g4954))|((~II10071));
assign g3769 = ((~g2548));
assign g6258 = ((~g5427));
assign g7079 = (g4259&g6677);
assign II12646 = ((~g6493));
assign g8901 = (g8804&g5631);
assign II12939 = ((~g7022));
assign II9034 = ((~g4317));
assign g4630 = ((~II8805));
assign II13493 = ((~g7132));
assign II12484 = ((~g6621));
assign g5545 = (g3617)|(g4824);
assign II8327 = ((~g2011))|((~II8326));
assign g5737 = ((~II10268));
assign g5956 = ((~II10582));
assign g5199 = ((~g4841));
assign g5812 = ((~II10469));
assign g6623 = ((~II11861));
assign II7987 = ((~g3528));
assign g1557 = ((~II5432));
assign g6262 = (g4074)|(g5334);
assign g6184 = ((~g875)&(~g5291));
assign g3681 = ((~g866))|((~g2368));
assign g4882 = ((~g4069));
assign II7486 = ((~g2989))|((~II7485));
assign II13628 = ((~g7248));
assign II7540 = ((~g1715))|((~II7538));
assign g6231 = ((~II11028));
assign g8765 = ((~g8524));
assign g5780 = ((~II10387));
assign g3914 = ((~II7532))|((~II7533));
assign g7456 = ((~g7174));
assign g2359 = ((~g1397));
assign g2330 = ((~II6134))|((~II6135));
assign II15231 = (g8701)|(g8715)|(g8730)|(g8720);
assign II13140 = ((~g6954));
assign g6123 = (g3617)|(g5556);
assign g6592 = ((~II11790));
assign II11443 = ((~g6038));
assign g4365 = (g237&g3097);
assign g6681 = ((~II11991));
assign g5568 = ((~g2044))|((~g4902))|((~g4320));
assign g6171 = (g5363&g4841);
assign II9425 = ((~g3917));
assign g6336 = ((~II11335));
assign g4228 = ((~g1408))|((~g2665));
assign g7534 = ((~II13782));
assign g7529 = ((~II13767));
assign II8205 = ((~g2655));
assign g6776 = ((~II12199));
assign g4491 = (g557&g2845);
assign II14831 = (g8483)|(g8464)|(g8514);
assign g3913 = ((~g2834));
assign g3678 = ((~II7173))|((~II7174));
assign g7263 = ((~II13231));
assign II12011 = ((~g5939));
assign g8296 = (g351&g7870);
assign g6179 = ((~II10896));
assign g9185 = ((~II15833));
assign g7522 = ((~II13746));
assign g8542 = (g661&g7887);
assign II11386 = ((~g5764));
assign II5577 = ((~g172));
assign g6798 = ((~II12265));
assign g1724 = ((~II5568));
assign II16046 = ((~g9288));
assign g6692 = ((~II12008));
assign g5207 = ((~g4673));
assign II12253 = ((~g6427));
assign g8965 = (g8739)|(g8742)|(g8914)|(g8847);
assign g9367 = ((~II16129));
assign g5219 = (g5065)|(g4394);
assign g1923 = ((~II5801));
assign g6056 = (g3760&g5286&g1695);
assign g6489 = ((~g5802)&(~g5769)&(~g5790));
assign II11215 = ((~g6156));
assign g5344 = ((~II9819));
assign g5164 = ((~II9618));
assign g2900 = ((~g2273));
assign g6901 = ((~g6525));
assign g6687 = ((~II12003));
assign g2728 = ((~g2256));
assign g2057 = ((~II5868));
assign g9387 = (g9349)|(g9384);
assign g4826 = (g1545&g4239);
assign II13365 = ((~g7267));
assign g8074 = (g855&g7616);
assign g7769 = ((~II14178));
assign g5050 = (g587&g3970);
assign II13512 = ((~g7138));
assign II12834 = ((~g6709))|((~II12832));
assign g5184 = ((~II9678));
assign g5794 = ((~II10421));
assign g3861 = ((~II7386));
assign II11488 = ((~g6034));
assign g7296 = ((~II13320));
assign g9299 = ((~II16023));
assign g4128 = (g98&g3693);
assign g6380 = ((~II11467));
assign g1869 = ((~g74));
assign g8699 = ((~g7658)&(~g8613)&(~g7634));
assign g3939 = ((~II7617))|((~II7618));
assign II13541 = ((~g7209));
assign II14732 = ((~g8155));
assign II12909 = ((~g7046));
assign II10976 = ((~g5726));
assign g4354 = ((~g1424)&(~g3541));
assign II9985 = ((~g4836))|((~g2096));
assign II15927 = ((~g9208));
assign g6107 = (g5478&g1849);
assign g4117 = (g2626&g2616);
assign g8381 = ((~II14603));
assign g8111 = ((~II14374));
assign g7159 = ((~II13051));
assign II10925 = ((~g2752))|((~II10923));
assign g9022 = (g8887&g5317);
assign II14022 = ((~g7443));
assign II13734 = ((~g7422));
assign II14397 = ((~g7686));
assign g7235 = (g6699&g7094);
assign g7101 = ((~II12891));
assign g1894 = ((~II5772));
assign g8861 = ((~g8493)&(~g8239)&(~II15169));
assign g8666 = ((~II14792));
assign gbuf50 = (g1163);
assign g6158 = ((~g3735))|((~g3716))|((~g5633))|((~g3754));
assign II15830 = ((~g9180));
assign II12561 = ((~g6449));
assign g5521 = ((~g4929));
assign g7038 = (g6466&g4841);
assign II6012 = ((~g384));
assign g8983 = (g8923)|(g8821);
assign II15423 = ((~g8894));
assign II10271 = ((~g5487));
assign g4714 = ((~g4344))|((~g4335))|((~g4328));
assign g6330 = ((~II11317));
assign g6295 = ((~II11212));
assign g2650 = ((~II6434));
assign g4379 = (g399&g3160);
assign g4677 = ((~II8932));
assign II6368 = ((~g20));
assign II11281 = ((~g5785));
assign g5488 = ((~II9910));
assign II7538 = ((~g2996))|((~g1715));
assign g6974 = (g3613&g6505);
assign II5545 = ((~g1276));
assign g9273 = (g4748&g9252);
assign g5152 = ((~II9582));
assign g9069 = ((~II15601));
assign g3932 = ((~II7595));
assign II8820 = ((~g3952));
assign g5734 = ((~II10259));
assign g4617 = ((~II8766));
assign g6190 = ((~II10933));
assign g4123 = (g2627&g2617);
assign g4169 = (II8052&II8053);
assign II8071 = (g2162&g2149&g2137&g2106);
assign II12391 = ((~g6744));
assign II12167 = ((~g5939));
assign II12078 = ((~g5988))|((~g5971));
assign g6312 = ((~II11263));
assign g4797 = (g3893&g1616);
assign g4724 = (g828&g4038);
assign g2618 = ((~g1566));
assign g8280 = (g114&g8111);
assign II14822 = ((~g8649));
assign II8617 = (g3430&g3398&g3359&g2106);
assign g2525 = ((~II6354));
assign II13915 = ((~g7360));
assign g2242 = ((~g985));
assign II15072 = (g7855)|(g7838)|(g7905)|(g7870);
assign g5714 = (g1532&g4733);
assign g4059 = (g1499&g2979);
assign g5060 = ((~II9422));
assign g8937 = (g4524&g8770);
assign g5824 = ((~II10497));
assign g8225 = ((~II14454));
assign g2695 = ((~g1672));
assign II11920 = ((~g5874));
assign g4187 = (II8078&II8079);
assign II15580 = ((~g8985));
assign g6657 = ((~II11951));
assign II8889 = ((~g4311));
assign II5377 = ((~g635));
assign g4548 = ((~II8636))|((~II8637));
assign II13403 = ((~g7269));
assign g7351 = ((~II13469));
assign II14789 = ((~g8544));
assign g8012 = ((~II14305));
assign g6357 = ((~II11398));
assign II7389 = ((~g3496));
assign II16154 = ((~g9370));
assign g8756 = ((~g8564));
assign II8574 = (g3316&g2057&g2020&g3238);
assign g3630 = ((~II7095));
assign g3852 = ((~II7359));
assign g8313 = (g4542&g7951);
assign II6232 = ((~g834))|((~g896));
assign II11251 = ((~g6152));
assign g5988 = ((~II10592));
assign g5744 = ((~II10289));
assign g9148 = (g9143)|(g9024);
assign g6645 = ((~II11917));
assign II12068 = ((~g5847));
assign II10180 = ((~g4721));
assign gbuf53 = (g1186);
assign g6984 = ((~II12725));
assign g4624 = ((~II8787));
assign g5576 = ((~g4894))|((~g4888))|((~g4884));
assign g1832 = ((~g763));
assign g7170 = (g6916)|(g6444);
assign II12181 = ((~g6163))|((~II12179));
assign g8903 = ((~II15315));
assign II11559 = ((~g6065));
assign g3187 = ((~II6860));
assign g8316 = (g513&g7966);
assign g6892 = ((~II12547));
assign g3770 = ((~g2551));
assign g6023 = ((~II10626))|((~II10627));
assign g2624 = ((~g1569));
assign II15850 = ((~g9154))|((~II15848));
assign g5265 = (g5126)|(g4491);
assign II12592 = ((~g1008));
assign g4001 = ((~g3160));
assign g2686 = ((~g1667));
assign g9000 = (g8940)|(g8845);
assign g9264 = (g9247)|(g6242);
assign II9419 = ((~g3916));
assign II10889 = ((~g5590))|((~II10888));
assign g8722 = (g2787&g8386);
assign g6400 = (g150&g6011);
assign g4305 = ((~g3712))|((~g3700))|((~g3732));
assign II10397 = ((~g5200));
assign II16100 = ((~g9338));
assign g7418 = ((~II13533));
assign g7338 = ((~II13432));
assign g5018 = (g232&g3930);
assign II7356 = ((~g2843));
assign g7081 = (g6172)|(g6629);
assign g2659 = ((~g1655));
assign II13873 = ((~g7342));
assign II5552 = ((~g1284));
assign II5359 = ((~g3839));
assign II15007 = ((~g8627));
assign g2870 = ((~g2225));
assign II7371 = ((~g3050));
assign g4599 = ((~II8712));
assign g9285 = (g9271)|(g6221);
assign II10608 = ((~g5701));
assign g2496 = ((~g942));
assign g3512 = ((~g1616));
assign g7241 = ((~II13185));
assign II8892 = ((~g4115));
assign g3993 = ((~g3192));
assign II14763 = ((~g7834));
assign g7229 = ((~g6938));
assign g9012 = (g8908&g8239);
assign g7494 = ((~g7260));
assign g6316 = ((~II11275));
assign g7211 = ((~II13147));
assign g6635 = ((~II11897));
assign II10256 = ((~g5401));
assign II10888 = ((~g5590))|((~g2259));
assign g5551 = ((~II9974));
assign g4684 = ((~II8949));
assign g6012 = ((~g5367));
assign g6957 = ((~II12672));
assign II9561 = ((~g4695));
assign g7044 = ((~g6543));
assign II12675 = ((~g6510));
assign g6555 = ((~II11729));
assign II12187 = ((~g5897));
assign g3539 = ((~g2424));
assign II13746 = ((~g7311));
assign g4386 = (g324&g3131);
assign II8537 = ((~g2506))|((~II8536));
assign g7577 = ((~II13876));
assign g6115 = (g3617)|(g5558);
assign II6363 = ((~g16));
assign II7504 = ((~g2498))|((~II7503));
assign g9121 = ((~II15747));
assign g4838 = (g4517&g1760);
assign g4146 = ((~II8011));
assign g6926 = (g6406)|(g6411);
assign II6457 = ((~g1886));
assign g4477 = ((~II8517));
assign g7097 = ((~II12881));
assign g6280 = ((~II11136))|((~II11137));
assign g4373 = ((~II8360));
assign II6437 = ((~g1784));
assign g2333 = ((~g985))|((~g990));
assign g5698 = (g5057)|(g5040);
assign g4420 = (g275&g3097);
assign g3533 = ((~g2397));
assign II10469 = ((~g5222));
assign g6877 = ((~II12502));
assign g8831 = (g423&g8564);
assign II15897 = ((~g9202))|((~g9203));
assign g9191 = ((~II15856))|((~II15857));
assign g5939 = ((~II10579));
assign g4552 = ((~g2890));
assign g3957 = ((~II7662));
assign II10169 = ((~g4873));
assign g7427 = (g1472&g7199);
assign g8742 = (g2973&g8493);
assign g2955 = ((~II6703));
assign g7601 = ((~g7450));
assign gbuf74 = (g911);
assign g9331 = ((~g9321));
assign g5724 = ((~g4969));
assign g4543 = ((~g2885));
assign g5057 = (g3939)|(g3925)|(g3915)|(g3907);
assign g4736 = (g4532)|(g4517)|(II9044);
assign g6795 = ((~II12256));
assign g2824 = ((~g1688));
assign g6277 = ((~II11123))|((~II11124));
assign II7640 = ((~g3062));
assign II11050 = ((~g5335));
assign g1718 = ((~II5562));
assign g7065 = ((~II12833))|((~II12834));
assign g3287 = ((~II6911));
assign g9042 = ((~II15530));
assign II5855 = ((~g71));
assign g2385 = ((~II6258))|((~II6259));
assign II12699 = ((~g6504));
assign II13131 = ((~g6951));
assign II12757 = ((~g6577));
assign II6523 = ((~g1919))|((~II6522));
assign g6148 = ((~II10807));
assign II13478 = ((~g7126));
assign II14780 = ((~g8284));
assign II8471 = ((~g2525))|((~II8470));
assign II9460 = ((~g3941));
assign g8460 = (g757&g8199);
assign g9318 = ((~g9304));
assign II11494 = ((~g6037));
assign g2367 = ((~II6202))|((~II6203));
assign g4393 = (g327&g3131);
assign g2944 = ((~g2363));
assign g4433 = (g278&g3097);
assign g3847 = ((~II7344));
assign g8325 = (g184&g8156);
assign II15714 = ((~g9077));
assign g2312 = ((~II6093));
assign g7983 = ((~II14294));
assign g1783 = ((~II5633));
assign g6033 = ((~g5384));
assign II9633 = ((~g4800));
assign II11157 = ((~g5482))|((~II11156));
assign g2262 = (g1384)|(g1385)|(g1386)|(g1387);
assign II10582 = ((~g5437));
assign II11110 = ((~g2734))|((~II11108));
assign II15510 = ((~g8969));
assign g5872 = ((~II10561));
assign g5417 = ((~g5006));
assign g9037 = (g8965&g5345);
assign g6366 = ((~II11425));
assign g4132 = (g2637&g2633);
assign g4643 = ((~II8844));
assign g5969 = (g5564&g2424);
assign g6810 = ((~II12301));
assign g7625 = (g7367&g4182);
assign II11163 = ((~g5469))|((~g3029));
assign II12145 = ((~g5971));
assign II8712 = ((~g4007));
assign II11461 = ((~g6094));
assign g5518 = (g4744)|(g4118);
assign g6567 = (g6265&g2424);
assign II11683 = ((~g5988));
assign II11550 = ((~g5984))|((~II11549));
assign II15043 = (g8363)|(g8342)|(g8407)|(g8386);
assign g3613 = ((~II7086))|((~II7087));
assign g4110 = ((~II7938))|((~II7939));
assign g7779 = ((~II14208));
assign g2105 = ((~g1444));
assign g6110 = ((~g5335));
assign g5622 = ((~g4938));
assign II15651 = ((~g9056));
assign II11929 = ((~g6190));
assign II11476 = ((~g6194));
assign g6993 = ((~II12731));
assign II8357 = ((~g1182));
assign g6352 = ((~II11383));
assign II10930 = ((~g5600));
assign II7931 = ((~g2780));
assign g3556 = ((~II7036));
assign II11945 = ((~g5874));
assign g2689 = ((~g1670));
assign g6076 = ((~g5287));
assign II7706 = ((~g2584));
assign II5945 = ((~g333));
assign g2633 = ((~g1577));
assign g4959 = (g376&g3898);
assign g1814 = ((~g630));
assign II12712 = ((~g6543));
assign II7599 = ((~g2734));
assign g8996 = (g8936)|(g8838);
assign g4341 = ((~II8308));
assign g3390 = ((~II6949));
assign II12763 = ((~g6686));
assign g8644 = ((~g4146)&(~g8128));
assign II7290 = ((~g2936));
assign g8303 = (g284&g7838);
assign II8412 = (g3430&g3398&g3359&g3341);
assign g1758 = ((~g1084));
assign g7253 = ((~g7049));
assign g7221 = ((~II13157));
assign II11359 = ((~g5810));
assign II7832 = ((~g2768));
assign g8943 = (g4560&g8781);
assign II11341 = ((~g5809));
assign g3014 = ((~II6767));
assign g7553 = (g7367&g4135);
assign II16180 = ((~g9387));
assign II14009 = ((~g7436));
assign II6956 = ((~g1907));
assign g8898 = ((~II15308));
assign g6506 = ((~II11680));
assign g5768 = ((~II10377));
assign g7554 = (g7367&g4139);
assign II9047 = (g4155)|(g4147)|(g4139);
assign g7175 = (g6893&g4841);
assign g7712 = ((~II14015));
assign g6562 = ((~II11736));
assign g9134 = ((~II15776));
assign g7834 = (g7724)|(g6762);
assign II8244 = ((~g2011))|((~II8243));
assign II13397 = ((~g1057))|((~II13395));
assign g7743 = ((~II14100));
assign g5684 = ((~II10183));
assign II10933 = ((~g5668));
assign II11696 = ((~g5971));
assign II11759 = ((~g6118))|((~II11757));
assign g6699 = (g6154)|(g5579);
assign g8931 = (g3867&g8761);
assign II13247 = ((~g6906));
assign g5067 = (g454&g3980);
assign g4158 = (II8033&II8034);
assign II15543 = ((~g9006));
assign II10770 = ((~g5441));
assign g3555 = ((~g2359)&(~g1398));
assign II7079 = ((~g2532));
assign II9999 = ((~g4839))|((~g1929));
assign g7313 = ((~II13369));
assign II12779 = ((~g6740));
assign II5520 = ((~g1087))|((~II5519));
assign II15010 = ((~g8584));
assign II14064 = ((~g7556));
assign II9258 = ((~g4249));
assign II10062 = ((~g2226))|((~II10060));
assign II14133 = ((~g7574));
assign g4310 = ((~g3666))|((~g2460));
assign II12918 = ((~g7013));
assign g7284 = ((~II13284));
assign II10708 = ((~g5545));
assign g4740 = (g2242&g4275);
assign II13583 = ((~g7252));
assign g8855 = ((~g7658)&(~g8613)&(~g7634));
assign g8067 = ((~II14342));
assign g5785 = ((~II10400));
assign II15285 = (g8709)|(g8713)|(g8803);
assign II8431 = (g3430&g3398&g3359&g3341);
assign g4080 = ((~II7867));
assign II10914 = ((~g5448));
assign g1704 = ((~II5548));
assign g2271 = ((~II6018));
assign g9272 = (g4748&g9248);
assign g6215 = ((~II10981))|((~II10982));
assign II13271 = ((~g7067));
assign g6181 = ((~II10907))|((~II10908));
assign g7304 = ((~II13344));
assign II10366 = ((~g5715));
assign II10151 = ((~g5007));
assign g4308 = ((~II8277));
assign II10494 = ((~g5232));
assign g1643 = ((~g1211));
assign II9837 = ((~g4781));
assign g2313 = ((~II6096));
assign g5638 = ((~g4748));
assign g3750 = ((~g2177));
assign II6752 = ((~g1494))|((~II6750));
assign II14674 = ((~g7788));
assign g7186 = (g6600&g7044);
assign g4434 = (g356&g3131);
assign g2664 = ((~II6463));
assign g6925 = (g6402)|(g6407);
assign g2901 = ((~g2284));
assign II11815 = ((~g6169));
assign g6446 = ((~II11591));
assign g3926 = ((~II7581));
assign II8955 = ((~g4246))|((~g1110));
assign g8443 = ((~g8015));
assign g4445 = (II8455&II8456);
assign g4334 = (g225&g3097);
assign g5223 = (g5069)|(g4398);
assign g2207 = ((~II5920));
assign g5806 = ((~II10451));
assign g9328 = (g9324&g6465);
assign g9107 = ((~II15711));
assign g5604 = ((~g4969));
assign g8332 = (g417&g7920);
assign II8736 = ((~g4008));
assign g8875 = ((~II15211));
assign g6160 = (g1504&g5718);
assign g6075 = ((~g5345));
assign g6914 = (g6483&g5246);
assign II7323 = ((~g2905));
assign g2867 = ((~g2222));
assign II6795 = ((~g1683));
assign II6856 = ((~g449));
assign g5621 = ((~g4748));
assign II10280 = ((~g5488));
assign g3577 = ((~g2372));
assign II5565 = ((~g1296));
assign g2294 = ((~II6065))|((~II6066));
assign g8798 = ((~g6984))|((~g8644));
assign II7728 = ((~g3675));
assign g6730 = ((~II12098));
assign g3081 = (g1682&g1616);
assign g1934 = ((~g154));
assign II15243 = (II15239)|(II15240)|(II15241)|(II15242);
assign g6307 = ((~II11248));
assign g8796 = (g8150)|(g8078)|(g8070)|(g8360);
assign II13646 = ((~g7245));
assign g4579 = ((~g2918));
assign g3497 = ((~g2185));
assign II14042 = ((~g7470));
assign g6253 = ((~g5403));
assign g3659 = ((~g2293));
assign g3904 = ((~g3160));
assign g3523 = ((~g2407));
assign II11299 = ((~g5786));
assign II11142 = ((~g5493))|((~g3062));
assign II6923 = ((~g1728))|((~g33));
assign g7653 = (g7480&g5754);
assign II11851 = ((~g6277));
assign g1888 = ((~g781));
assign g8304 = (g4523&g7905);
assign II14264 = ((~g7698));
assign II15616 = ((~g8997));
assign g7119 = ((~II12945));
assign II9692 = ((~g5096))|((~II9691));
assign II15110 = (g7855)|(g7838)|(g7905)|(g7870);
assign g4108 = (g782&g3655);
assign gbuf33 = (g1004);
assign II14378 = ((~g7691));
assign II14076 = ((~g7577));
assign g7547 = ((~II13825));
assign II10684 = ((~g5258));
assign g5704 = (g4936)|(g4334);
assign g3836 = ((~II7311));
assign g5108 = (g539&g4017);
assign g7632 = (g7445&g3548);
assign g1678 = ((~II5506))|((~II5507));
assign II12331 = ((~g6704));
assign II8483 = ((~g3641));
assign g4915 = ((~g4094));
assign II7610 = ((~g2471))|((~II7609));
assign g8658 = ((~g8199)&(~II14766)&(~II14767));
assign g7176 = ((~II13084));
assign g7511 = ((~II13713));
assign II6925 = ((~g33))|((~II6923));
assign II11227 = ((~g6130));
assign g1782 = ((~g624));
assign g5467 = ((~g4891));
assign g3970 = ((~g2845));
assign g2931 = ((~II6669));
assign II13698 = ((~g7348));
assign g2889 = (g1612&g1077);
assign g3561 = ((~II7041));
assign g1825 = ((~II5709));
assign II11576 = ((~g1122))|((~II11574));
assign g6910 = ((~g1011)&(~g1837)&(~g6559)&(~g1008));
assign g9114 = ((~II15732));
assign g6437 = (g859&g6050);
assign g8778 = ((~II14974));
assign g3771 = ((~g1853));
assign g2827 = (g1889&g1690);
assign II6054 = ((~g465));
assign II11556 = ((~g6065));
assign II8862 = ((~g3981));
assign II6834 = ((~g287));
assign g6809 = ((~II12298));
assign g6821 = ((~II12334));
assign g4679 = ((~II8939))|((~II8940));
assign g4058 = (g3656&g2407);
assign g6716 = (g6162)|(g5588);
assign g8564 = ((~g7951));
assign II10196 = ((~g4724))|((~g1958));
assign g3881 = ((~g2969));
assign II8811 = ((~g4022));
assign II6474 = ((~g1941));
assign g8524 = ((~g7855));
assign gbuf17 = (g1201);
assign g8648 = (g588&g8094);
assign II8006 = (g2074&g3287&g2020&g3238);
assign g8820 = (g261&g8524);
assign II15732 = ((~g9076));
assign g8784 = ((~g8545));
assign II12475 = ((~g6596));
assign g1562 = ((~g636));
assign II11874 = ((~g2543))|((~II11873));
assign g3994 = ((~g3192));
assign II13533 = ((~g7220));
assign g4537 = ((~g2878));
assign II7947 = ((~g3485));
assign g724 = ((~II5401));
assign g7425 = ((~II13550));
assign II8856 = ((~g3955));
assign II8781 = ((~g3932));
assign g1943 = ((~g1025));
assign g3784 = ((~g1768));
assign g7082 = ((~II12853))|((~II12854));
assign II13302 = ((~g7164));
assign II12921 = ((~g6993));
assign g5653 = ((~g4748));
assign II5371 = ((~g633));
assign II11413 = ((~g5871));
assign g6742 = ((~II12120));
assign g6876 = ((~II12499));
assign g8803 = ((~g8443)&(~g8421)&(~II15021));
assign g4453 = (g495&g3192);
assign g5287 = (g786&g4724);
assign g5345 = (g4736)|(g4734);
assign g4364 = (g2952)|(g1725);
assign g5364 = ((~g5124));
assign g8275 = (g4581&g7993);
assign g4427 = (II8431&II8432);
assign II12298 = ((~g6697));
assign II15084 = (g7951)|(g7920)|(g7983)|(g8181);
assign II11290 = ((~g5818));
assign g1804 = ((~II5664));
assign g6898 = ((~II12567));
assign g6441 = ((~II11586));
assign g9133 = ((~II15773));
assign g2972 = (g2397&g2407);
assign II9520 = ((~g3995));
assign g6481 = ((~II11641));
assign II9446 = ((~g3926));
assign II12725 = ((~g6565));
assign g5585 = (g4741&g4841);
assign g6457 = (g6196)|(g6209)|(g4937);
assign II12364 = ((~g6714));
assign g1576 = ((~g691));
assign g6703 = ((~II12041));
assign g5662 = ((~g5027));
assign g3965 = ((~II7676));
assign g2790 = ((~g1793));
assign II15645 = ((~g9043));
assign g6599 = ((~II11809));
assign II12853 = ((~g6701))|((~II12852));
assign g4802 = ((~II9129));
assign g4258 = ((~II8193));
assign II9964 = ((~g1938))|((~II9963));
assign II9826 = ((~g4729))|((~g1509));
assign II14467 = (g7993)|(g7966)|(g7793)|(g7811);
assign II10268 = ((~g5471));
assign II10545 = ((~g5259));
assign g8712 = (g2804&g8386);
assign II14753 = (g7993)|(g7966)|(g7793)|(g7811);
assign II15199 = ((~g8792));
assign II10298 = ((~g5461))|((~g2562));
assign II5842 = ((~g68));
assign g3656 = ((~II7139))|((~II7140));
assign II10259 = ((~g5362));
assign II6242 = ((~g1554));
assign g3732 = ((~g2533));
assign II7569 = ((~g3780))|((~II7567));
assign g7054 = ((~g6511));
assign g3944 = ((~II7635));
assign g8758 = (g8655)|(II14932)|(II14933);
assign g1638 = ((~g1092));
assign II9579 = ((~g4713));
assign g2267 = ((~II6006));
assign g8951 = (g8785&g6072);
assign II14097 = ((~g7595));
assign g7454 = ((~II13610));
assign g7951 = ((~II14288));
assign II7870 = ((~g2827));
assign g9332 = ((~g9322));
assign g5259 = (g5122)|(g4472);
assign g3093 = ((~g1686));
assign g3233 = ((~g1714)&(~g1459));
assign II9642 = ((~g4788));
assign g4264 = (g2490)|(g3315);
assign II13764 = ((~g7479));
assign II7864 = ((~g3812));
assign g6212 = ((~II10973));
assign g4489 = ((~g2826));
assign g9043 = ((~II15533));
assign g5618 = ((~g5015));
assign g2183 = ((~II5908));
assign g2539 = ((~II6363));
assign II13710 = ((~g7340));
assign g9112 = ((~II15726));
assign g7826 = (g4804)|(g7626);
assign g3505 = ((~g2263)&(~g1395));
assign II12597 = ((~g6582))|((~II12596));
assign g9288 = (g9272)|(g6235);
assign g4639 = ((~II8832));
assign g7233 = ((~g6940));
assign g2532 = ((~II6358));
assign g4779 = (g4176&g1760);
assign g3647 = ((~g2424));
assign g9306 = ((~II16036));
assign g8671 = ((~II14807));
assign g2921 = ((~g2312));
assign g4507 = (II8573&II8574);
assign II6299 = ((~g47));
assign II13879 = ((~g7332));
assign g2898 = ((~g2271));
assign g2214 = (g1376)|(g1377)|(g1378)|(g1379);
assign II12346 = ((~g6737));
assign g1917 = ((~II5795));
assign g1799 = ((~II5657));
assign II13084 = ((~g7071));
assign g2962 = ((~g2382));
assign g7518 = ((~II13734));
assign g8654 = (g570&g8094);
assign g6152 = ((~II10815));
assign g6885 = ((~II12526));
assign II7174 = ((~g2006))|((~II7172));
assign II14142 = ((~g7551));
assign g8613 = (g8082)|(g7616);
assign g5066 = (g395&g3978);
assign g4020 = ((~II7781));
assign g9201 = ((~g9183));
assign II8299 = (g3666&g3684&g3694&g3707);
assign g6405 = (g5956&g5494);
assign g5746 = ((~II10295));
assign II15507 = ((~g8968));
assign g2884 = ((~g2238));
assign g3679 = ((~II7180))|((~II7181));
assign II11233 = ((~g6147));
assign II11314 = ((~g5781));
assign g2402 = ((~g29));
assign II13810 = ((~g7312));
assign II8945 = ((~g4106));
assign II10277 = ((~g5472));
assign g5206 = ((~g4938));
assign II7574 = ((~g2999))|((~g1718));
assign g6708 = ((~g6250));
assign g6634 = ((~II11894));
assign II8089 = (g2162&g2149&g2137&g2106);
assign g5200 = (g5029)|(g4375);
assign II15933 = ((~g9210));
assign II9564 = ((~g4703));
assign II12214 = ((~g6507));
assign II12079 = ((~g5988))|((~II12078));
assign II10451 = ((~g5216));
assign g7142 = ((~II13012));
assign g9235 = ((~II15959));
assign II14683 = ((~g7825));
assign g5487 = ((~II9907));
assign g2810 = ((~g1922));
assign g9007 = (g8947)|(g8854);
assign g2221 = ((~II5936));
assign II11350 = ((~g5763));
assign g3237 = ((~g1444)&(~g1838)&(~g1454));
assign II12138 = ((~g5874));
assign II12445 = ((~g6568));
assign g9123 = (g8954)|(g9037);
assign g5084 = ((~g4477));
assign g5157 = ((~II9597));
assign g6415 = (g5988&g5367);
assign II7581 = ((~g3612));
assign II11793 = ((~g6188));
assign g2044 = ((~II5861));
assign II12948 = ((~g6919));
assign g1737 = ((~g597));
assign II14342 = ((~g7582));
assign II13565 = ((~g7181));
assign gbuf24 = (g1393);
assign g6083 = ((~II10702));
assign g1662 = ((~g1412));
assign g7507 = ((~II13701));
assign II11659 = ((~g5897));
assign g6346 = ((~II11365));
assign g8665 = ((~II14789));
assign g9039 = ((~II15527));
assign II13797 = ((~g7502));
assign II8480 = ((~g3640));
assign g7750 = ((~II14121));
assign g4616 = ((~II8763));
assign II8254 = ((~g2454))|((~II8253));
assign II7149 = ((~g799))|((~II7148));
assign g6651 = ((~II11933));
assign II12451 = ((~g6524));
assign g3835 = ((~II7308));
assign g4572 = ((~g2909));
assign g2241 = ((~II5984));
assign g2345 = ((~II6151));
assign II5670 = ((~g941));
assign g7102 = ((~II12894));
assign II8328 = ((~g2721))|((~II8326));
assign g5627 = ((~g4673));
assign g658 = ((~II5386));
assign g4784 = ((~II9095));
assign g4685 = ((~II8952));
assign II7749 = ((~g3692));
assign g7904 = ((~II14276));
assign II9502 = ((~g3972));
assign g3896 = ((~II7473));
assign II6428 = ((~g1818));
assign g8923 = (g4587&g8751);
assign g7488 = ((~g7225));
assign g7766 = ((~II14169));
assign g6286 = ((~II11178))|((~II11179));
assign g7048 = ((~II12810));
assign II13152 = ((~g6966));
assign II8582 = ((~g2498))|((~II8581));
assign II9196 = ((~g1652))|((~II9194));
assign II10334 = ((~g5462))|((~g2573));
assign g5030 = (g233&g3946);
assign II13103 = ((~g7055));
assign g5232 = (g5082)|(g4412);
assign II10899 = ((~g5520))|((~g2752));
assign II14276 = ((~g7720));
assign g6938 = ((~II12635));
assign g4072 = (g196)|(g2995);
assign g8860 = (g527&g8585);
assign g5192 = ((~g4841));
assign II8551 = (g3430&g3398&g3359&g2106);
assign g5261 = ((~g4748));
assign g6789 = ((~II12238));
assign II12289 = ((~g6702));
assign g8897 = (g8833)|(g8650);
assign g7755 = ((~II14136));
assign g8176 = (g7566)|(g1030)|(g6664)|(g6452);
assign g8738 = (g8619&g3338);
assign g6656 = ((~II11948));
assign g9279 = (g9255&g5665);
assign g8380 = (g681&g7887);
assign II8829 = ((~g4029));
assign g8836 = (g348&g8545);
assign g4282 = (g3549&g3568);
assign II10160 = ((~g5139));
assign g4823 = (g4238&g4230&g174);
assign g4194 = (II8089&II8090);
assign II11347 = ((~g5761));
assign II10506 = ((~g5236));
assign g4510 = ((~g2840));
assign g5840 = ((~II10535));
assign II8793 = ((~g3923));
assign g2485 = ((~g62));
assign g7724 = (g7337&g5938);
assign II11218 = ((~g6161));
assign II10406 = ((~g5203));
assign II5395 = ((~g698));
assign g7363 = (g7136)|(g6903);
assign II9618 = ((~g4742));
assign g7731 = ((~II14064));
assign II15773 = ((~g9126));
assign g4567 = ((~g2903));
assign II5353 = ((~g3833));
assign II11821 = ((~g6170));
assign g8582 = ((~g8094));
assign II11398 = ((~g5823));
assign II6103 = ((~g849))|((~II6102));
assign II15631 = ((~g9003));
assign II13656 = ((~g7228));
assign g3092 = ((~II6826));
assign II15598 = ((~g8991));
assign g7329 = ((~II13407));
assign g3002 = (g871&g1834);
assign g6224 = ((~II11011));
assign g2145 = ((~g1296));
assign g3466 = (g936&g2557);
assign g6980 = (g6745)|(g6028);
assign g8755 = ((~g8545));
assign g5127 = ((~II9525));
assign g4284 = (g3260&g3314);
assign II8835 = ((~g3954));
assign g1980 = ((~g1430)&(~g1431));
assign II14169 = ((~g7715));
assign g6766 = ((~II12167));
assign g6490 = ((~II11656));
assign g4923 = ((~g4112));
assign II5981 = ((~g459));
assign g7460 = ((~g7172));
assign II8932 = ((~g4096));
assign g5819 = ((~II10482));
assign g6752 = ((~II12131));
assign II13326 = ((~g7176));
assign g1745 = ((~g746));
assign g4881 = ((~g2460))|((~g4315));
assign g6462 = (g6215&g2424);
assign g9080 = (g9011&g5598);
assign II7216 = ((~g2091))|((~II7214));
assign g8059 = (g7682&g7032);
assign II10716 = ((~g5537));
assign II10463 = ((~g5220));
assign II11242 = ((~g6183));
assign g8605 = ((~II14680));
assign g9379 = ((~II16161));
assign g5441 = (g4870&g3497);
assign g7439 = ((~II13574));
assign II8802 = ((~g3963));
assign II12891 = ((~g6950));
assign g9073 = ((~II15613));
assign g8660 = (g1069&g8147);
assign g7467 = ((~g7236));
assign g1857 = ((~g889));
assign g3875 = ((~g2958));
assign g5158 = ((~II9600));
assign II9910 = ((~g4681));
assign g9212 = ((~II15912));
assign g7345 = ((~II13451));
assign II15481 = ((~g8913));
assign II8215 = ((~g3577));
assign II14049 = ((~g7493));
assign II13807 = ((~g7320));
assign II14302 = (g6664)|(g3492)|(g979);
assign g5078 = (g316&g3989);
assign II9222 = (g4041&g4044&g2584);
assign II8502 = ((~g2986))|((~g2038));
assign g6672 = ((~II11974));
assign II12397 = ((~g6764));
assign g3982 = ((~g3192));
assign II9979 = ((~g4880))|((~II9978));
assign II7009 = ((~g2295))|((~g2333));
assign g8661 = ((~II14777));
assign g1600 = ((~g976));
assign g1961 = ((~g1345));
assign g2495 = ((~g26));
assign g8719 = (g2821&g8443);
assign g1616 = ((~II5478));
assign g6967 = ((~II12696));
assign g6089 = ((~g5317));
assign g5397 = ((~g5076));
assign g9030 = ((~II15504));
assign g6777 = ((~II12202));
assign g8232 = ((~g8199)&(~II14479)&(~II14480));
assign II14810 = ((~g8481));
assign g5037 = ((~g4438));
assign g7208 = ((~II13140));
assign g3960 = ((~II7667));
assign g4744 = (g3525&g4296);
assign II10286 = ((~g5519));
assign g6797 = ((~II12262));
assign II11843 = ((~g6158))|((~II11841));
assign II10353 = ((~g5710));
assign II9547 = ((~g1952))|((~g4307));
assign II14175 = ((~g7718));
assign g8224 = ((~II14451));
assign II7335 = ((~g2910));
assign II14851 = ((~g8630));
assign g9377 = (g9371)|(g6757);
assign g4466 = (II8490&II8491);
assign II8607 = ((~g2764))|((~II8605));
assign g7708 = ((~II14005));
assign g6960 = ((~II12681));
assign II10842 = ((~g5701));
assign g4295 = (g2828)|(g2668);
assign II15265 = (II15261)|(II15262)|(II15263)|(II15264);
assign II14959 = (g8322)|(g8308)|(g8438)|(g8612);
assign g4738 = ((~II9050));
assign g5172 = ((~II9642));
assign g8611 = (g669&g7887);
assign g2562 = ((~g1652));
assign II9029 = (g4504)|(g4494)|(g4430);
assign g3706 = ((~g1556))|((~g2510));
assign II6791 = ((~g1967));
assign g6238 = ((~II11043));
assign II12737 = ((~g6460));
assign g3260 = ((~g1728)&(~g2490));
assign g8629 = ((~g6270)&(~g8009));
assign g2842 = ((~g2209));
assign g6790 = ((~II12241));
assign g2477 = ((~g25));
assign g9343 = (g9328&g1738);
assign g2374 = ((~II6220));
assign g9090 = ((~II15660));
assign II14028 = ((~g7501));
assign g7475 = ((~II13631));
assign g3359 = ((~II6946));
assign II11470 = ((~g6095));
assign II8511 = ((~g2517))|((~II8510));
assign II9892 = ((~g4879));
assign g7020 = (g3617)|(g6578);
assign II12586 = ((~g6643));
assign g7783 = (g4787)|(g7600);
assign g4737 = (g4135)|(g4529)|(g4514)|(II9047);
assign g7288 = ((~II13296));
assign g5831 = ((~II10516));
assign g8063 = ((~II14334));
assign II11967 = ((~g5971));
assign II14151 = ((~g7555));
assign II14127 = ((~g7594));
assign g9277 = (g9248&g5654);
assign II13779 = ((~g7406));
assign II14496 = (g7937)|(g7887)|(g8029)|(g8018);
assign g6713 = ((~II12065));
assign g2206 = (g1363)|(g1364)|(g1365)|(g1366);
assign g9302 = ((~g9281));
assign g7686 = ((~II13979));
assign g6807 = ((~II12292));
assign g8273 = (g185&g8156);
assign g5570 = (g1759&g4841);
assign g7509 = ((~II13707));
assign gbuf65 = (g530);
assign g4021 = ((~g3131));
assign II15811 = ((~g9151));
assign g3338 = ((~g1901));
assign g5672 = ((~g5056))|((~g5039))|((~g5023));
assign g6712 = ((~II12062));
assign g8912 = (g8796&g8239);
assign II5657 = ((~g921));
assign II6757 = ((~g186))|((~g1983));
assign g9056 = ((~II15562));
assign II10019 = ((~g2174))|((~II10017));
assign g9348 = (g9333&g6229);
assign g2185 = ((~II5914));
assign g6004 = ((~g5494));
assign g6686 = (g4068)|(g5970);
assign g9197 = ((~g9186));
assign II11710 = ((~g6098));
assign g5605 = ((~II10093))|((~II10094));
assign g8289 = (g348&g7870);
assign g3085 = ((~g1945));
assign g6471 = ((~II11627));
assign g8659 = ((~g8199)&(~II14771)&(~II14772));
assign II9271 = ((~g4263));
assign II13438 = ((~g7143));
assign II8157 = (g2686&g2689&g2692);
assign II15429 = ((~g8899));
assign II12379 = ((~g6768));
assign g8223 = ((~II14448));
assign II11392 = ((~g5800));
assign g6646 = ((~II11920));
assign II7461 = ((~g3815))|((~II7459));
assign II6045 = ((~g309));
assign II10436 = ((~g5213));
assign g2479 = ((~g32));
assign g4929 = ((~g4120));
assign II10359 = ((~g5552))|((~g1118));
assign g4397 = (g483&g3192);
assign g7470 = ((~g7253));
assign II13686 = ((~g1977))|((~II13685));
assign g7596 = (g7428&g7028);
assign II11434 = ((~g5789));
assign II11122 = ((~g5517))|((~g2712));
assign gbuf68 = (g890);
assign g5520 = ((~g4928));
assign g6888 = ((~II12535));
assign II12541 = ((~g6614));
assign g2920 = ((~II6652));
assign II13834 = ((~g7466));
assign II6770 = ((~g1590));
assign g9096 = ((~II15678));
assign g7360 = ((~II13496));
assign g3995 = ((~II7728));
assign g5071 = ((~g4438));
assign II9070 = ((~g4400))|((~II9069));
assign II13305 = ((~g7168));
assign II12352 = ((~g6752));
assign g9078 = ((~II15628));
assign g9219 = ((~II15933));
assign II8243 = ((~g2011))|((~g3506));
assign II14668 = ((~g7787));
assign g7614 = (g7367&g4176);
assign g2215 = ((~g1416));
assign g4018 = ((~II7775));
assign g8849 = (g513&g8585);
assign II14190 = ((~g7531));
assign g3047 = ((~g1736));
assign g4743 = (g3518&g4286);
assign g1987 = ((~II5842));
assign g2256 = ((~g1324));
assign g7277 = ((~II13267));
assign g3676 = ((~g2380));
assign g8610 = (g665&g7887);
assign g7751 = ((~II14124));
assign g6695 = ((~II12016))|((~II12017));
assign II15604 = ((~g8993));
assign gbuf12 = (g1195);
assign g2289 = ((~II6051));
assign g7037 = ((~g6525));
assign g7560 = ((~II13854));
assign g4633 = ((~II8814));
assign g6825 = ((~II12346));
assign g7772 = ((~II14187));
assign g7226 = ((~g6937));
assign II9819 = ((~g4691));
assign II13640 = ((~g7069))|((~II13638));
assign g9076 = ((~II15622));
assign g9089 = ((~II15657));
assign gbuf26 = (g1399);
assign II5535 = ((~g48));
assign II11838 = ((~g6281));
assign g6461 = ((~II11607));
assign II7453 = ((~g3226))|((~II7452));
assign g9154 = (g9142)|(g9021);
assign II10418 = ((~g5453));
assign g6788 = ((~II12235));
assign II5831 = ((~g1194));
assign g2237 = ((~II5972));
assign g1564 = ((~g642));
assign II6021 = ((~g495));
assign g7887 = ((~II14273));
assign II11848 = ((~g6159));
assign g5033 = (g393&g3953);
assign II7173 = ((~g1739))|((~II7172));
assign II15641 = ((~g9017));
assign II12190 = ((~g5918));
assign g8421 = ((~g8017));
assign g3999 = ((~II7738));
assign g4316 = ((~II8291));
assign II7480 = ((~g3808))|((~II7478));
assign II5936 = ((~g222));
assign II9129 = ((~g4475));
assign g8634 = (g6047)|(g8060);
assign II11704 = ((~g6076));
assign II5428 = ((~g49));
assign g5593 = (g4110&g4969);
assign II14416 = ((~g7727));
assign g8872 = ((~II15202));
assign II6431 = ((~g1825));
assign II14257 = ((~g7716));
assign g4904 = ((~g4085));
assign g4304 = (g2784&g3779);
assign II7262 = ((~g2514));
assign g6305 = ((~II11242));
assign g3097 = (g1746)|(g287);
assign g8612 = (g673&g7887);
assign II16072 = ((~g9303));
assign g4051 = ((~g3093));
assign g7698 = (g7367&g4483);
assign g5173 = ((~II9645));
assign g3980 = ((~g3192));
assign g4104 = ((~II7925));
assign g7543 = ((~II13813));
assign g5736 = ((~II10265));
assign g9227 = ((~II15947));
assign II15912 = ((~g9193));
assign g8290 = (g588&g8181);
assign II12505 = ((~g6612));
assign g6869 = ((~II12478));
assign g8889 = (II15283)|(II15284)|(II15285);
assign g7728 = ((~II14055));
assign II11248 = ((~g6149));
assign g6707 = (g6160)|(g5585);
assign g4793 = (g3887&g4202);
assign g8869 = ((~II15193));
assign g2161 = ((~g1454));
assign g8636 = ((~II14718));
assign II9366 = ((~g4350));
assign II8605 = ((~g2487))|((~g2764));
assign g5239 = ((~II9746))|((~II9747));
assign II13876 = ((~g7347));
assign g4656 = ((~II8883));
assign g4202 = ((~g2810));
assign g6516 = ((~g5897))|((~g5278));
assign g3643 = ((~g2453));
assign g7215 = (g6111&g6984);
assign II13454 = ((~g7147));
assign g2556 = ((~g1190));
assign g6469 = ((~g5918))|((~g5278));
assign g5708 = (g2889)|(g4699);
assign g3895 = ((~II7467))|((~II7468));
assign II15898 = ((~g9202))|((~II15897));
assign g4147 = (II8014&II8015);
assign g6639 = ((~g6198));
assign g8009 = (g3591)|(g7406)|(g7566)|(II14302);
assign g7721 = ((~g7344));
assign g8235 = ((~II14492));
assign II8727 = ((~g3944));
assign g4464 = ((~II8486));
assign g4907 = ((~g4087));
assign g2331 = ((~g933));
assign g8655 = ((~g8199)&(~II14753)&(~II14754));
assign g1708 = ((~II5552));
assign g6477 = ((~g5269))|((~g5918));
assign g4229 = ((~II8140));
assign II13234 = ((~g6898));
assign II10466 = ((~g5221));
assign II11014 = ((~g5621));
assign g6775 = ((~II12196));
assign g5224 = ((~g5114));
assign g3008 = ((~g1816));
assign g6170 = ((~II10874))|((~II10875));
assign g8859 = ((~g8493)&(~g8239)&(~II15165));
assign II14279 = ((~g7700));
assign II13063 = ((~g6973));
assign g6116 = (g5546)|(g4681);
assign g9236 = ((~II15962));
assign II6878 = ((~g1910))|((~II6876));
assign II11008 = ((~g5693));
assign g6153 = ((~II10819))|((~II10820));
assign II6974 = ((~g2528));
assign g8377 = (g507&g7966);
assign g6424 = ((~II11550))|((~II11551));
assign g6221 = ((~II11004));
assign II11506 = ((~g6189));
assign g6680 = ((~g5403))|((~g6252));
assign g6386 = ((~II11485));
assign II7867 = ((~g2818));
assign g5560 = (g3390&g5036);
assign II6419 = ((~g1799));
assign g3049 = (g2274&g1844);
assign II5633 = ((~g891));
assign g5644 = ((~g4748));
assign g8724 = (g3822&g8464);
assign g5264 = (g5125)|(g4490);
assign II12031 = ((~g5918))|((~g5897));
assign II12164 = ((~g5847));
assign II12051 = ((~g5956))|((~g5939));
assign g9352 = (g9343)|(g4526);
assign II8296 = (g3666&g3684&g3707);
assign II6751 = ((~g1733))|((~II6750));
assign g8774 = ((~II14964));
assign g5080 = (g396&g3991);
assign II5389 = ((~g690));
assign g5723 = ((~g4938));
assign II8538 = ((~g2798))|((~II8536));
assign g5031 = (g292&g3948);
assign g6242 = ((~II11047));
assign g5122 = (g436&g4030);
assign g7792 = ((~II14231));
assign g8737 = (g2992&g8493);
assign g5599 = (g4745&g4969);
assign g9300 = ((~II16026));
assign II10442 = ((~g5215));
assign g1671 = ((~g1494));
assign g4263 = ((~g3260))|((~g1435));
assign II5923 = ((~g252));
assign II8340 = ((~g1698))|((~II8338));
assign II5960 = ((~g187));
assign II9669 = ((~g4909));
assign II7893 = ((~g1499))|((~II7891));
assign II12552 = ((~g1462))|((~II12550));
assign g8966 = (g8741)|(g8745)|(g8912)|(g8850);
assign g1942 = ((~g828));
assign g6324 = ((~II11299));
assign g6068 = ((~II10687));
assign II11266 = ((~g5794));
assign g6449 = ((~II11596));
assign g4426 = ((~II8428));
assign g4912 = ((~II9277))|((~II9278));
assign g2131 = ((~g1300));
assign g5762 = ((~II10360))|((~II10361));
assign II13770 = ((~g7491));
assign II9603 = ((~g4719));
assign g3882 = ((~g2970));
assign g8156 = ((~II14394));
assign II9955 = ((~g4831))|((~II9953));
assign g6440 = (g6268)|(g5700);
assign g8808 = ((~II15062));
assign II8583 = ((~g2777))|((~II8581));
assign g3503 = ((~g2407));
assign g7540 = ((~II13801))|((~II13802));
assign g5873 = ((~g5367));
assign II13250 = ((~g7036));
assign g5678 = ((~II10169));
assign g7259 = ((~g7060));
assign g2233 = ((~II5960));
assign g6933 = (g6419)|(g6428);
assign g4081 = ((~II7870));
assign g7270 = ((~II13250));
assign g6973 = ((~II12708));
assign g3907 = ((~II7511))|((~II7512));
assign g9132 = ((~II15770));
assign II11942 = ((~g6015));
assign g8824 = (g264&g8524);
assign g7341 = ((~II13441));
assign II14311 = ((~g7566));
assign gbuf47 = (g1154);
assign II9235 = ((~g2180))|((~II9233));
assign g3956 = ((~g2845));
assign II15252 = (g8320)|(g8307)|(g8317)|(g8692);
assign g4254 = (g3583&g3568&g3549);
assign g4538 = ((~g2880));
assign g1570 = ((~g665));
assign II11809 = ((~g6285));
assign II6248 = ((~g411));
assign g4809 = ((~II9148));
assign II10627 = ((~g1514))|((~II10625));
assign II13527 = ((~g7217));
assign g2793 = ((~II6532));
assign g5094 = (g535&g4004);
assign g4788 = ((~II9103));
assign II12529 = ((~g6628));
assign II10952 = ((~g5565))|((~g2340));
assign g6187 = ((~g5633))|((~g3735))|((~g3716));
assign g7184 = (g6138&g7043);
assign II15196 = ((~g8778));
assign g8583 = ((~II14668));
assign II6233 = ((~g834))|((~II6232));
assign g7718 = ((~II14031));
assign II7847 = ((~g3798));
assign g5241 = (g5104)|(g4433);
assign II15635 = ((~g8976));
assign g5661 = ((~II10143))|((~II10144));
assign g4514 = (II8588&II8589);
assign g7151 = ((~II13035));
assign g2377 = ((~II6229));
assign g3962 = ((~g3131));
assign II7995 = (g2074&g3287&g2020&g3238);
assign g8607 = (g8154&g5616);
assign g5825 = ((~II10500));
assign g9192 = ((~II15863))|((~II15864));
assign g1913 = (g1528&g1532);
assign g1749 = ((~g371));
assign g5432 = (g1537&g4921);
assign II11172 = ((~g3038))|((~II11170));
assign g6574 = (g1045&g5984);
assign g5801 = ((~II10442));
assign II10061 = ((~g4910))|((~II10060));
assign II5507 = ((~g1528))|((~II5505));
assign II9195 = ((~g4252))|((~II9194));
assign II12731 = ((~g6579));
assign g1837 = ((~g1007));
assign g4299 = (g3233&g3358);
assign g8952 = (g8788&g6075);
assign II14082 = ((~g7539));
assign II12722 = ((~g6611));
assign II11875 = ((~g6187))|((~II11873));
assign g3665 = ((~II7157))|((~II7158));
assign g1788 = ((~g984));
assign g5139 = ((~II9543));
assign II8288 = (g3666&g3684&g3694);
assign II11936 = ((~g5918));
assign II9827 = ((~g4729))|((~II9826));
assign II14460 = ((~g7789));
assign II12334 = ((~g6713));
assign g6040 = (g1462&g5578);
assign II14136 = ((~g7633));
assign II5732 = ((~g859));
assign g4592 = ((~g2938));
assign g6311 = ((~II11260));
assign II5407 = ((~g4653));
assign g4517 = (II8593&II8594);
assign g3812 = ((~g1750));
assign g7303 = ((~II13341));
assign g9115 = ((~II15735));
assign g9025 = (g8889&g5317);
assign II13383 = ((~g7275));
assign II15577 = ((~g8984));
assign g2973 = ((~g1854));
assign g8323 = (g524&g7966);
assign g4532 = (II8617&II8618);
assign g3838 = ((~II7317));
assign II7765 = ((~g2595));
assign g7833 = (g6461&g7601);
assign g4250 = ((~II8177));
assign II10305 = ((~g5470))|((~g3019));
assign g4666 = ((~II8913));
assign g8626 = (g752&g8199);
assign g4877 = (g3746&g3723&g4288&g3764);
assign g2644 = ((~II6416));
assign g6802 = ((~II12277));
assign II6590 = ((~g2467));
assign g4521 = ((~g2866));
assign II11796 = ((~g6287));
assign II15241 = (g8269)|(g8314)|(g8309)|(g8695);
assign g8173 = ((~II14400));
assign g4808 = ((~II9145));
assign II12499 = ((~g6597));
assign II7326 = ((~g2940));
assign g7419 = (g7230&g3530);
assign g6408 = (g669&g6019);
assign g1667 = ((~g1481));
assign g8336 = (g420&g7920);
assign II12748 = ((~g6585));
assign g8331 = (g339&g7870);
assign g6038 = ((~II10649));
assign g5044 = (g234&g3959);
assign II10125 = ((~g5127));
assign g9106 = ((~II15708));
assign II7885 = ((~g2837));
assign II12158 = ((~g5956));
assign g6288 = ((~II11191));
assign II5356 = ((~g3837));
assign II14623 = ((~g7833));
assign II6081 = ((~g118));
assign g5220 = (g5066)|(g4395);
assign g8721 = (g2703&g8464);
assign II6192 = ((~g327));
assign g3545 = ((~g2344));
assign II8202 = ((~g3560));
assign II8491 = (g3316&g2057&g3264&g3238);
assign g5511 = (g4743)|(g4109);
assign II9202 = (g2605&g4044&g2584);
assign g4085 = ((~II7878));
assign II11185 = ((~g5474))|((~II11184));
assign g6438 = (g4829&g6051);
assign g5017 = (g211&g3928);
assign g7014 = ((~II12760));
assign II11818 = ((~g6276));
assign g6664 = ((~g5836)&(~g1901)&(~g1788));
assign II12101 = ((~g5971));
assign g7126 = ((~II12968));
assign II14199 = ((~g7704));
assign g3654 = ((~g2521));
assign II8363 = (g2655)|(g1163)|(g1160);
assign g699 = ((~II5395));
assign II7558 = ((~g2734));
assign II13716 = ((~g7331));
assign g1801 = ((~g618));
assign II8134 = ((~g1646))|((~II8132));
assign g7742 = ((~II14097));
assign g655 = ((~II5383));
assign g2546 = ((~II6368));
assign II7118 = ((~g2484));
assign g8793 = (g8637&g5622);
assign II13258 = ((~g6907));
assign II12669 = ((~g6477));
assign g3753 = ((~g2540));
assign g6210 = ((~II10969));
assign g6624 = ((~II11864));
assign II6189 = ((~g249));
assign II9393 = ((~g4266));
assign g7324 = ((~g7189)&(~g6994));
assign g2511 = ((~g1328));
assign g6315 = ((~II11272));
assign g5639 = ((~g4748));
assign g3949 = ((~II7644));
assign g8438 = (g649&g7793);
assign g3940 = ((~II7623));
assign g5014 = ((~II9344));
assign g4719 = ((~II9021));
assign g5793 = ((~II10418));
assign g8236 = ((~g8199)&(~II14495)&(~II14496));
assign II12223 = ((~g6655));
assign g2878 = ((~g2233));
assign II5598 = ((~g1481))|((~g1489));
assign g7420 = ((~II13537));
assign II12582 = ((~g6745));
assign g6342 = ((~II11353));
assign g5550 = ((~g1879))|((~g4830));
assign g5090 = (g317&g4000);
assign II7386 = ((~g3013));
assign II15678 = ((~g9060));
assign g5482 = ((~g4915));
assign II15208 = ((~g8810));
assign g7438 = (g7184)|(g6978);
assign g6784 = ((~II12223));
assign g3230 = ((~II6887));
assign g8442 = ((~II14623));
assign II12951 = ((~g7003))|((~g1467));
assign g5107 = (g478&g4016);
assign g5569 = ((~II10028));
assign II11884 = ((~g6091));
assign g7090 = ((~g6525));
assign II7811 = ((~g3019));
assign g7334 = ((~II13422));
assign g2932 = ((~g2329));
assign g3942 = ((~II7629));
assign II7939 = ((~g1138))|((~II7937));
assign II15681 = ((~g9063));
assign II16006 = ((~g9261));
assign g2909 = ((~g2291));
assign g3967 = ((~II7680));
assign g4038 = (g825&g2949);
assign II6446 = ((~g1812));
assign II10532 = ((~g5253));
assign g6019 = ((~g5367));
assign II13277 = ((~g7078));
assign g2490 = ((~II6326));
assign g8359 = (g642&g7793);
assign g1725 = (g1409&g1416);
assign g7098 = ((~g6525));
assign g2825 = ((~II6553));
assign II10295 = ((~g5523));
assign II15918 = ((~g9211));
assign II14234 = ((~g7614));
assign g3520 = ((~g1616));
assign II6814 = ((~g210))|((~II6813));
assign g1681 = ((~g929));
assign II7731 = ((~g3029));
assign g5428 = (g775&g4707);
assign g6911 = ((~II12597))|((~II12598));
assign g6165 = ((~II10855))|((~II10856));
assign g7583 = ((~II13894));
assign II12520 = ((~g6622));
assign II9081 = ((~g4357));
assign II5410 = ((~g8866));
assign g8852 = (g362&g8545);
assign g6582 = (g1122&g5894);
assign g7210 = ((~II13144));
assign g3978 = ((~g3160));
assign g6265 = ((~II11079))|((~II11080));
assign g4133 = (g2631&g2623);
assign g6432 = ((~II11569));
assign II13598 = ((~g2551))|((~g7244));
assign g5715 = (g4961)|(g4355);
assign II6171 = ((~g843))|((~II6170));
assign g4739 = ((~II9053));
assign g7083 = (g5448)|(g6267)|(g6710);
assign g3918 = ((~II7551));
assign g8174 = ((~II14403));
assign g6904 = ((~g6426));
assign g4878 = (g2573&g2562&II9222);
assign II12108 = ((~g5939));
assign g8969 = ((~II15411));
assign g3822 = ((~g1815));
assign g5917 = ((~g5412));
assign g4113 = ((~II7950));
assign II7204 = ((~g2520));
assign g8147 = (g1065&g7683);
assign g9127 = ((~II15759));
assign II12983 = ((~g6930));
assign II5984 = ((~g540));
assign g2634 = ((~g1578));
assign g5466 = ((~g4890));
assign g1817 = ((~II5689));
assign g6964 = (g6447)|(g6448);
assign g9031 = ((~II15507));
assign II9660 = ((~g4806));
assign g5654 = ((~g4748));
assign II8428 = ((~g3611));
assign II15017 = (g8131)|(g8111)|(g8042)|(g8156);
assign g6359 = ((~II11404));
assign II11861 = ((~g5747));
assign II7919 = ((~g3761));
assign II8432 = (g3316&g3287&g2020&g3238);
assign g3898 = ((~g3160));
assign g5722 = (g5001)|(g4361);
assign g8439 = (g699&g7811);
assign g5116 = (g355&g4021);
assign II10579 = ((~g5433));
assign g7336 = ((~II13428));
assign g2623 = ((~g1585));
assign g4588 = ((~g2929));
assign II7158 = ((~g929))|((~II7156));
assign II14531 = ((~g8178));
assign II8308 = ((~g3674));
assign g5132 = (II9534&II9535);
assign g7348 = ((~II13460));
assign II6451 = ((~g1895));
assign g8785 = (g8623)|(g8656)|(II14985);
assign II6102 = ((~g849))|((~g921));
assign II14970 = (g8457)|(g8383)|(g8626)|(g8233);
assign g9188 = ((~II15842));
assign g1670 = ((~g1489));
assign II13396 = ((~g7212))|((~II13395));
assign II13215 = ((~g7082))|((~II13213));
assign II6805 = ((~g1603));
assign II11627 = ((~g5874));
assign g3787 = ((~g1842));
assign II13416 = ((~g7165));
assign g2890 = ((~g2264));
assign II8024 = ((~g3076));
assign II6134 = ((~g846))|((~II6133));
assign II6130 = ((~g560));
assign g7239 = ((~g6945));
assign II6434 = ((~g1830));
assign II14485 = (g7937)|(g7887)|(g8029)|(g8018);
assign g8089 = (g840&g7658);
assign II15414 = ((~g8900));
assign g4570 = ((~g2907));
assign g9044 = ((~II15536));
assign II12538 = ((~g6606));
assign g1579 = ((~g703));
assign g4050 = ((~g3080));
assign g3981 = ((~II7706));
assign g6972 = (g5661&g6498);
assign II5605 = ((~g58));
assign g3790 = ((~g985)&(~g990)&(~g2295));
assign g6598 = ((~II11806));
assign g6875 = ((~II12496));
assign II9076 = ((~g4353));
assign g8514 = ((~g8040));
assign g3855 = ((~II7368));
assign II14121 = ((~g7587));
assign g8775 = ((~g8564));
assign g8265 = (g134&g8111);
assign II7085 = ((~g1753))|((~g1918));
assign g8604 = ((~II14677));
assign g6625 = ((~II11867));
assign II9181 = ((~g4231))|((~g2007));
assign g8713 = (g2777&g8421);
assign II16055 = ((~g9291));
assign II14766 = (g7993)|(g7966)|(g7793)|(g7811);
assign g7574 = ((~II13869));
assign g4303 = ((~II8268));
assign g3955 = ((~II7658));
assign II6723 = ((~g2052));
assign g8760 = ((~g8545));
assign g1588 = ((~g741));
assign II10060 = ((~g4910))|((~g2226));
assign II10528 = ((~g5245));
assign II12965 = ((~g6924));
assign g6341 = ((~II11350));
assign g5759 = ((~II10350));
assign g5740 = ((~II10277));
assign II15849 = ((~g9162))|((~II15848));
assign g8999 = (g8939)|(g8843);
assign g2843 = ((~II6571));
assign g6954 = (g5518&g6601);
assign g6840 = ((~II12391));
assign II15193 = ((~g8774));
assign g5299 = ((~II9804));
assign II12244 = ((~g6642));
assign g9140 = ((~II15784));
assign II13017 = ((~g6941))|((~II13016));
assign g6862 = ((~II12457));
assign g6566 = ((~II11740));
assign g8688 = (g3812&g8342);
assign g9321 = ((~g9311));
assign g4893 = ((~g2460))|((~g4312));
assign g2922 = ((~g2313));
assign II14091 = ((~g7589));
assign II10247 = ((~g5266));
assign II11206 = ((~g6133));
assign g1810 = ((~II5676));
assign II15814 = ((~g9154));
assign II9687 = ((~g4822));
assign g8306 = (g4525&g7951);
assign g5095 = ((~II9476))|((~II9477));
assign II5548 = ((~g1280));
assign g5677 = ((~II10166));
assign II8253 = ((~g2454))|((~g3825));
assign g8284 = ((~II14531));
assign g6274 = ((~II11102))|((~II11103));
assign g7232 = (g6694&g7091);
assign g2226 = ((~g1320));
assign g2902 = ((~g2285));
assign g9131 = (g9055&g5345);
assign II7911 = ((~g2767));
assign g6728 = (g6168)|(g5593);
assign g2958 = ((~g2377));
assign II7908 = ((~g3516));
assign g9171 = (g9146)|(g8962);
assign II15391 = ((~g8917));
assign g8407 = ((~g8013));
assign g3906 = ((~II7504))|((~II7505));
assign g3889 = ((~II7437))|((~II7438));
assign g2364 = ((~II6192));
assign g5100 = ((~II9484));
assign II6842 = ((~g205))|((~g2016));
assign g1975 = ((~g1253));
assign II6220 = ((~g126));
assign g5182 = ((~II9672));
assign g7692 = (g7367&g4430);
assign g5731 = ((~II10250));
assign g6816 = ((~II12319));
assign g2382 = ((~II6248));
assign II12017 = ((~g5847))|((~II12015));
assign g2487 = ((~II6323));
assign II11066 = ((~g5460));
assign II9069 = ((~g4400))|((~g1149));
assign II11686 = ((~g6076));
assign II11094 = ((~g5515))|((~g2734));
assign II8477 = ((~g3014));
assign g2746 = ((~g2259));
assign g8812 = ((~g8443)&(~g8421)&(~II15086));
assign g9065 = ((~II15589));
assign g3589 = ((~II7061));
assign II11428 = ((~g5813));
assign II10360 = ((~g5552))|((~II10359));
assign g4934 = ((~g4125));
assign g6636 = ((~II11900));
assign g6283 = ((~II11157))|((~II11158));
assign II10829 = ((~g5224));
assign g5613 = ((~g4748));
assign g9058 = ((~II15568));
assign g2344 = ((~II6148));
assign II12120 = ((~g5939));
assign g8649 = ((~II14743));
assign g4216 = (II8114&II8115);
assign g7565 = ((~II13865));
assign g2270 = ((~II6015));
assign II11800 = ((~g6164));
assign II7902 = ((~g2709));
assign II15592 = ((~g8989));
assign g6640 = ((~II11908));
assign g3530 = ((~g2185));
assign g8729 = (g2999&g8493);
assign g4490 = (g521&g3192);
assign g5841 = ((~II10538));
assign II13728 = ((~g7439));
assign g2677 = ((~g1664));
assign g8772 = ((~g8585));
assign g5029 = (g212&g3945);
assign g5516 = ((~g4924));
assign II8470 = ((~g2525))|((~g2821));
assign II13435 = ((~g7170));
assign g4573 = ((~g2911));
assign II11607 = ((~g5767));
assign g7118 = ((~II12942));
assign gbuf7 = (g1311);
assign g6794 = ((~II12253));
assign g2940 = ((~II6686));
assign II11666 = ((~g5772));
assign g4686 = ((~II8956))|((~II8957));
assign II9788 = ((~g4711));
assign II7479 = ((~g2502))|((~II7478));
assign g3865 = ((~g2944));
assign g8584 = (g8146&g7034);
assign g6052 = (g1049&g5604);
assign g8979 = (g8919)|(g8813);
assign g7411 = ((~g7202));
assign II7181 = ((~g795))|((~II7179));
assign g8082 = (g7654)|(g7628)|(g7611);
assign g3860 = ((~II7383));
assign II10433 = ((~g5212));
assign g8896 = (g8828)|(g8648);
assign g3849 = ((~II7350));
assign II10744 = ((~g5550))|((~II10743));
assign g3811 = ((~II7269))|((~II7270));
assign II13320 = ((~g7139));
assign g5697 = ((~g2044))|((~g5005));
assign g7060 = ((~g6654));
assign g6832 = ((~II12367));
assign II7588 = ((~g2584));
assign g8957 = ((~II15385));
assign g6498 = ((~II11666));
assign g7551 = ((~II13837));
assign g4272 = (g3233&g3286);
assign g5577 = ((~II10046));
assign g4525 = ((~g2870));
assign g2883 = ((~g2237));
assign II14985 = (g8341)|(g8384)|(g8542);
assign g2362 = ((~II6186));
assign II12400 = ((~g6767));
assign II12032 = ((~g5918))|((~II12031));
assign g6384 = ((~II11479));
assign II5709 = ((~g901));
assign g4107 = (g2625&g2615);
assign g5065 = (g374&g3977);
assign g2706 = ((~g1821));
assign g5772 = ((~g5428)&(~g1888));
assign II14709 = ((~g8198));
assign g8378 = (g677&g7887);
assign g7519 = ((~II13737));
assign g4638 = ((~II8829));
assign II15408 = ((~g8896));
assign II5682 = ((~g168));
assign g4118 = (g995&g3790);
assign g3074 = ((~II6800));
assign II15264 = (g8700)|(g8708)|(g8726)|(g8731);
assign II13854 = ((~g7327));
assign g6946 = ((~II12649));
assign II12179 = ((~g1961))|((~g6163));
assign II6087 = ((~g318));
assign g5189 = ((~II9692))|((~II9693));
assign g6476 = ((~g5939))|((~g5269));
assign g5799 = ((~II10436));
assign g9218 = ((~II15930));
assign II12148 = ((~g5988));
assign II11115 = ((~g5481))|((~g3062));
assign II15693 = ((~g9048));
assign II7011 = ((~g2333))|((~II7009));
assign g8071 = (g7540&g4969);
assign II15190 = ((~g8685));
assign g8730 = (g2863&g8407);
assign II9330 = (g2784&g2770&g2746);
assign II12277 = ((~g6681));
assign g4041 = ((~g2605));
assign g3938 = ((~II7610))|((~II7611));
assign g3802 = ((~g1832));
assign g8842 = (g429&g8564);
assign II15648 = ((~g9044));
assign g5818 = ((~II10479));
assign g7992 = ((~g7557));
assign g1563 = ((~g639));
assign II12062 = ((~g5988));
assign gbuf34 = (g1005);
assign g5286 = ((~g4714));
assign g7780 = ((~II14211));
assign II5568 = ((~g1409));
assign g3693 = ((~g2424));
assign g4820 = ((~II9170))|((~II9171));
assign II11790 = ((~g6282));
assign g6991 = (g5689&g6520);
assign g8878 = (g8777&g6106);
assign g6091 = (g5712&g5038);
assign II12412 = ((~g6404));
assign II6676 = ((~g1603));
assign g3158 = ((~II6853));
assign II9525 = ((~g4413));
assign gbuf41 = (g1146);
assign II6229 = ((~g486));
assign II12852 = ((~g6701))|((~g6695));
assign g8990 = (g8930)|(g8830);
assign g8868 = ((~II15190));
assign g4640 = ((~II8835));
assign g1800 = ((~g1477));
assign II11410 = ((~g5845));
assign g3642 = ((~II7118));
assign II13918 = ((~g7361));
assign II8496 = (g3316&g3287&g2020&g1987);
assign II12430 = ((~g6432));
assign g5442 = (g4679&g4202);
assign g6296 = ((~II11215));
assign g1757 = ((~g604));
assign g8685 = ((~II14851));
assign II12547 = ((~g6708));
assign II12409 = ((~g6398));
assign g7009 = ((~II12753));
assign g6205 = ((~g5628));
assign II12098 = ((~g5956));
assign g2454 = ((~II6294));
assign II15178 = ((~g8753));
assign g6774 = ((~II12193));
assign g9244 = ((~II15974));
assign II6036 = ((~g130));
assign g2459 = ((~II6299));
assign g2784 = ((~g2340));
assign g3878 = ((~g2962));
assign II10479 = ((~g5227));
assign g1661 = ((~g1405));
assign II11458 = ((~g6063));
assign g1694 = ((~g21));
assign II9171 = ((~g4244))|((~II9169));
assign g5719 = ((~II10236));
assign g6846 = ((~II12409));
assign II9965 = ((~g4869))|((~II9963));
assign g1006 = ((~II5410));
assign II8193 = ((~g3547));
assign g6778 = ((~II12205));
assign g8329 = (g527&g7966);
assign g2945 = ((~g2364));
assign g6137 = ((~II10776));
assign g8708 = (g3557&g8407);
assign g6347 = ((~II11368));
assign g8013 = ((~g7561));
assign II13885 = ((~g7351));
assign g7171 = ((~g7071));
assign g6289 = ((~II11194));
assign g6895 = ((~II12558));
assign g6003 = (g3716&g5633&II10597);
assign II5715 = ((~g896));
assign II6066 = ((~g883))|((~II6064));
assign g2311 = ((~II6090));
assign II11467 = ((~g6064));
assign II6686 = ((~g2246));
assign g4232 = ((~g1934)&(~g3591));
assign II11677 = ((~g6076));
assign II6839 = ((~g2185));
assign g6412 = (g158&g6024);
assign g6385 = ((~II11482));
assign g6591 = ((~II11787));
assign g6182 = (g1519&g5199);
assign g3705 = ((~II7204));
assign g6414 = (g673&g6025);
assign g8934 = (g3873&g8766);
assign g5314 = (g1509&g4729);
assign g6332 = ((~II11323));
assign II15953 = ((~g9215));
assign II8237 = (g2298&g2316&g2354);
assign gbuf19 = (g1204);
assign II6905 = ((~g2105))|((~II6904));
assign g4022 = ((~II7785));
assign g4887 = ((~II9234))|((~II9235));
assign II8730 = ((~g3987));
assign g7195 = (g6984&g4226);
assign II12044 = ((~g5847));
assign g8317 = (g547&g8181);
assign II8850 = ((~g4031));
assign II15824 = ((~g9157));
assign g3844 = ((~II7335));
assign g8040 = ((~g7699));
assign II13109 = ((~g7059));
assign g7581 = ((~II13888));
assign g7356 = ((~II13484));
assign II10011 = ((~g4821))|((~II10009));
assign g8866 = ((~II15184));
assign g1798 = ((~II5654));
assign g1701 = ((~II5545));
assign g7608 = (g7367&g4169);
assign g5155 = ((~II9591));
assign II7422 = ((~g2525))|((~II7421));
assign g7532 = ((~II13776));
assign g9314 = ((~II16058));
assign g7041 = (g6734&g5206);
assign g7526 = ((~II13758));
assign II10681 = ((~g5686));
assign II13290 = ((~g7158));
assign g4713 = ((~II9014));
assign g6059 = ((~g5317));
assign g9349 = (g9340&g5690);
assign g7443 = (g7192)|(g3158);
assign g9381 = ((~II16165));
assign II14103 = ((~g7584));
assign II12635 = ((~g6509));
assign g2911 = ((~g2292));
assign g5145 = ((~II9561));
assign II11491 = ((~g6010));
assign g4707 = (g812&g4062);
assign II10018 = ((~g4700))|((~II10017));
assign g4362 = ((~g2810));
assign g5811 = ((~II10466));
assign g7510 = ((~II13710));
assign II8523 = (g3430&g3398&g3359&g3341);
assign g7189 = ((~II13109));
assign g8908 = (g8079)|(g8066)|(g8855);
assign g4410 = (g408&g3160);
assign g6232 = ((~II11031));
assign g5559 = ((~g5132))|((~g1257));
assign II15109 = (g8131)|(g8111)|(g8042)|(g8156);
assign g6145 = (g1489&g5705);
assign g3258 = (g2298&g2316&g2334&g2354);
assign II7428 = ((~g3222))|((~g1541));
assign g7584 = ((~II13897));
assign g3935 = ((~II7602));
assign g7966 = ((~II14291));
assign gbuf54 = (g199);
assign II13676 = ((~g7256));
assign g4465 = ((~g3677));
assign g6763 = ((~II12158));
assign II8956 = ((~g4246))|((~II8955));
assign g6122 = ((~II10752));
assign g8014 = ((~g7564));
assign II6090 = ((~g390));
assign g3723 = ((~g2096));
assign g3358 = ((~II6940))|((~II6941));
assign II12577 = ((~g1049))|((~II12575));
assign g4604 = ((~II8727));
assign g8881 = ((~g8683));
assign g7042 = ((~g6543));
assign II9947 = ((~g2128))|((~II9946));
assign II7167 = ((~g2505));
assign g6132 = (g5436)|(g4793);
assign II9627 = ((~g4777));
assign g5163 = ((~II9615));
assign g5474 = ((~g4904));
assign II10617 = ((~g5677));
assign II16107 = ((~g9337));
assign g2324 = ((~II6115));
assign g5779 = ((~II10384));
assign g8274 = (g4580&g7951);
assign g4578 = ((~g2917));
assign g8267 = (g154&g8042);
assign g3917 = ((~II7548));
assign g4008 = ((~II7755));
assign g8692 = (g3462&g8363);
assign II7438 = ((~g3822))|((~II7436));
assign g5754 = ((~g5403));
assign II11011 = ((~g5693));
assign g3927 = ((~II7584));
assign II8354 = ((~g1163));
assign II10135 = ((~g4960));
assign g8297 = (g429&g7920);
assign g7631 = (g7367&g4187);
assign II7716 = ((~g3038));
assign II9760 = ((~g4838));
assign g6397 = ((~II11512));
assign g6689 = (g1519&g6239);
assign II13203 = ((~g7088));
assign II8150 = ((~g3229))|((~g38));
assign II8418 = (g3316&g3287&g3264&g3238);
assign II13758 = ((~g7414));
assign g2665 = ((~g1661));
assign g5440 = (g4790)|(g4786);
assign g6733 = (g685&g5873);
assign g7775 = ((~II14196));
assign g4034 = ((~II7811));
assign g5463 = ((~g5085));
assign g4377 = (g297&g3131);
assign g8094 = ((~g7705));
assign g6758 = ((~II12145));
assign g3011 = ((~II6751))|((~II6752));
assign g8076 = (g7690&g3521);
assign g7767 = ((~II14172));
assign II7953 = ((~g3542));
assign g2316 = ((~II6109));
assign II5392 = ((~g694));
assign II10739 = ((~g5572));
assign g6178 = ((~g2205))|((~g5568));
assign g9015 = (g8905&g8239);
assign g6025 = ((~g5367));
assign g4193 = (g145&g2727);
assign g4645 = ((~II8850));
assign g5212 = (g5047)|(g4387);
assign g5690 = ((~g4748));
assign II15102 = (II15098)|(II15099)|(II15100)|(II15101);
assign II8679 = ((~g2467))|((~II8678));
assign II12283 = ((~g6692));
assign g2006 = ((~g806));
assign g8832 = (g501&g8585);
assign II13749 = ((~g7313));
assign g7309 = ((~II13359));
assign II6646 = ((~g2246));
assign g8543 = (g706&g7887);
assign g1868 = ((~II5747));
assign g8839 = (g4050&g8581);
assign g8697 = (g3761&g8342);
assign g8150 = (g846&g7658);
assign II13299 = ((~g7163));
assign g9057 = ((~II15565));
assign II15546 = ((~g9007));
assign II7240 = ((~g1658))|((~II7239));
assign g7256 = ((~g7058));
assign II16043 = ((~g9285));
assign g4245 = ((~II8172));
assign II8121 = ((~g3220))|((~II8119));
assign II13410 = ((~g7274));
assign g7502 = ((~II13682));
assign g4653 = ((~II8874));
assign II6029 = ((~g1207));
assign II8041 = (g2074&g2057&g2020&g3238);
assign g1597 = ((~g973));
assign II9840 = ((~g4702));
assign g7737 = ((~II14082));
assign g8714 = (g2873&g8407);
assign g5034 = (g583&g3956);
assign g6306 = ((~II11245));
assign g7293 = ((~II13311));
assign g2872 = ((~II6590));
assign II5948 = ((~g378));
assign g6709 = ((~II12052))|((~II12053));
assign g3996 = ((~II7731));
assign II10482 = ((~g5228));
assign g3519 = ((~g2185));
assign g4015 = ((~g3160));
assign g2506 = ((~II6341));
assign g2350 = ((~II6166));
assign g6580 = (g6039)|(g6041);
assign II15553 = ((~g9009));
assign g2652 = ((~II6440));
assign II8315 = ((~g3691));
assign II6629 = ((~g2052));
assign g4013 = ((~g3131));
assign g7730 = ((~II14061));
assign II8078 = (g2162&g2149&g2137&g2106);
assign g9237 = ((~II15965));
assign g6154 = (g1499&g5713);
assign g4879 = ((~g2595))|((~g2584))|((~g4270))|((~g4281));
assign g4794 = (g954&g4574);
assign g2209 = ((~II5926));
assign g7172 = ((~g7092));
assign g1015 = ((~II5416));
assign II10144 = ((~g1916))|((~II10142));
assign g8637 = (g6057)|(g8071);
assign g2128 = ((~g1284));
assign g7741 = ((~II14094));
assign g1860 = ((~g162));
assign II9845 = ((~g4728));
assign g5079 = (g375&g3990);
assign g7046 = ((~II12806));
assign g4191 = ((~II8084));
assign II9828 = ((~g1509))|((~II9826));
assign II5747 = ((~g1260));
assign II10400 = ((~g5201));
assign g6474 = (g6203&g2424);
assign g7722 = ((~II14039));
assign II16119 = ((~g9351));
assign II16122 = ((~g9353));
assign g7091 = ((~g6525));
assign II5911 = ((~g216));
assign g5578 = ((~g4841));
assign II10953 = ((~g5565))|((~II10952));
assign II7180 = ((~g2351))|((~II7179));
assign g5064 = (g315&g3975);
assign g9046 = (g8744)|(g8749)|(g9016)|(g8862);
assign II15565 = ((~g8980));
assign II14374 = ((~g7693));
assign g5174 = ((~II9648));
assign II9539 = ((~g4018));
assign II9515 = ((~g4301));
assign g4905 = ((~g4282))|((~g3533));
assign II7778 = ((~g3019));
assign g4655 = ((~II8880));
assign g4906 = (g4320&g2728);
assign II13118 = ((~g7068));
assign II13161 = ((~g7080));
assign II13051 = ((~g6967));
assign g6826 = ((~II12349));
assign II9615 = ((~g4739));
assign II6578 = ((~g1603));
assign II12869 = ((~g2536))|((~g6618));
assign g8895 = (g8823)|(g8646);
assign g8674 = ((~II14816));
assign II9768 = ((~g4832))|((~II9767));
assign g8701 = (g2700&g8363);
assign II14677 = ((~g7791));
assign II9116 = ((~g4297));
assign II16090 = ((~g9336));
assign g1802 = ((~g628));
assign g9032 = ((~II15510));
assign g6370 = ((~II11437));
assign II7672 = ((~g3062));
assign g6348 = ((~II11371));
assign g2216 = ((~II5933));
assign g3780 = ((~g1847));
assign g6203 = ((~II10953))|((~II10954));
assign II11389 = ((~g5766));
assign g6482 = ((~g5269))|((~g5847));
assign g6965 = (g55&g6489);
assign g1672 = ((~g1499));
assign g6318 = ((~II11281));
assign g7832 = (g5343&g7599);
assign g7690 = (g4181)|(g7417);
assign g6611 = (g3390&g6249);
assign g5598 = ((~g4938));
assign g7697 = (g7419)|(g3187);
assign g4463 = ((~II8483));
assign g6683 = ((~g6237));
assign g7499 = ((~g7258));
assign II12328 = ((~g6760));
assign g6337 = ((~II11338));
assign II14643 = ((~g7837));
assign g4691 = (g4219&g1690);
assign g3691 = ((~II7195));
assign g8748 = (g2721&g8483);
assign g8177 = ((~II14410));
assign II5852 = ((~g1202));
assign g8656 = ((~g8199)&(~II14758)&(~II14759));
assign g4101 = (g108&g3649);
assign g4298 = ((~II8254))|((~II8255));
assign II10820 = ((~g2039))|((~II10818));
assign g5591 = ((~g4841));
assign g8635 = ((~g1034)&(~g8128));
assign II6877 = ((~g1967))|((~II6876));
assign g9371 = (g9352&g5917);
assign g4541 = ((~g2883));
assign g8828 = (g4573&g8541);
assign g1793 = ((~g626));
assign g5700 = (g1638&g4969);
assign II8282 = ((~g3515));
assign II15297 = (g8280)|(g8257)|(g8319)|(g8327);
assign g8234 = ((~II14489));
assign g6912 = (g4199)|(g6567);
assign g8754 = ((~g8524));
assign g5121 = ((~II9515));
assign II15082 = (g8131)|(g8111)|(g8042)|(g8156);
assign g6515 = ((~g6125));
assign II14112 = ((~g7560));
assign II8874 = ((~g3884));
assign II8618 = (g2074&g3287&g3264&g3238);
assign II12894 = ((~g7009));
assign II12436 = ((~g6635));
assign g5830 = (g5714)|(g5142);
assign g7710 = ((~II14009));
assign g7466 = ((~II13622));
assign g7050 = ((~g6618));
assign g2498 = ((~II6333));
assign g2007 = ((~g1223));
assign g5839 = ((~II10532));
assign g9014 = (g8906&g8239);
assign g5081 = (g455&g3993);
assign g1590 = ((~II5466));
assign gbuf61 = (g109);
assign g5032 = (g313&g3950);
assign g6463 = ((~g5918))|((~g5278));
assign g6880 = ((~II12511));
assign g1867 = ((~g878));
assign II8709 = ((~g4191));
assign II7498 = ((~g2752));
assign g2807 = ((~g1782));
assign g8833 = (g4583&g8562);
assign g6425 = ((~II11556));
assign g5561 = (g4168)|(g4797);
assign g4003 = ((~g3192));
assign g6088 = ((~II10708));
assign g8180 = ((~g7719));
assign II7044 = ((~g2402));
assign g8379 = (g691&g7793);
assign g5643 = ((~II10128));
assign g4504 = (II8568&II8569);
assign II12310 = ((~g6723));
assign II14015 = ((~g7440));
assign g3048 = ((~II6784));
assign g5437 = ((~g5041));
assign g9006 = (g8946)|(g8853);
assign g5671 = ((~II10160));
assign II13635 = ((~g7243));
assign II12340 = ((~g6725));
assign g6854 = ((~II12433));
assign g8627 = ((~g6232))|((~g8091));
assign II14838 = ((~g8660))|((~II14837));
assign g8694 = ((~g7658)&(~g8613)&(~g7634));
assign g8272 = (g158&g8042);
assign g9301 = ((~g9260));
assign g8963 = (g8891&g5317);
assign g7687 = (g6053)|(g7416);
assign g4928 = ((~g4119));
assign g5481 = ((~g4914));
assign II10183 = ((~g5129));
assign g5238 = (g5094)|(g4425);
assign II15152 = (g8483)|(g8464)|(g8514);
assign g9055 = (g8721)|(g8725)|(g9012)|(g8859);
assign II6711 = ((~g1726));
assign g3086 = ((~g1852));
assign g8929 = (g3865&g8759);
assign II5519 = ((~g1087))|((~g1098));
assign II15385 = ((~g8880));
assign II6952 = ((~g1896));
assign g6724 = ((~II12088));
assign g7287 = ((~II13293));
assign II15924 = ((~g9207));
assign g7627 = ((~II13956));
assign g4687 = ((~II8962));
assign II7214 = ((~g815))|((~g2091));
assign g1912 = ((~g1524));
assign g5592 = ((~g4969));
assign g6073 = ((~g5384));
assign g3988 = ((~g3097));
assign g5832 = ((~II10519));
assign II11021 = ((~g5627));
assign II12111 = ((~g5956));
assign g8922 = (g4586&g8750);
assign g4785 = (g1678&g4202);
assign II15501 = ((~g8975));
assign II12292 = ((~g6657));
assign g1877 = ((~g595));
assign g5606 = ((~g4748));
assign g3707 = ((~g2226));
assign g8493 = ((~g8041));
assign g6927 = (g6408)|(g6413);
assign g2996 = ((~g1828));
assign g7121 = ((~II12952))|((~II12953));
assign g6460 = (g6178&g2424);
assign g4632 = ((~II8811));
assign g5751 = ((~II10321))|((~II10322));
assign g7013 = ((~II12757));
assign g7125 = ((~II12965));
assign g6787 = ((~II12232));
assign g6647 = ((~II11923));
assign II8132 = ((~g3232))|((~g1646));
assign II7187 = ((~g2353))|((~II7186));
assign g7183 = (g6132&g7042);
assign II5664 = ((~g916));
assign II8547 = (g3316&g2057&g2020&g3238);
assign g1658 = ((~g1313));
assign g2376 = ((~II6226));
assign g5072 = ((~g4457));
assign g8761 = ((~g8564));
assign g3877 = ((~g2960));
assign g7033 = (g6716&g5190);
assign g5566 = (g3617)|(g4810);
assign g5169 = ((~II9633));
assign gbuf67 = (g646);
assign g6009 = ((~II10605));
assign g3677 = ((~g2485));
assign g4172 = (II8057&II8058);
assign II15041 = (g7855)|(g7838)|(g7905)|(g7870);
assign g6694 = (g6151)|(g5573);
assign g8911 = (g8798&g7688);
assign g6850 = ((~II12421));
assign g7150 = ((~g6952));
assign g2946 = ((~g2365));
assign g4286 = ((~g3790));
assign g4746 = ((~II9076));
assign II11278 = ((~g5780));
assign g5039 = ((~g3924)&(~g3914)&(~g3906)&(~g3899));
assign g7782 = (g4783)|(g7598);
assign g1816 = ((~g767));
assign g2629 = ((~g1574));
assign II15276 = (II15272)|(II15273)|(II15274)|(II15275);
assign g7029 = (g6433)|(g5765);
assign II8853 = ((~g4034));
assign g7773 = ((~II14190));
assign g2205 = ((~g13));
assign g2903 = ((~g2286));
assign g9088 = ((~II15654));
assign gbuf11 = (g1193);
assign g4486 = (II8528&II8529);
assign II11184 = ((~g5474))|((~g3029));
assign g1565 = ((~g649));
assign gbuf25 = (g1396);
assign g5735 = ((~II10262));
assign g6407 = (g5956&g5367);
assign g2467 = ((~II6305));
assign g8060 = (g7535&g4841);
assign g7361 = ((~II13499));
assign g7177 = (g7016&g5586);
assign II6669 = ((~g1698));
assign II16017 = ((~g9264));
assign g8291 = (g122&g8111);
assign g1742 = ((~g1486));
assign g1964 = ((~g1428)&(~g1429));
assign II7850 = ((~g2795));
assign II14118 = ((~g7565));
assign g5571 = ((~II10032));
assign g6166 = (g1509&g5725);
assign g7265 = ((~g7077));
assign II13199 = ((~g7025));
assign g7335 = ((~II13425));
assign II11353 = ((~g5788));
assign II9276 = ((~g2533))|((~g4313));
assign g7231 = ((~II13173));
assign g4079 = ((~II7864));
assign II8011 = ((~g3225));
assign II12427 = ((~g6553));
assign g3521 = ((~g2185));
assign g6039 = (g1037&g5574);
assign II8490 = (g3430&g3398&g3359&g3341);
assign II7568 = ((~g2481))|((~II7567));
assign II9496 = ((~g3971));
assign II9636 = ((~g4802));
assign g2517 = ((~II6348));
assign II13481 = ((~g7254));
assign g5118 = (g479&g4026);
assign II11757 = ((~g1758))|((~g6118));
assign g4568 = ((~g2904));
assign II14046 = ((~g7492));
assign g6906 = (g6715)|(g6726);
assign g9064 = ((~II15586));
assign g4270 = ((~g2573));
assign g4185 = (g2636&g2632);
assign g2877 = ((~g2232));
assign g2510 = ((~g58));
assign g6783 = ((~II12220));
assign g8873 = ((~II15205));
assign g8330 = (g261&g7838);
assign II14208 = ((~g7711));
assign g2238 = ((~II5975));
assign g4025 = ((~II7792));
assign g6834 = ((~II12373));
assign II11221 = ((~g6167));
assign g6188 = ((~II10924))|((~II10925));
assign g4872 = (g1924&g4225&g4224);
assign g6801 = ((~II12274));
assign g3657 = ((~II7145));
assign II8832 = ((~g3936));
assign g5285 = ((~g4841));
assign II13444 = ((~g7282));
assign g5162 = ((~II9612));
assign II12826 = ((~g6441));
assign g9322 = ((~g9313));
assign II10503 = ((~g5235));
assign II8635 = ((~g2481))|((~g2743));
assign II14857 = ((~g8657));
assign g2914 = ((~g2308));
assign gbuf31 = (g966);
assign g2986 = (g806&g1739);
assign II11955 = ((~g5988));
assign g5020 = (g579&g3937);
assign II15663 = ((~g9066));
assign g3528 = ((~g2343)&(~g1391));
assign g1558 = ((~II5435));
assign g5817 = (g5395&g3091);
assign g7353 = ((~II13475));
assign II13003 = ((~g7010))|((~II13002));
assign II15202 = ((~g8797));
assign g3868 = ((~g2948));
assign g3511 = ((~g1616));
assign II12702 = ((~g6497));
assign g2804 = ((~g1796));
assign g8794 = (g8153)|(g8074)|(g8069)|(g8523);
assign g8339 = (g345&g7870);
assign g7198 = ((~II13126));
assign g5205 = (g5034)|(g4380);
assign g4582 = ((~g2922));
assign g2291 = ((~II6057));
assign g6105 = (g5618&g2817);
assign g4577 = ((~g2914));
assign g4801 = ((~II9126));
assign g5427 = ((~g5115));
assign g9270 = (g4748&g9241);
assign g6251 = ((~II11060));
assign II13039 = ((~g6961));
assign g3941 = ((~II7626));
assign g6487 = (g5750&g4969);
assign g6058 = (g5561&g3501);
assign II10743 = ((~g5550))|((~g2100));
assign g9198 = ((~g9187));
assign II6815 = ((~g2052))|((~II6813));
assign g9282 = (g9270)|(g6238);
assign II9089 = ((~g4566));
assign g5796 = ((~II10427));
assign g4086 = (g103&g3629);
assign II7478 = ((~g2502))|((~g3808));
assign g8786 = ((~g8545));
assign g2234 = ((~II5963));
assign g2259 = ((~g1325));
assign g4476 = ((~II8511))|((~II8512));
assign g9105 = ((~II15705));
assign g1680 = ((~II5515));
assign g9187 = ((~II15839));
assign II15308 = ((~g8799));
assign g7920 = ((~II14282));
assign II10862 = ((~g5364));
assign g6732 = (g5874&g5367);
assign II6422 = ((~g1805));
assign g8818 = ((~g8443)&(~g8421)&(~II15102));
assign g1707 = ((~g955));
assign II13422 = ((~g7131));
assign II15985 = ((~g9237));
assign II6048 = ((~g387));
assign g3943 = ((~II7632));
assign g3968 = ((~II7683));
assign g6843 = ((~II12400));
assign II10424 = ((~g5209));
assign II15492 = ((~g8971));
assign g9312 = ((~II16052));
assign g7346 = ((~II13454));
assign II6186 = ((~g138));
assign g2269 = ((~II6012));
assign II7878 = ((~g2829));
assign g6448 = (g5918&g5384);
assign g4082 = (g1296&g3604);
assign g9116 = ((~II15738));
assign g2347 = ((~II6157));
assign II10262 = ((~g5551));
assign II8883 = ((~g4198));
assign g7541 = ((~II13807));
assign g2896 = ((~g2269));
assign II10387 = ((~g5194));
assign g7548 = ((~II13828));
assign g642 = ((~II5377));
assign II16176 = ((~g9385));
assign II8733 = ((~g3996));
assign II11729 = ((~g5772));
assign g7459 = ((~II13617));
assign g6675 = ((~II11981));
assign g9083 = ((~II15641));
assign g3870 = ((~g3466));
assign g4425 = (g536&g2845);
assign g5523 = ((~II9935));
assign II8090 = (g3316&g2057&g2020&g3238);
assign II15513 = ((~g8970));
assign II5649 = ((~g1389));
assign g8322 = (g4559&g7993);
assign II13930 = ((~g7405));
assign II12551 = ((~g6689))|((~II12550));
assign g8745 = (g2982&g8493);
assign g3231 = ((~g1889))|((~g1904));
assign II13924 = ((~g7365));
assign g5742 = ((~II10283));
assign g9340 = ((~II16090));
assign II15263 = (g8313)|(g8297)|(g8310)|(g8690);
assign g7036 = (g6728&g5197);
assign g5826 = ((~II10503));
assign g8858 = (g524&g8585);
assign g3582 = ((~g2407));
assign g5027 = ((~II9369));
assign g2557 = ((~g940));
assign g4590 = ((~g2932));
assign g5716 = (g4962)|(g4356);
assign g2285 = ((~II6039));
assign II5599 = ((~g1481))|((~II5598));
assign g5705 = ((~g4841));
assign g3850 = ((~II7353));
assign g5808 = ((~II10457));
assign II10643 = ((~g5267));
assign II14722 = ((~g8076));
assign g5091 = (g397&g4001);
assign g8810 = ((~II15068));
assign II15253 = (g8698)|(g8711)|(g8722)|(g8716);
assign g6323 = ((~II11296));
assign II13610 = ((~g7227));
assign II14424 = ((~g7652));
assign II14325 = ((~g7713));
assign II8196 = ((~g3654));
assign g8935 = (g3874&g8767);
assign g6573 = ((~g5868));
assign g3635 = ((~g1949));
assign II8560 = ((~g2790))|((~II8558));
assign g3500 = ((~g1616));
assign g6134 = ((~g5428));
assign II7061 = ((~g2457));
assign gbuf39 = (g1157);
assign g8809 = ((~II15065));
assign II7531 = ((~g2487))|((~g3787));
assign II13075 = ((~g6958));
assign g9329 = ((~g9317));
assign g7561 = (g7367&g4163);
assign g7086 = (g4101)|(g6464);
assign II7859 = ((~g2804));
assign II9505 = ((~g4300));
assign g2643 = ((~g1589));
assign g5800 = ((~II10439));
assign g4913 = ((~g4092));
assign g4539 = ((~g2881));
assign II11269 = ((~g5756));
assign II12286 = ((~g6696));
assign II8784 = ((~g3949));
assign II12117 = ((~g5918));
assign g4593 = ((~g2939));
assign g5732 = ((~II10253));
assign g5479 = (g5141&g5037);
assign II14479 = (g7993)|(g7966)|(g7793)|(g7811);
assign II11512 = ((~g5874));
assign g4351 = (g309&g3131);
assign g7719 = ((~g7475));
assign g6919 = (g6771)|(g6394);
assign g1775 = ((~II5620))|((~II5621));
assign II14031 = ((~g7448));
assign g1809 = ((~g759));
assign g6430 = (g5874&g5384);
assign II6946 = ((~g1887));
assign g1689 = ((~g855));
assign g5402 = ((~g5000));
assign II6143 = ((~g1217));
assign g4256 = ((~g3233))|((~g1444));
assign II11230 = ((~g6140));
assign II13617 = ((~g7276));
assign II9477 = ((~g1942))|((~II9475));
assign g4255 = (g3605&g3644&g3635&II8186);
assign g4163 = (II8040&II8041);
assign II12696 = ((~g6503));
assign II8817 = ((~g3935));
assign g7302 = ((~II13338));
assign II5963 = ((~g225));
assign g7007 = (g6627&g5072);
assign g1789 = ((~g1034));
assign II6317 = ((~g1339));
assign II10172 = ((~g4873));
assign II15684 = ((~g9067));
assign II14798 = ((~g8605));
assign g8512 = ((~g8094));
assign g7691 = (g7367&g4427);
assign g9141 = ((~g9129));
assign II15583 = ((~g8986));
assign g4935 = ((~g4202));
assign g4627 = ((~II8796));
assign g2584 = ((~g1646));
assign II6274 = ((~g840))|((~II6273));
assign II6843 = ((~g205))|((~II6842));
assign g2486 = ((~g959));
assign g6275 = ((~II11109))|((~II11110));
assign g7599 = ((~g7450));
assign g8305 = (g362&g7870);
assign II9170 = ((~g1935))|((~II9169));
assign g7607 = (g7325&g4969);
assign g5683 = ((~II10180));
assign g2617 = ((~g1565));
assign g4315 = (g3707&g3728&II8288);
assign g1815 = ((~g760));
assign II11137 = ((~g3052))|((~II11135));
assign II10597 = (g3769&g3754&g3735);
assign g7242 = (g7081&g6899);
assign g3934 = ((~II7599));
assign g6503 = ((~g5269))|((~g5897));
assign g2363 = ((~II6189));
assign g1585 = ((~g724));
assign g6041 = (g5189&g4969);
assign g3887 = ((~II7429))|((~II7430));
assign g1580 = ((~g706));
assign g2286 = ((~II6042));
assign g6106 = ((~g5345));
assign g4734 = (g4469)|(g4448)|(II9038);
assign II5775 = ((~g1240));
assign g5842 = ((~II10541));
assign g6326 = ((~II11305));
assign II6115 = ((~g134));
assign II10393 = ((~g5196));
assign g1732 = ((~g1439));
assign II11725 = ((~g6036));
assign g8128 = (g7566)|(g6910)|(g6452);
assign g8406 = ((~II14614));
assign g6793 = ((~II12250));
assign g3038 = ((~g2092));
assign g4936 = (g214&g3888);
assign g7087 = (g6440&g5311);
assign g6949 = (g5483&g6589);
assign II11903 = ((~g5939));
assign g7104 = ((~II12900));
assign g1919 = (g1098&g1087);
assign g7120 = ((~II12948));
assign II11908 = ((~g5918));
assign II11320 = ((~g5797));
assign g7260 = ((~g7064));
assign g4251 = ((~II8180));
assign II9194 = ((~g4252))|((~g1652));
assign II11897 = ((~g6141));
assign g1760 = ((~II5605));
assign g3557 = ((~g1773));
assign II6767 = ((~g1933));
assign g6637 = ((~II11903));
assign g4605 = ((~II8730));
assign II12912 = ((~g7006));
assign II9142 = ((~g4236));
assign II8119 = ((~g1904))|((~g3220));
assign II8360 = ((~g1186));
assign g8264 = (g105&g8131);
assign II6930 = ((~g1876));
assign g4831 = ((~g3635))|((~g3605))|((~g4220));
assign g8740 = (g2966&g8493);
assign g4070 = ((~II7847));
assign g4780 = ((~II9089));
assign g4727 = (g4417)|(g4172)|(g4163)|(II9029);
assign g3977 = ((~g3160));
assign II13428 = ((~g7167));
assign g5046 = (g314&g3962);
assign II11380 = ((~g5822));
assign II9935 = ((~g4812));
assign g8015 = ((~g7689));
assign g6381 = ((~II11470));
assign g6282 = ((~II11150))|((~II11151));
assign g3531 = ((~g1616));
assign g6727 = (g681&g5846);
assign g2957 = ((~g2376));
assign II5865 = ((~g1206));
assign g7006 = ((~II12748));
assign II12325 = ((~g6755));
assign g4589 = ((~g2930));
assign II11998 = ((~g5918));
assign g4090 = ((~II7892))|((~II7893));
assign g8092 = ((~g7634)&(~g7628)&(~g7616)&(~g7611));
assign g7099 = ((~II12885));
assign II15607 = ((~g8994));
assign g6641 = (g5939&g5494);
assign g2383 = ((~II6251));
assign II10236 = ((~g5014));
assign g2520 = ((~g41));
assign g6920 = (g6395)|(g6399);
assign g2325 = ((~II6118));
assign g6613 = ((~II11835));
assign g7255 = ((~II13209));
assign g6658 = ((~g6224));
assign g1824 = ((~II5706));
assign g4275 = ((~g3790));
assign g6051 = ((~g5246));
assign g7063 = ((~II12826));
assign g4547 = ((~g3466));
assign II8680 = ((~g2706))|((~II8678));
assign g8827 = (g498&g8585);
assign g7412 = (g7121&g4841);
assign g6018 = ((~g5494));
assign II12033 = ((~g5897))|((~II12031));
assign II15921 = ((~g9206));
assign g5213 = (g5048)|(g4388);
assign II7368 = ((~g3018));
assign g8958 = ((~II15388));
assign g8283 = (g267&g7838);
assign II7775 = ((~g3705));
assign g3225 = ((~g1021)&(~g1025)&(~g1889));
assign g6011 = ((~g5494));
assign g6932 = (g6417)|(g6423);
assign g8949 = (g4572&g8790);
assign II6170 = ((~g843))|((~g911));
assign g7437 = ((~II13570));
assign II10890 = ((~g2259))|((~II10888));
assign g6139 = ((~II10780));
assign g7349 = ((~II13463));
assign g9075 = ((~II15619));
assign II13353 = ((~g7231));
assign II14451 = ((~g8172));
assign g3604 = ((~g2407));
assign g5567 = ((~g1879))|((~g4883));
assign g9180 = ((~II15824));
assign II12247 = ((~g6646));
assign II6739 = ((~g195))|((~g1970));
assign II6135 = ((~g916))|((~II6133));
assign g6433 = (g778&g6134);
assign g6559 = ((~g5814))|((~g6109));
assign g8843 = (g507&g8585);
assign II11377 = ((~g5811));
assign II14160 = ((~g7549));
assign g1756 = ((~g533));
assign g3897 = ((~g3131));
assign II7511 = ((~g2992))|((~II7510));
assign g6565 = (g2396)|(g6131)|(g1603);
assign II6741 = ((~g1970))|((~II6739));
assign g8980 = (g8920)|(g8815);
assign II11864 = ((~g5753));
assign g4383 = (g222&g3097);
assign g2365 = ((~II6195));
assign II7139 = ((~g2404))|((~II7138));
assign g8723 = (g2706&g8421);
assign II7308 = ((~g3074));
assign g5115 = ((~II9505));
assign II5619 = ((~g1092))|((~g1130));
assign g9128 = ((~II15762));
assign g9165 = (g9159)|(g9023);
assign g7496 = ((~II13666));
assign g4718 = ((~II9018));
assign g1895 = ((~II5775));
assign II7892 = ((~g2979))|((~II7891));
assign II9476 = ((~g4038))|((~II9475));
assign g5458 = (g4686&g1616);
assign II5972 = ((~g356));
assign g8483 = ((~g8038));
assign g5267 = ((~II9785));
assign g2698 = ((~g1673));
assign g7276 = ((~II13264));
assign II7602 = ((~g2562));
assign II9588 = ((~g4704));
assign g4159 = (g1102&g3498);
assign g2404 = ((~g1276));
assign g6266 = (g1481&g5285);
assign g9294 = (g9274)|(g6230);
assign II7157 = ((~g2331))|((~II7156));
assign g2622 = ((~g1568));
assign g7776 = ((~II14199));
assign II10186 = ((~g5129));
assign g6264 = ((~g5403));
assign II13317 = ((~g7211));
assign g3825 = ((~g1826));
assign g5298 = (g1912&g4814);
assign g8088 = (g837&g7658);
assign II10377 = ((~g5188));
assign g3285 = ((~g1689));
assign g5686 = ((~g5132))|((~g1263));
assign II9132 = ((~g4284));
assign g7206 = ((~II13134));
assign g2979 = (g1494&g1733);
assign g2100 = ((~g1227));
assign g8763 = (g8232)|(II14941)|(II14942);
assign g3954 = ((~II7655));
assign II8808 = ((~g4014));
assign II13395 = ((~g7212))|((~g1057));
assign g3880 = ((~g2965));
assign II7592 = ((~g2712));
assign g4522 = ((~g2867));
assign g7337 = (g7278)|(g4546);
assign II12839 = ((~g6630));
assign II8986 = ((~g4552));
assign g7575 = (g7323)|(g7142);
assign g8917 = ((~II15337));
assign g9281 = ((~II16009));
assign g5558 = ((~II10000))|((~II10001));
assign g6861 = ((~II12454));
assign g6204 = (g5542&g5294);
assign II14366 = (g7566)|(g1030)|(g6664);
assign g4400 = (g1138&g3614);
assign g4569 = ((~g2906));
assign g4571 = ((~g2908));
assign g4921 = ((~g4202));
assign g6971 = (g6424&g4969);
assign g1904 = ((~g1021));
assign II12999 = ((~g7029));
assign II8001 = (g2074&g3287&g2020&g1987);
assign g6894 = ((~g6525));
assign g1878 = ((~g80));
assign g2635 = ((~g1579));
assign g8318 = (g183&g8156);
assign g5669 = ((~II10154));
assign g4475 = ((~g3818));
assign g7764 = ((~II14163));
assign II13599 = ((~g2551))|((~II13598));
assign g7247 = ((~II13199));
assign II12235 = ((~g6634));
assign g3310 = ((~g936)&(~g2557));
assign g9099 = ((~II15687));
assign g6868 = ((~II12475));
assign g7223 = ((~II13161));
assign g2276 = ((~II6029));
assign II10987 = ((~g5609));
assign g5221 = (g5067)|(g4396);
assign g6377 = ((~II11458));
assign II11984 = ((~g6246));
assign g6939 = ((~g6543));
assign g8222 = ((~II14445));
assign g5586 = ((~g4938));
assign g2170 = ((~g1229));
assign g4614 = ((~II8757));
assign g5918 = ((~II10574));
assign g4230 = (g2683&g3491&II8143);
assign II15478 = ((~g8910));
assign II10143 = ((~g4707))|((~II10142));
assign g8513 = (g718&g7937);
assign II11500 = ((~g6219));
assign g2895 = ((~g2268));
assign g4742 = ((~II9064));
assign g8606 = ((~II14683));
assign II14181 = ((~g7725));
assign g9045 = ((~II15539));
assign II15290 = (g8285)|(g8266)|(g8318)|(g8326);
assign II15218 = ((~g8801));
assign II8233 = ((~g3588));
assign g4654 = ((~II8877));
assign II15232 = (II15228)|(II15229)|(II15230)|(II15231);
assign g1808 = ((~g629));
assign g3722 = ((~II7215))|((~II7216));
assign II5763 = ((~g1207));
assign g8693 = (g3798&g8342);
assign II8452 = ((~g2816));
assign g3527 = ((~g1616));
assign g9313 = ((~II16055));
assign g7444 = ((~II13588))|((~II13589));
assign g8441 = (g746&g8018);
assign II11101 = ((~g5491))|((~g2712));
assign g4894 = ((~g4298)&(~g4575)&(~g4563));
assign g8544 = ((~II14657));
assign II12151 = ((~g5847));
assign II6904 = ((~g2105))|((~g1838));
assign gbuf51 = (g1160);
assign g7240 = (g6719&g6894);
assign II8101 = ((~g3259));
assign II6539 = ((~g2555))|((~II6538));
assign g9308 = ((~II16040));
assign g6177 = ((~II10889))|((~II10890));
assign g4370 = ((~II8351));
assign g5291 = ((~g4344))|((~g5002))|((~g4963));
assign II5692 = ((~g906));
assign II15696 = ((~g9050));
assign g4138 = (g2638&g2634);
assign g5810 = ((~II10463));
assign II9948 = ((~g4905))|((~II9946));
assign g1871 = ((~II5754));
assign g8851 = (g284&g8524);
assign g6688 = (g6145)|(g5570);
assign g6497 = ((~g5278))|((~g5847));
assign II9600 = ((~g4698));
assign g5278 = ((~II9794));
assign g9146 = (g9135&g6101);
assign II7377 = ((~g3189));
assign g6131 = ((~g5529));
assign g4555 = ((~g2894));
assign g7585 = ((~II13900));
assign II12806 = ((~g6602));
assign g4695 = ((~II8980));
assign g8298 = (g553&g8181);
assign II9794 = ((~g4778));
assign II11365 = ((~g5826));
assign II14837 = ((~g8660))|((~g1073));
assign II11095 = ((~g5515))|((~II11094));
assign g7527 = ((~II13761));
assign g6097 = ((~g5345));
assign g4131 = (g2630&g2622);
assign g5002 = ((~g4335));
assign g1780 = ((~g614));
assign II5975 = ((~g381));
assign II15839 = ((~g9168));
assign II12511 = ((~g6598));
assign gbuf8 = (g1312);
assign g3563 = ((~g2007));
assign II11109 = ((~g5522))|((~II11108));
assign g6121 = (g5425)|(g4785);
assign II12173 = ((~g5918));
assign II6163 = ((~g402));
assign II11638 = ((~g5847));
assign g7501 = ((~II13679));
assign g4192 = (g1126&g3531);
assign g7117 = ((~II12939));
assign II8351 = ((~g1160));
assign g4244 = ((~g3549))|((~g3533));
assign II15229 = (g8262)|(g8303)|(g8268)|(g8312);
assign g6823 = ((~II12340));
assign g3124 = ((~g1857));
assign g4106 = ((~II7931));
assign g2543 = ((~g1348));
assign II9767 = ((~g4832))|((~g1114));
assign II15101 = (g8363)|(g8342)|(g8407)|(g8386);
assign g4352 = (g387&g3160);
assign II6258 = ((~g837))|((~II6257));
assign g8880 = ((~II15218));
assign g8867 = ((~II15187));
assign g5970 = (g5605&g2424);
assign II15504 = ((~g8967));
assign II13767 = ((~g7486));
assign II13009 = ((~g6935));
assign g4122 = ((~II7973));
assign II13134 = ((~g7017));
assign g7308 = ((~II13356));
assign g4704 = ((~II9001));
assign g8857 = (g446&g8564);
assign II14433 = ((~g8061));
assign g5146 = ((~II9564));
assign g6193 = ((~g1926)&(~g5310));
assign g5473 = ((~g4903));
assign g7286 = ((~II13290));
assign g4391 = (g249&g3097);
assign g2970 = ((~g2394));
assign g6062 = ((~II10675));
assign II7755 = ((~g3019));
assign g6903 = ((~II12582));
assign II8971 = ((~g4464));
assign g2235 = ((~II5966));
assign g6024 = ((~g5494));
assign g2919 = ((~g2311));
assign II8589 = (g2074&g3287&g3264&g3238);
assign II6065 = ((~g852))|((~II6064));
assign g4175 = (g1110&g3502);
assign g3916 = ((~II7545));
assign g4962 = (g457&g3905);
assign g1776 = ((~g608));
assign g4646 = ((~II8853));
assign g2641 = ((~g1587));
assign gbuf27 = (g1402);
assign g7310 = ((~II13362));
assign g2011 = ((~II5847));
assign g4119 = ((~II7964));
assign g6740 = (g4100)|(g6022);
assign g6955 = ((~II12666));
assign g3071 = ((~g1948));
assign II7296 = ((~g2915));
assign g9026 = ((~II15492));
assign g6092 = ((~g5317));
assign g5614 = ((~g3002)&(~g1590)&(~g4714));
assign g2868 = ((~g2223));
assign g6945 = ((~II12646));
assign II5812 = ((~g1243));
assign g8900 = (g8840)|(g8653);
assign g6338 = ((~II11341));
assign g8974 = ((~II15426));
assign g6590 = (g3617)|(g6153);
assign g6714 = ((~II12068));
assign g8989 = (g8929)|(g8829);
assign g3632 = ((~II7101));
assign II15172 = (g8483)|(g8464)|(g8514);
assign g5611 = ((~g4969));
assign II11116 = ((~g5481))|((~II11115));
assign g4005 = ((~II7746));
assign g5334 = (g4887&g2424);
assign II15222 = ((~g8834));
assign g7294 = ((~II13314));
assign g3692 = ((~II7198));
assign gbuf20 = (g1205);
assign g5257 = ((~II9768))|((~II9769));
assign g2310 = ((~II6087));
assign II5542 = ((~g1272));
assign II14804 = ((~g8563));
assign g7217 = (g1142&g6941);
assign II13801 = ((~g7429))|((~II13800));
assign g4870 = (g4154)|(g3081);
assign II15516 = ((~g8977));
assign g4455 = ((~g3811));
assign g9222 = ((~II15940));
assign g9020 = ((~II15484));
assign II6636 = ((~g1704));
assign II13692 = ((~g7343));
assign g6759 = ((~II12148));
assign II9151 = ((~g3883))|((~g1649));
assign g7109 = ((~II12915));
assign g6297 = ((~II11218));
assign II10454 = ((~g5217));
assign II6499 = ((~g1913))|((~g1537));
assign g6159 = ((~II10835))|((~II10836));
assign g8707 = ((~g7658)&(~g8613)&(~g7634));
assign II10071 = ((~g4954))|((~g2253));
assign g3083 = ((~II6814))|((~II6815));
assign gbuf42 = (g1147);
assign g3495 = ((~g1616));
assign II8636 = ((~g2481))|((~II8635));
assign II12382 = ((~g6772));
assign g4692 = ((~II8971));
assign II12180 = ((~g1961))|((~II12179));
assign g8879 = (g8782&g6108);
assign g5150 = ((~II9576));
assign II12460 = ((~g6674));
assign II6864 = ((~g2528));
assign g5156 = ((~II9594));
assign II11778 = ((~g6180));
assign g4888 = ((~g4548)&(~g4528)&(~g4513)&(~g4502));
assign II15394 = ((~g8916));
assign g8776 = ((~g8585));
assign g1970 = ((~II5831));
assign g5008 = (g231&g3920);
assign II14969 = (g8315)|(g8377)|(g8359)|(g8611);
assign g9139 = (g8879)|(g9120);
assign g6069 = ((~II10690));
assign II11718 = ((~g6115));
assign II14442 = ((~g8065));
assign II13743 = ((~g7454));
assign II9057 = ((~g4059))|((~g1504));
assign g8328 = (g4571&g7993);
assign g9370 = ((~II16138));
assign II5374 = ((~g634));
assign g8813 = (g255&g8524);
assign II7734 = ((~g2595));
assign g6773 = ((~II12190));
assign II16145 = ((~g9367));
assign g6908 = (g6478&g5246);
assign II16138 = ((~g9358));
assign g8266 = (g2157&g8042);
assign II15909 = ((~g9201));
assign g7301 = ((~II13335));
assign g2092 = ((~g1225));
assign II6202 = ((~g831))|((~II6201));
assign g7829 = ((~II14251));
assign II15051 = (g8131)|(g8111)|(g8042)|(g8156);
assign II6532 = ((~g1694));
assign g6413 = (g5939&g5367);
assign II12958 = ((~g6920));
assign II10780 = ((~g5445));
assign g9063 = ((~II15583));
assign g5631 = ((~g4938));
assign II6121 = ((~g321));
assign II14484 = (g7993)|(g7966)|(g7793)|(g7811);
assign II16023 = ((~g9267));
assign II11362 = ((~g5821));
assign g1830 = ((~II5718));
assign g8829 = (g267&g8524);
assign g7993 = ((~II14298));
assign II10412 = ((~g5205));
assign II11591 = ((~g5814));
assign g9334 = (g9318&g6205);
assign II9621 = ((~g4732));
assign II13813 = ((~g7314));
assign II8939 = ((~g4239))|((~II8938));
assign II8063 = (g2162&g2149&g2137&g2106);
assign II14318 = ((~g7657));
assign g6525 = (g6112)|(g5547);
assign II12065 = ((~g5897));
assign g4910 = ((~g2460))|((~g4314));
assign II15536 = ((~g9004));
assign g1955 = (g1189)|(g16);
assign II8565 = ((~g3071));
assign g6723 = ((~II12085));
assign g5005 = (g2728&g4320&II9330);
assign II12367 = ((~g6754));
assign g7563 = ((~II13861));
assign II8790 = ((~g4020));
assign II15762 = ((~g9039));
assign II9645 = ((~g4900));
assign II13800 = ((~g7429))|((~g1061));
assign II13605 = ((~g7197));
assign II10786 = ((~g5452));
assign g5082 = (g476&g3994);
assign g8759 = ((~g8524));
assign g7068 = ((~g6556));
assign g6445 = (g6105)|(g6107);
assign II14904 = ((~g8629));
assign g2640 = ((~g1584));
assign g8744 = (g3802&g8464);
assign g4437 = (g540&g2845);
assign II11744 = ((~g6120));
assign g6936 = ((~II12629));
assign g3846 = ((~II7341));
assign g6921 = (g6396)|(g6401);
assign g4688 = (g4193)|(g3190);
assign g6257 = ((~g5685));
assign g4563 = ((~II8659))|((~II8660));
assign g4252 = ((~g2276))|((~g3313));
assign g8840 = (g4590&g8582);
assign g6249 = (g4066)|(g5313);
assign g6806 = ((~II12289));
assign II7532 = ((~g2487))|((~II7531));
assign g4483 = (II8523&II8524);
assign II12038 = ((~g5847));
assign g6756 = ((~II12141));
assign g1834 = (g933&g929);
assign g6996 = (g3678&g6552);
assign g8029 = ((~II14318));
assign g3501 = ((~g2185));
assign II8880 = ((~g4303));
assign g6632 = ((~II11890));
assign II12690 = ((~g6467));
assign g1688 = ((~II5535));
assign II8940 = ((~g1545))|((~II8938));
assign II8569 = (g3316&g2057&g2020&g1987);
assign g3648 = ((~g2424));
assign II7891 = ((~g2979))|((~g1499));
assign g6510 = ((~g5278))|((~g5874));
assign II10574 = ((~g5426));
assign g2642 = ((~g1588));
assign II6018 = ((~g462));
assign g1786 = ((~g623));
assign g4813 = ((~II9162));
assign II11401 = ((~g5828));
assign g6169 = ((~II10867))|((~II10868));
assign g5600 = ((~g5128));
assign g7611 = (g7367&g4507);
assign g8181 = ((~II14420));
assign g8216 = ((~II14427));
assign g7434 = ((~II13565));
assign g5626 = ((~g4748));
assign g2349 = ((~II6163));
assign g4591 = ((~g2937));
assign g3462 = ((~g1743));
assign g7579 = ((~II13882));
assign g1572 = ((~g673));
assign II10193 = ((~g4670));
assign II10766 = ((~g5674));
assign g6496 = ((~II11662));
assign g2795 = ((~g1801));
assign II11787 = ((~g6273));
assign g1908 = ((~g812));
assign II10605 = ((~g5440));
assign g4741 = ((~II9058))|((~II9059));
assign g5016 = ((~II9350));
assign II10649 = ((~g5657));
assign II14728 = ((~g8152));
assign II12810 = ((~g6607));
assign g7422 = ((~II13541));
assign II13072 = ((~g6969));
assign g5243 = (g5106)|(g4435);
assign II7623 = ((~g3631));
assign g6630 = ((~II11884));
assign II8898 = ((~g4089));
assign g5092 = (g456&g4002);
assign g4087 = ((~II7882));
assign g8312 = (g365&g7870);
assign g5403 = ((~g5088));
assign g6700 = ((~g6244));
assign g4200 = ((~II8105));
assign g2966 = ((~g1856));
assign g6851 = ((~II12424));
assign g6897 = ((~II12564));
assign II11497 = ((~g6014));
assign g7182 = (g6902&g4969);
assign g5438 = (g1545&g4932);
assign g9323 = ((~g9315));
assign II14388 = ((~g7605));
assign g2817 = ((~g1849));
assign II15262 = (g8293)|(g8283)|(g8304)|(g8289);
assign g9130 = (g9054&g5345);
assign II15982 = ((~g9236));
assign g5137 = ((~II9539));
assign g8822 = (g417&g8564);
assign g6237 = ((~II11040));
assign II10010 = ((~g1949))|((~II10009));
assign g4474 = ((~II8503))|((~II8504));
assign II15181 = ((~g8734));
assign II13378 = ((~g1472))|((~II13376));
assign II9058 = ((~g4059))|((~II9057));
assign II10761 = ((~g5302));
assign II5422 = ((~g1234));
assign g5749 = ((~g5207));
assign g8308 = (g510&g7966);
assign g4130 = ((~II7987));
assign II12211 = ((~g6502));
assign II11047 = ((~g5653));
assign g6508 = ((~II11686));
assign II11515 = ((~g5897));
assign II8868 = ((~g4035));
assign II8980 = ((~g4535));
assign g2424 = ((~g1329));
assign g9117 = ((~II15741));
assign g2654 = ((~II6446));
assign II7978 = ((~g3574));
assign II13865 = ((~g7333));
assign II6203 = ((~g891))|((~II6201));
assign g8321 = (g446&g7920);
assign g5652 = ((~II10135));
assign g6615 = ((~II11842))|((~II11843));
assign g4271 = (g3666&g3684);
assign g3653 = ((~g2459));
assign g6317 = ((~II11278));
assign g7749 = ((~II14118));
assign II11616 = ((~g1519))|((~II11614));
assign g4806 = ((~II9139));
assign g5657 = ((~g5021))|((~g4381));
assign g8791 = ((~g8585));
assign g6907 = (g6727)|(g6732);
assign II10313 = ((~g5484))|((~g1041));
assign g8271 = (g130&g8111);
assign g9388 = ((~II16180));
assign g6163 = ((~g5633))|((~g3716));
assign g3518 = ((~II6997))|((~II6998));
assign g4036 = ((~g3192));
assign g9209 = ((~g9199));
assign g9104 = ((~II15702));
assign II10954 = ((~g2340))|((~II10952));
assign g3617 = ((~g1655));
assign II9443 = ((~g4564));
assign II11575 = ((~g5894))|((~II11574));
assign g8700 = (g3784&g8342);
assign II13425 = ((~g7166));
assign II7320 = ((~g2927));
assign II10343 = ((~g5704));
assign g2904 = ((~g2287));
assign g7166 = (g6437)|(g6914);
assign g2470 = ((~g42));
assign g8609 = (g7828&g4969);
assign II7632 = ((~g3634));
assign g3853 = ((~II7362));
assign g2352 = ((~II6171))|((~II6172));
assign g9071 = ((~II15607));
assign g4026 = ((~g3192));
assign g5480 = ((~g4913));
assign II5600 = ((~g1489))|((~II5598));
assign g2649 = ((~II6431));
assign g8334 = (g264&g7838);
assign g6603 = ((~II11815));
assign II14073 = ((~g7627));
assign II8766 = ((~g3960));
assign g6800 = ((~II12271));
assign g5426 = ((~g5013));
assign g6087 = ((~II10705));
assign g2905 = ((~II6629));
assign g6216 = ((~II10987));
assign II16168 = ((~g9381));
assign g7032 = ((~g6525));
assign II7010 = ((~g2295))|((~II7009));
assign g1726 = ((~g158));
assign g5769 = ((~II10380));
assign g7332 = ((~II13416));
assign II10522 = ((~g5243));
assign g8146 = (g6045)|(g7597);
assign g2514 = ((~g1330));
assign g4319 = (g3728&g3694&g3750&II8296);
assign II13189 = ((~g7002));
assign g3096 = ((~II6834));
assign g5161 = ((~II9609));
assign g2985 = ((~II6733));
assign g5096 = (g1149&g4400);
assign g4452 = (g437&g3160);
assign II7800 = ((~g2605));
assign g6734 = (g6176)|(g5599);
assign II10625 = ((~g5314))|((~g1514));
assign g8964 = (g8915)|(g8863)|(II15400);
assign II13332 = ((~g7241));
assign g4694 = ((~II8977));
assign g5214 = (g5049)|(g4389);
assign g6737 = ((~II12111));
assign g6782 = ((~II12217));
assign g1911 = ((~II5789));
assign II7517 = ((~g3578));
assign g6036 = ((~II10643));
assign g5114 = ((~II9502));
assign g7092 = ((~II12866));
assign II6270 = ((~g492));
assign g4594 = ((~g2941));
assign II12358 = ((~g6761));
assign II6072 = ((~g1211));
assign g3947 = ((~II7640));
assign II14334 = ((~g7578));
assign g2231 = ((~II5954));
assign g7311 = ((~II13365));
assign g6820 = ((~II12331));
assign g4375 = (g219&g3097);
assign II12813 = ((~g6607));
assign II10818 = ((~g5567))|((~g2039));
assign g5204 = (g5033)|(g4379);
assign g5311 = ((~g4938));
assign II13580 = ((~g7208));
assign g4829 = (g863)|(g4051);
assign g8042 = ((~II14325));
assign g6917 = (g6743)|(g6753);
assign g2621 = ((~g1567));
assign II7551 = ((~g2712));
assign g9102 = ((~II15696));
assign g4297 = (g3617)|(g3602);
assign g3547 = ((~g2345));
assign g639 = ((~II5374));
assign g3909 = ((~II7520));
assign g8585 = ((~g7993));
assign g6674 = ((~II11978));
assign II13787 = ((~g1477))|((~II13785));
assign II9889 = ((~g4819));
assign II14219 = (g979)|(g7566)|(g1865);
assign g2264 = ((~II5997));
assign g8154 = (g6054)|(g7607);
assign g9362 = ((~II16122));
assign g8971 = ((~II15417));
assign II10157 = ((~g5109));
assign g4032 = ((~II7807));
assign II5847 = ((~g1360));
assign II13559 = ((~g7177));
assign II15495 = ((~g8973));
assign g4424 = (g489&g3192);
assign II10867 = ((~g5480))|((~II10866));
assign g5572 = (g5051)|(g1236);
assign II11482 = ((~g6117));
assign II5861 = ((~g1313));
assign g1686 = ((~II5531));
assign II11078 = ((~g5697))|((~g2511));
assign II10361 = ((~g1118))|((~II10359));
assign g7436 = (g7183)|(g6975);
assign g5042 = ((~II9396));
assign g1582 = ((~g714));
assign g8819 = ((~g8443)&(~g8421)&(~II15113));
assign II6057 = ((~g518));
assign II5697 = ((~g1524))|((~II5695));
assign g6947 = ((~II12652));
assign g5021 = (g943)|(g4501);
assign II13048 = ((~g6956));
assign II6695 = ((~g2246));
assign g4868 = (g4227&g4160);
assign g9094 = ((~II15672));
assign II9009 = ((~g4591));
assign II10962 = ((~g5719));
assign II10000 = ((~g4839))|((~II9999));
assign II12472 = ((~g6591));
assign g7035 = ((~g6543));
assign g3605 = ((~g1938));
assign g3831 = ((~II7296));
assign g5579 = (g4090&g4841);
assign g8179 = ((~II14416));
assign g2395 = ((~II6274))|((~II6275));
assign g7688 = ((~g7406));
assign II10789 = ((~g5512))|((~g2170));
assign g9304 = ((~g9298));
assign II6740 = ((~g195))|((~II6739));
assign g2346 = ((~II6154));
assign g2210 = ((~g1326));
assign g8231 = ((~II14473))|((~II14474));
assign g5237 = (g5093)|(g4424);
assign g3567 = ((~g2407));
assign II9585 = ((~g4697));
assign g5538 = ((~g5132))|((~g1266));
assign II10300 = ((~g2562))|((~II10298));
assign g7058 = ((~g6649));
assign g1603 = ((~II5471));
assign g9205 = ((~II15898))|((~II15899));
assign g7594 = ((~II13927));
assign II15484 = ((~g8918));
assign g3573 = ((~g2424));
assign II11124 = ((~g2712))|((~II11122));
assign g8928 = (g4595&g8757);
assign gbuf62 = (g287);
assign g3890 = ((~II7444))|((~II7445));
assign g5362 = ((~II9823));
assign II12681 = ((~g6469));
assign g4023 = ((~II7788));
assign II9534 = (g3019&g3029&g3038&g3052);
assign g7689 = (g7367&g4417);
assign g8913 = ((~II15329));
assign g5522 = ((~g4930));
assign g4190 = (g1122&g3527);
assign II13472 = ((~g7266));
assign II12936 = ((~g7015));
assign g5897 = ((~II10569));
assign II12544 = ((~g6617));
assign g3674 = ((~II7164));
assign g6648 = ((~II11926));
assign II9025 = ((~g4462));
assign II11479 = ((~g6201));
assign g9217 = ((~II15927));
assign g6244 = ((~g5670));
assign g636 = ((~II5371));
assign g9372 = ((~II16142));
assign II10380 = ((~g5448));
assign g4357 = ((~g3679));
assign II7069 = ((~g1639))|((~II7068));
assign g2284 = ((~II6036));
assign g7279 = ((~II13271));
assign g3588 = ((~g2379));
assign g6143 = ((~II10796));
assign g8799 = ((~II15007));
assign g1901 = ((~II5781));
assign g6303 = ((~II11236));
assign II10040 = ((~g2202))|((~II10038));
assign II8401 = (g3316&g3287&g3264&g3238);
assign II6151 = ((~g12));
assign II8568 = (g3430&g3398&g3359&g3341);
assign II14157 = ((~g7547));
assign II8019 = (g3430&g3398&g3359&g2106);
assign II12609 = ((~g6571));
assign g1819 = ((~II5696))|((~II5697));
assign II15261 = (g8256)|(g8271)|(g8267)|(g8286);
assign g7281 = ((~II13277));
assign g7323 = (g4065&g7171);
assign II6326 = ((~g1443));
assign g7318 = ((~g7185)&(~g6979));
assign II8928 = ((~g4153));
assign g6696 = ((~II12022));
assign g8906 = (g8088)|(g8062)|(g8699);
assign g8847 = ((~g8493)&(~g8239)&(~II15147));
assign g2292 = ((~II6060));
assign II15610 = ((~g8995));
assign g6367 = ((~II11428));
assign II9609 = ((~g4780));
assign g5781 = ((~II10390));
assign g8299 = (g591&g8181);
assign II13518 = ((~g7141));
assign II11656 = ((~g5772));
assign g6652 = ((~II11936));
assign g6291 = ((~II11200));
assign gbuf14 = (g1197);
assign g5587 = ((~g4938));
assign II10369 = ((~g5716));
assign g6008 = ((~g5367));
assign II12307 = ((~g6712));
assign g5833 = ((~II10522));
assign II11732 = ((~g6076));
assign g6786 = ((~II12229));
assign g4444 = ((~II8452));
assign II8245 = ((~g3506))|((~II8243));
assign g8993 = (g8933)|(g8835);
assign g4776 = ((~II9081));
assign II11191 = ((~g6155));
assign g3900 = ((~II7486))|((~II7487));
assign g6760 = ((~II12151));
assign II9570 = ((~g4696));
assign II8593 = (g3430&g3398&g3359&g2106);
assign II5817 = ((~g1081));
assign II16026 = ((~g9267));
assign II15842 = ((~g9171));
assign g8910 = ((~II15324));
assign g3997 = ((~II7734));
assign II16132 = ((~g9356));
assign II9834 = ((~g4782));
assign II8143 = (g2674&g2677&g2680);
assign g7124 = ((~g6896));
assign g5168 = ((~II9630));
assign g7770 = ((~II14181));
assign g7493 = ((~II13659));
assign g6928 = (g6409)|(g6415);
assign II8180 = ((~g3529));
assign g6596 = ((~II11800));
assign II7140 = ((~g2397))|((~II7138));
assign g5843 = ((~g5367));
assign g8632 = ((~II14712));
assign g4580 = ((~g2919));
assign g5580 = ((~g4938));
assign g9138 = (g8878)|(g9119);
assign II14792 = ((~g8583));
assign g4626 = ((~II8793));
assign II10488 = ((~g5230));
assign II14637 = ((~g8012));
assign II9850 = ((~g4798));
assign II15113 = (II15109)|(II15110)|(II15111)|(II15112);
assign g2821 = ((~g1786));
assign g7790 = ((~II14227));
assign II11641 = ((~g5918));
assign II13311 = ((~g7162));
assign g5086 = ((~II9460));
assign g5648 = ((~g4748));
assign II15595 = ((~g8990));
assign g8752 = ((~g8564));
assign g7704 = ((~II14001));
assign II15817 = ((~g9151))|((~g9148));
assign g2880 = ((~g2234));
assign g1673 = ((~g1504));
assign g8715 = (g2761&g8386);
assign g8286 = (g180&g8156);
assign g6855 = ((~II12436));
assign g5190 = ((~g4938));
assign g9067 = ((~II15595));
assign g4269 = (g2354&g3563&II8209);
assign g2327 = ((~II6124));
assign g7130 = ((~II12976));
assign g1897 = ((~g789));
assign II6876 = ((~g1967))|((~g1910));
assign g8459 = (g655&g7793);
assign g7447 = ((~II13599))|((~II13600));
assign g2501 = ((~g27));
assign II10509 = ((~g5237));
assign II8841 = ((~g3979));
assign II7510 = ((~g2992))|((~g1711));
assign II10592 = ((~g5444));
assign g8259 = (g4538&g7855);
assign II12424 = ((~g6446));
assign g9238 = (g4748&g9223);
assign II11335 = ((~g5839));
assign g6835 = ((~II12376));
assign g4016 = ((~g3192));
assign g7789 = ((~II14224));
assign II8503 = ((~g2986))|((~II8502));
assign g2871 = ((~II6587));
assign g9350 = ((~II16100));
assign g6467 = ((~g5956))|((~g5269));
assign g8292 = (g181&g8156);
assign g2862 = ((~II6578));
assign g6717 = (g4082)|(g6005);
assign II5416 = ((~g8868));
assign g6677 = ((~II11987));
assign g6473 = ((~g5269))|((~g5988));
assign g7476 = ((~g7229));
assign g5597 = ((~g4969));
assign g6010 = ((~II10608));
assign g4389 = (g480&g3192);
assign II14687 = ((~g7826));
assign g4748 = ((~g4465));
assign II10497 = ((~g5233));
assign g3641 = ((~II7115));
assign II14473 = ((~g8147))|((~II14472));
assign g6020 = ((~g5367));
assign g4014 = ((~II7769));
assign g4302 = (g3086&g3659&g3124);
assign II13002 = ((~g7010))|((~g1053));
assign g4102 = ((~II7919));
assign g4735 = (g4427)|(g4414)|(g4403)|(II9041);
assign g6047 = (g1477&g5596);
assign gbuf21 = (g1271);
assign II5969 = ((~g303));
assign II15899 = ((~g9203))|((~II15897));
assign g4078 = (g3753&g3732&g3712&g3700);
assign g8080 = (g7467&g7634);
assign II8919 = ((~g4196));
assign g4280 = (II8224)|(II8225);
assign II12945 = ((~g7066));
assign II12632 = ((~g6514));
assign II10448 = ((~g5335));
assign g3987 = ((~II7716));
assign II13666 = ((~g7238));
assign g6682 = ((~II11994));
assign II6917 = ((~g2360))|((~II6916));
assign g4745 = ((~II9070))|((~II9071));
assign II10998 = ((~g5672));
assign g9082 = ((~II15638));
assign II12256 = ((~g6647));
assign g1639 = ((~g1207));
assign II7667 = ((~g3052));
assign g9003 = (g8943)|(g8849);
assign g6881 = ((~II12514));
assign g4074 = (g137&g3573);
assign g5615 = ((~g4714)&(~g3002));
assign g2764 = ((~g1802));
assign II10500 = ((~g5234));
assign II12316 = ((~g6736));
assign II13164 = ((~g7086));
assign g7736 = ((~II14079));
assign g8078 = (g7463&g7634);
assign g4676 = ((~g3885)&(~g3094));
assign g7479 = ((~II13635));
assign g4369 = (g580&g2845);
assign II12564 = ((~g6720));
assign g4909 = ((~II9271));
assign g5124 = ((~II9520));
assign g5590 = ((~g2044))|((~g4906));
assign II7468 = ((~g1704))|((~II7466));
assign g9005 = (g8945)|(g8852);
assign g8178 = ((~II14413));
assign g2893 = ((~II6615));
assign II8799 = ((~g3951));
assign II10614 = ((~g5302));
assign II11455 = ((~g6087));
assign g5056 = ((~g3556)&(~g2872)&(~g3938));
assign g8887 = (II15265)|(g8819);
assign g9190 = ((~II15849))|((~II15850));
assign II7738 = ((~g3038));
assign g4791 = (g949&g4562);
assign II6657 = ((~g1701));
assign II14001 = ((~g7433));
assign g5827 = ((~II10506));
assign g2528 = ((~g1260));
assign g6387 = ((~II11488));
assign II13752 = ((~g7315));
assign g4528 = ((~II8606))|((~II8607));
assign II6471 = ((~g1923));
assign g5710 = (g4958)|(g4351);
assign II11245 = ((~g6143));
assign g5871 = ((~II10558));
assign g8217 = ((~II14430));
assign g6597 = ((~II11803));
assign II13956 = ((~g7499));
assign g9051 = ((~II15553));
assign g6944 = ((~II12643));
assign II15298 = (g8332)|(g8333)|(g8686)|(g8702);
assign g7765 = ((~II14166));
assign g2326 = ((~II6121));
assign g6290 = ((~II11197));
assign II7429 = ((~g3222))|((~II7428));
assign II13088 = ((~g7045));
assign g8073 = ((~g7658)&(~g7654));
assign II9963 = ((~g1938))|((~g4869));
assign g1855 = ((~g866));
assign g8973 = ((~II15423));
assign g4523 = ((~g2868));
assign g6422 = (g714&g6033);
assign II10320 = ((~g5459))|((~g2573));
assign g6452 = ((~g6270)&(~g2245));
assign g1805 = ((~II5667));
assign g8706 = ((~g7658)&(~g8613)&(~g7634));
assign g9178 = ((~II15814));
assign g5448 = ((~g5137));
assign g5556 = ((~II9986))|((~II9987));
assign g5764 = ((~II10369));
assign g6410 = ((~II11533));
assign II10307 = ((~g3019))|((~II10305));
assign II13574 = ((~g7205));
assign g4384 = (g246&g3097);
assign g8992 = (g8932)|(g8832);
assign II6257 = ((~g837))|((~g901));
assign g7700 = (g7367&g4494);
assign g4320 = (g3728&g3750&g3768&II8299);
assign g8732 = (g3808&g8464);
assign II6294 = ((~g1330));
assign g6095 = ((~II10719));
assign g8016 = ((~II14311));
assign II6788 = ((~g1681));
assign II11923 = ((~g5939));
assign g7703 = (g7367&g4504);
assign II15589 = ((~g8988));
assign g6661 = ((~II11961));
assign g6267 = ((~II11086));
assign g7582 = ((~II13891));
assign II6015 = ((~g437));
assign g4408 = (g330&g3131);
assign g4099 = (g117&g3647);
assign g6585 = (g3617)|(g6119);
assign g5284 = ((~g4344))|((~g4335))|((~g4963));
assign g4902 = (g4304&g2770&g2746&g2728);
assign g5175 = ((~II9651));
assign g4668 = ((~II8919));
assign g4673 = ((~II8928));
assign II6538 = ((~g2555))|((~g2557));
assign II15699 = ((~g9061));
assign g2502 = ((~II6337));
assign g6520 = ((~II11704));
assign II11747 = ((~g6123));
assign II14758 = (g7993)|(g7966)|(g7793)|(g7811);
assign g8691 = (g3805&g8342);
assign g4142 = (II8005&II8006);
assign g7057 = ((~g6644));
assign g1770 = ((~g606));
assign g2573 = ((~g1649));
assign g6098 = (g5681&g1247);
assign g5790 = ((~II10415));
assign g2840 = ((~g2207));
assign g5180 = ((~II9666));
assign II8152 = ((~g38))|((~II8150));
assign g1017 = ((~II5419));
assign II10946 = ((~g5563));
assign g6979 = (g5095&g6511);
assign II16148 = ((~g9368));
assign g9143 = (g9122&g6089);
assign g4281 = ((~g2562));
assign II10299 = ((~g5461))|((~II10298));
assign II5419 = ((~g1603));
assign g4360 = ((~II8333));
assign g5685 = ((~II10186));
assign II10796 = ((~g5397));
assign g1864 = ((~g162));
assign g3964 = ((~g3160));
assign II15978 = ((~g9235));
assign g6538 = ((~II11714));
assign g9303 = ((~g9301));
assign II9791 = ((~g4779));
assign II10094 = ((~g2177))|((~II10092));
assign g4125 = ((~II7978));
assign g4055 = (g187)|(g3012);
assign II8528 = (g3430&g3398&g3359&g2106);
assign II5386 = ((~g648));
assign II13506 = ((~g7148));
assign g2452 = ((~g23));
assign II15272 = (g8237)|(g8300)|(g8261)|(g8282);
assign g3808 = ((~g1827));
assign II5795 = ((~g1236));
assign g6867 = ((~II12472));
assign g4885 = ((~g4070));
assign II12672 = ((~g6473));
assign II11648 = ((~g6028));
assign g6722 = ((~II12079))|((~II12080));
assign g9333 = ((~g9323));
assign g5557 = ((~II9993))|((~II9994));
assign g5187 = ((~II9687));
assign II10991 = ((~g5632))|((~g2389));
assign II8108 = (g2162&g2149&g2137&g2106);
assign II12973 = ((~g6927));
assign II12993 = ((~g6933));
assign II9980 = ((~g2092))|((~II9978));
assign II14680 = ((~g7810));
assign g8864 = ((~II15178));
assign g3818 = ((~II7278))|((~II7279));
assign g7266 = ((~II13238));
assign g4651 = ((~II8868));
assign g5784 = ((~II10397));
assign g1739 = (g803&g799);
assign g1779 = ((~g612));
assign g8230 = ((~g8199)&(~II14467)&(~II14468));
assign g9358 = (g9279)|(g9348);
assign g3959 = ((~g3097));
assign g8220 = ((~II14439));
assign g3591 = ((~g1789));
assign g8221 = ((~II14442));
assign g7530 = ((~II13770));
assign g9383 = ((~g9380));
assign II7362 = ((~g2933));
assign g6027 = ((~g5384));
assign g5730 = ((~II10247));
assign g4641 = ((~II8838));
assign g8386 = ((~g8014));
assign g4367 = (g240&g3097);
assign g6378 = ((~II11461));
assign II9691 = ((~g5096))|((~g1037));
assign II6680 = ((~g1558));
assign g6735 = (g4091)|(g6013);
assign g2942 = ((~g2350));
assign g6353 = ((~II11386));
assign g2949 = (g822&g1753);
assign g6983 = ((~II12722));
assign g3524 = ((~g2306));
assign g9017 = ((~II15475));
assign g6959 = ((~II12678));
assign g1781 = ((~g622));
assign g2782 = ((~g1616));
assign II12717 = ((~g6543));
assign II15021 = (II15017)|(II15018)|(II15019)|(II15020);
assign g3510 = ((~g2185));
assign II11404 = ((~g5834));
assign g6042 = (g1041&g5581);
assign g7128 = (g6926&g3047);
assign II9095 = ((~g4283));
assign g7016 = (g6042)|(g6487);
assign g4554 = ((~g2892));
assign II8057 = (g3430&g3398&g3359&g3341);
assign g7524 = ((~II13752));
assign g2947 = ((~II6695));
assign II8642 = (g3430&g3398&g3359&g2106);
assign g8155 = (g7632)|(g3219);
assign g7504 = ((~II13692));
assign gbuf52 = (g1182);
assign gbuf57 = (g92);
assign II14430 = ((~g7836));
assign II8588 = (g3430&g3398&g3359&g3341);
assign g9162 = (g9158)|(g9022);
assign II6006 = ((~g306));
assign II15239 = (g8264)|(g8260)|(g8277)|(g8301);
assign g6218 = ((~II10992))|((~II10993));
assign g7187 = ((~II13103));
assign g2927 = ((~II6663));
assign g6916 = (g727&g6515);
assign g6120 = (g3617)|(g5555);
assign II14813 = ((~g8640));
assign gbuf1 = (g1240);
assign g4729 = (g1504&g4059);
assign g8440 = (g714&g7937);
assign g8269 = (g4569&g7951);
assign II14282 = ((~g7709));
assign g5013 = ((~II9341));
assign II7922 = ((~g3462));
assign g9258 = (g9227&g5628);
assign g8683 = ((~g8235));
assign II6109 = ((~g1214));
assign II11615 = ((~g6239))|((~II11614));
assign II8659 = ((~g2471))|((~II8658));
assign g4313 = ((~g3712))|((~g3700));
assign g3587 = ((~g1964));
assign g9315 = ((~II16061));
assign g4544 = ((~g2886));
assign II10079 = ((~g4911))|((~II10078));
assign gbuf32 = (g963);
assign g7445 = (g4192)|(g7193);
assign g4647 = ((~II8856));
assign g4963 = ((~g4328));
assign g6791 = ((~II12244));
assign gbuf48 = (g1155);
assign g4576 = ((~g2913));
assign g9255 = ((~II15985));
assign II10565 = ((~g5402));
assign II11752 = ((~g1486))|((~II11750));
assign g2952 = (g2474&g2215);
assign g5795 = ((~II10424));
assign g7034 = ((~g6525));
assign g1747 = ((~g599));
assign g6180 = ((~II10900))|((~II10901));
assign g1866 = ((~g71));
assign g7739 = ((~II14088));
assign II9166 = (g4041&g2595&g2584);
assign g9010 = (g8950)|(g8860);
assign g6394 = (g5988&g5494);
assign II15717 = ((~g9051));
assign g9368 = ((~II16132));
assign g4968 = (g4403&g1760);
assign g4705 = (g190&g3986);
assign II13725 = ((~g7437));
assign gbuf28 = (g1403);
assign g5701 = ((~g5120));
assign g5484 = (g1037&g5096);
assign g9019 = ((~II15481));
assign II6774 = ((~g2386))|((~g1134));
assign II12575 = ((~g6574))|((~g1049));
assign g8545 = ((~g7905));
assign g2521 = ((~g65)&(~g62));
assign g4390 = (g560&g2845);
assign g9248 = ((~II15978));
assign g2309 = ((~II6084));
assign g7343 = ((~II13447));
assign g3937 = ((~g2845));
assign g6478 = ((~II11638));
assign g6761 = ((~II12154));
assign g8734 = ((~II14904));
assign g5255 = (g5118)|(g4453);
assign II6663 = ((~g2246));
assign g4711 = (g190&g4072);
assign II12742 = ((~g6590));
assign II13255 = ((~g7057));
assign g5755 = ((~g5494));
assign II14743 = ((~g8174));
assign g2628 = ((~g1573));
assign g8739 = (g3780&g8464);
assign g8835 = (g270&g8524);
assign II13308 = ((~g7169));
assign g2263 = ((~g1394));
assign II9145 = ((~g4264));
assign g8888 = (II15276)|(g8807);
assign II9657 = ((~g4784));
assign g7273 = ((~II13255));
assign g2287 = ((~II6045));
assign II7156 = ((~g2331))|((~g929));
assign II14294 = ((~g7553));
assign g2869 = ((~g2224));
assign II8020 = (g2074&g3287&g2020&g1987);
assign II10558 = ((~g5264));
assign g5266 = ((~II9782));
assign g9220 = ((~g9205));
assign II11549 = ((~g5984))|((~g1045));
assign g4105 = ((~II7928));
assign g5461 = ((~g4885));
assign II14055 = ((~g7495));
assign g1879 = ((~II5763));
assign II10472 = ((~g5223));
assign g3226 = (g1102&g1919);
assign II15776 = ((~g9127));
assign g6399 = (g5971&g5494);
assign g3700 = ((~g2514));
assign II14990 = (g8337)|(g8379)|(g8543);
assign g2378 = ((~II6233))|((~II6234));
assign g7225 = ((~g6936));
assign II5872 = ((~g77));
assign II5754 = ((~g966));
assign II9782 = ((~g4720));
assign II12952 = ((~g7003))|((~II12951));
assign g1246 = ((~II5425));
assign II9573 = ((~g4701));
assign g3079 = ((~g1603));
assign g3574 = ((~g1771));
assign II9475 = ((~g4038))|((~g1942));
assign II14381 = ((~g7596));
assign g4841 = ((~g4250));
assign g4154 = (g1098&g3495);
assign II12496 = ((~g6592));
assign g5229 = (g5079)|(g4409);
assign II10541 = ((~g5256));
assign g2240 = ((~II5981));
assign II15044 = (II15040)|(II15041)|(II15042)|(II15043);
assign g3264 = ((~II6900));
assign g7216 = ((~II13152));
assign II9675 = ((~g4807));
assign g4814 = (g150&g4265);
assign g7545 = ((~II13819));
assign g6149 = ((~II10810));
assign II15498 = ((~g8974));
assign g6403 = ((~II11522));
assign II6172 = ((~g911))|((~II6170));
assign II12053 = ((~g5939))|((~II12051));
assign g8311 = (g4540&g7905);
assign g7134 = ((~II12986));
assign g3461 = ((~II6959));
assign g3316 = ((~II6930));
assign g7291 = ((~II13305));
assign g5007 = ((~II9336));
assign II8164 = ((~g1943))|((~g3231));
assign II15753 = ((~g9080));
assign g7248 = (g7079)|(g5652);
assign II9994 = ((~g4871))|((~II9992));
assign II9277 = ((~g2533))|((~II9276));
assign g1843 = ((~g771));
assign g6860 = ((~II12451));
assign II7564 = ((~g2752));
assign II13837 = ((~g7324));
assign g2636 = ((~g1580));
assign II11951 = ((~g5847));
assign II10327 = ((~g5467))|((~g2562));
assign g7558 = ((~II13850));
assign g1646 = ((~g1214));
assign II6733 = ((~g1718));
assign g7758 = ((~II14145));
assign g8463 = ((~g8094));
assign g8773 = (II14959)|(II14960);
assign g1715 = ((~II5559));
assign g6273 = ((~II11095))|((~II11096));
assign II13825 = ((~g7318));
assign g2639 = ((~g1583));
assign g6814 = ((~II12313));
assign g5023 = ((~g3894)&(~g3889)&(~g3886)&(~g4359));
assign g5739 = ((~II10274));
assign g8948 = (g4570&g8789);
assign II13496 = ((~g7133));
assign II13407 = ((~g7271));
assign g2478 = ((~g31));
assign II7635 = ((~g3052));
assign II9774 = ((~g4678));
assign g9336 = ((~II16084));
assign g8326 = (g258&g7838);
assign II9148 = ((~g4354));
assign g4098 = (g985&g3790);
assign g1952 = ((~g1333));
assign g691 = ((~II5389));
assign g8675 = ((~II14819));
assign g2471 = ((~II6309));
assign II6759 = ((~g1983))|((~II6757));
assign II9183 = ((~g2007))|((~II9181));
assign g7557 = (g7367&g4147);
assign g3953 = ((~g3160));
assign g5144 = ((~II9558));
assign g6002 = (g5539&g2407);
assign g7280 = ((~II13274));
assign g4615 = ((~II8760));
assign g3746 = ((~g2100));
assign II6764 = ((~g1955));
assign g7088 = (g6638)|(g6641);
assign g8686 = (g3819&g8342);
assign g2937 = ((~g2346));
assign g6627 = ((~II11874))|((~II11875));
assign g7261 = ((~II13225));
assign II10847 = ((~g5490))|((~g2595));
assign II12271 = ((~g6663));
assign g4296 = ((~g3790));
assign g3061 = ((~II6795));
assign g5195 = (g5019)|(g4368);
assign g4231 = ((~g2276))|((~g3258));
assign II6844 = ((~g2016))|((~II6842));
assign g2699 = ((~g1674));
assign II10046 = ((~g4840));
assign II12241 = ((~g6640));
assign g6339 = ((~II11344));
assign gbuf59 = (g99);
assign g1812 = ((~II5682));
assign g6223 = ((~II11008));
assign g4955 = (g215&g3891);
assign II14298 = ((~g7678));
assign II7359 = ((~g2871));
assign g5063 = (g294&g3974);
assign II10166 = ((~g5016));
assign II7875 = ((~g3819));
assign g6887 = ((~II12532));
assign g3222 = (g1537&g1913);
assign II11419 = ((~g5835));
assign g8464 = ((~g8039));
assign II12942 = ((~g7023));
assign g4301 = ((~II8264));
assign g6278 = ((~II11129));
assign II8536 = ((~g2506))|((~g2798));
assign g8405 = (g741&g8018);
assign g7415 = (g7222&g5603);
assign g4781 = (g4182&g1760);
assign g6103 = ((~g5317));
assign II7115 = ((~g2547));
assign g8950 = (g4582&g8791);
assign g2457 = ((~g24));
assign g4696 = ((~II8983));
assign g5019 = (g312&g3933);
assign g7405 = ((~II13518));
assign g2380 = ((~II6242));
assign g6343 = ((~II11356));
assign II9946 = ((~g2128))|((~g4905));
assign g1823 = ((~g768));
assign II6443 = ((~g1774));
assign II15888 = ((~g9192))|((~II15887));
assign g2963 = ((~g2383));
assign g2828 = ((~g1980));
assign II7548 = ((~g3590));
assign II10032 = ((~g1236));
assign g8263 = (g4555&g7905);
assign II7138 = ((~g2404))|((~g2397));
assign g9047 = ((~II15543));
assign II6060 = ((~g580));
assign g4167 = (g2783&g1616);
assign gbuf6 = (g1310);
assign g7740 = ((~II14091));
assign II6831 = ((~g2185));
assign g3888 = ((~g3097));
assign g6948 = ((~II12655));
assign II6154 = ((~g122));
assign g2148 = ((~g1304));
assign g3976 = ((~II7697));
assign g6054 = (g1057&g5611);
assign II12596 = ((~g6582))|((~g1126));
assign II13761 = ((~g7418));
assign g6607 = ((~II11827));
assign g4279 = ((~g3340));
assign g8894 = (g8817)|(g8645);
assign g6001 = (g5540&g2407);
assign g7694 = (g7367&g4448);
assign g6285 = ((~II11171))|((~II11172));
assign II12980 = ((~g6929));
assign g9033 = ((~II15513));
assign g6638 = (g174&g5755);
assign II14474 = ((~g1069))|((~II14472));
assign g8145 = ((~II14381));
assign g9126 = ((~II15756));
assign g2886 = ((~g2240));
assign II11900 = ((~g5847));
assign g4937 = (g3086&g4309);
assign II13441 = ((~g7146));
assign g6811 = ((~II12304));
assign g3832 = ((~II7299));
assign g8939 = (g3879&g8772);
assign g6874 = ((~II12493));
assign II10080 = ((~g2256))|((~II10078));
assign II10937 = ((~g5560));
assign g6254 = ((~g5683));
assign II6354 = ((~g1357));
assign II8261 = ((~g3643));
assign g7116 = ((~II12936));
assign g4836 = ((~g4288))|((~g1879));
assign g2660 = ((~II6451));
assign g8770 = ((~g8545));
assign g2348 = ((~II6160));
assign II7595 = ((~g2573));
assign II15254 = (II15250)|(II15251)|(II15252)|(II15253);
assign g1945 = ((~g1081));
assign II11485 = ((~g6137));
assign g6195 = ((~II10940));
assign g3924 = ((~II7568))|((~II7569));
assign II10336 = ((~g2573))|((~II10334));
assign II9746 = ((~g4826))|((~II9745));
assign g2360 = ((~g1435));
assign g4586 = ((~g2926));
assign g7103 = ((~II12897));
assign g6726 = (g5897&g5367);
assign g2397 = ((~g1272));
assign g2801 = ((~II6539))|((~II6540));
assign II15112 = (g8363)|(g8342)|(g8407)|(g8386);
assign g703 = ((~II5398));
assign g6570 = ((~II11751))|((~II11752));
assign II7107 = ((~g2480));
assign II7758 = ((~g2605));
assign g6642 = ((~II11912));
assign II8962 = ((~g4553));
assign g8726 = (g2795&g8386);
assign g4083 = (g125&g3610);
assign g8093 = ((~II14370));
assign g7413 = ((~II13524));
assign g6501 = ((~II11669));
assign g8300 = (g126&g8111);
assign II11260 = ((~g5779));
assign g5717 = ((~g4969));
assign II8748 = ((~g3997));
assign II6239 = ((~g8));
assign II12753 = ((~g6445));
assign II9752 = ((~g4705));
assign g6998 = (g4474&g6555);
assign g2616 = ((~g1564));
assign g4876 = (g4159)|(g4167);
assign II5478 = ((~g1148));
assign g6071 = ((~II10694));
assign II8273 = ((~g2976));
assign II9594 = ((~g4718));
assign g3863 = ((~II7392));
assign g5699 = (g1667&g4841);
assign g4621 = ((~II8778));
assign g5493 = ((~g4920));
assign g4344 = ((~g3124));
assign II10548 = ((~g5260));
assign g4139 = (II8000&II8001);
assign g7517 = ((~II13731));
assign g7077 = ((~g6676));
assign g5089 = (g273&g3998);
assign g4497 = (II8551&II8552);
assign g7715 = ((~II14022));
assign g2224 = ((~II5945));
assign g5109 = ((~II9493));
assign II14214 = ((~g7576));
assign II12760 = ((~g6685));
assign II14085 = ((~g7583));
assign II13466 = ((~g7122));
assign g2353 = ((~g871));
assign II7473 = ((~g3546));
assign g5104 = (g274&g4010);
assign II11806 = ((~g6275));
assign g7580 = ((~II13885));
assign II12385 = ((~g6397));
assign II11917 = ((~g5897));
assign g4037 = ((~g2845));
assign g4807 = ((~II9142));
assign g7748 = ((~II14115));
assign g5425 = (g1528&g4916);
assign g7406 = ((~g7191)&(~g1600));
assign g3485 = ((~g1737));
assign II13356 = ((~g7221));
assign g3655 = ((~g1844));
assign gbuf16 = (g1200);
assign II14079 = ((~g7579));
assign g7165 = (g6434)|(g6908);
assign g5633 = ((~g4895));
assign II6024 = ((~g544));
assign II11374 = ((~g5844));
assign g8337 = (g498&g7966);
assign g9103 = ((~II15699));
assign g9101 = ((~II15693));
assign g5581 = ((~g4969));
assign g8270 = (g110&g8131);
assign II12361 = ((~g6765));
assign gbuf37 = (g1081);
assign g7333 = ((~II13419));
assign II6440 = ((~g1806));
assign g3546 = ((~II7029));
assign II8678 = ((~g2467))|((~g2706));
assign II16116 = ((~g9350));
assign II15379 = ((~g8882));
assign g8792 = ((~II14996));
assign g7837 = (g6470&g7610);
assign g6161 = ((~II10842));
assign g9226 = (g9220&g5403);
assign II8268 = ((~g2801));
assign g2912 = (g1080&g1945);
assign g2965 = ((~g2384));
assign g2873 = ((~g1779));
assign g8871 = ((~II15199));
assign g6061 = (g5257&g1616);
assign II14267 = ((~g7695));
assign g4318 = ((~g3681)&(~g1590));
assign II14454 = ((~g8177));
assign g6836 = ((~II12379));
assign g7448 = ((~II13605));
assign II10314 = ((~g5484))|((~II10313));
assign g4007 = ((~II7752));
assign g5335 = ((~g4677));
assign g6769 = ((~II12176));
assign g3652 = ((~II7132));
assign II10321 = ((~g5459))|((~II10320));
assign g7325 = ((~II13396))|((~II13397));
assign II15791 = ((~g9140));
assign g8237 = (g89&g8131);
assign II13238 = ((~g6900));
assign II13023 = ((~g7040));
assign g1685 = ((~II5528));
assign g1727 = ((~g596));
assign II13909 = ((~g7339));
assign g5453 = ((~g4680));
assign II16009 = ((~g9261));
assign g9216 = ((~II15924));
assign g2879 = ((~II6597));
assign g4376 = (g243&g3097);
assign g6037 = ((~II10646));
assign g3509 = (g1637&g1616);
assign II11356 = ((~g5799));
assign g4077 = (g1284&g3582);
assign II7792 = ((~g3038));
assign II12280 = ((~g6684));
assign g9159 = (g9138&g6074);
assign g2935 = (g1612&g1077);
assign g7300 = ((~II13332));
assign II9123 = ((~g4455));
assign g2648 = ((~II6428));
assign II9014 = ((~g3864));
assign g3948 = ((~g3131));
assign g8853 = (g365&g8545);
assign g6164 = ((~II10848))|((~II10849));
assign II11987 = ((~g6278));
assign g3526 = ((~g2185));
assign g3640 = ((~II7112));
assign g6852 = ((~II12427));
assign II10868 = ((~g2605))|((~II10866));
assign g9280 = ((~II16006));
assign II10626 = ((~g5314))|((~II10625));
assign g5113 = ((~II9499));
assign g4462 = ((~II8480));
assign II15628 = ((~g9001));
assign II11867 = ((~g6286));
assign g6466 = ((~II11615))|((~II11616));
assign II15747 = ((~g9042));
assign g2401 = ((~g22));
assign g9380 = ((~g9379));
assign II10427 = ((~g5210));
assign II12059 = ((~g5874));
assign II11395 = ((~g5812));
assign II11407 = ((~g5841));
assign g9208 = ((~g9198));
assign II13274 = ((~g6917));
assign g6552 = ((~II11722));
assign II8094 = ((~g2976));
assign g6578 = (g6218&g3913);
assign g3908 = ((~II7517));
assign g9079 = ((~II15631));
assign g1652 = ((~g1220));
assign g3830 = ((~II7293));
assign g1910 = ((~g1435))|((~g1439));
assign g8153 = (g852&g7658);
assign g6918 = ((~II12609));
assign II12930 = ((~g7019));
assign II16129 = ((~g9355));
assign II9325 = ((~g4242));
assign II6084 = ((~g240));
assign II10804 = ((~g5526));
assign g5573 = (g3011&g4841);
assign g4084 = ((~II7875));
assign II14960 = (g8621)|(g8622)|(g8628)|(g8230);
assign II11586 = ((~g6256));
assign g8816 = (g336&g8545);
assign II13126 = ((~g6949));
assign II12768 = ((~g6718));
assign g1787 = ((~g625));
assign II15741 = ((~g9083));
assign g5625 = ((~g2044))|((~g4957));
assign II13782 = ((~g7498));
assign g1807 = ((~g619));
assign g2394 = ((~II6270));
assign g9137 = (g8877)|(g9118);
assign g5022 = ((~g4438));
assign g3872 = ((~g2954));
assign g8199 = ((~II14424));
assign g9024 = (g8884&g5317);
assign g4423 = (g465&g3192);
assign g6245 = ((~g5690));
assign II15068 = ((~g8638));
assign II10415 = ((~g5397));
assign g4562 = ((~g3466));
assign g9196 = ((~g9185));
assign g2894 = ((~g2267));
assign g8320 = (g4557&g7951);
assign g8743 = ((~g8524));
assign g7433 = ((~II13562));
assign g7429 = (g1057&g7212);
assign g3430 = ((~II6956));
assign g9179 = ((~II15818))|((~II15819));
assign g6935 = (g6429)|(g6431);
assign g1687 = ((~g10));
assign g6633 = (g5526&g5987);
assign g6702 = ((~II12038));
assign g3961 = ((~g3131));
assign II12265 = ((~g6660));
assign g4911 = ((~g4320))|((~g2044));
assign g8805 = ((~g8443)&(~g8421)&(~II15033));
assign g7133 = ((~II12983));
assign II15687 = ((~g9071));
assign g1566 = ((~g652));
assign g2888 = ((~II6608));
assign II14130 = ((~g7592));
assign II9666 = ((~g4931));
assign g9145 = ((~II15791));
assign II5679 = ((~g911));
assign II12493 = ((~g6587));
assign II12439 = ((~g6566));
assign II12448 = ((~g6569));
assign g6934 = (g6422)|(g6430);
assign II14718 = ((~g8068));
assign g4253 = ((~g2734));
assign g5083 = ((~g4457));
assign II10826 = ((~g5434));
assign II11981 = ((~g6246));
assign II14205 = ((~g7710));
assign II5766 = ((~g1254));
assign g6889 = ((~II12538));
assign g9070 = ((~II15604));
assign g5093 = (g477&g4003);
assign II9745 = ((~g4826))|((~g1549));
assign II13819 = ((~g7426));
assign g7870 = ((~II14270));
assign II6245 = ((~g142));
assign II9234 = ((~g4310))|((~II9233));
assign g7578 = ((~II13879));
assign g4201 = (II8108&II8109);
assign II8637 = ((~g2743))|((~II8635));
assign II7617 = ((~g3008))|((~II7616));
assign g3666 = ((~g2134));
assign g9324 = ((~II16072));
assign g7258 = (g7083)|(g5403)|(II13220);
assign g4535 = ((~g2876));
assign g5240 = ((~II9752));
assign g8825 = (g342&g8545);
assign II11680 = ((~g5939));
assign g5802 = ((~II10445));
assign II7723 = ((~g3052));
assign II8072 = (g3316&g3287&g2020&g3238);
assign g3131 = (g1749)|(g368);
assign g4635 = ((~II8820));
assign g7421 = (g6745)|(g7202);
assign g6631 = ((~II11887));
assign II9278 = ((~g4313))|((~II9276));
assign g4665 = ((~II8910));
assign g2960 = ((~g2381));
assign g1571 = ((~g669));
assign II13447 = ((~g7261));
assign II12532 = ((~g6594));
assign II6195 = ((~g405));
assign g4088 = ((~II7885));
assign g8955 = ((~II15379));
assign II12961 = ((~g6921));
assign II7844 = ((~g3784));
assign II9612 = ((~g4776));
assign II6597 = ((~g1970));
assign g1898 = (g959&g955);
assign II10705 = ((~g5463));
assign g7717 = ((~II14028));
assign g7515 = ((~II13725));
assign g1811 = ((~II5679));
assign II8218 = ((~g3002));
assign g4392 = (g303&g3131);
assign II15562 = ((~g8979));
assign II15337 = ((~g8802));
assign g9278 = (g9252&g5658);
assign II12394 = ((~g6759));
assign g2655 = ((~g1611));
assign g2283 = ((~II6033));
assign g3839 = ((~II7320));
assign II10306 = ((~g5470))|((~II10305));
assign g1666 = ((~g1472));
assign g4089 = ((~II7888));
assign II12523 = ((~g6624));
assign g9118 = (g9046&g5345);
assign g1777 = ((~g611));
assign g9066 = ((~II15592));
assign II11102 = ((~g5491))|((~II11101));
assign g2794 = ((~g2185));
assign g4473 = (g518&g3192);
assign g6256 = ((~II11069));
assign II13377 = ((~g7199))|((~II13376));
assign g2236 = ((~II5969));
assign II7503 = ((~g2498))|((~g3802));
assign g5688 = ((~II10193));
assign II12208 = ((~g6496));
assign II8594 = (g3316&g2057&g2020&g1987);
assign g3879 = ((~g2963));
assign g7127 = ((~g6974));
assign g1587 = ((~g734));
assign II14463 = ((~g8072));
assign II7299 = ((~g2961));
assign g1674 = ((~g1514));
assign g5036 = (g4047)|(g2972);
assign g8751 = ((~g8545));
assign g7123 = ((~II12961));
assign II8660 = ((~g2724))|((~II8658));
assign g8285 = (g118&g8111);
assign g4721 = ((~II9025));
assign II11108 = ((~g5522))|((~g2734));
assign g6891 = ((~II12544));
assign g3590 = ((~II7064));
assign g5645 = ((~g4748));
assign g8893 = (g8814)|(g8643);
assign g7720 = ((~II14035));
assign II8989 = ((~g4537));
assign g5043 = (g213&g3958);
assign g6808 = ((~II12295));
assign g6409 = (g706&g6020);
assign g2481 = ((~II6317));
assign g8482 = ((~g8094));
assign g453 = ((~II5362));
assign II15930 = ((~g9209));
assign II6916 = ((~g2360))|((~g1732));
assign g2615 = ((~g1563));
assign II9059 = ((~g1504))|((~II9057));
assign g6718 = (g4083)|(g6006);
assign g4176 = (II8063&II8064);
assign II13057 = ((~g6968));
assign g2225 = ((~II5948));
assign g2761 = ((~g1820));
assign g8258 = (g142&g8111);
assign g4052 = (g1276&g3522);
assign g2536 = ((~g1354));
assign g5844 = ((~II10545));
assign II14844 = ((~g8641));
assign g4268 = (g2216&g2655);
assign g4073 = (g1300&g3567);
assign g6856 = ((~II12439));
assign g4747 = (g3984)|(g2912);
assign g2180 = ((~g1318));
assign II11338 = ((~g5798));
assign g6785 = ((~II12226));
assign II10204 = ((~g5060));
assign II14109 = ((~g7590));
assign g4011 = ((~II7762));
assign II8910 = ((~g4200));
assign g6246 = ((~II11055));
assign g9002 = (g8942)|(g8848);
assign g7788 = (g4794)|(g7604);
assign g7015 = ((~II12763));
assign g6211 = ((~g5645));
assign g5472 = ((~II9892));
assign g9239 = (g7653)|(g9226);
assign II8255 = ((~g3825))|((~II8253));
assign g7738 = ((~II14085));
assign g5123 = (g516&g4033);
assign g8079 = (g831&g7658);
assign II7658 = ((~g2562));
assign g3492 = ((~II6970));
assign g1849 = ((~II5732));
assign g9004 = (g8944)|(g8851);
assign g5789 = ((~II10412));
assign II11437 = ((~g5801));
assign g1856 = ((~g774));
assign g4792 = ((~II9111));
assign g4890 = ((~g4075));
assign g6517 = ((~II11701));
assign g4448 = (II8460&II8461);
assign g4581 = ((~g2921));
assign II7467 = ((~g2982))|((~II7466));
assign II13042 = ((~g6963));
assign g5055 = ((~g4477));
assign II10896 = ((~g5475));
assign g6325 = ((~II11302));
assign g6046 = (g1073&g5592);
assign II10142 = ((~g4707))|((~g1916));
assign g6676 = ((~II11984));
assign g6418 = (g5897&g5494);
assign II11416 = ((~g5829));
assign g4407 = (g252&g3097);
assign g8771 = ((~g8564));
assign g2668 = ((~g1662));
assign II12322 = ((~g6751));
assign g8008 = ((~g7559));
assign g6831 = ((~II12364));
assign g6096 = ((~g5317));
assign II8559 = ((~g2502))|((~II8558));
assign II8393 = ((~g2949))|((~II8392));
assign g2863 = ((~g1778));
assign g4693 = ((~II8974));
assign g4317 = (g878&g3086&g1857&g3659);
assign g6423 = (g5897&g5384);
assign g9353 = ((~II16107));
assign g8633 = ((~g8176))|((~g6232));
assign II9084 = ((~g4358));
assign II9241 = ((~g2540))|((~g4305));
assign g4092 = ((~II7899));
assign II7148 = ((~g799))|((~g1974));
assign g7705 = (g7367&g4514);
assign II12202 = ((~g6481));
assign g7699 = (g7367&g4486);
assign g8988 = (g8928)|(g8827);
assign II12274 = ((~g6672));
assign II13031 = ((~g6984));
assign g7735 = ((~II14076));
assign g4368 = (g318&g3131);
assign g6383 = ((~II11476));
assign g8038 = ((~g7694));
assign g6595 = ((~g6083));
assign II14061 = ((~g7546));
assign II15937 = ((~g9212));
assign II10535 = ((~g5254));
assign II9107 = (g4133)|(g4145)|(g4138)|(g4132);
assign g1795 = ((~II5649));
assign g7652 = (g7367&g4194);
assign II12418 = ((~g6572));
assign g4918 = ((~g4103));
assign g5126 = (g556&g4037);
assign g6963 = ((~II12690));
assign g6781 = ((~II12214));
assign II14783 = ((~g8324));
assign g5483 = (g4740)|(g4098);
assign gbuf45 = (g1167);
assign II14495 = (g7993)|(g7966)|(g7793)|(g7811);
assign gbuf69 = (g878);
assign g5167 = ((~II9627));
assign g4787 = (g953&g4547);
assign g4024 = ((~g3160));
assign II15165 = (g8483)|(g8464)|(g8514);
assign II14238 = ((~g7608));
assign g4602 = ((~II8721));
assign II13900 = ((~g7356));
assign g7027 = (g3390&g6698);
assign g4891 = ((~g4076));
assign II6813 = ((~g210))|((~g2052));
assign g9077 = ((~II15625));
assign g3974 = ((~g3131));
assign g4810 = ((~II9152))|((~II9153));
assign gbuf13 = (g1196);
assign II8838 = ((~g3967));
assign II11031 = ((~g5335));
assign II7746 = ((~g3591));
assign g3602 = ((~II7069))|((~II7070));
assign II12514 = ((~g6605));
assign II11117 = ((~g3062))|((~II11115));
assign II8938 = ((~g4239))|((~g1545));
assign g9204 = ((~II15894));
assign II5839 = ((~g1198));
assign g7435 = (g6052)|(g7182);
assign II14154 = ((~g7558));
assign II13707 = ((~g7420));
assign g1938 = ((~g1288));
assign g1612 = ((~II5475));
assign g7793 = ((~II14234));
assign g7340 = ((~II13438));
assign g5153 = ((~II9585));
assign II6750 = ((~g1733))|((~g1494));
assign g5674 = ((~g5042));
assign g9247 = (g4748&g9227);
assign g8914 = (g8795&g8239);
assign g7366 = ((~II13512));
assign g3675 = ((~II7167));
assign g6649 = ((~II11929));
assign g6209 = ((~g2332)&(~g5305));
assign g7220 = (g1304)|(g7062);
assign g5679 = ((~II10172));
assign g6711 = ((~II12059));
assign g6470 = (g5817)|(g2934);
assign g7059 = ((~g6538));
assign g8279 = ((~g7658)&(~g7616)&(~g8082)&(~g7634));
assign II10350 = ((~g5707));
assign g5236 = (g5092)|(g4423);
assign g9059 = ((~II15571));
assign g7322 = ((~g7188)&(~g6991));
assign g2232 = ((~II5957));
assign II13685 = ((~g1977))|((~g7237));
assign g6304 = ((~II11239));
assign g9373 = ((~II16145));
assign II8658 = ((~g2471))|((~g2724));
assign II9535 = (g3062&g2712&g4253&g2752);
assign g7564 = (g7367&g4172);
assign II8172 = ((~g3524));
assign g3050 = ((~II6788));
assign II12022 = ((~g5874));
assign g7811 = ((~II14238));
assign g7271 = (g6436&g6922);
assign g4926 = ((~g4202));
assign g7155 = ((~II13039));
assign II11284 = ((~g5795));
assign g5176 = ((~II9654));
assign g7727 = ((~II14052));
assign II7095 = ((~g2539));
assign g6653 = ((~II11939));
assign g5834 = ((~II10525));
assign II16052 = ((~g9291));
assign gbuf38 = (g1156);
assign g9110 = ((~II15720));
assign II7454 = ((~g1106))|((~II7452));
assign II7068 = ((~g1639))|((~g1643));
assign g4697 = ((~II8986));
assign II5620 = ((~g1092))|((~II5619));
assign II13157 = ((~g6997));
assign g5539 = ((~II9947))|((~II9948));
assign II12008 = ((~g5897));
assign g6007 = ((~g5494));
assign g4689 = ((~II8966));
assign g7319 = ((~g7124));
assign II11079 = ((~g5697))|((~II11078));
assign g8608 = ((~II14687));
assign g7471 = ((~g7233));
assign II13502 = ((~g7135));
assign II11123 = ((~g5517))|((~II11122));
assign II13451 = ((~g7262));
assign II6000 = ((~g202));
assign g7031 = (g3390&g6717);
assign g7762 = ((~II14157));
assign g7152 = ((~g6253)&(~g7083)&(~g5418));
assign g5015 = ((~II9347));
assign g4243 = ((~II8165))|((~II8166));
assign g4618 = ((~II8769));
assign g3712 = ((~g1952));
assign g4288 = (g3563&g3579&g3603&II8240);
assign II6093 = ((~g468));
assign g3339 = (g1424)|(g2014);
assign g8458 = (g756&g8199);
assign II12421 = ((~g6486));
assign g4198 = ((~II8101));
assign g5384 = ((~II9837));
assign II12897 = ((~g6962));
assign g5868 = ((~II10555));
assign g8942 = (g4522&g8780);
assign II9350 = ((~g4503));
assign g4469 = (II8495&II8496);
assign g6292 = ((~II11203));
assign II15240 = (g8259)|(g8294)|(g8263)|(g8305);
assign g3078 = ((~g1603));
assign II5914 = ((~g1097));
assign g5658 = ((~g4748));
assign II14251 = ((~g7541));
assign II13843 = ((~g7326));
assign g6602 = (g6058)|(g3092);
assign g1909 = ((~g998));
assign g4659 = ((~II8892));
assign g5588 = (g3028&g4969);
assign II15613 = ((~g8996));
assign g7771 = ((~II14184));
assign g4358 = ((~g3680));
assign II10776 = ((~g5576));
assign g8927 = (g4594&g8756);
assign g8625 = ((~g1000)&(~g6573)&(~g1860)&(~g8009));
assign II5654 = ((~g921));
assign II7882 = ((~g2700));
assign II11693 = ((~g6076));
assign g4903 = ((~g4084));
assign g4799 = (g951&g4596);
assign g3764 = ((~g2039));
assign g5517 = ((~g4925));
assign II13600 = ((~g7244))|((~II13598));
assign II12454 = ((~g6581));
assign II7561 = ((~g2562));
assign II13659 = ((~g7232));
assign g8865 = ((~II15181));
assign g5809 = ((~II10460));
assign g7040 = (g6439)|(g5783);
assign gbuf40 = (g1159);
assign g9161 = ((~II15803));
assign g3018 = ((~II6770));
assign g5073 = ((~g4477));
assign g7525 = ((~II13755));
assign II5398 = ((~g702));
assign g5783 = (g1897&g5287);
assign g7559 = (g7367&g4155);
assign II13028 = ((~g7087));
assign g6873 = ((~II12490));
assign II8957 = ((~g1110))|((~II8955));
assign II10409 = ((~g5204));
assign g7272 = (g6182)|(g7038);
assign II15887 = ((~g9192))|((~g9191));
assign II10078 = ((~g4911))|((~g2256));
assign g8650 = (g591&g8094);
assign II10356 = ((~g5711));
assign g7503 = ((~II13686))|((~II13687));
assign g2308 = ((~II6081));
assign g4892 = ((~II9250));
assign g2837 = ((~g1780));
assign II15574 = ((~g8983));
assign g4652 = ((~II8871));
assign II9111 = ((~g4232));
assign g6146 = ((~II10801));
assign g8769 = (II14951)|(II14952);
assign II13891 = ((~g7336));
assign II7437 = ((~g2517))|((~II7436));
assign g2928 = ((~g2326));
assign g6026 = ((~g5384));
assign g5753 = ((~II10335))|((~II10336));
assign gbuf58 = (g94);
assign g4642 = ((~II8841));
assign II13144 = ((~g7031));
assign g6772 = ((~II12187));
assign II10289 = ((~g5569));
assign II9044 = (g4150)|(g4142)|(g4549);
assign g8811 = ((~g8443)&(~g8421)&(~II15075));
assign g5549 = (g2935)|(g4712);
assign II13537 = ((~g7152));
assign g4869 = ((~g4254))|((~g3533));
assign g3694 = ((~g2174));
assign g4648 = ((~II8859));
assign g3525 = ((~II7010))|((~II7011));
assign g7446 = ((~II13595));
assign g6235 = ((~II11034));
assign II14025 = ((~g7500));
assign g7550 = ((~II13834));
assign II12232 = ((~g6662));
assign g3819 = ((~g1748));
assign gbuf29 = (g1404);
assign II8974 = ((~g3871));
assign II11103 = ((~g2712))|((~II11101));
assign II13264 = ((~g7061));
assign II10017 = ((~g4700))|((~g2174));
assign g9359 = (g4748&g9340);
assign II7400 = ((~g3075));
assign II7421 = ((~g2525))|((~g2703));
assign II15175 = (g8483)|(g8464)|(g8514);
assign II16183 = ((~g9388));
assign II15675 = ((~g9058));
assign g5490 = ((~g4917));
assign g1649 = ((~g1217));
assign II11329 = ((~g5825));
assign g2674 = ((~g1675));
assign g4728 = (g190&g4179);
assign II10177 = ((~g4721));
assign g3614 = (g1134&g2386);
assign II12666 = ((~g6476));
assign g2480 = ((~g44));
assign g6882 = ((~II12517));
assign g9182 = ((~g9178));
assign g5235 = (g5091)|(g4422);
assign g6060 = (g1065&g5623);
assign g6990 = (g799&g6517);
assign g4027 = ((~g2845));
assign g7463 = ((~g7239));
assign II12433 = ((~g6632));
assign II13888 = ((~g7335));
assign g3798 = ((~g1757));
assign II7676 = ((~g2584));
assign II8417 = (g3430&g3398&g3359&g2106);
assign II7702 = ((~g3062));
assign g6612 = ((~II11832));
assign g5616 = ((~g4938));
assign II6775 = ((~g2386))|((~II6774));
assign II8028 = (g3430&g3398&g3359&g3341);
assign II7329 = ((~g2920));
assign g4153 = ((~II8024));
assign g1753 = (g819&g815);
assign gbuf22 = (g1270);
assign g4121 = ((~II7970));
assign g6762 = (g5847&g5412);
assign g4242 = ((~II8161));
assign g5469 = ((~g4898));
assign g9356 = (g9277)|(g9346);
assign g1974 = ((~g803));
assign g1748 = ((~g601));
assign g8961 = (g8885&g5317);
assign g1778 = ((~g613));
assign g7267 = ((~II13241));
assign g4969 = (g4362&g2216);
assign II6251 = ((~g489));
assign II12903 = ((~g6905));
assign II13940 = ((~g7355));
assign g6502 = ((~II11672));
assign g8733 = (g2996&g8493);
assign g5000 = ((~II9325));
assign g8624 = (g754&g8199);
assign II10907 = ((~g5492))|((~II10906));
assign g9018 = ((~II15478));
assign g3843 = ((~II7332));
assign g4359 = ((~II8327))|((~II8328));
assign g3866 = ((~g2945));
assign g5542 = ((~g5061));
assign g5761 = ((~II10356));
assign II11090 = ((~g1000));
assign g3899 = ((~II7479))|((~II7480));
assign g9291 = (g9273)|(g6216);
assign II10949 = ((~g5513));
assign g4235 = ((~g1415))|((~g2668));
assign g4350 = ((~II8315));
assign g4822 = ((~II9177));
assign g6194 = ((~II10937));
assign II6587 = ((~g1708));
assign II11371 = ((~g5840));
assign g9085 = ((~II15645));
assign g4867 = ((~II9209));
assign g7355 = ((~II13481));
assign g2910 = ((~II6636));
assign II9974 = ((~g4676));
assign g8838 = (g504&g8585);
assign g8268 = (g4568&g7905);
assign g8933 = (g4511&g8765);
assign g4908 = ((~g4088));
assign II11824 = ((~g6283));
assign II15053 = (g7951)|(g7920)|(g7983)|(g8181);
assign II15065 = ((~g8636));
assign II6341 = ((~g1351));
assign II11707 = ((~g5988));
assign II6302 = ((~g1313));
assign II12176 = ((~g5939));
assign g6833 = ((~II12370));
assign g8705 = (g2798&g8421);
assign g6372 = ((~II11443));
assign II7956 = ((~g2810));
assign g6349 = ((~II11374));
assign g8731 = (g2743&g8421);
assign g8746 = ((~g8524));
assign g6369 = ((~II11434));
assign g5760 = ((~II10353));
assign g5254 = (g5117)|(g4452);
assign II11464 = ((~g6088));
assign g8886 = (g8727)|(g8812)|(II15254);
assign g2976 = ((~II6728));
assign II15770 = ((~g9121));
assign g2149 = ((~II5894));
assign II12953 = ((~g1467))|((~II12951));
assign g7590 = ((~II13915));
assign II8949 = ((~g4116));
assign II10403 = ((~g5202));
assign II11446 = ((~g6062));
assign II6348 = ((~g1354));
assign g5471 = ((~II9889));
assign II15029 = (g8131)|(g8111)|(g8042)|(g8156);
assign g8218 = ((~II14433));
assign g8987 = (g8927)|(g8826);
assign II15273 = (g8287)|(g8334)|(g8295)|(g8339);
assign g9016 = (g8904&g8239);
assign g5596 = ((~g4841));
assign g6950 = ((~II12659));
assign g5564 = ((~II10018))|((~II10019));
assign g4529 = (II8612&II8613);
assign g5401 = ((~II9845));
assign g1771 = ((~g609));
assign II10038 = ((~g4893))|((~g2202));
assign g6978 = ((~II12717));
assign g1806 = ((~II5670));
assign II6906 = ((~g1838))|((~II6904));
assign g8696 = (g3743&g8342);
assign g6411 = (g5918&g5494);
assign g3634 = ((~II7107));
assign II6039 = ((~g207));
assign g2540 = ((~g1339));
assign g6393 = ((~II11506));
assign II14166 = ((~g7702));
assign II14406 = ((~g7681));
assign g3012 = ((~II6758))|((~II6759));
assign II6564 = ((~g2073));
assign g3801 = ((~II7262));
assign g9346 = (g9331&g6222);
assign g3910 = ((~II7523));
assign II14819 = ((~g8647));
assign g7292 = ((~II13308));
assign II8871 = ((~g3869));
assign g2841 = ((~g2208));
assign g6626 = ((~II11870));
assign II5506 = ((~g1532))|((~II5505));
assign g4224 = (g2680&g2683&II8127);
assign II13547 = ((~g1170));
assign II14187 = ((~g7728));
assign g6138 = (g5438)|(g5442);
assign g7827 = (g7575&g7173);
assign g6721 = ((~g6257));
assign g6813 = ((~II12310));
assign g5555 = ((~II9979))|((~II9980));
assign II8151 = ((~g3229))|((~II8150));
assign II10328 = ((~g5467))|((~II10327));
assign II8058 = (g2074&g2057&g2020&g1987);
assign g3856 = ((~II7371));
assign II15032 = (g8363)|(g8342)|(g8407)|(g8386);
assign g4927 = (g4318)|(g1590);
assign g6905 = ((~II12586));
assign g2245 = ((~g999));
assign II12885 = ((~g6946));
assign g3219 = ((~II6872));
assign g6671 = ((~II11971));
assign g2948 = ((~g2366));
assign II15947 = ((~g9221));
assign II6371 = ((~g33));
assign g1863 = ((~g68));
assign II8520 = ((~g3652));
assign II8109 = (g2074&g3287&g3264&g3238);
assign g6344 = ((~II11359));
assign II11672 = ((~g5971));
assign II11177 = ((~g5466))|((~g3019));
assign g9050 = ((~II15550));
assign g7025 = (g6541)|(g3095);
assign g5798 = ((~II10433));
assign II14394 = ((~g7536));
assign g6953 = ((~g6745));
assign g6390 = ((~II11497));
assign II10675 = ((~g5662));
assign II9153 = ((~g1649))|((~II9151));
assign II11040 = ((~g5299));
assign g6586 = ((~II11778));
assign II6460 = ((~g2104));
assign g7106 = ((~II12906));
assign II7967 = ((~g2787));
assign II9651 = ((~g4805));
assign g3998 = ((~g3097));
assign g5188 = (g5008)|(g4365);
assign II13731 = ((~g7441));
assign g4886 = ((~g4071));
assign g5154 = ((~II9588));
assign g8039 = ((~g7696));
assign g8229 = (g8180&g5680);
assign II12349 = ((~g6742));
assign II14839 = ((~g1073))|((~II14837));
assign II13016 = ((~g6941))|((~g1142));
assign g2700 = ((~g1744));
assign g4124 = (g2641&g2640);
assign II8097 = ((~g3237));
assign II10687 = ((~g5674));
assign g6090 = ((~g5529));
assign II15864 = ((~g9171))|((~II15862));
assign II10819 = ((~g5567))|((~II10818));
assign II10093 = ((~g4881))|((~II10092));
assign g6331 = ((~II11320));
assign g1738 = ((~g741));
assign g3975 = ((~g3131));
assign g6104 = ((~g5345));
assign g7605 = (g7435&g5607);
assign g4710 = ((~II9009));
assign g6999 = (g815&g6556);
assign II9372 = ((~g3902));
assign g7416 = (g7140&g4969);
assign II12015 = ((~g5874))|((~g5847));
assign g4361 = (g471&g3192);
assign II5897 = ((~g173));
assign g6328 = ((~II11311));
assign II5555 = ((~g1288));
assign II11933 = ((~g5847));
assign II11209 = ((~g6139));
assign g6053 = (g1053&g5608);
assign g2885 = ((~g2239));
assign g6606 = ((~II11824));
assign g9195 = ((~II15871));
assign g7209 = ((~g1789)&(~g146)&(~g6984));
assign g6043 = (g1069&g5582);
assign II15184 = ((~g8684));
assign g7299 = ((~II13329));
assign g7350 = ((~II13466));
assign g5665 = ((~g4748));
assign g8907 = (g8081)|(g8064)|(g8707);
assign g4612 = ((~II8751));
assign g2381 = ((~II6245));
assign g7262 = ((~II13228));
assign g2458 = ((~g30));
assign II6157 = ((~g246));
assign II15965 = ((~g9219));
assign g7693 = (g7367&g4445);
assign g6725 = ((~II12091));
assign II10855 = ((~g5521))|((~II10854));
assign g4300 = ((~II8261));
assign g6220 = ((~II11001));
assign II5879 = ((~g1267));
assign g5718 = ((~g4841));
assign II6333 = ((~g1345));
assign II7129 = ((~g2495));
assign II5889 = ((~g83));
assign g9189 = ((~II15845));
assign g8360 = ((~g7658)&(~g7616)&(~g8082)&(~g7634));
assign g8956 = ((~II15382));
assign g5181 = ((~II9669));
assign g5317 = (g4727)|(g4737)|(g4735);
assign II13244 = ((~g7033));
assign g8672 = ((~II14810));
assign g6428 = (g5874&g5494);
assign g4938 = ((~II9310));
assign II13722 = ((~g7442));
assign g2361 = ((~II6183));
assign II7762 = ((~g3029));
assign II12016 = ((~g5874))|((~II12015));
assign g8262 = (g4554&g7855);
assign g2162 = ((~II5901));
assign g6354 = ((~II11389));
assign g7542 = ((~II13810));
assign II12370 = ((~g6758));
assign g6072 = ((~g5345));
assign g2637 = ((~g1581));
assign II5475 = ((~g1084));
assign g6509 = ((~II11689));
assign II5966 = ((~g278));
assign II7188 = ((~g1834))|((~II7186));
assign II7029 = ((~g2392));
assign g6643 = (g1860&g5868);
assign g2829 = ((~g1785));
assign g5470 = ((~g4899));
assign II5894 = ((~g86));
assign g7516 = ((~II13728));
assign II7533 = ((~g3787))|((~II7531));
assign g7760 = ((~II14151));
assign g6757 = (g5874&g5412);
assign II10335 = ((~g5462))|((~II10334));
assign g4049 = (g141&g3514);
assign g2770 = ((~g2210));
assign g4782 = (g4187&g1760);
assign II14834 = (g8483)|(g8464)|(g8514);
assign g4629 = ((~II8802));
assign g4273 = ((~II8215));
assign g4587 = ((~g2928));
assign g9260 = ((~II15990));
assign g7597 = (g7316&g4841);
assign II10253 = ((~g5240));
assign g5707 = (g4956)|(g4343);
assign II10552 = ((~g5396));
assign II11662 = ((~g5956));
assign g4166 = (II8045&II8046);
assign II15003 = ((~g8633));
assign II7644 = ((~g2584));
assign II9407 = ((~g4232));
assign g6922 = ((~g6525));
assign g5494 = ((~II9918));
assign g5938 = ((~g5412));
assign g8725 = (g3008&g8493);
assign g5215 = (g5050)|(g4390);
assign g7028 = ((~g6525));
assign g6284 = ((~II11164))|((~II11165));
assign II15568 = ((~g8981));
assign g6805 = ((~II12286));
assign II9064 = ((~g4302));
assign II7781 = ((~g2605));
assign II11569 = ((~g6279));
assign g7257 = ((~II13214))|((~II13215));
assign g5088 = ((~II9466));
assign g4033 = ((~g3192));
assign g1926 = ((~g874));
assign g6270 = (g1000)|(g5335)|(g1909);
assign g7414 = ((~II13527));
assign g5828 = ((~II10509));
assign II10516 = ((~g5241));
assign g1865 = ((~g1013));
assign II15971 = ((~g9233));
assign II5435 = ((~g1461));
assign II7150 = ((~g1974))|((~II7148));
assign II8209 = (g2298&g2316&g2334);
assign g4438 = ((~II8446));
assign II8120 = ((~g1904))|((~II8119));
assign g2522 = ((~g1342));
assign g1944 = ((~II5817));
assign II15940 = ((~g9213));
assign II12906 = ((~g6918));
assign II6042 = ((~g237));
assign g7774 = ((~II14193));
assign II9416 = ((~g4273));
assign II15819 = ((~g9148))|((~II15817));
assign g8070 = (g863&g7616);
assign II14224 = ((~g7722));
assign II6776 = ((~g1134))|((~II6774));
assign g5756 = ((~II10343));
assign g3925 = ((~II7575))|((~II7576));
assign g2605 = ((~g1639));
assign g7122 = ((~II12958));
assign g6997 = ((~II12737));
assign g2396 = ((~g1033));
assign g7061 = ((~g6650));
assign II5772 = ((~g1240));
assign II7769 = ((~g3038));
assign g8404 = (g710&g7937);
assign II12708 = ((~g6482));
assign g6320 = ((~II11287));
assign II14614 = ((~g7832));
assign g9241 = ((~II15971));
assign g9221 = ((~II15937));
assign g4620 = ((~II8775));
assign II9050 = ((~g3881));
assign II14445 = ((~g8067));
assign g9097 = ((~II15681));
assign g8870 = ((~II15196));
assign II11473 = ((~g6069));
assign g8920 = (g4578&g8746);
assign g6388 = ((~II11491));
assign II8778 = ((~g3922));
assign g6404 = ((~II11525));
assign II15848 = ((~g9162))|((~g9154));
assign g7716 = ((~II14025));
assign g1818 = ((~II5692));
assign g7196 = ((~II13122));
assign g8841 = (g351&g8545);
assign g8848 = (g281&g8524);
assign g6581 = ((~II11773));
assign g7491 = ((~II13653));
assign g9144 = (g9123&g6096);
assign II14067 = ((~g7550));
assign g3919 = ((~II7554));
assign g2266 = ((~II6003));
assign II6133 = ((~g846))|((~g916));
assign g8684 = ((~II14848));
assign g8062 = (g7476&g7634);
assign g6719 = (g6166)|(g6171);
assign g4557 = ((~g2896));
assign II10745 = ((~g2100))|((~II10743));
assign g3952 = ((~II7651));
assign g7245 = ((~II13193));
assign g3739 = ((~g2536));
assign II15654 = ((~g9057));
assign g2661 = ((~II6454));
assign g7278 = (g6965&g1745);
assign II8925 = ((~g4482));
assign g4398 = (g567&g2845);
assign g8991 = (g8931)|(g8831);
assign g2074 = ((~II5872));
assign g6375 = ((~II11452));
assign g4381 = ((~g3466));
assign g7838 = ((~II14264));
assign g1792 = ((~g616));
assign g7533 = ((~II13779));
assign g6929 = (g6412)|(g6418);
assign II15527 = ((~g9020));
assign II13284 = ((~g7156));
assign II10810 = ((~g5403));
assign II14942 = (g8439)|(g8440)|(g8405)|(g8460);
assign g8457 = (g724&g7811);
assign II11302 = ((~g5796));
assign g6845 = ((~II12406));
assign gbuf70 = (g891);
assign g6202 = ((~II10949));
assign g2630 = ((~g1575));
assign g4199 = (g93&g2769);
assign g8481 = ((~II14637));
assign II7380 = ((~g3461));
assign g4112 = ((~II7947));
assign II14767 = (g7937)|(g7887)|(g8029)|(g8018);
assign II6517 = ((~g1687));
assign II5695 = ((~g1513))|((~g1524));
assign II6223 = ((~g330));
assign II11308 = ((~g5759));
assign g4182 = (II8071&II8072);
assign II15959 = ((~g9217));
assign g7498 = ((~II13672));
assign g6119 = ((~II10744))|((~II10745));
assign g4069 = ((~II7844));
assign g2938 = ((~g2347));
assign II10848 = ((~g5490))|((~II10847));
assign g1714 = (g1454&g1450);
assign g1844 = (g792&g795);
assign g6129 = ((~II10758));
assign g6610 = (g4180)|(g6061);
assign g7181 = (g6124&g7039);
assign g3979 = ((~II7702));
assign g9335 = (g9320&g6206);
assign g4000 = ((~g3131));
assign II8994 = ((~g4565));
assign g5194 = (g5018)|(g4367);
assign g8687 = (g3488&g8363);
assign g2783 = ((~II6523))|((~II6524));
assign II8718 = ((~g3909));
assign g6819 = ((~II12328));
assign g3062 = ((~g2100));
assign g2638 = ((~g1582));
assign g8307 = (g432&g7920);
assign g7759 = ((~II14148));
assign II10225 = ((~g4895))|((~II10223));
assign g4680 = ((~II8945));
assign II15075 = (II15071)|(II15072)|(II15073)|(II15074);
assign II5751 = ((~g963));
assign g9389 = ((~II16183));
assign g6360 = ((~II11407));
assign II13927 = ((~g7366));
assign g5024 = ((~II9360));
assign g8968 = ((~II15408));
assign g7179 = (g6121&g7035);
assign II7691 = ((~g3651));
assign II9457 = ((~g3940));
assign II14771 = (g7993)|(g7966)|(g7793)|(g7811);
assign g5367 = ((~II9834));
assign g8947 = (g4558&g8787);
assign II9261 = (g3777&g3764&g3746);
assign II15014 = ((~g8607));
assign g3774 = ((~g1770));
assign g8919 = (g4567&g8743);
assign g7089 = (g4128)|(g6474);
endmodule
