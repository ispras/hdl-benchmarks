//NOTE: no-implementation module stub

module ejtag_setclr (
    output wire SETQ,
    output wire CLRQ,
    input wire SET,
    input wire CLR,
    input wire SETCLK,
    input wire SETRST_N,
    input wire CLRCLK,
    input wire CLRRST_N
);

endmodule
