//NOTE: no-implementation module stub

module obj_q (
    input wire DATA14,
    input wire DATA13,
    input wire CLKSOURCE1,
    input wire VXI2C,
    input wire VXI2D,
    input wire VXI2E,
    input wire DATA12,
    input wire CLKSOURCE0,
    input wire DATA15,
    input wire [15:0] DATA0,
    input wire [15:0] DATA1,
    input wire [15:0] DATA2,
    input wire [15:0] DATA3,
    input wire [15:0] DATA4,
    input wire [15:0] DATA5,
    input wire [15:0] DATA6,
    input wire [15:0] DATA7,
    inout wire [31:0] DATA08,
    inout wire [7:0] WEC1,
    input wire [5:1] DATA10,
    output wire DATA29,
    output wire DATA19,
    output wire DATA24,
    output wire DATA20,
    output wire WEC2,
    output wire WEC3,
    output wire WEC8,
    output wire WEC6,
    output wire WEC7,
    output wire DATA18,
    output wire [3:0] WEC4,
    output wire [7:0] WEC5,
    output wire [31:0] vxi2a,
    output wire [31:0] vxi2b,
    output wire [19:0] pr4
);

endmodule
