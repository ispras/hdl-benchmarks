//NOTE: no-implementation module stub

module lmi_iram (
    input wire CLK,
    input wire TMODE,
    input wire RESET_D1_R_N,
    input wire INVALIDATE,
    input wire MEMSEQUENTIAL,
    input wire MEMZEROFIRST,
    input wire CFG_IRAMISROM,
    input wire EXT_IWREQRAM_R,
    input wire IW_GNTRAM_R,
    output wire IW_DATAOE,
    output wire IW_LBCOE,
    input wire NEXTADDR,
    input wire RDOP_N,
    output wire IS_VAL,
    output wire IW_VAL,
    output wire X_HALT_R,
    output wire IW_ACK,
    output wire IW_MISS_R,
    output wire IW_MISS_P,
    output wire IW_HALT_S_R,
    input wire IW_VALINDEX,
    input wire IWR_VALRD,
    input wire IW_VALWR,
    input wire IW_VALWE,
    input wire IW_VALWEN,
    input wire IW_VALRE,
    input wire IW_VALREN,
    input wire IW_VALCS,
    input wire IW_VALCSN,
    input wire IW_DATAINDEX,
    input wire IW_DATAWE,
    input wire IW_DATAWEN,
    input wire IW_DATARE,
    input wire IW_DATAREN,
    input wire IW_DATACS,
    input wire IW_DATACSN,
    input wire CONFIGBASE,
    input wire CONFIGTOP
);

endmodule
