//NOTE: no-implementation module stub

module MAbufx (
    input [13:0] CMAin,
    output [13:0] CMAinx
);

endmodule
