module Mod_7 ( constr__0___3__constr_inst1851__0___3__cp_sub_out , impl__0___0__I_546__0___0__o
 , constr__0___0__wp_test__0__in2[7:0]  , constr__0___0__wp_test__0__in1[7:0] 
 , constr__0___0__wp_test__0__in4[7:0]  , constr__0___0__wp_test__0__in3[7:0] ,
himanshu_clock	
 ) ;
 input himanshu_clock;
 output  [7:0]  constr__0___3__constr_inst1851__0___3__cp_sub_out ;
 output  [7:0]  impl__0___0__I_546__0___0__o ;
 input    [7:0]  constr__0___0__wp_test__0__in2  ;
 input    [7:0]  constr__0___0__wp_test__0__in1  ;
 input    [7:0]  constr__0___0__wp_test__0__in4  ;
 input    [7:0]  constr__0___0__wp_test__0__in3  ;
 wire  [7:0] impl__0___0__r71672__0___0 ;
 wire  [11:0] impl__0___0__r7__0___0 ;
 wire  [11:0] impl__0___0__E_13481704__0___0 ;
 wire    [6:0] impl__0___0__E_1348__0___0 ;
 wire  [0:0] E_1878__0___0 ;
 wire    [5:0] impl__0___0__r1__0___0 ;
 wire  [5:0] impl__0___0__in21663__0___0 ;
 wire  [7:0] constr__0___0__constr_inst1861__0___0__ce1821__3___0 ;
 wire    [7:0] constr__0___0__ce_test__0__in2__0___0  ;
assign constr__0___0__ce_test__0__in2__0___0  = constr__0___0__wp_test__0__in2[7:0]  ;
 wire  [5:0] impl__0___0__in11662__0___0 ;
 wire  [7:0] spec__0___0__E_68__0___0 ;
 wire    [7:0] constr__0___0__ce_test__0__in1__0___0  ;
assign constr__0___0__ce_test__0__in1__0___0  = constr__0___0__wp_test__0__in1[7:0]  ;
 wire  [11:0] impl__0___0__E_13471703__0___0 ;
 wire  [9:0] impl__0___0__E_1347__0___0 ;
 wire  [1:0] E_1876__0___0 ;
 wire  [11:0] impl__0___0__E_13281701__0___0 ;
 wire    [10:0] impl__0___0__r6__0___0 ;
 wire    [10:0] impl__0___0__r6_inp13601774__0___0 ;
 wire  [10:0] impl__0___0__r6_inp1360__0___0 ;
 wire  [10:0] impl__0___0__E_13691717__0___0 ;
 wire    [7:0] impl__0___0__r3__0___0 ;
 wire  [7:0] impl__0___0__E_1411__0___0 ;
 wire  [7:0] constr__0___0__constr_inst1857__0___0__ce1821__5___0 ;
 wire    [7:0] constr__0___0__ce_test__0__in4__0___0  ;
assign constr__0___0__ce_test__0__in4__0___0  = constr__0___0__wp_test__0__in4[7:0]  ;
 wire    [6:0] impl__0___0__r2__0___0 ;
 wire  [6:0] impl__0___0__in31664__0___0 ;
 wire  [7:0] constr__0___0__constr_inst1859__0___0__ce1821__4___0 ;
 wire    [7:0] constr__0___0__ce_test__0__in3__0___0  ;
assign constr__0___0__ce_test__0__in3__0___0  = constr__0___0__wp_test__0__in3[7:0]  ;
 wire  [6:0] impl__0___0__E_141016791729__0___0 ;
 wire  [7:0] impl__0___0__E_13891719__0___0 ;
 wire  [10:0] impl__0___0__E_13681716__0___0 ;
 wire    [10:0] impl__0___0__r613431773__0___0 ;
 wire    [6:0] impl__0___0__r61343__0___0 ;
 wire impl__0___0__r6_inp__0___0 ;
 wire  [7:0] impl__0___0__E_1362__0___0 ;
 wire  [7:0] impl__0___0__eq_s_s_9eq_s_s_9_output1720__0___0  ;
 wire impl__0___0__eq_s_s_9eq_s_s_9_output__0___0  ;
 wire  [8:0] impl__0___0__E_1413__0___0 ;
 wire impl__0___0__E_1421__0___0 ;
 wire  [0:0] impl__0___0__mul_s_s_9t1_inp1722__0___0  ;
 wire  [0:0] E_1879__0___0 ;
 wire  [0:8] impl__0___0__mul_s_s_9in0_inp__0___0  ;
 wire  [7:0] impl__0___0__mul_s_s_9in0_inp1681__0___0  ;
 wire  [8:0] impl__0___0__E_1412__0___0 ;
 wire impl__0___0__E_1419__0___0 ;
 wire impl__0___0__E_1426__0___0 ;
 wire  [0:8] impl__0___0__r4__0___0 ;
 wire  [0:8] impl__0___0__mul_s_s_9mul_s_s_9_output__0___0  ;
 wire  [0:8] impl__0___0__mul_s_s_9mul_s_s_9_output_inp14331772__0___0  ;
 wire  [8:0] impl__0___0__mul_s_s_9mul_s_s_9_output_inp1433__0___0  ;
 wire  [0:8] impl__0___0__mul_s_s_9t3__0___0  ;
 wire    [2:8] impl__0___0__mul_s_s_9t2__0___0  ;
 wire    [2:8] impl__0___0__mul_s_s_9t2_inp14411771__0___0  ;
 wire    [6:0] impl__0___0__mul_s_s_9t2_inp1441__0___0  ;
 wire  [0:8] impl__0___0__mul_s_s_9in1_inp__0___0  ;
 wire    [2:8] impl__0___0__mul_s_s_9in1_inp1770__0___0  ;
 wire  [0:0] impl__0___0__mul_s_s_9t2_inp1723__0___0  ;
 wire  [0:8] impl__0___0__mul_s_s_9t1__0___0  ;
 wire  [0:8] impl__0___0__mul_s_s_9t1_inp14391769__0___0  ;
 wire  [8:0] impl__0___0__mul_s_s_9t1_inp1439__0___0  ;
 wire impl__0___0__mul_s_s_9mul_s_s_9_output_inp__0___0  ;
 wire  [7:0] impl__0___0__eq_s_s_9in0_inp1680__0___0  ;
 wire  [7:0] impl__0___0__E_1323__0___0 ;
 wire  [7:0] impl__0___0__E_13281666__0___0 ;
 wire  [7:0] impl__0___0__r5__0___0 ;
 wire  [7:0] impl__0___0__r5_inp__0___0 ;
 wire  [7:0] impl__0___0__E_13871718__0___0 ;
 wire  [7:0] impl__0___0__r5_inp1371__0___0 ;
 wire  [7:0] impl__0___0__r31653__0___0 ;
 wire  [7:0] constr__0___3__constr_inst1851__0___3__ce1824__3___3 ;
assign constr__0___3__constr_inst1851__0___3__cp_sub_out = constr__0___3__constr_inst1851__0___3__ce1824__3___3 ;
 wire  [7:0] constr__0___3__constr_inst1849__0___3__ce1821__7___3 ;
 wire    [7:0] spec__0___0__out2_inp__0___0 ;
 wire  [7:0] spec__0___0__r71779__0___0 ;
 wire  [8:0] spec__0___0__r7__0___0 ;
 wire  [8:0] spec__0___0__E_521789__0___0 ;
 wire    [6:0] spec__0___0__E_52__0___0 ;
 wire  [0:0] E_1881__0___0 ;
 wire    [5:0] spec__0___0__r1__0___0 ;
 wire  [5:0] spec__0___0__in21776__0___0 ;
 wire  [5:0] spec__0___0__in11775__0___0 ;
 wire  [8:0] spec__0___0__E_51__0___0 ;
 wire  [1:0] E_1880__0___0 ;
 wire  [10:0] spec__0___0__r6__0___0 ;
 wire  [10:0] spec__0___0__r6_inp60__0___0 ;
 wire  [10:0] spec__0___0__E_651791__0___0 ;
 wire    [7:0] spec__0___0__r3__0___0 ;
 wire  [7:0] spec__0___0__E_77__0___0 ;
 wire    [6:0] spec__0___0__r2__0___0 ;
 wire  [6:0] spec__0___0__in31777__0___0 ;
 wire  [6:0] spec__0___0__E_7617811802__0___0 ;
 wire  [7:0] spec__0___0__E_721796__0___0 ;
 wire  [10:0] spec__0___0__E_661793__0___0 ;
 wire  [10:0] spec__0___0__r6_inp61__0___0 ;
 wire spec__0___0__r6_inp__0___0 ;
 wire  [7:0] spec__0___0__E_62__0___0 ;
 wire  [7:0] spec__0___0__E_671794__0___0 ;
 wire spec__0___0__E_67__0___0 ;
 wire    [8:0] spec__0___0__r4__0___0 ;
 wire  [8:0] spec__0___0__E_78__0___0 ;
 wire  [7:0] spec__0___0__E_43__0___0 ;
 wire  [7:0] spec__0___0__r61780__0___0 ;
 wire  [7:0] spec__0___0__r5__0___0 ;
 wire  [7:0] spec__0___0__r5_inp__0___0 ;
 wire  [7:0] spec__0___0__E_701795__0___0 ;
 wire  [7:0] spec__0___0__r5_inp63__0___0 ;
  assign /* un  8-bit */  impl__0___0__I_546__0___0__o = impl__0___0__E_1323__0___0 & impl__0___0__r71672__0___0 ;
  assign /* un  8-bit */  impl__0___0__r71672__0___0 = impl__0___0__r7__0___0 ;
  assign /* un 12-bit */  impl__0___0__r7__0___0 = impl__0___0__E_13471703__0___0 | impl__0___0__E_13481704__0___0 ;
  assign /* un 12-bit */  impl__0___0__E_13481704__0___0 = impl__0___0__E_1348__0___0 ;
  assign /*     7-bit */  impl__0___0__E_1348__0___0 = impl__0___0__r1__0___0 << E_1878__0___0 ;
  assign /* un  1-bit */  E_1878__0___0 = 1'h1;
  assign /*     6-bit */  impl__0___0__r1__0___0 = impl__0___0__in11662__0___0 + impl__0___0__in21663__0___0 ;
  assign /* un  6-bit */  impl__0___0__in21663__0___0 = constr__0___0__constr_inst1861__0___0__ce1821__3___0 ;
  assign /* un  8-bit */  constr__0___0__constr_inst1861__0___0__ce1821__3___0 = constr__0___0__ce_test__0__in2__0___0  ;
  assign /* un  6-bit */  impl__0___0__in11662__0___0 = spec__0___0__E_68__0___0 ;
  assign /* un  8-bit */  spec__0___0__E_68__0___0 = constr__0___0__ce_test__0__in1__0___0  ;
  assign /* un 12-bit */  impl__0___0__E_13471703__0___0 = impl__0___0__E_1347__0___0 ;
  assign /* un 10-bit */  impl__0___0__E_1347__0___0 = impl__0___0__E_13281701__0___0 >> E_1876__0___0 ;
  assign /* un  2-bit */  E_1876__0___0 = 2'h2;
  assign /* un 12-bit */  impl__0___0__E_13281701__0___0 = impl__0___0__r6__0___0 ;
  assign /*    11-bit */  impl__0___0__r6__0___0 = impl__0___0__r6_inp__0___0 ? impl__0___0__r6_inp13601774__0___0 : impl__0___0__r613431773__0___0 ;
  assign /*    11-bit */  impl__0___0__r6_inp13601774__0___0 = impl__0___0__r6_inp1360__0___0 ;
  assign /* un 11-bit */  impl__0___0__r6_inp1360__0___0 = impl__0___0__E_13681716__0___0 | impl__0___0__E_13691717__0___0 ;
  assign /* un 11-bit */  impl__0___0__E_13691717__0___0 = impl__0___0__r3__0___0 ;
  assign /*     8-bit */  impl__0___0__r3__0___0 = impl__0___0__E_13891719__0___0 ^ impl__0___0__E_1411__0___0 ;
wire  [7:0]  impl__0___0__r2__0___01936 = impl__0___0__r2__0___0; /* sign-extend */ 
  assign /* un  8-bit */  impl__0___0__E_1411__0___0 = impl__0___0__r2__0___01936 - constr__0___0__constr_inst1857__0___0__ce1821__5___0 ;
  assign /* un  8-bit */  constr__0___0__constr_inst1857__0___0__ce1821__5___0 = constr__0___0__ce_test__0__in4__0___0  ;
  assign /*     7-bit */  impl__0___0__r2__0___0 = impl__0___0__E_141016791729__0___0 | impl__0___0__in31664__0___0 ;
  assign /* un  7-bit */  impl__0___0__in31664__0___0 = constr__0___0__constr_inst1859__0___0__ce1821__4___0 ;
  assign /* un  8-bit */  constr__0___0__constr_inst1859__0___0__ce1821__4___0 = constr__0___0__ce_test__0__in3__0___0  ;
  assign /* un  7-bit */  impl__0___0__E_141016791729__0___0 = impl__0___0__r1__0___0 ;
  assign /* un  8-bit */  impl__0___0__E_13891719__0___0 = impl__0___0__r1__0___0 ;
  assign /* un 11-bit */  impl__0___0__E_13681716__0___0 = impl__0___0__r2__0___0 ;
  assign /*    11-bit */  impl__0___0__r613431773__0___0 = impl__0___0__r61343__0___0 ;
  assign /*     7-bit */  impl__0___0__r61343__0___0 = ~impl__0___0__r2__0___0 ;
  assign /* un    bit */  impl__0___0__r6_inp__0___0 = |impl__0___0__E_1362__0___0 ;
  assign /* un  8-bit */  impl__0___0__E_1362__0___0 = impl__0___0__eq_s_s_9eq_s_s_9_output1720__0___0  | spec__0___0__E_68__0___0 ;
  assign /* un  8-bit */  impl__0___0__eq_s_s_9eq_s_s_9_output1720__0___0  = impl__0___0__eq_s_s_9eq_s_s_9_output__0___0  ;
  assign /* un    bit */  impl__0___0__eq_s_s_9eq_s_s_9_output__0___0  = impl__0___0__E_1412__0___0 == impl__0___0__E_1413__0___0 ;
  assign /* un  9-bit */  impl__0___0__E_1413__0___0 = { impl__0___0__E_1421__0___0 , impl__0___0__mul_s_s_9in0_inp1681__0___0  };
  assign /* un    bit */  impl__0___0__E_1421__0___0 = ~impl__0___0__mul_s_s_9t1_inp1722__0___0  ;
  assign /* un  1-bit */  impl__0___0__mul_s_s_9t1_inp1722__0___0  = impl__0___0__mul_s_s_9in0_inp__0___0  [ 1'h0 : 1'h0 ] ; 
  assign /* un  1-bit */  E_1879__0___0 = 1'h0;
  assign /* un  9-bit */  impl__0___0__mul_s_s_9in0_inp__0___0  = impl__0___0__r3__0___0 ;
  assign /* un  8-bit */  impl__0___0__mul_s_s_9in0_inp1681__0___0  = impl__0___0__mul_s_s_9in0_inp__0___0  ;
  assign /* un  9-bit */  impl__0___0__E_1412__0___0 = { impl__0___0__E_1419__0___0 , impl__0___0__eq_s_s_9in0_inp1680__0___0  };
  assign /* un    bit */  impl__0___0__E_1419__0___0 = ~impl__0___0__E_1426__0___0 ;
  assign /* un    bit */  impl__0___0__E_1426__0___0 = impl__0___0__r4__0___0 [ 1'h0 : 1'h0 ] ; 
wire  [8:0]  impl__0___0__r2__0___01937 = impl__0___0__r2__0___0; /* sign-extend */ 
  assign /* un  9-bit */  impl__0___0__r4__0___0 = impl__0___0__mul_s_s_9mul_s_s_9_output__0___0  + impl__0___0__r2__0___01937 ;
  assign /* un  9-bit */  impl__0___0__mul_s_s_9mul_s_s_9_output__0___0  = impl__0___0__mul_s_s_9mul_s_s_9_output_inp__0___0  ? impl__0___0__mul_s_s_9mul_s_s_9_output_inp14331772__0___0  : impl__0___0__mul_s_s_9t3__0___0  ;
  assign /* un  9-bit */  impl__0___0__mul_s_s_9mul_s_s_9_output_inp14331772__0___0  = impl__0___0__mul_s_s_9mul_s_s_9_output_inp1433__0___0  ;
  assign /* un  9-bit */  impl__0___0__mul_s_s_9mul_s_s_9_output_inp1433__0___0  = -impl__0___0__mul_s_s_9t3__0___0  ;
wire  [8:0]  impl__0___0__mul_s_s_9t2__0___01938  = impl__0___0__mul_s_s_9t2__0___0 ; /* sign-extend */ 
  assign /* un  9-bit */  impl__0___0__mul_s_s_9t3__0___0  = impl__0___0__mul_s_s_9t1__0___0  * impl__0___0__mul_s_s_9t2__0___01938  ;
  assign /*     7-bit */  impl__0___0__mul_s_s_9t2__0___0  = impl__0___0__mul_s_s_9t2_inp1723__0___0  ? impl__0___0__mul_s_s_9t2_inp14411771__0___0  : impl__0___0__mul_s_s_9in1_inp1770__0___0  ;
  assign /*     7-bit */  impl__0___0__mul_s_s_9t2_inp14411771__0___0  = impl__0___0__mul_s_s_9t2_inp1441__0___0  ;
  assign /*     7-bit */  impl__0___0__mul_s_s_9t2_inp1441__0___0  = -impl__0___0__mul_s_s_9in1_inp__0___0  ;
  assign /* un  9-bit */  impl__0___0__mul_s_s_9in1_inp__0___0  = impl__0___0__r1__0___0 ;
  assign /*     7-bit */  impl__0___0__mul_s_s_9in1_inp1770__0___0  = impl__0___0__mul_s_s_9in1_inp__0___0  ;
  assign /* un  1-bit */  impl__0___0__mul_s_s_9t2_inp1723__0___0  = impl__0___0__mul_s_s_9in1_inp__0___0  [ 1'h0 : 1'h0 ] ; 
  assign /* un  9-bit */  impl__0___0__mul_s_s_9t1__0___0  = impl__0___0__mul_s_s_9t1_inp1722__0___0  ? impl__0___0__mul_s_s_9t1_inp14391769__0___0  : impl__0___0__mul_s_s_9in0_inp__0___0  ;
  assign /* un  9-bit */  impl__0___0__mul_s_s_9t1_inp14391769__0___0  = impl__0___0__mul_s_s_9t1_inp1439__0___0  ;
  assign /* un  9-bit */  impl__0___0__mul_s_s_9t1_inp1439__0___0  = -impl__0___0__mul_s_s_9in0_inp__0___0  ;
  assign /* un    bit */  impl__0___0__mul_s_s_9mul_s_s_9_output_inp__0___0  = impl__0___0__mul_s_s_9t1_inp1722__0___0  ^ impl__0___0__mul_s_s_9t2_inp1723__0___0  ;
  assign /* un  8-bit */  impl__0___0__eq_s_s_9in0_inp1680__0___0  = impl__0___0__r4__0___0 ;
  assign /* un  8-bit */  impl__0___0__E_1323__0___0 = impl__0___0__r5__0___0 + impl__0___0__E_13281666__0___0 ;
  assign /* un  8-bit */  impl__0___0__E_13281666__0___0 = impl__0___0__r6__0___0 ;
  assign /* un  8-bit */  impl__0___0__r5__0___0 = impl__0___0__r6_inp__0___0 ? impl__0___0__r5_inp__0___0 : impl__0___0__r5_inp1371__0___0 ;
  assign /* un  8-bit */  impl__0___0__r5_inp__0___0 = impl__0___0__E_13891719__0___0 ^ impl__0___0__E_13871718__0___0 ;
  assign /* un  8-bit */  impl__0___0__E_13871718__0___0 = impl__0___0__r2__0___0 ;
wire  [7:0]  impl__0___0__r1__0___01939 = impl__0___0__r1__0___0; /* sign-extend */ 
  assign /* un  8-bit */  impl__0___0__r5_inp1371__0___0 = impl__0___0__r31653__0___0 + impl__0___0__r1__0___01939 ;
  assign /* un  8-bit */  impl__0___0__r31653__0___0 = impl__0___0__r3__0___0 ;
  assign /* un  8-bit */  constr__0___3__constr_inst1851__0___3__ce1824__3___3 = constr__0___3__constr_inst1849__0___3__ce1821__7___3 ;
  assign /* un  8-bit */  constr__0___3__constr_inst1849__0___3__ce1821__7___3 = spec__0___0__out2_inp__0___0 ;
  assign /*     8-bit */  spec__0___0__out2_inp__0___0 = spec__0___0__E_43__0___0 & spec__0___0__r71779__0___0 ;
  assign /* un  8-bit */  spec__0___0__r71779__0___0 = spec__0___0__r7__0___0 ;
  assign /* un  9-bit */  spec__0___0__r7__0___0 = spec__0___0__E_51__0___0 | spec__0___0__E_521789__0___0 ;
  assign /* un  9-bit */  spec__0___0__E_521789__0___0 = spec__0___0__E_52__0___0 ;
  assign /*     7-bit */  spec__0___0__E_52__0___0 = spec__0___0__r1__0___0 <<< E_1881__0___0 ;
  assign /* un  1-bit */  E_1881__0___0 = 1'h1;
  assign /*     6-bit */  spec__0___0__r1__0___0 = spec__0___0__in11775__0___0 + spec__0___0__in21776__0___0 ;
  assign /* un  6-bit */  spec__0___0__in21776__0___0 = constr__0___0__ce_test__0__in2__0___0  ;
  assign /* un  6-bit */  spec__0___0__in11775__0___0 = constr__0___0__ce_test__0__in1__0___0  ;
  assign /* un  9-bit */  spec__0___0__E_51__0___0 = spec__0___0__r6__0___0 >> E_1880__0___0 ;
  assign /* un  2-bit */  E_1880__0___0 = 2'h2;
  assign /* un 11-bit */  spec__0___0__r6__0___0 = spec__0___0__r6_inp__0___0 ? spec__0___0__r6_inp60__0___0 : spec__0___0__r6_inp61__0___0 ;
  assign /* un 11-bit */  spec__0___0__r6_inp60__0___0 = spec__0___0__E_661793__0___0 | spec__0___0__E_651791__0___0 ;
  assign /* un 11-bit */  spec__0___0__E_651791__0___0 = spec__0___0__r3__0___0 ;
  assign /*     8-bit */  spec__0___0__r3__0___0 = spec__0___0__E_721796__0___0 ^ spec__0___0__E_77__0___0 ;
  assign /* un  8-bit */  spec__0___0__E_77__0___0 = spec__0___0__r2__0___0 - constr__0___0__ce_test__0__in4__0___0  ;
  assign /*     7-bit */  spec__0___0__r2__0___0 = spec__0___0__E_7617811802__0___0 | spec__0___0__in31777__0___0 ;
  assign /* un  7-bit */  spec__0___0__in31777__0___0 = constr__0___0__ce_test__0__in3__0___0  ;
  assign /* un  7-bit */  spec__0___0__E_7617811802__0___0 = spec__0___0__r1__0___0 ;
  assign /* un  8-bit */  spec__0___0__E_721796__0___0 = spec__0___0__r1__0___0 ;
  assign /* un 11-bit */  spec__0___0__E_661793__0___0 = spec__0___0__r2__0___0 ;
  assign /* un 11-bit */  spec__0___0__r6_inp61__0___0 = ~spec__0___0__E_661793__0___0 ;
  assign /* un    bit */  spec__0___0__r6_inp__0___0 = |spec__0___0__E_62__0___0 ;
  assign /* un  8-bit */  spec__0___0__E_62__0___0 = spec__0___0__E_671794__0___0 | spec__0___0__E_68__0___0 ;
  assign /* un  8-bit */  spec__0___0__E_671794__0___0 = spec__0___0__E_67__0___0 ;
  assign /* un    bit */  spec__0___0__E_67__0___0 = spec__0___0__r4__0___0 == spec__0___0__r3__0___0 ;
wire  [8:0]  spec__0___0__r2__0___01940 = spec__0___0__r2__0___0; /* sign-extend */ 
  assign /*     9-bit */  spec__0___0__r4__0___0 = spec__0___0__E_78__0___0 + spec__0___0__r2__0___01940 ;
  assign /* un  9-bit */  spec__0___0__E_78__0___0 = spec__0___0__r3__0___0 * spec__0___0__r1__0___0 ;
  assign /* un  8-bit */  spec__0___0__E_43__0___0 = spec__0___0__r5__0___0 + spec__0___0__r61780__0___0 ;
  assign /* un  8-bit */  spec__0___0__r61780__0___0 = spec__0___0__r6__0___0 ;
  assign /* un  8-bit */  spec__0___0__r5__0___0 = spec__0___0__r6_inp__0___0 ? spec__0___0__r5_inp__0___0 : spec__0___0__r5_inp63__0___0 ;
  assign /* un  8-bit */  spec__0___0__r5_inp__0___0 = spec__0___0__E_721796__0___0 ^ spec__0___0__E_701795__0___0 ;
  assign /* un  8-bit */  spec__0___0__E_701795__0___0 = spec__0___0__r2__0___0 ;
  assign /* un  8-bit */  spec__0___0__r5_inp63__0___0 = spec__0___0__r3__0___0 + spec__0___0__r1__0___0 ;
endmodule

