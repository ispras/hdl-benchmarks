//NOTE: no-implementation module stub

module GTECH_NOR3 (
    input wire A,
    input wire B,
    input wire C,
    output wire Z
);

endmodule
