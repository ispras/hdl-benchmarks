module top ( g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 , g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 );
input g0 , g1 , g2 , g3 , g4 , g5 , g6 , g7 , g8 , g9 , g10 , g11 , g12 , g13 , g14 , g15 , g16 , g17 , g18 , g19 , g20 , g21 , g22 , g23 , g24 , g25 , g26 , g27 , g28 , g29 , g30 , g31 , g32 , g33 , g34 , g35 , g36 , g37 , g38 , g39 , g40 , g41 , g42 , g43 , g44 , g45 , g46 , g47 , g48 , g49 , g50 , g51 , g52 , g53 , g54 , g55 , g56 , g57 , g58 , g59 , g60 , g61 , g62 , g63 , g64 , g65 , g66 , g67 , g68 , g69 , g70 , g71 , g72 , g73 , g74 , g75 , g76 , g77 , g78 , g79 , g80 , g81 , g82 , g83 , g84 , g85 , g86 , g87 , g88 , g89 , g90 , g91 , g92 , g93 , g94 , g95 , g96 , g97 , g98 , g99 , g100 , g101 , g102 , g103 , g104 , g105 , g106 , g107 , g108 , g109 , g110 , g111 , g112 , g113 , g114 , g115 , g116 , g117 , g118 , g119 , g120 , g121 , g122 , g123 , g124 , g125 , g126 , g127 , g128 , g129 , g130 , g131 , g132 , g133 , g134 , g135 , g136 , g137 , g138 , g139 , g140 , g141 , g142 , g143 , g144 , g145 , g146 , g147 , g148 , g149 , g150 , g151 , g152 , g153 , g154 , g155 , g156 , g157 , g158 , g159 , g160 , g161 , g162 , g163 , g164 , g165 , g166 , g167 , g168 , g169 , g170 , g171 , g172 , g173 , g174 , g175 , g176 , g177 , g178 , g179 , g180 , g181 , g182 , g183 , g184 , g185 , g186 , g187 , g188 , g189 , g190 , g191 , g192 , g193 , g194 , g195 , g196 , g197 , g198 , g199 , g200 , g201 , g202 , g203 , g204 , g205 , g206 ;
output g207 , g208 , g209 , g210 , g211 , g212 , g213 , g214 , g215 , g216 , g217 , g218 , g219 , g220 , g221 , g222 , g223 , g224 , g225 , g226 , g227 , g228 , g229 , g230 ;

wire n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , 
     n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , 
     n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , 
     n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , 
     n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , 
     n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , 
     n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , 
     n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , 
     n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , 
     n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , 
     n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , 
     n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , 
     n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , 
     n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , 
     n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , 
     n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , 
     n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , 
     n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , 
     n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , 
     n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , 
     n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , 
     n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , 
     n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , 
     n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , 
     n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , 
     n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , 
     n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , 
     n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , 
     n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , 
     n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , 
     n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , 
     n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , 
     n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , 
     n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , 
     n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , 
     n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , 
     n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , 
     n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , 
     n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , 
     n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , 
     n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , 
     n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , 
     n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , 
     n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , 
     n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , 
     n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , 
     n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , 
     n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , 
     n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , 
     n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , 
     n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , 
     n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , 
     n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , 
     n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , 
     n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , 
     n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , 
     n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , 
     n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , 
     n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , 
     n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , 
     n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , 
     n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , 
     n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , 
     n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , 
     n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , 
     n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , 
     n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , 
     n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , 
     n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , 
     n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , 
     n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , 
     n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , 
     n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , 
     n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , 
     n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , 
     n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , 
     n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , 
     n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , 
     n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , 
     n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , 
     n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , 
     n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , 
     n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , 
     n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , 
     n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , 
     n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , 
     n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , 
     n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , 
     n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , 
     n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , 
     n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , 
     n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , 
     n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , 
     n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , 
     n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , 
     n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , 
     n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , 
     n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , 
     n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , 
     n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , 
     n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , 
     n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , 
     n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , 
     n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , 
     n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , 
     n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , 
     n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , 
     n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , 
     n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , 
     n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , 
     n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , 
     n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , 
     n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , 
     n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , 
     n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , 
     n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , 
     n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , 
     n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , 
     n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , 
     n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , 
     n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , 
     n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , 
     n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , 
     n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , 
     n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , 
     n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , 
     n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , 
     n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , 
     n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , 
     n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , 
     n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , 
     n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , 
     n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , 
     n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , 
     n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , 
     n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , 
     n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , 
     n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , 
     n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , 
     n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , 
     n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , 
     n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , 
     n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , 
     n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , 
     n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , 
     n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , 
     n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , 
     n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , 
     n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , 
     n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , 
     n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , 
     n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , 
     n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , 
     n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , 
     n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , 
     n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , 
     n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , 
     n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , 
     n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , 
     n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , 
     n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , 
     n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , 
     n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , 
     n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , 
     n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , 
     n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , 
     n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , 
     n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , 
     n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , 
     n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 ;
buf ( n1 , g0 );
buf ( n2 , g1 );
buf ( n3 , g2 );
buf ( n4 , g3 );
buf ( n5 , g4 );
buf ( n6 , g5 );
buf ( n7 , g6 );
buf ( n8 , g7 );
buf ( n9 , g8 );
buf ( n10 , g9 );
buf ( n11 , g10 );
buf ( n12 , g11 );
buf ( n13 , g12 );
buf ( n14 , g13 );
buf ( n15 , g14 );
buf ( n16 , g15 );
buf ( n17 , g16 );
buf ( n18 , g17 );
buf ( n19 , g18 );
buf ( n20 , g19 );
buf ( n21 , g20 );
buf ( n22 , g21 );
buf ( n23 , g22 );
buf ( n24 , g23 );
buf ( n25 , g24 );
buf ( n26 , g25 );
buf ( n27 , g26 );
buf ( n28 , g27 );
buf ( n29 , g28 );
buf ( n30 , g29 );
buf ( n31 , g30 );
buf ( n32 , g31 );
buf ( n33 , g32 );
buf ( n34 , g33 );
buf ( n35 , g34 );
buf ( n36 , g35 );
buf ( n37 , g36 );
buf ( n38 , g37 );
buf ( n39 , g38 );
buf ( n40 , g39 );
buf ( n41 , g40 );
buf ( n42 , g41 );
buf ( n43 , g42 );
buf ( n44 , g43 );
buf ( n45 , g44 );
buf ( n46 , g45 );
buf ( n47 , g46 );
buf ( n48 , g47 );
buf ( n49 , g48 );
buf ( n50 , g49 );
buf ( n51 , g50 );
buf ( n52 , g51 );
buf ( n53 , g52 );
buf ( n54 , g53 );
buf ( n55 , g54 );
buf ( n56 , g55 );
buf ( n57 , g56 );
buf ( n58 , g57 );
buf ( n59 , g58 );
buf ( n60 , g59 );
buf ( n61 , g60 );
buf ( n62 , g61 );
buf ( n63 , g62 );
buf ( n64 , g63 );
buf ( n65 , g64 );
buf ( n66 , g65 );
buf ( n67 , g66 );
buf ( n68 , g67 );
buf ( n69 , g68 );
buf ( n70 , g69 );
buf ( n71 , g70 );
buf ( n72 , g71 );
buf ( n73 , g72 );
buf ( n74 , g73 );
buf ( n75 , g74 );
buf ( n76 , g75 );
buf ( n77 , g76 );
buf ( n78 , g77 );
buf ( n79 , g78 );
buf ( n80 , g79 );
buf ( n81 , g80 );
buf ( n82 , g81 );
buf ( n83 , g82 );
buf ( n84 , g83 );
buf ( n85 , g84 );
buf ( n86 , g85 );
buf ( n87 , g86 );
buf ( n88 , g87 );
buf ( n89 , g88 );
buf ( n90 , g89 );
buf ( n91 , g90 );
buf ( n92 , g91 );
buf ( n93 , g92 );
buf ( n94 , g93 );
buf ( n95 , g94 );
buf ( n96 , g95 );
buf ( n97 , g96 );
buf ( n98 , g97 );
buf ( n99 , g98 );
buf ( n100 , g99 );
buf ( n101 , g100 );
buf ( n102 , g101 );
buf ( n103 , g102 );
buf ( n104 , g103 );
buf ( n105 , g104 );
buf ( n106 , g105 );
buf ( n107 , g106 );
buf ( n108 , g107 );
buf ( n109 , g108 );
buf ( n110 , g109 );
buf ( n111 , g110 );
buf ( n112 , g111 );
buf ( n113 , g112 );
buf ( n114 , g113 );
buf ( n115 , g114 );
buf ( n116 , g115 );
buf ( n117 , g116 );
buf ( n118 , g117 );
buf ( n119 , g118 );
buf ( n120 , g119 );
buf ( n121 , g120 );
buf ( n122 , g121 );
buf ( n123 , g122 );
buf ( n124 , g123 );
buf ( n125 , g124 );
buf ( n126 , g125 );
buf ( n127 , g126 );
buf ( n128 , g127 );
buf ( n129 , g128 );
buf ( n130 , g129 );
buf ( n131 , g130 );
buf ( n132 , g131 );
buf ( n133 , g132 );
buf ( n134 , g133 );
buf ( n135 , g134 );
buf ( n136 , g135 );
buf ( n137 , g136 );
buf ( n138 , g137 );
buf ( n139 , g138 );
buf ( n140 , g139 );
buf ( n141 , g140 );
buf ( n142 , g141 );
buf ( n143 , g142 );
buf ( n144 , g143 );
buf ( n145 , g144 );
buf ( n146 , g145 );
buf ( n147 , g146 );
buf ( n148 , g147 );
buf ( n149 , g148 );
buf ( n150 , g149 );
buf ( n151 , g150 );
buf ( n152 , g151 );
buf ( n153 , g152 );
buf ( n154 , g153 );
buf ( n155 , g154 );
buf ( n156 , g155 );
buf ( n157 , g156 );
buf ( n158 , g157 );
buf ( n159 , g158 );
buf ( n160 , g159 );
buf ( n161 , g160 );
buf ( n162 , g161 );
buf ( n163 , g162 );
buf ( n164 , g163 );
buf ( n165 , g164 );
buf ( n166 , g165 );
buf ( n167 , g166 );
buf ( n168 , g167 );
buf ( n169 , g168 );
buf ( n170 , g169 );
buf ( n171 , g170 );
buf ( n172 , g171 );
buf ( n173 , g172 );
buf ( n174 , g173 );
buf ( n175 , g174 );
buf ( n176 , g175 );
buf ( n177 , g176 );
buf ( n178 , g177 );
buf ( n179 , g178 );
buf ( n180 , g179 );
buf ( n181 , g180 );
buf ( n182 , g181 );
buf ( n183 , g182 );
buf ( n184 , g183 );
buf ( n185 , g184 );
buf ( n186 , g185 );
buf ( n187 , g186 );
buf ( n188 , g187 );
buf ( n189 , g188 );
buf ( n190 , g189 );
buf ( n191 , g190 );
buf ( n192 , g191 );
buf ( n193 , g192 );
buf ( n194 , g193 );
buf ( n195 , g194 );
buf ( n196 , g195 );
buf ( n197 , g196 );
buf ( n198 , g197 );
buf ( n199 , g198 );
buf ( n200 , g199 );
buf ( n201 , g200 );
buf ( n202 , g201 );
buf ( n203 , g202 );
buf ( n204 , g203 );
buf ( n205 , g204 );
buf ( n206 , g205 );
buf ( n207 , g206 );
buf ( g207 , n208 );
buf ( g208 , n209 );
buf ( g209 , n210 );
buf ( g210 , n211 );
buf ( g211 , n212 );
buf ( g212 , n213 );
buf ( g213 , n214 );
buf ( g214 , n215 );
buf ( g215 , n216 );
buf ( g216 , n217 );
buf ( g217 , n218 );
buf ( g218 , n219 );
buf ( g219 , n220 );
buf ( g220 , n221 );
buf ( g221 , n222 );
buf ( g222 , n223 );
buf ( g223 , n224 );
buf ( g224 , n225 );
buf ( g225 , n226 );
buf ( g226 , n227 );
buf ( g227 , n228 );
buf ( g228 , n229 );
buf ( g229 , n230 );
buf ( g230 , n231 );
buf ( n208 , n1699 );
buf ( n209 , n1331 );
buf ( n210 , n1457 );
buf ( n211 , n932 );
buf ( n212 , n1660 );
buf ( n213 , n1291 );
buf ( n214 , n1114 );
buf ( n215 , n1000 );
buf ( n216 , n1414 );
buf ( n217 , n1484 );
buf ( n218 , n1081 );
buf ( n219 , n1367 );
buf ( n220 , n1386 );
buf ( n221 , n1025 );
buf ( n222 , n1548 );
buf ( n223 , n1643 );
buf ( n224 , n1572 );
buf ( n225 , n1591 );
buf ( n226 , n1610 );
buf ( n227 , n1690 );
buf ( n228 , n1401 );
buf ( n229 , n1620 );
buf ( n230 , n1528 );
buf ( n231 , n478 );
not ( n234 , n177 );
not ( n235 , n2 );
nand ( n236 , n235 , n178 );
nand ( n237 , n234 , n236 );
or ( n238 , n181 , n182 );
and ( n239 , n237 , n238 );
not ( n240 , n239 );
not ( n241 , n196 );
not ( n242 , n241 );
nand ( n243 , n184 , n185 );
not ( n244 , n243 );
or ( n245 , n242 , n244 );
or ( n246 , n243 , n241 );
not ( n247 , n197 );
nand ( n248 , n246 , n247 );
nand ( n249 , n245 , n248 );
not ( n250 , n187 );
nand ( n251 , n189 , n186 , n188 );
nand ( n252 , n250 , n251 );
nor ( n253 , n184 , n185 );
nor ( n254 , n196 , n197 );
nor ( n255 , n253 , n254 );
not ( n256 , n186 );
nand ( n257 , n188 , n189 );
nand ( n258 , n256 , n257 );
nand ( n259 , n252 , n255 , n258 );
and ( n260 , n249 , n259 );
not ( n261 , n195 );
nor ( n262 , n261 , n2 );
or ( n263 , n262 , n194 );
nand ( n264 , n263 , n235 );
nor ( n265 , n260 , n264 );
and ( n266 , n262 , n194 );
or ( n267 , n265 , n266 );
or ( n268 , n192 , n193 );
nand ( n269 , n267 , n268 );
nand ( n270 , n235 , n192 , n193 );
nand ( n271 , n269 , n270 );
or ( n272 , n190 , n191 );
nand ( n273 , n271 , n272 );
nand ( n274 , n235 , n190 , n191 );
and ( n275 , n273 , n274 );
nor ( n276 , n202 , n203 );
nor ( n277 , n204 , n205 );
or ( n278 , n276 , n277 );
nor ( n279 , n275 , n278 );
nor ( n280 , n179 , n180 );
nor ( n281 , n167 , n168 );
nor ( n282 , n280 , n281 );
not ( n283 , n169 );
not ( n284 , n170 );
nand ( n285 , n283 , n284 );
nand ( n286 , n282 , n285 );
nor ( n287 , n173 , n174 );
nor ( n288 , n286 , n287 );
or ( n289 , n171 , n172 );
nand ( n290 , n288 , n289 );
not ( n291 , n290 );
or ( n292 , n159 , n160 );
nand ( n293 , n291 , n292 );
nor ( n294 , n163 , n164 );
nor ( n295 , n165 , n166 );
nor ( n296 , n294 , n295 );
not ( n297 , n296 );
nor ( n298 , n155 , n156 );
nor ( n299 , n297 , n298 );
or ( n300 , n157 , n158 );
or ( n301 , n151 , n152 );
nand ( n302 , n300 , n301 );
not ( n303 , n302 );
not ( n304 , n153 );
not ( n305 , n154 );
nand ( n306 , n304 , n305 );
nand ( n307 , n303 , n306 );
nor ( n308 , n161 , n162 );
nor ( n309 , n198 , n199 );
or ( n310 , n308 , n309 );
nor ( n311 , n307 , n310 );
nand ( n312 , n299 , n311 );
nor ( n313 , n200 , n201 );
nor ( n314 , n312 , n313 );
not ( n315 , n314 );
nor ( n316 , n293 , n315 );
nand ( n317 , n279 , n316 );
not ( n318 , n2 );
nand ( n319 , n318 , n200 , n201 );
not ( n320 , n319 );
nand ( n321 , n198 , n199 );
nor ( n322 , n321 , n2 );
nor ( n323 , n320 , n322 );
nor ( n324 , n312 , n323 );
not ( n325 , n324 );
nand ( n326 , n235 , n204 , n205 );
or ( n327 , n326 , n276 );
nand ( n328 , n235 , n202 , n203 );
nand ( n329 , n327 , n328 );
nand ( n330 , n314 , n329 );
nand ( n331 , n325 , n330 );
not ( n332 , n293 );
and ( n333 , n331 , n332 );
nand ( n334 , n235 , n171 , n172 );
not ( n335 , n334 );
and ( n336 , n288 , n335 );
nand ( n337 , n169 , n170 );
nor ( n338 , n337 , n2 );
nand ( n339 , n167 , n168 );
nor ( n340 , n339 , n2 );
nor ( n341 , n338 , n340 );
not ( n342 , n282 );
or ( n343 , n341 , n342 );
not ( n344 , n2 );
nand ( n345 , n344 , n181 , n182 );
nand ( n346 , n343 , n345 );
nor ( n347 , n336 , n346 );
not ( n348 , n180 );
not ( n349 , n179 );
or ( n350 , n348 , n349 );
nand ( n351 , n173 , n174 );
or ( n352 , n286 , n351 );
nand ( n353 , n350 , n352 );
nand ( n354 , n353 , n235 );
nand ( n355 , n347 , n354 );
nor ( n356 , n333 , n355 );
nand ( n357 , n235 , n155 , n156 );
not ( n358 , n357 );
not ( n359 , n158 );
not ( n360 , n157 );
or ( n361 , n359 , n360 );
and ( n362 , n153 , n154 );
and ( n363 , n151 , n152 );
nor ( n364 , n362 , n363 );
or ( n365 , n302 , n364 );
nand ( n366 , n361 , n365 );
nand ( n367 , n366 , n235 );
not ( n368 , n367 );
or ( n369 , n358 , n368 );
nand ( n370 , n369 , n299 );
not ( n371 , n2 );
nand ( n372 , n371 , n165 , n166 );
not ( n373 , n372 );
not ( n374 , n294 );
and ( n375 , n373 , n374 );
nand ( n376 , n161 , n162 );
nand ( n377 , n163 , n164 );
and ( n378 , n376 , n377 );
nor ( n379 , n378 , n2 );
nor ( n380 , n375 , n379 );
and ( n381 , n370 , n380 );
nor ( n382 , n381 , n308 );
and ( n383 , n235 , n159 , n160 );
or ( n384 , n382 , n383 );
nand ( n385 , n384 , n332 );
nand ( n386 , n317 , n356 , n385 );
not ( n387 , n386 );
or ( n388 , n240 , n387 );
and ( n389 , n235 , n175 );
nand ( n390 , n389 , n176 );
not ( n391 , n236 );
nand ( n392 , n391 , n177 );
nand ( n393 , n390 , n392 );
not ( n394 , n393 );
nand ( n395 , n388 , n394 );
not ( n396 , n2 );
nand ( n397 , n396 , n115 );
not ( n398 , n397 );
not ( n399 , n398 );
not ( n400 , n183 );
and ( n401 , n399 , n400 );
nor ( n402 , n389 , n176 );
nor ( n403 , n401 , n402 );
and ( n404 , n395 , n403 );
and ( n405 , n398 , n183 );
nor ( n406 , n404 , n405 );
not ( n407 , n207 );
and ( n408 , n406 , n407 );
not ( n409 , n406 );
and ( n410 , n409 , n207 );
nor ( n411 , n408 , n410 );
not ( n412 , n117 );
nor ( n413 , n412 , n150 );
or ( n414 , n413 , n126 );
not ( n415 , n82 );
and ( n416 , n415 , n126 );
nor ( n417 , n416 , n2 );
and ( n418 , n117 , n82 );
not ( n419 , n117 );
and ( n420 , n419 , n116 );
nor ( n421 , n418 , n420 );
nand ( n422 , n414 , n417 , n421 );
nand ( n423 , n411 , n422 );
nand ( n424 , n235 , n206 );
not ( n425 , n424 );
and ( n426 , n423 , n425 );
not ( n427 , n423 );
and ( n428 , n427 , n424 );
nor ( n429 , n426 , n428 );
or ( n430 , n429 , n67 );
not ( n431 , n3 );
nor ( n432 , n431 , n2 );
buf ( n433 , n432 );
nand ( n434 , n433 , n4 );
and ( n435 , n434 , n1 );
not ( n436 , n435 );
nor ( n437 , n19 , n28 );
nor ( n438 , n23 , n24 );
nor ( n439 , n16 , n26 );
nand ( n440 , n437 , n438 , n439 );
nor ( n441 , n17 , n25 );
nor ( n442 , n18 , n31 );
nand ( n443 , n441 , n442 );
nor ( n444 , n440 , n443 );
nor ( n445 , n13 , n15 );
not ( n446 , n12 );
nand ( n447 , n445 , n446 );
not ( n448 , n20 );
nor ( n449 , n21 , n27 );
nand ( n450 , n448 , n449 );
nor ( n451 , n447 , n450 );
nor ( n452 , n8 , n11 );
nor ( n453 , n9 , n14 );
nand ( n454 , n452 , n453 );
nor ( n455 , n22 , n29 );
nor ( n456 , n10 , n30 );
nand ( n457 , n455 , n456 );
nor ( n458 , n454 , n457 );
nand ( n459 , n444 , n451 , n458 );
not ( n460 , n459 );
nor ( n461 , n7 , n5 , n6 );
and ( n462 , n460 , n461 );
not ( n463 , n2 );
nand ( n464 , n463 , n3 );
buf ( n465 , n464 );
nor ( n466 , n462 , n465 );
nor ( n467 , n466 , n2 );
not ( n468 , n467 );
or ( n469 , n436 , n468 );
not ( n470 , n434 );
not ( n471 , n466 );
not ( n472 , n471 );
or ( n473 , n470 , n472 );
not ( n474 , n1 );
nand ( n475 , n473 , n474 );
nand ( n476 , n469 , n475 );
nand ( n477 , n476 , n67 );
nand ( n478 , n430 , n477 );
or ( n479 , n432 , n17 );
not ( n480 , n479 );
nor ( n481 , n22 , n26 );
nor ( n482 , n18 , n21 );
nor ( n483 , n24 , n27 );
nand ( n484 , n481 , n482 , n483 );
nor ( n485 , n23 , n25 );
not ( n486 , n20 );
nand ( n487 , n485 , n486 );
nor ( n488 , n484 , n487 );
buf ( n489 , n488 );
nor ( n490 , n16 , n17 , n19 );
nand ( n491 , n489 , n490 );
not ( n492 , n491 );
nor ( n493 , n480 , n492 );
nand ( n494 , n432 , n16 );
not ( n495 , n494 );
not ( n496 , n19 );
not ( n497 , n496 );
not ( n498 , n488 );
or ( n499 , n497 , n498 );
nand ( n500 , n499 , n432 );
not ( n501 , n500 );
or ( n502 , n495 , n501 );
nand ( n503 , n502 , n17 );
nand ( n504 , n493 , n503 );
not ( n505 , n47 );
and ( n506 , n504 , n505 );
not ( n507 , n504 );
and ( n508 , n507 , n47 );
nor ( n509 , n506 , n508 );
not ( n510 , n509 );
not ( n511 , n27 );
not ( n512 , n2 );
nand ( n513 , n512 , n3 );
not ( n514 , n513 );
not ( n515 , n514 );
nor ( n516 , n511 , n515 );
not ( n517 , n516 );
nor ( n518 , n23 , n22 , n25 );
nor ( n519 , n20 , n21 );
not ( n520 , n24 );
nand ( n521 , n518 , n519 , n520 );
not ( n522 , n521 );
or ( n523 , n517 , n522 );
not ( n524 , n3 );
nor ( n525 , n524 , n2 );
not ( n526 , n525 );
not ( n527 , n27 );
and ( n528 , n526 , n527 );
not ( n529 , n487 );
nor ( n530 , n21 , n24 );
nor ( n531 , n22 , n27 );
nand ( n532 , n530 , n531 );
not ( n533 , n532 );
and ( n534 , n529 , n533 );
nor ( n535 , n528 , n534 );
nand ( n536 , n523 , n535 );
not ( n537 , n536 );
not ( n538 , n537 );
not ( n539 , n40 );
or ( n540 , n538 , n539 );
not ( n541 , n22 );
not ( n542 , n513 );
not ( n543 , n542 );
or ( n544 , n541 , n543 );
not ( n545 , n23 );
not ( n546 , n545 );
not ( n547 , n519 );
or ( n548 , n546 , n547 );
nand ( n549 , n548 , n542 );
nand ( n550 , n544 , n549 );
not ( n551 , n25 );
and ( n552 , n550 , n551 );
not ( n553 , n550 );
and ( n554 , n553 , n25 );
nor ( n555 , n552 , n554 );
not ( n556 , n555 );
and ( n557 , n556 , n42 );
nand ( n558 , n519 , n518 );
nand ( n559 , n558 , n525 , n24 );
nand ( n560 , n515 , n520 );
nand ( n561 , n559 , n521 , n560 );
not ( n562 , n561 );
and ( n563 , n562 , n39 );
nor ( n564 , n557 , n563 );
not ( n565 , n564 );
not ( n566 , n549 );
and ( n567 , n566 , n22 );
not ( n568 , n566 );
not ( n569 , n22 );
and ( n570 , n568 , n569 );
nor ( n571 , n567 , n570 );
not ( n572 , n571 );
not ( n573 , n41 );
nor ( n574 , n572 , n573 );
not ( n575 , n37 );
or ( n576 , n20 , n21 );
nand ( n577 , n576 , n3 );
xor ( n578 , n577 , n23 );
not ( n579 , n578 );
not ( n580 , n579 );
or ( n581 , n575 , n580 );
and ( n582 , n37 , n23 );
not ( n583 , n37 );
and ( n584 , n583 , n545 );
or ( n585 , n582 , n584 );
not ( n586 , n585 );
not ( n587 , n3 );
nor ( n588 , n20 , n21 );
nor ( n589 , n587 , n588 );
not ( n590 , n589 );
or ( n591 , n586 , n590 );
or ( n592 , n589 , n585 );
nand ( n593 , n591 , n592 );
and ( n594 , n20 , n38 );
not ( n595 , n594 );
xor ( n596 , n36 , n21 );
nand ( n597 , n3 , n20 );
not ( n598 , n597 );
xor ( n599 , n596 , n598 );
not ( n600 , n599 );
or ( n601 , n595 , n600 );
not ( n602 , n597 );
not ( n603 , n21 );
not ( n604 , n603 );
and ( n605 , n602 , n604 );
and ( n606 , n597 , n603 );
nor ( n607 , n605 , n606 );
nand ( n608 , n607 , n36 );
nand ( n609 , n601 , n608 );
nand ( n610 , n593 , n609 );
nand ( n611 , n581 , n610 );
or ( n612 , n574 , n611 );
not ( n613 , n571 );
nand ( n614 , n613 , n573 );
nand ( n615 , n612 , n614 );
not ( n616 , n615 );
not ( n617 , n42 );
not ( n618 , n555 );
or ( n619 , n617 , n618 );
or ( n620 , n555 , n42 );
nand ( n621 , n619 , n620 );
nand ( n622 , n616 , n621 );
not ( n623 , n622 );
or ( n624 , n565 , n623 );
not ( n625 , n40 );
and ( n626 , n536 , n625 );
not ( n627 , n536 );
and ( n628 , n627 , n40 );
nor ( n629 , n626 , n628 );
not ( n630 , n39 );
nand ( n631 , n630 , n561 );
and ( n632 , n629 , n631 );
nand ( n633 , n624 , n632 );
nand ( n634 , n540 , n633 );
not ( n635 , n634 );
nor ( n636 , n500 , n16 );
not ( n637 , n636 );
nand ( n638 , n500 , n16 );
nand ( n639 , n637 , n638 );
xnor ( n640 , n43 , n639 );
not ( n641 , n640 );
not ( n642 , n26 );
not ( n643 , n642 );
not ( n644 , n533 );
not ( n645 , n529 );
or ( n646 , n644 , n645 );
nand ( n647 , n646 , n525 );
not ( n648 , n647 );
or ( n649 , n643 , n648 );
not ( n650 , n647 );
nand ( n651 , n650 , n26 );
nand ( n652 , n649 , n651 );
xnor ( n653 , n45 , n652 );
not ( n654 , n46 );
nor ( n655 , n23 , n25 , n20 );
nand ( n656 , n533 , n655 );
nor ( n657 , n656 , n26 );
nor ( n658 , n657 , n515 );
and ( n659 , n658 , n18 );
not ( n660 , n658 );
not ( n661 , n18 );
and ( n662 , n660 , n661 );
nor ( n663 , n659 , n662 );
not ( n664 , n663 );
xor ( n665 , n654 , n664 );
nor ( n666 , n488 , n464 );
and ( n667 , n666 , n19 );
not ( n668 , n666 );
and ( n669 , n668 , n496 );
nor ( n670 , n667 , n669 );
xor ( n671 , n44 , n670 );
and ( n672 , n653 , n665 , n671 );
and ( n673 , n641 , n672 );
not ( n674 , n673 );
or ( n675 , n635 , n674 );
and ( n676 , n654 , n664 );
not ( n677 , n652 );
nand ( n678 , n677 , n45 );
or ( n679 , n676 , n678 );
and ( n680 , n658 , n18 );
not ( n681 , n658 );
and ( n682 , n681 , n661 );
nor ( n683 , n680 , n682 );
nand ( n684 , n683 , n46 );
nand ( n685 , n679 , n684 );
and ( n686 , n685 , n671 );
and ( n687 , n44 , n670 );
nor ( n688 , n686 , n687 );
not ( n689 , n688 );
and ( n690 , n689 , n641 );
and ( n691 , n639 , n43 );
nor ( n692 , n690 , n691 );
nand ( n693 , n675 , n692 );
not ( n694 , n693 );
or ( n695 , n510 , n694 );
not ( n696 , n504 );
nand ( n697 , n696 , n47 );
nand ( n698 , n695 , n697 );
and ( n699 , n432 , n28 );
not ( n700 , n699 );
not ( n701 , n491 );
or ( n702 , n700 , n701 );
not ( n703 , n28 );
not ( n704 , n703 );
not ( n705 , n465 );
or ( n706 , n704 , n705 );
nor ( n707 , n16 , n22 );
nor ( n708 , n25 , n27 );
and ( n709 , n438 , n437 , n707 , n708 );
nor ( n710 , n26 , n17 , n18 );
and ( n711 , n588 , n710 );
nand ( n712 , n709 , n711 );
nand ( n713 , n706 , n712 );
not ( n714 , n713 );
nand ( n715 , n702 , n714 );
xor ( n716 , n715 , n48 );
buf ( n717 , n716 );
not ( n718 , n717 );
nand ( n719 , n698 , n718 );
not ( n720 , n719 );
not ( n721 , n467 );
nand ( n722 , n721 , n4 );
not ( n723 , n4 );
nand ( n724 , n723 , n471 );
and ( n725 , n722 , n724 , n67 );
and ( n726 , n725 , n476 );
buf ( n727 , n726 );
buf ( n728 , n727 );
not ( n729 , n49 );
and ( n730 , n712 , n432 );
and ( n731 , n730 , n29 );
not ( n732 , n730 );
not ( n733 , n29 );
and ( n734 , n732 , n733 );
nor ( n735 , n731 , n734 );
not ( n736 , n735 );
not ( n737 , n736 );
or ( n738 , n729 , n737 );
or ( n739 , n49 , n736 );
nand ( n740 , n738 , n739 );
buf ( n741 , n740 );
not ( n742 , n741 );
and ( n743 , n728 , n742 );
nand ( n744 , n720 , n743 );
not ( n745 , n698 );
not ( n746 , n718 );
or ( n747 , n745 , n746 );
not ( n748 , n742 );
nand ( n749 , n748 , n727 );
and ( n750 , n491 , n699 );
nor ( n751 , n750 , n713 );
and ( n752 , n751 , n48 );
nor ( n753 , n749 , n752 );
nand ( n754 , n747 , n753 );
and ( n755 , n58 , n556 );
not ( n756 , n58 );
and ( n757 , n756 , n555 );
nor ( n758 , n755 , n757 );
not ( n759 , n758 );
nand ( n760 , n20 , n54 );
not ( n761 , n760 );
and ( n762 , n607 , n761 );
and ( n763 , n761 , n52 );
nor ( n764 , n762 , n763 );
nand ( n765 , n607 , n52 );
and ( n766 , n764 , n765 );
not ( n767 , n766 );
not ( n768 , n578 );
not ( n769 , n53 );
or ( n770 , n768 , n769 );
or ( n771 , n578 , n53 );
nand ( n772 , n770 , n771 );
nand ( n773 , n767 , n772 );
not ( n774 , n57 );
not ( n775 , n571 );
or ( n776 , n774 , n775 );
nand ( n777 , n579 , n53 );
nand ( n778 , n776 , n777 );
not ( n779 , n778 );
and ( n780 , n773 , n779 );
buf ( n781 , n571 );
nor ( n782 , n781 , n57 );
nor ( n783 , n780 , n782 );
not ( n784 , n783 );
or ( n785 , n759 , n784 );
nand ( n786 , n670 , n60 );
nand ( n787 , n663 , n62 );
and ( n788 , n786 , n787 );
not ( n789 , n788 );
nand ( n790 , n556 , n58 );
nand ( n791 , n677 , n61 );
nand ( n792 , n537 , n56 );
nand ( n793 , n562 , n55 );
nand ( n794 , n790 , n791 , n792 , n793 );
nor ( n795 , n789 , n794 );
nand ( n796 , n785 , n795 );
not ( n797 , n56 );
and ( n798 , n536 , n797 );
nand ( n799 , n791 , n787 , n798 );
not ( n800 , n799 );
xor ( n801 , n670 , n60 );
not ( n802 , n801 );
or ( n803 , n800 , n802 );
buf ( n804 , n786 );
buf ( n805 , n804 );
nand ( n806 , n803 , n805 );
not ( n807 , n793 );
not ( n808 , n55 );
not ( n809 , n808 );
not ( n810 , n562 );
or ( n811 , n809 , n810 );
or ( n812 , n562 , n808 );
nand ( n813 , n811 , n812 );
nor ( n814 , n807 , n813 );
nand ( n815 , n814 , n804 , n791 );
nand ( n816 , n787 , n792 );
nor ( n817 , n815 , n816 );
not ( n818 , n59 );
and ( n819 , n639 , n818 );
not ( n820 , n639 );
and ( n821 , n820 , n59 );
nor ( n822 , n819 , n821 );
nor ( n823 , n817 , n822 );
xnor ( n824 , n62 , n664 );
not ( n825 , n824 );
not ( n826 , n61 );
xor ( n827 , n647 , n26 );
nand ( n828 , n826 , n827 );
not ( n829 , n828 );
or ( n830 , n825 , n829 );
nand ( n831 , n830 , n788 );
nand ( n832 , n796 , n806 , n823 , n831 );
not ( n833 , n504 );
nand ( n834 , n833 , n63 );
nand ( n835 , n751 , n64 );
nand ( n836 , n639 , n59 );
and ( n837 , n834 , n835 , n836 );
nand ( n838 , n832 , n837 );
nor ( n839 , n833 , n63 );
and ( n840 , n835 , n839 );
not ( n841 , n835 );
not ( n842 , n64 );
not ( n843 , n715 );
or ( n844 , n842 , n843 );
not ( n845 , n64 );
nand ( n846 , n845 , n751 );
nand ( n847 , n844 , n846 );
nor ( n848 , n841 , n847 );
nor ( n849 , n840 , n848 );
nand ( n850 , n838 , n849 );
not ( n851 , n736 );
xor ( n852 , n65 , n851 );
not ( n853 , n852 );
and ( n854 , n850 , n853 );
not ( n855 , n850 );
and ( n856 , n855 , n852 );
nor ( n857 , n854 , n856 );
nand ( n858 , n724 , n722 );
not ( n859 , n858 );
nor ( n860 , n477 , n859 );
buf ( n861 , n860 );
buf ( n862 , n861 );
nand ( n863 , n857 , n862 );
not ( n864 , n7 );
not ( n865 , n864 );
not ( n866 , n460 );
or ( n867 , n865 , n866 );
nand ( n868 , n867 , n433 );
or ( n869 , n6 , n868 );
not ( n870 , n6 );
nor ( n871 , n870 , n2 );
nand ( n872 , n868 , n871 );
nand ( n873 , n869 , n872 );
nor ( n874 , n16 , n29 );
nand ( n875 , n481 , n874 );
nor ( n876 , n875 , n450 );
nor ( n877 , n17 , n23 );
nor ( n878 , n24 , n25 );
nand ( n879 , n877 , n878 );
nor ( n880 , n18 , n19 );
nor ( n881 , n28 , n31 );
nand ( n882 , n880 , n881 );
nor ( n883 , n879 , n882 );
nand ( n884 , n876 , n883 );
not ( n885 , n884 );
not ( n886 , n30 );
nand ( n887 , n885 , n886 );
or ( n888 , n454 , n447 );
or ( n889 , n887 , n888 );
nand ( n890 , n889 , n10 );
and ( n891 , n864 , n890 );
not ( n892 , n10 );
not ( n893 , n465 );
or ( n894 , n892 , n893 );
nand ( n895 , n433 , n7 );
or ( n896 , n895 , n460 );
nand ( n897 , n894 , n896 );
nor ( n898 , n891 , n897 );
and ( n899 , n873 , n898 );
not ( n900 , n6 );
not ( n901 , n433 );
or ( n902 , n900 , n901 );
nand ( n903 , n902 , n868 );
and ( n904 , n903 , n5 );
not ( n905 , n903 );
nand ( n906 , n235 , n5 );
and ( n907 , n905 , n906 );
nor ( n908 , n904 , n907 );
nand ( n909 , n899 , n908 );
nand ( n910 , n909 , n858 );
not ( n911 , n910 );
not ( n912 , n476 );
not ( n913 , n67 );
nor ( n914 , n913 , n2 );
and ( n915 , n911 , n912 , n914 );
and ( n916 , n915 , n75 );
nor ( n917 , n476 , n913 );
and ( n918 , n910 , n917 );
not ( n919 , n918 );
not ( n920 , n851 );
or ( n921 , n919 , n920 );
not ( n922 , n726 );
not ( n923 , n922 );
not ( n924 , n752 );
nor ( n925 , n924 , n741 );
and ( n926 , n923 , n925 );
and ( n927 , n235 , n913 );
and ( n928 , n927 , n76 );
nor ( n929 , n926 , n928 );
nand ( n930 , n921 , n929 );
nor ( n931 , n916 , n930 );
nand ( n932 , n744 , n754 , n863 , n931 );
not ( n933 , n31 );
nor ( n934 , n465 , n933 );
not ( n935 , n934 );
not ( n936 , n712 );
nand ( n937 , n936 , n733 );
not ( n938 , n937 );
or ( n939 , n935 , n938 );
not ( n940 , n884 );
and ( n941 , n464 , n933 );
nor ( n942 , n940 , n941 );
nand ( n943 , n939 , n942 );
xnor ( n944 , n943 , n50 );
buf ( n945 , n944 );
nor ( n946 , n749 , n945 );
nand ( n947 , n720 , n946 );
not ( n948 , n943 );
not ( n949 , n66 );
and ( n950 , n948 , n949 );
and ( n951 , n943 , n66 );
nor ( n952 , n950 , n951 );
buf ( n953 , n952 );
not ( n954 , n953 );
not ( n955 , n838 );
and ( n956 , n849 , n852 );
not ( n957 , n956 );
or ( n958 , n955 , n957 );
nand ( n959 , n735 , n65 );
nand ( n960 , n958 , n959 );
not ( n961 , n960 );
or ( n962 , n954 , n961 );
or ( n963 , n960 , n953 );
nand ( n964 , n962 , n963 );
nand ( n965 , n964 , n862 );
nand ( n966 , n476 , n725 );
buf ( n967 , n966 );
nand ( n968 , n735 , n49 );
nand ( n969 , n945 , n968 , n924 );
nor ( n970 , n967 , n969 );
nand ( n971 , n719 , n970 );
or ( n972 , n945 , n742 , n924 );
nand ( n973 , n740 , n944 );
not ( n974 , n973 );
and ( n975 , n945 , n968 );
not ( n976 , n945 );
not ( n977 , n968 );
and ( n978 , n976 , n977 );
nor ( n979 , n975 , n978 );
or ( n980 , n974 , n979 );
nand ( n981 , n972 , n980 );
and ( n982 , n981 , n727 );
and ( n983 , n927 , n90 );
nor ( n984 , n982 , n983 );
not ( n985 , n984 );
not ( n986 , n911 );
buf ( n987 , n986 );
not ( n988 , n987 );
not ( n989 , n988 );
not ( n990 , n943 );
not ( n991 , n990 );
and ( n992 , n989 , n991 );
buf ( n993 , n918 );
not ( n994 , n993 );
and ( n995 , n917 , n235 );
nand ( n996 , n995 , n89 );
and ( n997 , n994 , n996 );
nor ( n998 , n992 , n997 );
nor ( n999 , n985 , n998 );
nand ( n1000 , n947 , n965 , n971 , n999 );
not ( n1001 , n847 );
not ( n1002 , n834 );
and ( n1003 , n832 , n836 );
not ( n1004 , n1003 );
or ( n1005 , n1002 , n1004 );
not ( n1006 , n839 );
nand ( n1007 , n1005 , n1006 );
not ( n1008 , n1007 );
or ( n1009 , n1001 , n1008 );
or ( n1010 , n847 , n1007 );
nand ( n1011 , n1009 , n1010 );
nand ( n1012 , n1011 , n862 );
and ( n1013 , n698 , n718 );
not ( n1014 , n698 );
and ( n1015 , n1014 , n717 );
nor ( n1016 , n1013 , n1015 );
nand ( n1017 , n1016 , n728 );
and ( n1018 , n915 , n101 );
not ( n1019 , n751 );
not ( n1020 , n918 );
or ( n1021 , n1019 , n1020 );
nand ( n1022 , n927 , n102 );
nand ( n1023 , n1021 , n1022 );
nor ( n1024 , n1018 , n1023 );
nand ( n1025 , n1012 , n1017 , n1024 );
not ( n1026 , n861 );
buf ( n1027 , n822 );
not ( n1028 , n1027 );
not ( n1029 , n791 );
nor ( n1030 , n1029 , n816 );
not ( n1031 , n1030 );
buf ( n1032 , n813 );
not ( n1033 , n1032 );
nand ( n1034 , n773 , n779 );
not ( n1035 , n1034 );
nor ( n1036 , n556 , n58 );
nor ( n1037 , n1036 , n782 );
not ( n1038 , n1037 );
or ( n1039 , n1035 , n1038 );
nand ( n1040 , n1039 , n790 );
not ( n1041 , n1040 );
or ( n1042 , n1033 , n1041 );
nand ( n1043 , n1042 , n793 );
xor ( n1044 , n536 , n797 );
nand ( n1045 , n1043 , n1044 );
not ( n1046 , n1045 );
or ( n1047 , n1031 , n1046 );
nand ( n1048 , n824 , n828 );
buf ( n1049 , n787 );
nand ( n1050 , n1048 , n1049 );
buf ( n1051 , n801 );
and ( n1052 , n1050 , n1051 );
nand ( n1053 , n1047 , n1052 );
nand ( n1054 , n1053 , n805 );
not ( n1055 , n1054 );
or ( n1056 , n1028 , n1055 );
or ( n1057 , n1054 , n1027 );
nand ( n1058 , n1056 , n1057 );
not ( n1059 , n1058 );
or ( n1060 , n1026 , n1059 );
and ( n1061 , n915 , n95 );
not ( n1062 , n993 );
not ( n1063 , n639 );
or ( n1064 , n1062 , n1063 );
not ( n1065 , n641 );
not ( n1066 , n632 );
nand ( n1067 , n622 , n564 );
not ( n1068 , n1067 );
or ( n1069 , n1066 , n1068 );
nand ( n1070 , n537 , n40 );
nand ( n1071 , n1069 , n1070 );
nand ( n1072 , n1071 , n672 );
nand ( n1073 , n1072 , n688 );
not ( n1074 , n1073 );
xor ( n1075 , n1065 , n1074 );
and ( n1076 , n1075 , n923 );
and ( n1077 , n927 , n96 );
nor ( n1078 , n1076 , n1077 );
nand ( n1079 , n1064 , n1078 );
nor ( n1080 , n1061 , n1079 );
nand ( n1081 , n1060 , n1080 );
and ( n1082 , n1045 , n792 );
nand ( n1083 , n1082 , n791 );
not ( n1084 , n1048 );
nand ( n1085 , n1083 , n1084 );
nand ( n1086 , n1085 , n1049 );
not ( n1087 , n861 );
not ( n1088 , n1087 );
nand ( n1089 , n1088 , n1051 );
or ( n1090 , n1086 , n1089 );
not ( n1091 , n665 );
not ( n1092 , n653 );
nand ( n1093 , n633 , n1070 );
not ( n1094 , n1093 );
or ( n1095 , n1092 , n1094 );
nand ( n1096 , n1095 , n678 );
not ( n1097 , n1096 );
or ( n1098 , n1091 , n1097 );
nand ( n1099 , n1098 , n684 );
xnor ( n1100 , n1099 , n671 );
not ( n1101 , n1100 );
not ( n1102 , n967 );
and ( n1103 , n1101 , n1102 );
not ( n1104 , n87 );
not ( n1105 , n915 );
or ( n1106 , n1104 , n1105 );
and ( n1107 , n918 , n670 );
and ( n1108 , n927 , n88 );
nor ( n1109 , n1107 , n1108 );
nand ( n1110 , n1106 , n1109 );
nor ( n1111 , n1103 , n1110 );
nor ( n1112 , n1087 , n1051 );
nand ( n1113 , n1086 , n1112 );
nand ( n1114 , n1090 , n1111 , n1113 );
nor ( n1115 , n464 , n886 );
not ( n1116 , n1115 );
not ( n1117 , n884 );
or ( n1118 , n1116 , n1117 );
nand ( n1119 , n465 , n886 );
nand ( n1120 , n1118 , n1119 );
not ( n1121 , n1120 );
nand ( n1122 , n1121 , n887 );
and ( n1123 , n35 , n1122 );
not ( n1124 , n35 );
not ( n1125 , n1122 );
and ( n1126 , n1124 , n1125 );
nor ( n1127 , n1123 , n1126 );
and ( n1128 , n883 , n876 , n886 );
not ( n1129 , n1128 );
nand ( n1130 , n1129 , n433 );
not ( n1131 , n1130 );
not ( n1132 , n446 );
and ( n1133 , n1131 , n1132 );
not ( n1134 , n12 );
and ( n1135 , n1130 , n1134 );
nor ( n1136 , n1133 , n1135 );
not ( n1137 , n1136 );
not ( n1138 , n1137 );
not ( n1139 , n69 );
and ( n1140 , n1138 , n1139 );
and ( n1141 , n1137 , n69 );
nor ( n1142 , n1140 , n1141 );
nor ( n1143 , n1127 , n1142 );
not ( n1144 , n1143 );
not ( n1145 , n509 );
nor ( n1146 , n973 , n1145 , n716 , n640 );
not ( n1147 , n1146 );
not ( n1148 , n1073 );
or ( n1149 , n1147 , n1148 );
and ( n1150 , n944 , n977 );
and ( n1151 , n990 , n50 );
nor ( n1152 , n1150 , n1151 );
not ( n1153 , n1152 );
not ( n1154 , n716 );
nand ( n1155 , n1154 , n509 , n691 );
not ( n1156 , n697 );
not ( n1157 , n716 );
and ( n1158 , n1156 , n1157 );
nor ( n1159 , n1158 , n752 );
and ( n1160 , n1155 , n1159 );
nor ( n1161 , n1160 , n973 );
nor ( n1162 , n1153 , n1161 );
nand ( n1163 , n1149 , n1162 );
not ( n1164 , n1163 );
or ( n1165 , n1144 , n1164 );
nand ( n1166 , n1125 , n35 );
or ( n1167 , n1142 , n1166 );
nand ( n1168 , n1165 , n1167 );
not ( n1169 , n1168 );
not ( n1170 , n13 );
not ( n1171 , n433 );
or ( n1172 , n1170 , n1171 );
not ( n1173 , n446 );
not ( n1174 , n1128 );
or ( n1175 , n1173 , n1174 );
nand ( n1176 , n1175 , n525 );
nand ( n1177 , n1172 , n1176 );
and ( n1178 , n1177 , n15 );
not ( n1179 , n1177 );
not ( n1180 , n15 );
and ( n1181 , n1179 , n1180 );
nor ( n1182 , n1178 , n1181 );
and ( n1183 , n1182 , n81 );
not ( n1184 , n80 );
xor ( n1185 , n1176 , n13 );
not ( n1186 , n1185 );
or ( n1187 , n1184 , n1186 );
or ( n1188 , n80 , n1185 );
nand ( n1189 , n1187 , n1188 );
and ( n1190 , n1136 , n69 );
nand ( n1191 , n1189 , n1190 );
not ( n1192 , n1185 );
nand ( n1193 , n1192 , n80 );
and ( n1194 , n1191 , n1193 );
nor ( n1195 , n1182 , n81 );
nor ( n1196 , n1194 , n1195 );
nor ( n1197 , n1183 , n1196 );
not ( n1198 , n887 );
not ( n1199 , n447 );
and ( n1200 , n1198 , n1199 );
nor ( n1201 , n1200 , n465 );
and ( n1202 , n1201 , n14 );
not ( n1203 , n1201 );
not ( n1204 , n14 );
and ( n1205 , n1203 , n1204 );
nor ( n1206 , n1202 , n1205 );
not ( n1207 , n79 );
and ( n1208 , n1206 , n1207 );
not ( n1209 , n1206 );
and ( n1210 , n1209 , n79 );
nor ( n1211 , n1208 , n1210 );
nor ( n1212 , n966 , n1211 );
and ( n1213 , n1197 , n1212 );
nand ( n1214 , n1169 , n1213 );
nand ( n1215 , n726 , n1211 );
not ( n1216 , n1189 );
or ( n1217 , n1216 , n1195 );
or ( n1218 , n1215 , n1217 );
not ( n1219 , n1218 );
nand ( n1220 , n1219 , n1168 );
not ( n1221 , n66 );
nor ( n1222 , n1221 , n943 );
not ( n1223 , n1222 );
and ( n1224 , n959 , n1223 );
nand ( n1225 , n837 , n1224 );
and ( n1226 , n1192 , n84 );
and ( n1227 , n1136 , n70 );
nor ( n1228 , n1226 , n1227 );
nand ( n1229 , n1182 , n85 );
not ( n1230 , n70 );
nand ( n1231 , n1230 , n1137 );
nand ( n1232 , n1231 , n1125 , n51 );
nand ( n1233 , n1228 , n1229 , n1232 );
nor ( n1234 , n1225 , n1233 );
not ( n1235 , n1234 );
not ( n1236 , n832 );
or ( n1237 , n1235 , n1236 );
nor ( n1238 , n1222 , n63 );
nand ( n1239 , n1238 , n959 , n835 , n504 );
nand ( n1240 , n952 , n1223 );
and ( n1241 , n1239 , n1240 );
nand ( n1242 , n848 , n959 , n1223 );
nor ( n1243 , n934 , n1221 );
and ( n1244 , n942 , n1243 );
not ( n1245 , n730 );
and ( n1246 , n1245 , n29 );
nor ( n1247 , n1244 , n1246 );
and ( n1248 , n730 , n733 );
nor ( n1249 , n1248 , n65 );
not ( n1250 , n937 );
nand ( n1251 , n1250 , n884 , n66 );
nand ( n1252 , n1247 , n1249 , n1251 );
not ( n1253 , n51 );
nand ( n1254 , n1253 , n1122 );
and ( n1255 , n1252 , n1231 , n1254 );
nand ( n1256 , n1241 , n1242 , n1255 );
not ( n1257 , n1233 );
and ( n1258 , n1256 , n1257 );
or ( n1259 , n1182 , n85 );
not ( n1260 , n85 );
not ( n1261 , n1182 );
or ( n1262 , n1260 , n1261 );
nor ( n1263 , n1192 , n84 );
nand ( n1264 , n1262 , n1263 );
nand ( n1265 , n1259 , n1264 );
nor ( n1266 , n1258 , n1265 );
nand ( n1267 , n1237 , n1266 );
not ( n1268 , n83 );
and ( n1269 , n1267 , n1268 );
not ( n1270 , n1267 );
and ( n1271 , n1270 , n83 );
nor ( n1272 , n1269 , n1271 );
nor ( n1273 , n1087 , n1206 );
and ( n1274 , n1272 , n1273 );
not ( n1275 , n1206 );
not ( n1276 , n986 );
or ( n1277 , n1275 , n1276 );
nand ( n1278 , n235 , n82 );
or ( n1279 , n1278 , n986 );
nand ( n1280 , n1277 , n1279 );
and ( n1281 , n1280 , n917 );
and ( n1282 , n927 , n86 );
nor ( n1283 , n1281 , n1282 );
nand ( n1284 , n1197 , n1212 , n1217 );
or ( n1285 , n1197 , n1215 );
nand ( n1286 , n1283 , n1284 , n1285 );
nor ( n1287 , n1274 , n1286 );
not ( n1288 , n1272 );
and ( n1289 , n862 , n1206 );
nand ( n1290 , n1288 , n1289 );
nand ( n1291 , n1214 , n1220 , n1287 , n1290 );
not ( n1292 , n1127 );
and ( n1293 , n1163 , n1292 );
nand ( n1294 , n1142 , n1166 );
nor ( n1295 , n1293 , n1294 );
nor ( n1296 , n1295 , n967 );
not ( n1297 , n1168 );
nand ( n1298 , n1296 , n1297 );
and ( n1299 , n1125 , n51 );
not ( n1300 , n1299 );
not ( n1301 , n1227 );
nand ( n1302 , n1231 , n1301 );
not ( n1303 , n1302 );
nand ( n1304 , n1300 , n861 , n1303 );
not ( n1305 , n1304 );
not ( n1306 , n1225 );
not ( n1307 , n1306 );
not ( n1308 , n832 );
or ( n1309 , n1307 , n1308 );
and ( n1310 , n1241 , n1242 , n1252 );
nand ( n1311 , n1309 , n1310 );
not ( n1312 , n1311 );
or ( n1313 , n1305 , n1312 );
not ( n1314 , n1254 );
nor ( n1315 , n1087 , n1303 , n1314 );
or ( n1316 , n1311 , n1315 );
nand ( n1317 , n1313 , n1316 );
nand ( n1318 , n995 , n71 );
and ( n1319 , n994 , n1318 );
and ( n1320 , n987 , n1137 );
nor ( n1321 , n1319 , n1320 );
not ( n1322 , n72 );
not ( n1323 , n927 );
or ( n1324 , n1322 , n1323 );
and ( n1325 , n1303 , n1314 );
and ( n1326 , n1302 , n1299 );
nor ( n1327 , n1325 , n1326 );
or ( n1328 , n1087 , n1327 );
nand ( n1329 , n1324 , n1328 );
nor ( n1330 , n1321 , n1329 );
nand ( n1331 , n1298 , n1317 , n1330 );
not ( n1332 , n1256 );
not ( n1333 , n1332 );
nand ( n1334 , n832 , n1306 );
not ( n1335 , n1334 );
or ( n1336 , n1333 , n1335 );
and ( n1337 , n1232 , n1301 );
nand ( n1338 , n1336 , n1337 );
not ( n1339 , n84 );
not ( n1340 , n1192 );
not ( n1341 , n1340 );
or ( n1342 , n1339 , n1341 );
or ( n1343 , n1340 , n84 );
nand ( n1344 , n1342 , n1343 );
nor ( n1345 , n1344 , n1087 );
and ( n1346 , n1338 , n1345 );
and ( n1347 , n910 , n1340 );
not ( n1348 , n1347 );
and ( n1349 , n995 , n97 );
and ( n1350 , n1348 , n1349 );
nor ( n1351 , n1346 , n1350 );
nor ( n1352 , n967 , n1216 , n1190 );
nand ( n1353 , n1297 , n1352 );
nor ( n1354 , n966 , n1189 );
buf ( n1355 , n1354 );
and ( n1356 , n1355 , n1168 );
nand ( n1357 , n861 , n1344 );
or ( n1358 , n1338 , n1357 );
not ( n1359 , n1347 );
nand ( n1360 , n1359 , n918 );
and ( n1361 , n1354 , n1190 );
and ( n1362 , n927 , n98 );
nor ( n1363 , n1361 , n1362 );
and ( n1364 , n1360 , n1363 );
nand ( n1365 , n1358 , n1364 );
nor ( n1366 , n1356 , n1365 );
nand ( n1367 , n1351 , n1353 , n1366 );
and ( n1368 , n1085 , n824 );
not ( n1369 , n828 );
nor ( n1370 , n1369 , n1084 );
and ( n1371 , n1083 , n1370 );
nor ( n1372 , n1368 , n1371 );
not ( n1373 , n862 );
or ( n1374 , n1372 , n1373 );
not ( n1375 , n665 );
xor ( n1376 , n1096 , n1375 );
or ( n1377 , n1376 , n967 );
nand ( n1378 , n927 , n100 );
nand ( n1379 , n1377 , n1378 );
not ( n1380 , n99 );
not ( n1381 , n915 );
or ( n1382 , n1380 , n1381 );
nand ( n1383 , n993 , n683 );
nand ( n1384 , n1382 , n1383 );
nor ( n1385 , n1379 , n1384 );
nand ( n1386 , n1374 , n1385 );
and ( n1387 , n386 , n238 );
and ( n1388 , n1387 , n237 );
nor ( n1389 , n1388 , n393 );
nor ( n1390 , n1389 , n402 );
and ( n1391 , n397 , n183 );
nor ( n1392 , n397 , n183 );
nor ( n1393 , n1391 , n1392 );
xor ( n1394 , n1390 , n1393 );
nand ( n1395 , n422 , n913 );
or ( n1396 , n1394 , n1395 );
and ( n1397 , n859 , n67 );
nor ( n1398 , n422 , n67 );
and ( n1399 , n1398 , n398 );
nor ( n1400 , n1397 , n1399 );
nand ( n1401 , n1396 , n1400 );
nand ( n1402 , n834 , n1006 );
xor ( n1403 , n1003 , n1402 );
nand ( n1404 , n1403 , n862 );
nand ( n1405 , n915 , n91 );
and ( n1406 , n993 , n833 );
and ( n1407 , n927 , n92 );
nor ( n1408 , n1406 , n1407 );
and ( n1409 , n693 , n509 );
not ( n1410 , n693 );
and ( n1411 , n1410 , n1145 );
nor ( n1412 , n1409 , n1411 );
nand ( n1413 , n1412 , n728 );
nand ( n1414 , n1404 , n1405 , n1408 , n1413 );
and ( n1415 , n1163 , n1127 );
not ( n1416 , n1163 );
and ( n1417 , n1416 , n1292 );
nor ( n1418 , n1415 , n1417 );
nor ( n1419 , n1418 , n967 );
not ( n1420 , n34 );
not ( n1421 , n915 );
or ( n1422 , n1420 , n1421 );
and ( n1423 , n993 , n1125 );
and ( n1424 , n927 , n68 );
nor ( n1425 , n1423 , n1424 );
nand ( n1426 , n1422 , n1425 );
nor ( n1427 , n1419 , n1426 );
not ( n1428 , n861 );
xor ( n1429 , n1044 , n1043 );
not ( n1430 , n1429 );
or ( n1431 , n1428 , n1430 );
not ( n1432 , n629 );
not ( n1433 , n1432 );
and ( n1434 , n39 , n562 );
not ( n1435 , n39 );
and ( n1436 , n1435 , n561 );
nor ( n1437 , n1434 , n1436 );
not ( n1438 , n1437 );
nand ( n1439 , n42 , n556 );
nand ( n1440 , n1439 , n622 );
not ( n1441 , n1440 );
or ( n1442 , n1438 , n1441 );
nand ( n1443 , n562 , n39 );
nand ( n1444 , n1442 , n1443 );
not ( n1445 , n1444 );
or ( n1446 , n1433 , n1445 );
or ( n1447 , n1444 , n1432 );
nand ( n1448 , n1446 , n1447 );
and ( n1449 , n1448 , n923 );
and ( n1450 , n917 , n537 );
nor ( n1451 , n1449 , n1450 );
nand ( n1452 , n1431 , n1451 );
nand ( n1453 , n988 , n912 );
nand ( n1454 , n1452 , n1453 );
nand ( n1455 , n73 , n915 );
nand ( n1456 , n927 , n74 );
nand ( n1457 , n1454 , n1455 , n1456 );
xor ( n1458 , n1093 , n653 );
and ( n1459 , n859 , n1458 );
not ( n1460 , n859 );
not ( n1461 , n1082 );
not ( n1462 , n61 );
not ( n1463 , n652 );
or ( n1464 , n1462 , n1463 );
or ( n1465 , n652 , n61 );
nand ( n1466 , n1464 , n1465 );
and ( n1467 , n1461 , n1466 );
not ( n1468 , n1461 );
not ( n1469 , n1466 );
and ( n1470 , n1468 , n1469 );
nor ( n1471 , n1467 , n1470 );
and ( n1472 , n1460 , n1471 );
nor ( n1473 , n1459 , n1472 );
or ( n1474 , n1473 , n477 );
and ( n1475 , n915 , n93 );
not ( n1476 , n94 );
not ( n1477 , n927 );
or ( n1478 , n1476 , n1477 );
buf ( n1479 , n918 );
not ( n1480 , n1479 );
or ( n1481 , n1480 , n652 );
nand ( n1482 , n1478 , n1481 );
nor ( n1483 , n1475 , n1482 );
nand ( n1484 , n1474 , n1483 );
not ( n1485 , n402 );
not ( n1486 , n1395 );
nand ( n1487 , n1485 , n1389 , n1486 );
or ( n1488 , n278 , n326 );
nand ( n1489 , n1488 , n328 , n319 );
or ( n1490 , n279 , n1489 );
not ( n1491 , n315 );
nand ( n1492 , n1490 , n1491 );
not ( n1493 , n307 );
nand ( n1494 , n1493 , n322 );
and ( n1495 , n367 , n1494 );
nor ( n1496 , n1495 , n298 );
not ( n1497 , n379 );
nand ( n1498 , n1497 , n372 , n357 );
or ( n1499 , n1496 , n1498 );
not ( n1500 , n296 );
not ( n1501 , n379 );
and ( n1502 , n1500 , n1501 );
nor ( n1503 , n1502 , n308 );
nand ( n1504 , n1499 , n1503 );
and ( n1505 , n1492 , n1504 );
not ( n1506 , n332 );
nor ( n1507 , n1505 , n1506 );
not ( n1508 , n383 );
and ( n1509 , n334 , n1508 );
nor ( n1510 , n1509 , n290 );
or ( n1511 , n1507 , n1510 );
not ( n1512 , n402 );
nand ( n1513 , n1512 , n390 );
and ( n1514 , n1486 , n239 , n1513 );
nand ( n1515 , n1511 , n1514 );
nand ( n1516 , n908 , n67 );
not ( n1517 , n338 );
or ( n1518 , n1517 , n286 );
not ( n1519 , n340 );
or ( n1520 , n1519 , n280 );
nand ( n1521 , n1518 , n1520 , n354 );
and ( n1522 , n1514 , n1521 );
nand ( n1523 , n392 , n345 );
and ( n1524 , n1513 , n1523 , n237 );
and ( n1525 , n1486 , n1524 );
and ( n1526 , n1398 , n389 );
nor ( n1527 , n1522 , n1525 , n1526 );
nand ( n1528 , n1487 , n1515 , n1516 , n1527 );
not ( n1529 , n1479 );
not ( n1530 , n966 );
not ( n1531 , n38 );
and ( n1532 , n1530 , n1531 );
not ( n1533 , n54 );
and ( n1534 , n861 , n1533 );
nor ( n1535 , n1532 , n1534 );
nand ( n1536 , n1529 , n1535 );
nand ( n1537 , n1536 , n20 );
nand ( n1538 , n915 , n103 );
and ( n1539 , n927 , n104 );
not ( n1540 , n966 );
not ( n1541 , n38 );
not ( n1542 , n1541 );
and ( n1543 , n1540 , n1542 );
and ( n1544 , n861 , n54 );
nor ( n1545 , n1543 , n1544 );
nor ( n1546 , n1545 , n20 );
nor ( n1547 , n1539 , n1546 );
nand ( n1548 , n1537 , n1538 , n1547 );
buf ( n1549 , n993 );
not ( n1550 , n1549 );
buf ( n1551 , n781 );
not ( n1552 , n1551 );
or ( n1553 , n1550 , n1552 );
nor ( n1554 , n1453 , n913 );
nand ( n1555 , n1554 , n107 );
and ( n1556 , n57 , n1552 );
not ( n1557 , n57 );
and ( n1558 , n1557 , n1551 );
nor ( n1559 , n1556 , n1558 );
not ( n1560 , n1559 );
nand ( n1561 , n773 , n777 );
not ( n1562 , n1561 );
or ( n1563 , n1560 , n1562 );
or ( n1564 , n1561 , n1559 );
nand ( n1565 , n1563 , n1564 );
and ( n1566 , n861 , n1565 );
and ( n1567 , n927 , n108 );
xor ( n1568 , n41 , n1551 );
xor ( n1569 , n1568 , n611 );
and ( n1570 , n1569 , n726 );
nor ( n1571 , n1566 , n1567 , n1570 );
nand ( n1572 , n1553 , n1555 , n1571 );
or ( n1573 , n1550 , n578 );
nand ( n1574 , n1554 , n109 );
buf ( n1575 , n772 );
not ( n1576 , n1575 );
not ( n1577 , n766 );
or ( n1578 , n1576 , n1577 );
or ( n1579 , n1575 , n766 );
nand ( n1580 , n1578 , n1579 );
and ( n1581 , n861 , n1580 );
and ( n1582 , n913 , n110 );
not ( n1583 , n609 );
not ( n1584 , n1583 );
not ( n1585 , n593 );
or ( n1586 , n1584 , n1585 );
or ( n1587 , n593 , n1583 );
nand ( n1588 , n1586 , n1587 );
and ( n1589 , n726 , n1588 );
nor ( n1590 , n1581 , n1582 , n1589 );
nand ( n1591 , n1573 , n1574 , n1590 );
not ( n1592 , n607 );
or ( n1593 , n1550 , n1592 );
nand ( n1594 , n1554 , n111 );
not ( n1595 , n760 );
not ( n1596 , n52 );
not ( n1597 , n1592 );
or ( n1598 , n1596 , n1597 );
or ( n1599 , n1592 , n52 );
nand ( n1600 , n1598 , n1599 );
not ( n1601 , n1600 );
or ( n1602 , n1595 , n1601 );
or ( n1603 , n1600 , n760 );
nand ( n1604 , n1602 , n1603 );
and ( n1605 , n861 , n1604 );
and ( n1606 , n927 , n112 );
xor ( n1607 , n599 , n594 );
and ( n1608 , n726 , n1607 );
nor ( n1609 , n1605 , n1606 , n1608 );
nand ( n1610 , n1593 , n1594 , n1609 );
nand ( n1611 , n237 , n392 );
and ( n1612 , n1387 , n1611 );
nor ( n1613 , n1387 , n1611 );
nor ( n1614 , n1612 , n1613 );
or ( n1615 , n1614 , n1395 );
not ( n1616 , n873 );
or ( n1617 , n913 , n1616 );
not ( n1618 , n1398 );
or ( n1619 , n236 , n1618 );
nand ( n1620 , n1615 , n1617 , n1619 );
not ( n1621 , n105 );
not ( n1622 , n915 );
or ( n1623 , n1621 , n1622 );
not ( n1624 , n556 );
not ( n1625 , n1479 );
or ( n1626 , n1624 , n1625 );
not ( n1627 , n621 );
not ( n1628 , n1627 );
not ( n1629 , n615 );
not ( n1630 , n1629 );
or ( n1631 , n1628 , n1630 );
or ( n1632 , n1629 , n1627 );
nand ( n1633 , n1631 , n1632 );
nand ( n1634 , n923 , n1633 );
nand ( n1635 , n1626 , n1634 );
xor ( n1636 , n783 , n758 );
not ( n1637 , n1636 );
not ( n1638 , n861 );
or ( n1639 , n1637 , n1638 );
nand ( n1640 , n927 , n106 );
nand ( n1641 , n1639 , n1640 );
nor ( n1642 , n1635 , n1641 );
nand ( n1643 , n1623 , n1642 );
not ( n1644 , n77 );
not ( n1645 , n915 );
or ( n1646 , n1644 , n1645 );
not ( n1647 , n562 );
not ( n1648 , n993 );
or ( n1649 , n1647 , n1648 );
xor ( n1650 , n1440 , n1437 );
nand ( n1651 , n727 , n1650 );
nand ( n1652 , n1649 , n1651 );
xor ( n1653 , n1040 , n1032 );
not ( n1654 , n1653 );
not ( n1655 , n861 );
or ( n1656 , n1654 , n1655 );
nand ( n1657 , n927 , n78 );
nand ( n1658 , n1656 , n1657 );
nor ( n1659 , n1652 , n1658 );
nand ( n1660 , n1646 , n1659 );
not ( n1661 , n44 );
and ( n1662 , n32 , n465 );
not ( n1663 , n32 );
and ( n1664 , n1663 , n433 );
nor ( n1665 , n1662 , n1664 );
not ( n1666 , n1665 );
or ( n1667 , n1661 , n1666 );
and ( n1668 , n94 , n106 , n100 , n108 );
nand ( n1669 , n1668 , n74 , n78 );
and ( n1670 , n1669 , n88 );
nor ( n1671 , n1669 , n88 );
nor ( n1672 , n1670 , n1671 );
or ( n1673 , n1665 , n1672 );
nand ( n1674 , n1667 , n1673 );
and ( n1675 , n33 , n433 );
not ( n1676 , n33 );
and ( n1677 , n1676 , n465 );
nor ( n1678 , n1675 , n1677 );
and ( n1679 , n1674 , n1678 );
nand ( n1680 , n1665 , n114 );
not ( n1681 , n1665 );
nand ( n1682 , n1681 , n60 );
and ( n1683 , n1680 , n1682 );
nor ( n1684 , n1683 , n1678 );
nor ( n1685 , n1679 , n1684 );
not ( n1686 , n909 );
nand ( n1687 , n1686 , n67 );
or ( n1688 , n1685 , n1687 );
nand ( n1689 , n1687 , n235 , n113 );
nand ( n1690 , n1688 , n1689 );
and ( n1691 , n51 , n1122 );
not ( n1692 , n51 );
and ( n1693 , n1692 , n1125 );
nor ( n1694 , n1691 , n1693 );
xor ( n1695 , n1311 , n1694 );
not ( n1696 , n1695 );
not ( n1697 , n862 );
or ( n1698 , n1696 , n1697 );
nand ( n1699 , n1698 , n1427 );
endmodule

