//NOTE: no-implementation module stub

module mfa (
    input  wire S,
    input  wire C,
    input  wire P,
    output wire Q,
    output wire R
);

endmodule
