module pipeKuz(
    input [127:0] block,
    input [255:0] key,
    input clk,
    output reg [127:0] enc);

  reg [127:0] key3; reg [127:0] key4; reg [127:0] key5; reg [127:0] key6;
  reg [127:0] key7; reg [127:0] key8; reg [127:0] key9; reg [127:0] key10;
  
  //-------------------------------------------------------------------------------------------------------------------------------------------//
  // TABLES AND CONSTS
  //-------------------------------------------------------------------------------------------------------------------------------------------//
  
  // S BLOCK
  reg [7:0] sTab [255:0];
  `define C(ind, val) assign sTab[ind] = 8'd``val
    `C(0, 252); `C(1, 238); `C(2, 221); `C(3, 17); `C(4, 207); `C(5, 110); `C(6, 49);  `C(7, 22); `C(8, 251); `C(9, 196); `C(10, 250); `C(11, 218);
    `C(12, 35); `C(13, 197); `C(14, 4); `C(15, 77); `C(16, 233); `C(17, 119); `C(18, 240); `C(19, 219); `C(20, 147); `C(21, 46); `C(22, 153); `C(23, 186);
    `C(24, 23); `C(25, 54); `C(26, 241); `C(27, 187); `C(28, 20); `C(29, 205); `C(30, 95); `C(31, 193); `C(32, 249); `C(33, 24); `C(34, 101); `C(35, 90);
    `C(36, 226); `C(37, 92); `C(38, 239); `C(39, 33); `C(40, 129); `C(41, 28); `C(42, 60); `C(43, 66); `C(44, 139); `C(45, 1); `C(46, 142); `C(47, 79);
    `C(48, 5); `C(49, 132); `C(50, 2); `C(51, 174); `C(52, 227); `C(53, 106); `C(54, 143); `C(55, 160); `C(56, 6); `C(57, 11); `C(58, 237); `C(59, 152);
    `C(60, 127); `C(61, 212); `C(62, 211); `C(63, 31); `C(64, 235); `C(65, 52); `C(66, 44); `C(67, 81); `C(68, 234); `C(69, 200); `C(70, 72); `C(71, 171);
    `C(72, 242); `C(73, 42); `C(74, 104); `C(75, 162); `C(76, 253); `C(77, 58); `C(78, 206); `C(79, 204); `C(80, 181); `C(81, 112); `C(82, 14); `C(83, 86);
    `C(84, 8);  `C(85, 12); `C(86, 118); `C(87, 18); `C(88, 191); `C(89, 114); `C(90, 19); `C(91, 71); `C(92, 156); `C(93, 183); `C(94, 93); `C(95, 135);
    `C(96, 21); `C(97, 161); `C(98, 150); `C(99, 41); `C(100, 16); `C(101, 123); `C(102, 154); `C(103, 199); `C(104, 243); `C(105, 145); `C(106, 120);
    `C(107, 111); `C(108, 157); `C(109, 158); `C(110, 178); `C(111, 177); `C(112, 50); `C(113, 117); `C(114, 25); `C(115, 61); `C(116, 255);
    `C(117, 53); `C(118, 138); `C(119, 126); `C(120, 109); `C(121, 84); `C(122, 198); `C(123, 128); `C(124, 195); `C(125, 189); `C(126, 13);
    `C(127, 87); `C(128, 223); `C(129, 245); `C(130, 36); `C(131, 169); `C(132, 62); `C(133, 168); `C(134, 67); `C(135, 201); `C(136, 215);
    `C(137, 121); `C(138, 214); `C(139, 246); `C(140, 124); `C(141, 34); `C(142, 185); `C(143, 3); `C(144, 224); `C(145, 15); `C(146, 236);
    `C(147, 222); `C(148, 122); `C(149, 148); `C(150, 176); `C(151, 188); `C(152, 220); `C(153, 232); `C(154, 40); `C(155, 80); `C(156, 78);
    `C(157, 51); `C(158, 10); `C(159, 74); `C(160, 167); `C(161, 151); `C(162, 96); `C(163, 115); `C(164, 30); `C(165, 0); `C(166, 98);
    `C(167, 68); `C(168, 26); `C(169, 184); `C(170, 56); `C(171, 130); `C(172, 100); `C(173, 159); `C(174, 38); `C(175, 65); `C(176, 173);
    `C(177, 69); `C(178, 70); `C(179, 146); `C(180, 39); `C(181, 94); `C(182, 85); `C(183, 47); `C(184, 140); `C(185, 163); `C(186, 165);
    `C(187, 125); `C(188, 105); `C(189, 213); `C(190, 149); `C(191, 59); `C(192, 7); `C(193, 88); `C(194, 179); `C(195, 64); `C(196, 134);
    `C(197, 172); `C(198, 29); `C(199, 247); `C(200, 48); `C(201, 55); `C(202, 107); `C(203, 228); `C(204, 136); `C(205, 217); `C(206, 231);
    `C(207, 137); `C(208, 225); `C(209, 27); `C(210, 131); `C(211, 73); `C(212, 76); `C(213, 63); `C(214, 248); `C(215, 254); `C(216, 141);
    `C(217, 83); `C(218, 170); `C(219, 144); `C(220, 202); `C(221, 216); `C(222, 133); `C(223, 97); `C(224, 32); `C(225, 113); `C(226, 103);
    `C(227, 164); `C(228, 45); `C(229, 43); `C(230, 9); `C(231, 91); `C(232, 203); `C(233, 155); `C(234, 37); `C(235, 208); `C(236, 190);
    `C(237, 229); `C(238, 108); `C(239, 82); `C(240, 89); `C(241, 166); `C(242, 116); `C(243, 210); `C(244, 230); `C(245, 244); `C(246, 180);
    `C(247, 192); `C(248, 209); `C(249, 102); `C(250, 175); `C(251, 194); `C(252, 57); `C(253, 75); `C(254, 99); `C(255, 182);
  
  function automatic [127:0] sBlock;
    input [127:0] in;
    begin
      sBlock[7:0] = sTab[in[7:0]]; sBlock[15:8] = sTab[in[15:8]]; sBlock[23:16] = sTab[in[23:16]]; sBlock[31:24] = sTab[in[31:24]];
      sBlock[39:32] = sTab[in[39:32]]; sBlock[47:40] = sTab[in[47:40]]; sBlock[55:48] = sTab[in[55:48]]; sBlock[63:56] = sTab[in[63:56]];
      sBlock[71:64] = sTab[in[71:64]]; sBlock[79:72] = sTab[in[79:72]]; sBlock[87:80] = sTab[in[87:80]]; sBlock[95:88] = sTab[in[95:88]];
      sBlock[103:96] = sTab[in[103:96]]; sBlock[111:104] = sTab[in[111:104]]; sBlock[119:112] = sTab[in[119:112]]; sBlock[127:120] = sTab[in[127:120]];
    end
  endfunction
  
  // L BLOCK
  `define LC(name, ind, val) assign name[ind] = 8'd``val
  reg [7:0] l94 [255:0]; reg [7:0] l20 [255:0]; reg [7:0] l85 [255:0]; reg [7:0] l10 [255:0];
  reg [7:0] lC2 [255:0]; reg [7:0] lC0 [255:0]; reg [7:0] lFB [255:0];
    `LC(l94, 0, 0); `LC(l94, 1, 148); `LC(l94, 2, 235); `LC(l94, 3, 127); `LC(l94, 4, 21); `LC(l94, 5, 129); `LC(l94, 6, 254); `LC(l94, 7, 106); `LC(l94, 8, 42); `LC(l94, 9, 190);
    `LC(l94, 10, 193); `LC(l94, 11, 85); `LC(l94, 12, 63); `LC(l94, 13, 171); `LC(l94, 14, 212); `LC(l94, 15, 64); `LC(l94, 16, 84); `LC(l94, 17, 192); `LC(l94, 18, 191);
    `LC(l94, 19, 43); `LC(l94, 20, 65); `LC(l94, 21, 213); `LC(l94, 22, 170); `LC(l94, 23, 62); `LC(l94, 24, 126); `LC(l94, 25, 234); `LC(l94, 26, 149); `LC(l94, 27, 1);
    `LC(l94, 28, 107); `LC(l94, 29, 255); `LC(l94, 30, 128); `LC(l94, 31, 20); `LC(l94, 32, 168); `LC(l94, 33, 60); `LC(l94, 34, 67); `LC(l94, 35, 215); `LC(l94, 36, 189);
    `LC(l94, 37, 41); `LC(l94, 38, 86); `LC(l94, 39, 194); `LC(l94, 40, 130); `LC(l94, 41, 22); `LC(l94, 42, 105); `LC(l94, 43, 253); `LC(l94, 44, 151); `LC(l94, 45, 3);
    `LC(l94, 46, 124); `LC(l94, 47, 232); `LC(l94, 48, 252); `LC(l94, 49, 104); `LC(l94, 50, 23); `LC(l94, 51, 131); `LC(l94, 52, 233); `LC(l94, 53, 125); `LC(l94, 54, 2);
    `LC(l94, 55, 150); `LC(l94, 56, 214); `LC(l94, 57, 66); `LC(l94, 58, 61); `LC(l94, 59, 169); `LC(l94, 60, 195); `LC(l94, 61, 87); `LC(l94, 62, 40); `LC(l94, 63, 188);
    `LC(l94, 64, 147); `LC(l94, 65, 7); `LC(l94, 66, 120); `LC(l94, 67, 236); `LC(l94, 68, 134); `LC(l94, 69, 18); `LC(l94, 70, 109); `LC(l94, 71, 249); `LC(l94, 72, 185);
    `LC(l94, 73, 45); `LC(l94, 74, 82); `LC(l94, 75, 198); `LC(l94, 76, 172); `LC(l94, 77, 56); `LC(l94, 78, 71); `LC(l94, 79, 211); `LC(l94, 80, 199); `LC(l94, 81, 83);
    `LC(l94, 82, 44); `LC(l94, 83, 184); `LC(l94, 84, 210); `LC(l94, 85, 70); `LC(l94, 86, 57); `LC(l94, 87, 173); `LC(l94, 88, 237); `LC(l94, 89, 121); `LC(l94, 90, 6);
    `LC(l94, 91, 146); `LC(l94, 92, 248); `LC(l94, 93, 108); `LC(l94, 94, 19); `LC(l94, 95, 135); `LC(l94, 96, 59); `LC(l94, 97, 175); `LC(l94, 98, 208); `LC(l94, 99, 68);
    `LC(l94, 100, 46); `LC(l94, 101, 186); `LC(l94, 102, 197); `LC(l94, 103, 81); `LC(l94, 104, 17); `LC(l94, 105, 133); `LC(l94, 106, 250); `LC(l94, 107, 110); `LC(l94, 108, 4);
    `LC(l94, 109, 144); `LC(l94, 110, 239); `LC(l94, 111, 123); `LC(l94, 112, 111); `LC(l94, 113, 251); `LC(l94, 114, 132); `LC(l94, 115, 16); `LC(l94, 116, 122); `LC(l94, 117, 238);
    `LC(l94, 118, 145); `LC(l94, 119, 5); `LC(l94, 120, 69); `LC(l94, 121, 209); `LC(l94, 122, 174); `LC(l94, 123, 58); `LC(l94, 124, 80); `LC(l94, 125, 196); `LC(l94, 126, 187);
    `LC(l94, 127, 47); `LC(l94, 128, 229); `LC(l94, 129, 113); `LC(l94, 130, 14); `LC(l94, 131, 154); `LC(l94, 132, 240); `LC(l94, 133, 100); `LC(l94, 134, 27); `LC(l94, 135, 143);
    `LC(l94, 136, 207); `LC(l94, 137, 91); `LC(l94, 138, 36); `LC(l94, 139, 176); `LC(l94, 140, 218); `LC(l94, 141, 78); `LC(l94, 142, 49); `LC(l94, 143, 165); `LC(l94, 144, 177);
    `LC(l94, 145, 37); `LC(l94, 146, 90); `LC(l94, 147, 206); `LC(l94, 148, 164); `LC(l94, 149, 48); `LC(l94, 150, 79); `LC(l94, 151, 219); `LC(l94, 152, 155); `LC(l94, 153, 15);
    `LC(l94, 154, 112); `LC(l94, 155, 228); `LC(l94, 156, 142); `LC(l94, 157, 26); `LC(l94, 158, 101); `LC(l94, 159, 241); `LC(l94, 160, 77); `LC(l94, 161, 217); `LC(l94, 162, 166);
    `LC(l94, 163, 50); `LC(l94, 164, 88); `LC(l94, 165, 204); `LC(l94, 166, 179); `LC(l94, 167, 39); `LC(l94, 168, 103); `LC(l94, 169, 243); `LC(l94, 170, 140); `LC(l94, 171, 24);
    `LC(l94, 172, 114); `LC(l94, 173, 230); `LC(l94, 174, 153); `LC(l94, 175, 13); `LC(l94, 176, 25); `LC(l94, 177, 141); `LC(l94, 178, 242); `LC(l94, 179, 102); `LC(l94, 180, 12);
    `LC(l94, 181, 152); `LC(l94, 182, 231); `LC(l94, 183, 115); `LC(l94, 184, 51); `LC(l94, 185, 167); `LC(l94, 186, 216); `LC(l94, 187, 76); `LC(l94, 188, 38); `LC(l94, 189, 178);
    `LC(l94, 190, 205); `LC(l94, 191, 89); `LC(l94, 192, 118); `LC(l94, 193, 226); `LC(l94, 194, 157); `LC(l94, 195, 9); `LC(l94, 196, 99); `LC(l94, 197, 247); `LC(l94, 198, 136);
    `LC(l94, 199, 28); `LC(l94, 200, 92); `LC(l94, 201, 200); `LC(l94, 202, 183); `LC(l94, 203, 35); `LC(l94, 204, 73); `LC(l94, 205, 221); `LC(l94, 206, 162); `LC(l94, 207, 54);
    `LC(l94, 208, 34); `LC(l94, 209, 182); `LC(l94, 210, 201); `LC(l94, 211, 93); `LC(l94, 212, 55); `LC(l94, 213, 163); `LC(l94, 214, 220); `LC(l94, 215, 72); `LC(l94, 216, 8);
    `LC(l94, 217, 156); `LC(l94, 218, 227); `LC(l94, 219, 119); `LC(l94, 220, 29); `LC(l94, 221, 137); `LC(l94, 222, 246); `LC(l94, 223, 98); `LC(l94, 224, 222); `LC(l94, 225, 74);
    `LC(l94, 226, 53); `LC(l94, 227, 161); `LC(l94, 228, 203); `LC(l94, 229, 95); `LC(l94, 230, 32); `LC(l94, 231, 180); `LC(l94, 232, 244); `LC(l94, 233, 96); `LC(l94, 234, 31);
    `LC(l94, 235, 139); `LC(l94, 236, 225); `LC(l94, 237, 117); `LC(l94, 238, 10); `LC(l94, 239, 158); `LC(l94, 240, 138); `LC(l94, 241, 30); `LC(l94, 242, 97); `LC(l94, 243, 245);
    `LC(l94, 244, 159); `LC(l94, 245, 11); `LC(l94, 246, 116); `LC(l94, 247, 224); `LC(l94, 248, 160); `LC(l94, 249, 52); `LC(l94, 250, 75); `LC(l94, 251, 223); `LC(l94, 252, 181);
    `LC(l94, 253, 33); `LC(l94, 254, 94); `LC(l94, 255, 202);
    `LC(l20, 0, 0); `LC(l20, 1, 32); `LC(l20, 2, 64); `LC(l20, 3, 96); `LC(l20, 4, 128); `LC(l20, 5, 160); `LC(l20, 6, 192); `LC(l20, 7, 224); `LC(l20, 8, 195); `LC(l20, 9, 227);
    `LC(l20, 10, 131); `LC(l20, 11, 163); `LC(l20, 12, 67); `LC(l20, 13, 99); `LC(l20, 14, 3); `LC(l20, 15, 35); `LC(l20, 16, 69); `LC(l20, 17, 101); `LC(l20, 18, 5); `LC(l20, 19, 37);
    `LC(l20, 20, 197); `LC(l20, 21, 229); `LC(l20, 22, 133); `LC(l20, 23, 165); `LC(l20, 24, 134); `LC(l20, 25, 166); `LC(l20, 26, 198); `LC(l20, 27, 230); `LC(l20, 28, 6);
    `LC(l20, 29, 38); `LC(l20, 30, 70); `LC(l20, 31, 102); `LC(l20, 32, 138); `LC(l20, 33, 170); `LC(l20, 34, 202); `LC(l20, 35, 234); `LC(l20, 36, 10); `LC(l20, 37, 42);
    `LC(l20, 38, 74); `LC(l20, 39, 106); `LC(l20, 40, 73); `LC(l20, 41, 105); `LC(l20, 42, 9); `LC(l20, 43, 41); `LC(l20, 44, 201); `LC(l20, 45, 233); `LC(l20, 46, 137);
    `LC(l20, 47, 169); `LC(l20, 48, 207); `LC(l20, 49, 239); `LC(l20, 50, 143); `LC(l20, 51, 175); `LC(l20, 52, 79); `LC(l20, 53, 111); `LC(l20, 54, 15); `LC(l20, 55, 47);
    `LC(l20, 56, 12); `LC(l20, 57, 44); `LC(l20, 58, 76); `LC(l20, 59, 108); `LC(l20, 60, 140); `LC(l20, 61, 172); `LC(l20, 62, 204); `LC(l20, 63, 236); `LC(l20, 64, 215);
    `LC(l20, 65, 247); `LC(l20, 66, 151); `LC(l20, 67, 183); `LC(l20, 68, 87); `LC(l20, 69, 119); `LC(l20, 70, 23); `LC(l20, 71, 55); `LC(l20, 72, 20); `LC(l20, 73, 52);
    `LC(l20, 74, 84); `LC(l20, 75, 116); `LC(l20, 76, 148); `LC(l20, 77, 180); `LC(l20, 78, 212); `LC(l20, 79, 244); `LC(l20, 80, 146); `LC(l20, 81, 178); `LC(l20, 82, 210);
    `LC(l20, 83, 242); `LC(l20, 84, 18); `LC(l20, 85, 50); `LC(l20, 86, 82); `LC(l20, 87, 114); `LC(l20, 88, 81); `LC(l20, 89, 113); `LC(l20, 90, 17); `LC(l20, 91, 49);
    `LC(l20, 92, 209); `LC(l20, 93, 241); `LC(l20, 94, 145); `LC(l20, 95, 177); `LC(l20, 96, 93); `LC(l20, 97, 125); `LC(l20, 98, 29); `LC(l20, 99, 61); `LC(l20, 100, 221);
    `LC(l20, 101, 253); `LC(l20, 102, 157); `LC(l20, 103, 189); `LC(l20, 104, 158); `LC(l20, 105, 190); `LC(l20, 106, 222); `LC(l20, 107, 254); `LC(l20, 108, 30); `LC(l20, 109, 62);
    `LC(l20, 110, 94); `LC(l20, 111, 126); `LC(l20, 112, 24); `LC(l20, 113, 56); `LC(l20, 114, 88); `LC(l20, 115, 120); `LC(l20, 116, 152); `LC(l20, 117, 184); `LC(l20, 118, 216);
    `LC(l20, 119, 248); `LC(l20, 120, 219); `LC(l20, 121, 251); `LC(l20, 122, 155); `LC(l20, 123, 187); `LC(l20, 124, 91); `LC(l20, 125, 123); `LC(l20, 126, 27); `LC(l20, 127, 59);
    `LC(l20, 128, 109); `LC(l20, 129, 77); `LC(l20, 130, 45); `LC(l20, 131, 13); `LC(l20, 132, 237); `LC(l20, 133, 205); `LC(l20, 134, 173); `LC(l20, 135, 141);
    `LC(l20, 136, 174); `LC(l20, 137, 142); `LC(l20, 138, 238); `LC(l20, 139, 206); `LC(l20, 140, 46); `LC(l20, 141, 14); `LC(l20, 142, 110); `LC(l20, 143, 78); `LC(l20, 144, 40);
    `LC(l20, 145, 8); `LC(l20, 146, 104); `LC(l20, 147, 72); `LC(l20, 148, 168); `LC(l20, 149, 136); `LC(l20, 150, 232); `LC(l20, 151, 200); `LC(l20, 152, 235); `LC(l20, 153, 203);
    `LC(l20, 154, 171); `LC(l20, 155, 139); `LC(l20, 156, 107); `LC(l20, 157, 75); `LC(l20, 158, 43); `LC(l20, 159, 11); `LC(l20, 160, 231); `LC(l20, 161, 199); `LC(l20, 162, 167);
    `LC(l20, 163, 135); `LC(l20, 164, 103); `LC(l20, 165, 71); `LC(l20, 166, 39); `LC(l20, 167, 7); `LC(l20, 168, 36); `LC(l20, 169, 4); `LC(l20, 170, 100);
    `LC(l20, 171, 68); `LC(l20, 172, 164); `LC(l20, 173, 132); `LC(l20, 174, 228); `LC(l20, 175, 196); `LC(l20, 176, 162); `LC(l20, 177, 130); `LC(l20, 178, 226); `LC(l20, 179, 194);
    `LC(l20, 180, 34); `LC(l20, 181, 2); `LC(l20, 182, 98); `LC(l20, 183, 66); `LC(l20, 184, 97); `LC(l20, 185, 65); `LC(l20, 186, 33); `LC(l20, 187, 1); `LC(l20, 188, 225);
    `LC(l20, 189, 193); `LC(l20, 190, 161); `LC(l20, 191, 129); `LC(l20, 192, 186); `LC(l20, 193, 154); `LC(l20, 194, 250); `LC(l20, 195, 218); `LC(l20, 196, 58); `LC(l20, 197, 26);
    `LC(l20, 198, 122); `LC(l20, 199, 90); `LC(l20, 200, 121); `LC(l20, 201, 89); `LC(l20, 202, 57); `LC(l20, 203, 25); `LC(l20, 204, 249); `LC(l20, 205, 217);
    `LC(l20, 206, 185); `LC(l20, 207, 153); `LC(l20, 208, 255); `LC(l20, 209, 223); `LC(l20, 210, 191); `LC(l20, 211, 159); `LC(l20, 212, 127); `LC(l20, 213, 95); `LC(l20, 214, 63);
    `LC(l20, 215, 31); `LC(l20, 216, 60); `LC(l20, 217, 28); `LC(l20, 218, 124); `LC(l20, 219, 92); `LC(l20, 220, 188); `LC(l20, 221, 156); `LC(l20, 222, 252); `LC(l20, 223, 220);
    `LC(l20, 224, 48); `LC(l20, 225, 16); `LC(l20, 226, 112); `LC(l20, 227, 80); `LC(l20, 228, 176); `LC(l20, 229, 144); `LC(l20, 230, 240);
    `LC(l20, 231, 208); `LC(l20, 232, 243); `LC(l20, 233, 211); `LC(l20, 234, 179); `LC(l20, 235, 147); `LC(l20, 236, 115); `LC(l20, 237, 83); `LC(l20, 238, 51); `LC(l20, 239, 19);
    `LC(l20, 240, 117); `LC(l20, 241, 85); `LC(l20, 242, 53); `LC(l20, 243, 21); `LC(l20, 244, 245); `LC(l20, 245, 213); `LC(l20, 246, 181); `LC(l20, 247, 149); `LC(l20, 248, 182);
    `LC(l20, 249, 150); `LC(l20, 250, 246); `LC(l20, 251, 214); `LC(l20, 252, 54); `LC(l20, 253, 22); `LC(l20, 254, 118); `LC(l20, 255, 86);
    `LC(l85, 0, 0); `LC(l85, 1, 133); `LC(l85, 2, 201); `LC(l85, 3, 76); `LC(l85, 4, 81); `LC(l85, 5, 212); `LC(l85, 6, 152); `LC(l85, 7, 29); `LC(l85, 8, 162); `LC(l85, 9, 39);
    `LC(l85, 10, 107); `LC(l85, 11, 238); `LC(l85, 12, 243); `LC(l85, 13, 118); `LC(l85, 14, 58); `LC(l85, 15, 191); `LC(l85, 16, 135); `LC(l85, 17, 2); `LC(l85, 18, 78);
    `LC(l85, 19, 203); `LC(l85, 20, 214); `LC(l85, 21, 83); `LC(l85, 22, 31); `LC(l85, 23, 154); `LC(l85, 24, 37); `LC(l85, 25, 160); `LC(l85, 26, 236); `LC(l85, 27, 105);
    `LC(l85, 28, 116); `LC(l85, 29, 241); `LC(l85, 30, 189); `LC(l85, 31, 56); `LC(l85, 32, 205); `LC(l85, 33, 72); `LC(l85, 34, 4); `LC(l85, 35, 129); `LC(l85, 36, 156);
    `LC(l85, 37, 25); `LC(l85, 38, 85); `LC(l85, 39, 208); `LC(l85, 40, 111); `LC(l85, 41, 234); `LC(l85, 42, 166); `LC(l85, 43, 35); `LC(l85, 44, 62); `LC(l85, 45, 187);
    `LC(l85, 46, 247); `LC(l85, 47, 114); `LC(l85, 48, 74); `LC(l85, 49, 207); `LC(l85, 50, 131); `LC(l85, 51, 6); `LC(l85, 52, 27); `LC(l85, 53, 158); `LC(l85, 54, 210);
    `LC(l85, 55, 87); `LC(l85, 56, 232); `LC(l85, 57, 109); `LC(l85, 58, 33); `LC(l85, 59, 164); `LC(l85, 60, 185); `LC(l85, 61, 60); `LC(l85, 62, 112); `LC(l85, 63, 245);
    `LC(l85, 64, 89); `LC(l85, 65, 220); `LC(l85, 66, 144); `LC(l85, 67, 21); `LC(l85, 68, 8); `LC(l85, 69, 141); `LC(l85, 70, 193); `LC(l85, 71, 68); `LC(l85, 72, 251);
    `LC(l85, 73, 126); `LC(l85, 74, 50); `LC(l85, 75, 183); `LC(l85, 76, 170); `LC(l85, 77, 47); `LC(l85, 78, 99); `LC(l85, 79, 230); `LC(l85, 80, 222); `LC(l85, 81, 91);
    `LC(l85, 82, 23); `LC(l85, 83, 146); `LC(l85, 84, 143); `LC(l85, 85, 10); `LC(l85, 86, 70); `LC(l85, 87, 195); `LC(l85, 88, 124); `LC(l85, 89, 249); `LC(l85, 90, 181);
    `LC(l85, 91, 48); `LC(l85, 92, 45); `LC(l85, 93, 168); `LC(l85, 94, 228); `LC(l85, 95, 97); `LC(l85, 96, 148); `LC(l85, 97, 17); `LC(l85, 98, 93); `LC(l85, 99, 216);
    `LC(l85, 100, 197); `LC(l85, 101, 64); `LC(l85, 102, 12); `LC(l85, 103, 137); `LC(l85, 104, 54); `LC(l85, 105, 179); `LC(l85, 106, 255); `LC(l85, 107, 122); `LC(l85, 108, 103);
    `LC(l85, 109, 226); `LC(l85, 110, 174); `LC(l85, 111, 43); `LC(l85, 112, 19); `LC(l85, 113, 150); `LC(l85, 114, 218); `LC(l85, 115, 95); `LC(l85, 116, 66); `LC(l85, 117, 199);
    `LC(l85, 118, 139); `LC(l85, 119, 14); `LC(l85, 120, 177); `LC(l85, 121, 52); `LC(l85, 122, 120); `LC(l85, 123, 253); `LC(l85, 124, 224); `LC(l85, 125, 101); `LC(l85, 126, 41);
    `LC(l85, 127, 172); `LC(l85, 128, 178); `LC(l85, 129, 55); `LC(l85, 130, 123); `LC(l85, 131, 254); `LC(l85, 132, 227); `LC(l85, 133, 102); `LC(l85, 134, 42); `LC(l85, 135, 175);
    `LC(l85, 136, 16); `LC(l85, 137, 149); `LC(l85, 138, 217); `LC(l85, 139, 92); `LC(l85, 140, 65); `LC(l85, 141, 196); `LC(l85, 142, 136); `LC(l85, 143, 13); `LC(l85, 144, 53);
    `LC(l85, 145, 176); `LC(l85, 146, 252); `LC(l85, 147, 121); `LC(l85, 148, 100); `LC(l85, 149, 225); `LC(l85, 150, 173); `LC(l85, 151, 40); `LC(l85, 152, 151); `LC(l85, 153, 18);
    `LC(l85, 154, 94); `LC(l85, 155, 219); `LC(l85, 156, 198); `LC(l85, 157, 67); `LC(l85, 158, 15); `LC(l85, 159, 138); `LC(l85, 160, 127); `LC(l85, 161, 250); `LC(l85, 162, 182);
    `LC(l85, 163, 51); `LC(l85, 164, 46); `LC(l85, 165, 171); `LC(l85, 166, 231); `LC(l85, 167, 98); `LC(l85, 168, 221); `LC(l85, 169, 88); `LC(l85, 170, 20); `LC(l85, 171, 145);
    `LC(l85, 172, 140); `LC(l85, 173, 9); `LC(l85, 174, 69); `LC(l85, 175, 192); `LC(l85, 176, 248); `LC(l85, 177, 125); `LC(l85, 178, 49); `LC(l85, 179, 180); `LC(l85, 180, 169);
    `LC(l85, 181, 44); `LC(l85, 182, 96); `LC(l85, 183, 229); `LC(l85, 184, 90); `LC(l85, 185, 223); `LC(l85, 186, 147); `LC(l85, 187, 22); `LC(l85, 188, 11); `LC(l85, 189, 142);
    `LC(l85, 190, 194); `LC(l85, 191, 71); `LC(l85, 192, 235); `LC(l85, 193, 110); `LC(l85, 194, 34); `LC(l85, 195, 167); `LC(l85, 196, 186); `LC(l85, 197, 63); `LC(l85, 198, 115);
    `LC(l85, 199, 246); `LC(l85, 200, 73); `LC(l85, 201, 204); `LC(l85, 202, 128); `LC(l85, 203, 5); `LC(l85, 204, 24); `LC(l85, 205, 157); `LC(l85, 206, 209); `LC(l85, 207, 84);
    `LC(l85, 208, 108); `LC(l85, 209, 233); `LC(l85, 210, 165); `LC(l85, 211, 32); `LC(l85, 212, 61); `LC(l85, 213, 184); `LC(l85, 214, 244); `LC(l85, 215, 113); `LC(l85, 216, 206);
    `LC(l85, 217, 75); `LC(l85, 218, 7); `LC(l85, 219, 130); `LC(l85, 220, 159); `LC(l85, 221, 26); `LC(l85, 222, 86); `LC(l85, 223, 211); `LC(l85, 224, 38); `LC(l85, 225, 163);
    `LC(l85, 226, 239); `LC(l85, 227, 106); `LC(l85, 228, 119); `LC(l85, 229, 242); `LC(l85, 230, 190); `LC(l85, 231, 59); `LC(l85, 232, 132); `LC(l85, 233, 1); `LC(l85, 234, 77);
    `LC(l85, 235, 200); `LC(l85, 236, 213); `LC(l85, 237, 80); `LC(l85, 238, 28); `LC(l85, 239, 153); `LC(l85, 240, 161); `LC(l85, 241, 36); `LC(l85, 242, 104); `LC(l85, 243, 237);
    `LC(l85, 244, 240); `LC(l85, 245, 117); `LC(l85, 246, 57); `LC(l85, 247, 188); `LC(l85, 248, 3); `LC(l85, 249, 134); `LC(l85, 250, 202);
    `LC(l85, 251, 79); `LC(l85, 252, 82); `LC(l85, 253, 215); `LC(l85, 254, 155); `LC(l85, 255, 30);
    `LC(l10, 0, 0); `LC(l10, 1, 16); `LC(l10, 2, 32); `LC(l10, 3, 48); `LC(l10, 4, 64); `LC(l10, 5, 80); `LC(l10, 6, 96); `LC(l10, 7, 112); `LC(l10, 8, 128); `LC(l10, 9, 144);
    `LC(l10, 10, 160); `LC(l10, 11, 176); `LC(l10, 12, 192); `LC(l10, 13, 208); `LC(l10, 14, 224); `LC(l10, 15, 240); `LC(l10, 16, 195); `LC(l10, 17, 211); `LC(l10, 18, 227);
    `LC(l10, 19, 243); `LC(l10, 20, 131); `LC(l10, 21, 147); `LC(l10, 22, 163); `LC(l10, 23, 179); `LC(l10, 24, 67); `LC(l10, 25, 83); `LC(l10, 26, 99); `LC(l10, 27, 115);
    `LC(l10, 28, 3); `LC(l10, 29, 19); `LC(l10, 30, 35); `LC(l10, 31, 51); `LC(l10, 32, 69); `LC(l10, 33, 85); `LC(l10, 34, 101); `LC(l10, 35, 117); `LC(l10, 36, 5); `LC(l10, 37, 21);
    `LC(l10, 38, 37); `LC(l10, 39, 53); `LC(l10, 40, 197); `LC(l10, 41, 213); `LC(l10, 42, 229); `LC(l10, 43, 245); `LC(l10, 44, 133); `LC(l10, 45, 149); `LC(l10, 46, 165);
    `LC(l10, 47, 181); `LC(l10, 48, 134); `LC(l10, 49, 150); `LC(l10, 50, 166); `LC(l10, 51, 182); `LC(l10, 52, 198); `LC(l10, 53, 214); `LC(l10, 54, 230); `LC(l10, 55, 246);
    `LC(l10, 56, 6); `LC(l10, 57, 22); `LC(l10, 58, 38); `LC(l10, 59, 54); `LC(l10, 60, 70); `LC(l10, 61, 86); `LC(l10, 62, 102); `LC(l10, 63, 118); `LC(l10, 64, 138);
    `LC(l10, 65, 154); `LC(l10, 66, 170); `LC(l10, 67, 186); `LC(l10, 68, 202); `LC(l10, 69, 218); `LC(l10, 70, 234); `LC(l10, 71, 250); `LC(l10, 72, 10); `LC(l10, 73, 26);
    `LC(l10, 74, 42); `LC(l10, 75, 58); `LC(l10, 76, 74); `LC(l10, 77, 90); `LC(l10, 78, 106); `LC(l10, 79, 122); `LC(l10, 80, 73); `LC(l10, 81, 89); `LC(l10, 82, 105);
    `LC(l10, 83, 121); `LC(l10, 84, 9); `LC(l10, 85, 25); `LC(l10, 86, 41); `LC(l10, 87, 57); `LC(l10, 88, 201); `LC(l10, 89, 217); `LC(l10, 90, 233); `LC(l10, 91, 249);
    `LC(l10, 92, 137); `LC(l10, 93, 153); `LC(l10, 94, 169); `LC(l10, 95, 185); `LC(l10, 96, 207); `LC(l10, 97, 223); `LC(l10, 98, 239); `LC(l10, 99, 255); `LC(l10, 100, 143);
    `LC(l10, 101, 159); `LC(l10, 102, 175); `LC(l10, 103, 191); `LC(l10, 104, 79); `LC(l10, 105, 95); `LC(l10, 106, 111); `LC(l10, 107, 127); `LC(l10, 108, 15); `LC(l10, 109, 31);
    `LC(l10, 110, 47); `LC(l10, 111, 63); `LC(l10, 112, 12); `LC(l10, 113, 28); `LC(l10, 114, 44); `LC(l10, 115, 60); `LC(l10, 116, 76); `LC(l10, 117, 92); `LC(l10, 118, 108);
    `LC(l10, 119, 124); `LC(l10, 120, 140); `LC(l10, 121, 156); `LC(l10, 122, 172); `LC(l10, 123, 188); `LC(l10, 124, 204); `LC(l10, 125, 220); `LC(l10, 126, 236); `LC(l10, 127, 252);
    `LC(l10, 128, 215); `LC(l10, 129, 199); `LC(l10, 130, 247); `LC(l10, 131, 231); `LC(l10, 132, 151); `LC(l10, 133, 135); `LC(l10, 134, 183); `LC(l10, 135, 167); `LC(l10, 136, 87);
    `LC(l10, 137, 71); `LC(l10, 138, 119); `LC(l10, 139, 103); `LC(l10, 140, 23); `LC(l10, 141, 7); `LC(l10, 142, 55); `LC(l10, 143, 39); `LC(l10, 144, 20); `LC(l10, 145, 4);
    `LC(l10, 146, 52); `LC(l10, 147, 36); `LC(l10, 148, 84); `LC(l10, 149, 68); `LC(l10, 150, 116); `LC(l10, 151, 100); `LC(l10, 152, 148); `LC(l10, 153, 132); `LC(l10, 154, 180);
    `LC(l10, 155, 164); `LC(l10, 156, 212); `LC(l10, 157, 196); `LC(l10, 158, 244); `LC(l10, 159, 228); `LC(l10, 160, 146); `LC(l10, 161, 130); `LC(l10, 162, 178);
    `LC(l10, 163, 162); `LC(l10, 164, 210); `LC(l10, 165, 194); `LC(l10, 166, 242); `LC(l10, 167, 226); `LC(l10, 168, 18); `LC(l10, 169, 2); `LC(l10, 170, 50); `LC(l10, 171, 34);
    `LC(l10, 172, 82); `LC(l10, 173, 66); `LC(l10, 174, 114); `LC(l10, 175, 98); `LC(l10, 176, 81); `LC(l10, 177, 65); `LC(l10, 178, 113); `LC(l10, 179, 97); `LC(l10, 180, 17);
    `LC(l10, 181, 1); `LC(l10, 182, 49); `LC(l10, 183, 33); `LC(l10, 184, 209); `LC(l10, 185, 193); `LC(l10, 186, 241); `LC(l10, 187, 225); `LC(l10, 188, 145); `LC(l10, 189, 129);
    `LC(l10, 190, 177); `LC(l10, 191, 161); `LC(l10, 192, 93); `LC(l10, 193, 77); `LC(l10, 194, 125); `LC(l10, 195, 109); `LC(l10, 196, 29); `LC(l10, 197, 13); `LC(l10, 198, 61);
    `LC(l10, 199, 45); `LC(l10, 200, 221); `LC(l10, 201, 205); `LC(l10, 202, 253); `LC(l10, 203, 237); `LC(l10, 204, 157); `LC(l10, 205, 141); `LC(l10, 206, 189); `LC(l10, 207, 173);
    `LC(l10, 208, 158); `LC(l10, 209, 142); `LC(l10, 210, 190); `LC(l10, 211, 174); `LC(l10, 212, 222); `LC(l10, 213, 206); `LC(l10, 214, 254); `LC(l10, 215, 238); `LC(l10, 216, 30);
    `LC(l10, 217, 14); `LC(l10, 218, 62); `LC(l10, 219, 46); `LC(l10, 220, 94); `LC(l10, 221, 78); `LC(l10, 222, 126); `LC(l10, 223, 110); `LC(l10, 224, 24); `LC(l10, 225, 8);
    `LC(l10, 226, 56); `LC(l10, 227, 40); `LC(l10, 228, 88); `LC(l10, 229, 72); `LC(l10, 230, 120); `LC(l10, 231, 104); `LC(l10, 232, 152); `LC(l10, 233, 136); `LC(l10, 234, 184);
    `LC(l10, 235, 168); `LC(l10, 236, 216); `LC(l10, 237, 200); `LC(l10, 238, 248); `LC(l10, 239, 232); `LC(l10, 240, 219); `LC(l10, 241, 203); `LC(l10, 242, 251);
    `LC(l10, 243, 235); `LC(l10, 244, 155); `LC(l10, 245, 139); `LC(l10, 246, 187); `LC(l10, 247, 171); `LC(l10, 248, 91); `LC(l10, 249, 75); `LC(l10, 250, 123); `LC(l10, 251, 107);
    `LC(l10, 252, 27); `LC(l10, 253, 11); `LC(l10, 254, 59); `LC(l10, 255, 43);
    `LC(lC2, 0, 0); `LC(lC2, 1, 194); `LC(lC2, 2, 71); `LC(lC2, 3, 133); `LC(lC2, 4, 142); `LC(lC2, 5, 76); `LC(lC2, 6, 201); `LC(lC2, 7, 11); `LC(lC2, 8, 223); `LC(lC2, 9, 29);
    `LC(lC2, 10, 152); `LC(lC2, 11, 90); `LC(lC2, 12, 81); `LC(lC2, 13, 147); `LC(lC2, 14, 22); `LC(lC2, 15, 212); `LC(lC2, 16, 125); `LC(lC2, 17, 191); `LC(lC2, 18, 58);
    `LC(lC2, 19, 248); `LC(lC2, 20, 243); `LC(lC2, 21, 49); `LC(lC2, 22, 180); `LC(lC2, 23, 118); `LC(lC2, 24, 162); `LC(lC2, 25, 96); `LC(lC2, 26, 229); `LC(lC2, 27, 39);
    `LC(lC2, 28, 44); `LC(lC2, 29, 238); `LC(lC2, 30, 107); `LC(lC2, 31, 169); `LC(lC2, 32, 250); `LC(lC2, 33, 56); `LC(lC2, 34, 189); `LC(lC2, 35, 127); `LC(lC2, 36, 116);
    `LC(lC2, 37, 182); `LC(lC2, 38, 51); `LC(lC2, 39, 241); `LC(lC2, 40, 37); `LC(lC2, 41, 231); `LC(lC2, 42, 98); `LC(lC2, 43, 160); `LC(lC2, 44, 171); `LC(lC2, 45, 105);
    `LC(lC2, 46, 236); `LC(lC2, 47, 46); `LC(lC2, 48, 135); `LC(lC2, 49, 69); `LC(lC2, 50, 192); `LC(lC2, 51, 2); `LC(lC2, 52, 9); `LC(lC2, 53, 203); `LC(lC2, 54, 78);
    `LC(lC2, 55, 140); `LC(lC2, 56, 88); `LC(lC2, 57, 154); `LC(lC2, 58, 31); `LC(lC2, 59, 221); `LC(lC2, 60, 214); `LC(lC2, 61, 20); `LC(lC2, 62, 145); `LC(lC2, 63, 83);
    `LC(lC2, 64, 55); `LC(lC2, 65, 245); `LC(lC2, 66, 112); `LC(lC2, 67, 178); `LC(lC2, 68, 185); `LC(lC2, 69, 123); `LC(lC2, 70, 254); `LC(lC2, 71, 60); `LC(lC2, 72, 232);
    `LC(lC2, 73, 42); `LC(lC2, 74, 175); `LC(lC2, 75, 109); `LC(lC2, 76, 102); `LC(lC2, 77, 164); `LC(lC2, 78, 33); `LC(lC2, 79, 227); `LC(lC2, 80, 74); `LC(lC2, 81, 136);
    `LC(lC2, 82, 13); `LC(lC2, 83, 207); `LC(lC2, 84, 196); `LC(lC2, 85, 6); `LC(lC2, 86, 131); `LC(lC2, 87, 65); `LC(lC2, 88, 149); `LC(lC2, 89, 87); `LC(lC2, 90, 210);
    `LC(lC2, 91, 16); `LC(lC2, 92, 27); `LC(lC2, 93, 217); `LC(lC2, 94, 92); `LC(lC2, 95, 158); `LC(lC2, 96, 205); `LC(lC2, 97, 15); `LC(lC2, 98, 138); `LC(lC2, 99, 72);
    `LC(lC2, 100, 67); `LC(lC2, 101, 129); `LC(lC2, 102, 4); `LC(lC2, 103, 198); `LC(lC2, 104, 18); `LC(lC2, 105, 208); `LC(lC2, 106, 85); `LC(lC2, 107, 151); `LC(lC2, 108, 156);
    `LC(lC2, 109, 94); `LC(lC2, 110, 219); `LC(lC2, 111, 25); `LC(lC2, 112, 176); `LC(lC2, 113, 114); `LC(lC2, 114, 247); `LC(lC2, 115, 53); `LC(lC2, 116, 62); `LC(lC2, 117, 252);
    `LC(lC2, 118, 121); `LC(lC2, 119, 187); `LC(lC2, 120, 111); `LC(lC2, 121, 173); `LC(lC2, 122, 40); `LC(lC2, 123, 234); `LC(lC2, 124, 225); `LC(lC2, 125, 35); `LC(lC2, 126, 166);
    `LC(lC2, 127, 100); `LC(lC2, 128, 110); `LC(lC2, 129, 172); `LC(lC2, 130, 41); `LC(lC2, 131, 235); `LC(lC2, 132, 224); `LC(lC2, 133, 34); `LC(lC2, 134, 167); `LC(lC2, 135, 101);
    `LC(lC2, 136, 177); `LC(lC2, 137, 115); `LC(lC2, 138, 246); `LC(lC2, 139, 52); `LC(lC2, 140, 63); `LC(lC2, 141, 253); `LC(lC2, 142, 120); `LC(lC2, 143, 186); `LC(lC2, 144, 19);
    `LC(lC2, 145, 209); `LC(lC2, 146, 84); `LC(lC2, 147, 150); `LC(lC2, 148, 157); `LC(lC2, 149, 95); `LC(lC2, 150, 218); `LC(lC2, 151, 24); `LC(lC2, 152, 204); `LC(lC2, 153, 14);
    `LC(lC2, 154, 139); `LC(lC2, 155, 73); `LC(lC2, 156, 66); `LC(lC2, 157, 128); `LC(lC2, 158, 5); `LC(lC2, 159, 199); `LC(lC2, 160, 148); `LC(lC2, 161, 86); `LC(lC2, 162, 211);
    `LC(lC2, 163, 17); `LC(lC2, 164, 26); `LC(lC2, 165, 216); `LC(lC2, 166, 93); `LC(lC2, 167, 159); `LC(lC2, 168, 75); `LC(lC2, 169, 137); `LC(lC2, 170, 12); `LC(lC2, 171, 206);
    `LC(lC2, 172, 197); `LC(lC2, 173, 7); `LC(lC2, 174, 130); `LC(lC2, 175, 64); `LC(lC2, 176, 233); `LC(lC2, 177, 43); `LC(lC2, 178, 174); `LC(lC2, 179, 108); `LC(lC2, 180, 103);
    `LC(lC2, 181, 165); `LC(lC2, 182, 32); `LC(lC2, 183, 226); `LC(lC2, 184, 54); `LC(lC2, 185, 244); `LC(lC2, 186, 113); `LC(lC2, 187, 179); `LC(lC2, 188, 184); `LC(lC2, 189, 122);
    `LC(lC2, 190, 255); `LC(lC2, 191, 61); `LC(lC2, 192, 89); `LC(lC2, 193, 155); `LC(lC2, 194, 30); `LC(lC2, 195, 220); `LC(lC2, 196, 215); `LC(lC2, 197, 21); `LC(lC2, 198, 144);
    `LC(lC2, 199, 82); `LC(lC2, 200, 134); `LC(lC2, 201, 68); `LC(lC2, 202, 193); `LC(lC2, 203, 3); `LC(lC2, 204, 8); `LC(lC2, 205, 202); `LC(lC2, 206, 79); `LC(lC2, 207, 141);
    `LC(lC2, 208, 36); `LC(lC2, 209, 230); `LC(lC2, 210, 99); `LC(lC2, 211, 161); `LC(lC2, 212, 170); `LC(lC2, 213, 104); `LC(lC2, 214, 237); `LC(lC2, 215, 47); `LC(lC2, 216, 251);
    `LC(lC2, 217, 57); `LC(lC2, 218, 188); `LC(lC2, 219, 126); `LC(lC2, 220, 117); `LC(lC2, 221, 183); `LC(lC2, 222, 50); `LC(lC2, 223, 240); `LC(lC2, 224, 163); `LC(lC2, 225, 97);
    `LC(lC2, 226, 228); `LC(lC2, 227, 38); `LC(lC2, 228, 45); `LC(lC2, 229, 239); `LC(lC2, 230, 106); `LC(lC2, 231, 168); `LC(lC2, 232, 124); `LC(lC2, 233, 190); `LC(lC2, 234, 59);
    `LC(lC2, 235, 249); `LC(lC2, 236, 242); `LC(lC2, 237, 48); `LC(lC2, 238, 181); `LC(lC2, 239, 119); `LC(lC2, 240, 222); `LC(lC2, 241, 28); `LC(lC2, 242, 153); `LC(lC2, 243, 91);
    `LC(lC2, 244, 80); `LC(lC2, 245, 146); `LC(lC2, 246, 23); `LC(lC2, 247, 213); `LC(lC2, 248, 1); `LC(lC2, 249, 195); `LC(lC2, 250, 70); `LC(lC2, 251, 132); `LC(lC2, 252, 143);
    `LC(lC2, 253, 77); `LC(lC2, 254, 200); `LC(lC2, 255, 10);
    `LC(lC0, 0, 0); `LC(lC0, 1, 192); `LC(lC0, 2, 67); `LC(lC0, 3, 131); `LC(lC0, 4, 134); `LC(lC0, 5, 70); `LC(lC0, 6, 197); `LC(lC0, 7, 5); `LC(lC0, 8, 207); `LC(lC0, 9, 15);
    `LC(lC0, 10, 140); `LC(lC0, 11, 76); `LC(lC0, 12, 73); `LC(lC0, 13, 137); `LC(lC0, 14, 10); `LC(lC0, 15, 202); `LC(lC0, 16, 93); `LC(lC0, 17, 157); `LC(lC0, 18, 30);
    `LC(lC0, 19, 222); `LC(lC0, 20, 219); `LC(lC0, 21, 27); `LC(lC0, 22, 152); `LC(lC0, 23, 88); `LC(lC0, 24, 146); `LC(lC0, 25, 82); `LC(lC0, 26, 209); `LC(lC0, 27, 17);
    `LC(lC0, 28, 20); `LC(lC0, 29, 212); `LC(lC0, 30, 87); `LC(lC0, 31, 151); `LC(lC0, 32, 186); `LC(lC0, 33, 122); `LC(lC0, 34, 249); `LC(lC0, 35, 57); `LC(lC0, 36, 60);
    `LC(lC0, 37, 252); `LC(lC0, 38, 127); `LC(lC0, 39, 191); `LC(lC0, 40, 117); `LC(lC0, 41, 181); `LC(lC0, 42, 54); `LC(lC0, 43, 246); `LC(lC0, 44, 243); `LC(lC0, 45, 51);
    `LC(lC0, 46, 176); `LC(lC0, 47, 112); `LC(lC0, 48, 231); `LC(lC0, 49, 39); `LC(lC0, 50, 164); `LC(lC0, 51, 100); `LC(lC0, 52, 97); `LC(lC0, 53, 161); `LC(lC0, 54, 34);
    `LC(lC0, 55, 226); `LC(lC0, 56, 40); `LC(lC0, 57, 232); `LC(lC0, 58, 107); `LC(lC0, 59, 171); `LC(lC0, 60, 174); `LC(lC0, 61, 110); `LC(lC0, 62, 237); `LC(lC0, 63, 45);
    `LC(lC0, 64, 183); `LC(lC0, 65, 119); `LC(lC0, 66, 244); `LC(lC0, 67, 52); `LC(lC0, 68, 49); `LC(lC0, 69, 241); `LC(lC0, 70, 114); `LC(lC0, 71, 178); `LC(lC0, 72, 120);
    `LC(lC0, 73, 184); `LC(lC0, 74, 59); `LC(lC0, 75, 251); `LC(lC0, 76, 254); `LC(lC0, 77, 62); `LC(lC0, 78, 189); `LC(lC0, 79, 125); `LC(lC0, 80, 234); `LC(lC0, 81, 42);
    `LC(lC0, 82, 169); `LC(lC0, 83, 105); `LC(lC0, 84, 108); `LC(lC0, 85, 172); `LC(lC0, 86, 47); `LC(lC0, 87, 239); `LC(lC0, 88, 37); `LC(lC0, 89, 229); `LC(lC0, 90, 102);
    `LC(lC0, 91, 166); `LC(lC0, 92, 163); `LC(lC0, 93, 99); `LC(lC0, 94, 224); `LC(lC0, 95, 32); `LC(lC0, 96, 13); `LC(lC0, 97, 205); `LC(lC0, 98, 78); `LC(lC0, 99, 142);
    `LC(lC0, 100, 139); `LC(lC0, 101, 75); `LC(lC0, 102, 200); `LC(lC0, 103, 8); `LC(lC0, 104, 194); `LC(lC0, 105, 2); `LC(lC0, 106, 129); `LC(lC0, 107, 65); `LC(lC0, 108, 68);
    `LC(lC0, 109, 132); `LC(lC0, 110, 7); `LC(lC0, 111, 199); `LC(lC0, 112, 80); `LC(lC0, 113, 144); `LC(lC0, 114, 19); `LC(lC0, 115, 211); `LC(lC0, 116, 214); `LC(lC0, 117, 22);
    `LC(lC0, 118, 149); `LC(lC0, 119, 85); `LC(lC0, 120, 159); `LC(lC0, 121, 95); `LC(lC0, 122, 220); `LC(lC0, 123, 28); `LC(lC0, 124, 25); `LC(lC0, 125, 217); `LC(lC0, 126, 90);
    `LC(lC0, 127, 154); `LC(lC0, 128, 173); `LC(lC0, 129, 109); `LC(lC0, 130, 238); `LC(lC0, 131, 46); `LC(lC0, 132, 43); `LC(lC0, 133, 235); `LC(lC0, 134, 104); `LC(lC0, 135, 168);
    `LC(lC0, 136, 98); `LC(lC0, 137, 162); `LC(lC0, 138, 33); `LC(lC0, 139, 225); `LC(lC0, 140, 228); `LC(lC0, 141, 36); `LC(lC0, 142, 167); `LC(lC0, 143, 103); `LC(lC0, 144, 240);
    `LC(lC0, 145, 48); `LC(lC0, 146, 179); `LC(lC0, 147, 115); `LC(lC0, 148, 118); `LC(lC0, 149, 182); `LC(lC0, 150, 53); `LC(lC0, 151, 245); `LC(lC0, 152, 63); `LC(lC0, 153, 255);
    `LC(lC0, 154, 124); `LC(lC0, 155, 188); `LC(lC0, 156, 185); `LC(lC0, 157, 121); `LC(lC0, 158, 250); `LC(lC0, 159, 58); `LC(lC0, 160, 23); `LC(lC0, 161, 215); `LC(lC0, 162, 84);
    `LC(lC0, 163, 148); `LC(lC0, 164, 145); `LC(lC0, 165, 81); `LC(lC0, 166, 210); `LC(lC0, 167, 18); `LC(lC0, 168, 216); `LC(lC0, 169, 24); `LC(lC0, 170, 155); `LC(lC0, 171, 91);
    `LC(lC0, 172, 94); `LC(lC0, 173, 158); `LC(lC0, 174, 29); `LC(lC0, 175, 221); `LC(lC0, 176, 74); `LC(lC0, 177, 138); `LC(lC0, 178, 9); `LC(lC0, 179, 201); `LC(lC0, 180, 204);
    `LC(lC0, 181, 12); `LC(lC0, 182, 143); `LC(lC0, 183, 79); `LC(lC0, 184, 133); `LC(lC0, 185, 69); `LC(lC0, 186, 198); `LC(lC0, 187, 6); `LC(lC0, 188, 3); `LC(lC0, 189, 195);
    `LC(lC0, 190, 64); `LC(lC0, 191, 128); `LC(lC0, 192, 26); `LC(lC0, 193, 218); `LC(lC0, 194, 89); `LC(lC0, 195, 153); `LC(lC0, 196, 156); `LC(lC0, 197, 92); `LC(lC0, 198, 223);
    `LC(lC0, 199, 31); `LC(lC0, 200, 213); `LC(lC0, 201, 21); `LC(lC0, 202, 150); `LC(lC0, 203, 86); `LC(lC0, 204, 83); `LC(lC0, 205, 147); `LC(lC0, 206, 16); `LC(lC0, 207, 208);
    `LC(lC0, 208, 71); `LC(lC0, 209, 135); `LC(lC0, 210, 4); `LC(lC0, 211, 196); `LC(lC0, 212, 193); `LC(lC0, 213, 1); `LC(lC0, 214, 130); `LC(lC0, 215, 66); `LC(lC0, 216, 136);
    `LC(lC0, 217, 72); `LC(lC0, 218, 203); `LC(lC0, 219, 11); `LC(lC0, 220, 14); `LC(lC0, 221, 206); `LC(lC0, 222, 77); `LC(lC0, 223, 141); `LC(lC0, 224, 160); `LC(lC0, 225, 96);
    `LC(lC0, 226, 227); `LC(lC0, 227, 35); `LC(lC0, 228, 38); `LC(lC0, 229, 230); `LC(lC0, 230, 101); `LC(lC0, 231, 165); `LC(lC0, 232, 111); `LC(lC0, 233, 175); `LC(lC0, 234, 44);
    `LC(lC0, 235, 236); `LC(lC0, 236, 233); `LC(lC0, 237, 41); `LC(lC0, 238, 170); `LC(lC0, 239, 106); `LC(lC0, 240, 253); `LC(lC0, 241, 61); `LC(lC0, 242, 190); `LC(lC0, 243, 126);
    `LC(lC0, 244, 123); `LC(lC0, 245, 187); `LC(lC0, 246, 56); `LC(lC0, 247, 248); `LC(lC0, 248, 50); `LC(lC0, 249, 242); `LC(lC0, 250, 113); `LC(lC0, 251, 177); `LC(lC0, 252, 180);
    `LC(lC0, 253, 116); `LC(lC0, 254, 247); `LC(lC0, 255, 55);
    `LC(lFB, 0, 0); `LC(lFB, 1, 251); `LC(lFB, 2, 53); `LC(lFB, 3, 206); `LC(lFB, 4, 106); `LC(lFB, 5, 145); `LC(lFB, 6, 95); `LC(lFB, 7, 164); `LC(lFB, 8, 212); `LC(lFB, 9, 47);
    `LC(lFB, 10, 225); `LC(lFB, 11, 26); `LC(lFB, 12, 190); `LC(lFB, 13, 69); `LC(lFB, 14, 139); `LC(lFB, 15, 112); `LC(lFB, 16, 107); `LC(lFB, 17, 144); `LC(lFB, 18, 94);
    `LC(lFB, 19, 165); `LC(lFB, 20, 1); `LC(lFB, 21, 250); `LC(lFB, 22, 52); `LC(lFB, 23, 207); `LC(lFB, 24, 191); `LC(lFB, 25, 68); `LC(lFB, 26, 138); `LC(lFB, 27, 113);
    `LC(lFB, 28, 213); `LC(lFB, 29, 46); `LC(lFB, 30, 224); `LC(lFB, 31, 27); `LC(lFB, 32, 214); `LC(lFB, 33, 45); `LC(lFB, 34, 227); `LC(lFB, 35, 24); `LC(lFB, 36, 188);
    `LC(lFB, 37, 71); `LC(lFB, 38, 137); `LC(lFB, 39, 114); `LC(lFB, 40, 2); `LC(lFB, 41, 249); `LC(lFB, 42, 55); `LC(lFB, 43, 204); `LC(lFB, 44, 104); `LC(lFB, 45, 147);
    `LC(lFB, 46, 93); `LC(lFB, 47, 166); `LC(lFB, 48, 189); `LC(lFB, 49, 70); `LC(lFB, 50, 136); `LC(lFB, 51, 115); `LC(lFB, 52, 215); `LC(lFB, 53, 44); `LC(lFB, 54, 226);
    `LC(lFB, 55, 25); `LC(lFB, 56, 105); `LC(lFB, 57, 146); `LC(lFB, 58, 92); `LC(lFB, 59, 167); `LC(lFB, 60, 3); `LC(lFB, 61, 248); `LC(lFB, 62, 54); `LC(lFB, 63, 205);
    `LC(lFB, 64, 111); `LC(lFB, 65, 148); `LC(lFB, 66, 90); `LC(lFB, 67, 161); `LC(lFB, 68, 5); `LC(lFB, 69, 254); `LC(lFB, 70, 48); `LC(lFB, 71, 203); `LC(lFB, 72, 187);
    `LC(lFB, 73, 64); `LC(lFB, 74, 142); `LC(lFB, 75, 117); `LC(lFB, 76, 209); `LC(lFB, 77, 42); `LC(lFB, 78, 228); `LC(lFB, 79, 31); `LC(lFB, 80, 4); `LC(lFB, 81, 255);
    `LC(lFB, 82, 49); `LC(lFB, 83, 202); `LC(lFB, 84, 110); `LC(lFB, 85, 149); `LC(lFB, 86, 91); `LC(lFB, 87, 160); `LC(lFB, 88, 208); `LC(lFB, 89, 43); `LC(lFB, 90, 229);
    `LC(lFB, 91, 30); `LC(lFB, 92, 186); `LC(lFB, 93, 65); `LC(lFB, 94, 143); `LC(lFB, 95, 116); `LC(lFB, 96, 185); `LC(lFB, 97, 66); `LC(lFB, 98, 140); `LC(lFB, 99, 119);
    `LC(lFB, 100, 211); `LC(lFB, 101, 40); `LC(lFB, 102, 230); `LC(lFB, 103, 29); `LC(lFB, 104, 109); `LC(lFB, 105, 150); `LC(lFB, 106, 88); `LC(lFB, 107, 163); `LC(lFB, 108, 7);
    `LC(lFB, 109, 252); `LC(lFB, 110, 50); `LC(lFB, 111, 201); `LC(lFB, 112, 210); `LC(lFB, 113, 41); `LC(lFB, 114, 231); `LC(lFB, 115, 28); `LC(lFB, 116, 184); `LC(lFB, 117, 67);
    `LC(lFB, 118, 141); `LC(lFB, 119, 118); `LC(lFB, 120, 6); `LC(lFB, 121, 253); `LC(lFB, 122, 51); `LC(lFB, 123, 200); `LC(lFB, 124, 108); `LC(lFB, 125, 151); `LC(lFB, 126, 89);
    `LC(lFB, 127, 162); `LC(lFB, 128, 222); `LC(lFB, 129, 37); `LC(lFB, 130, 235); `LC(lFB, 131, 16); `LC(lFB, 132, 180); `LC(lFB, 133, 79); `LC(lFB, 134, 129); `LC(lFB, 135, 122);
    `LC(lFB, 136, 10); `LC(lFB, 137, 241); `LC(lFB, 138, 63); `LC(lFB, 139, 196); `LC(lFB, 140, 96); `LC(lFB, 141, 155); `LC(lFB, 142, 85); `LC(lFB, 143, 174); `LC(lFB, 144, 181);
    `LC(lFB, 145, 78); `LC(lFB, 146, 128); `LC(lFB, 147, 123); `LC(lFB, 148, 223); `LC(lFB, 149, 36); `LC(lFB, 150, 234); `LC(lFB, 151, 17); `LC(lFB, 152, 97); `LC(lFB, 153, 154);
    `LC(lFB, 154, 84); `LC(lFB, 155, 175); `LC(lFB, 156, 11); `LC(lFB, 157, 240); `LC(lFB, 158, 62); `LC(lFB, 159, 197); `LC(lFB, 160, 8); `LC(lFB, 161, 243); `LC(lFB, 162, 61);
    `LC(lFB, 163, 198); `LC(lFB, 164, 98); `LC(lFB, 165, 153); `LC(lFB, 166, 87); `LC(lFB, 167, 172); `LC(lFB, 168, 220); `LC(lFB, 169, 39); `LC(lFB, 170, 233); `LC(lFB, 171, 18);
    `LC(lFB, 172, 182); `LC(lFB, 173, 77); `LC(lFB, 174, 131); `LC(lFB, 175, 120); `LC(lFB, 176, 99); `LC(lFB, 177, 152); `LC(lFB, 178, 86); `LC(lFB, 179, 173); `LC(lFB, 180, 9);
    `LC(lFB, 181, 242); `LC(lFB, 182, 60); `LC(lFB, 183, 199); `LC(lFB, 184, 183); `LC(lFB, 185, 76); `LC(lFB, 186, 130); `LC(lFB, 187, 121); `LC(lFB, 188, 221); `LC(lFB, 189, 38);
    `LC(lFB, 190, 232); `LC(lFB, 191, 19); `LC(lFB, 192, 177); `LC(lFB, 193, 74); `LC(lFB, 194, 132); `LC(lFB, 195, 127); `LC(lFB, 196, 219); `LC(lFB, 197, 32); `LC(lFB, 198, 238);
    `LC(lFB, 199, 21); `LC(lFB, 200, 101); `LC(lFB, 201, 158); `LC(lFB, 202, 80); `LC(lFB, 203, 171); `LC(lFB, 204, 15); `LC(lFB, 205, 244); `LC(lFB, 206, 58); `LC(lFB, 207, 193);
    `LC(lFB, 208, 218); `LC(lFB, 209, 33); `LC(lFB, 210, 239); `LC(lFB, 211, 20); `LC(lFB, 212, 176); `LC(lFB, 213, 75); `LC(lFB, 214, 133); `LC(lFB, 215, 126); `LC(lFB, 216, 14);
    `LC(lFB, 217, 245); `LC(lFB, 218, 59); `LC(lFB, 219, 192); `LC(lFB, 220, 100); `LC(lFB, 221, 159); `LC(lFB, 222, 81); `LC(lFB, 223, 170); `LC(lFB, 224, 103); `LC(lFB, 225, 156);
    `LC(lFB, 226, 82); `LC(lFB, 227, 169); `LC(lFB, 228, 13); `LC(lFB, 229, 246); `LC(lFB, 230, 56); `LC(lFB, 231, 195); `LC(lFB, 232, 179); `LC(lFB, 233, 72); `LC(lFB, 234, 134);
    `LC(lFB, 235, 125); `LC(lFB, 236, 217); `LC(lFB, 237, 34); `LC(lFB, 238, 236); `LC(lFB, 239, 23); `LC(lFB, 240, 12); `LC(lFB, 241, 247); `LC(lFB, 242, 57); `LC(lFB, 243, 194);
    `LC(lFB, 244, 102); `LC(lFB, 245, 157); `LC(lFB, 246, 83); `LC(lFB, 247, 168); `LC(lFB, 248, 216); `LC(lFB, 249, 35); `LC(lFB, 250, 237); `LC(lFB, 251, 22); `LC(lFB, 252, 178);
    `LC(lFB, 253, 73); `LC(lFB, 254, 135); `LC(lFB, 255, 124);
  
  function automatic [127:0] lBlock;
    input [127:0] in;
    reg [127:0] R1; reg [127:0] R2; reg [127:0] R3; reg [127:0] R4; reg [127:0] R5; reg [127:0] R6; reg [127:0] R7; reg [127:0] R8;
    reg [127:0] R9; reg [127:0] R10; reg [127:0] R11; reg [127:0] R12; reg [127:0] R13; reg [127:0] R14; reg [127:0] R15;
    begin
      R1[119:0] = in[127:8];
      R1[127:120] = in[7:0] ^ l94[in[15:8]] ^ l20[in[23:16]] ^ l85[in[31:24]] ^ l10[in[39:32]] ^ lC2[in[47:40]] ^ lC0[in[55:48]] ^ in[63:56] ^ lFB[in[71:64]] ^
                    in[79:72] ^ lC0[in[87:80]] ^ lC2[in[95:88]] ^ l10[in[103:96]] ^ l85[in[111:104]] ^ l20[in[119:112]] ^ l94[in[127:120]];
      R2[119:0] = R1[127:8];
      R2[127:120] = R1[7:0] ^ l94[R1[15:8]] ^ l20[R1[23:16]] ^ l85[R1[31:24]] ^ l10[R1[39:32]] ^ lC2[R1[47:40]] ^ lC0[R1[55:48]] ^ R1[63:56] ^ lFB[R1[71:64]] ^
                    R1[79:72] ^ lC0[R1[87:80]] ^ lC2[R1[95:88]] ^ l10[R1[103:96]] ^ l85[R1[111:104]] ^ l20[R1[119:112]] ^ l94[R1[127:120]];
      R3[119:0] = R2[127:8];
      R3[127:120] = R2[7:0] ^ l94[R2[15:8]] ^ l20[R2[23:16]] ^ l85[R2[31:24]] ^ l10[R2[39:32]] ^ lC2[R2[47:40]] ^ lC0[R2[55:48]] ^ R2[63:56] ^ lFB[R2[71:64]] ^
                    R2[79:72] ^ lC0[R2[87:80]] ^ lC2[R2[95:88]] ^ l10[R2[103:96]] ^ l85[R2[111:104]] ^ l20[R2[119:112]] ^ l94[R2[127:120]];
      R4[119:0] = R3[127:8];
      R4[127:120] = R3[7:0] ^ l94[R3[15:8]] ^ l20[R3[23:16]] ^ l85[R3[31:24]] ^ l10[R3[39:32]] ^ lC2[R3[47:40]] ^ lC0[R3[55:48]] ^ R3[63:56] ^ lFB[R3[71:64]] ^
                    R3[79:72] ^ lC0[R3[87:80]] ^ lC2[R3[95:88]] ^ l10[R3[103:96]] ^ l85[R3[111:104]] ^ l20[R3[119:112]] ^ l94[R3[127:120]];
      R5[119:0] = R4[127:8];
      R5[127:120] = R4[7:0] ^ l94[R4[15:8]] ^ l20[R4[23:16]] ^ l85[R4[31:24]] ^ l10[R4[39:32]] ^ lC2[R4[47:40]] ^ lC0[R4[55:48]] ^ R4[63:56] ^ lFB[R4[71:64]] ^
                    R4[79:72] ^ lC0[R4[87:80]] ^ lC2[R4[95:88]] ^ l10[R4[103:96]] ^ l85[R4[111:104]] ^ l20[R4[119:112]] ^ l94[R4[127:120]];
      R6[119:0] = R5[127:8];
      R6[127:120] = R5[7:0] ^ l94[R5[15:8]] ^ l20[R5[23:16]] ^ l85[R5[31:24]] ^ l10[R5[39:32]] ^ lC2[R5[47:40]] ^ lC0[R5[55:48]] ^ R5[63:56] ^ lFB[R5[71:64]] ^
                    R5[79:72] ^ lC0[R5[87:80]] ^ lC2[R5[95:88]] ^ l10[R5[103:96]] ^ l85[R5[111:104]] ^ l20[R5[119:112]] ^ l94[R5[127:120]];
      R7[119:0] = R6[127:8];
      R7[127:120] = R6[7:0] ^ l94[R6[15:8]] ^ l20[R6[23:16]] ^ l85[R6[31:24]] ^ l10[R6[39:32]] ^ lC2[R6[47:40]] ^ lC0[R6[55:48]] ^ R6[63:56] ^ lFB[R6[71:64]] ^
                    R6[79:72] ^ lC0[R6[87:80]] ^ lC2[R6[95:88]] ^ l10[R6[103:96]] ^ l85[R6[111:104]] ^ l20[R6[119:112]] ^ l94[R6[127:120]];
      R8[119:0] = R7[127:8];
      R8[127:120] = R7[7:0] ^ l94[R7[15:8]] ^ l20[R7[23:16]] ^ l85[R7[31:24]] ^ l10[R7[39:32]] ^ lC2[R7[47:40]] ^ lC0[R7[55:48]] ^ R7[63:56] ^ lFB[R7[71:64]] ^
                    R7[79:72] ^ lC0[R7[87:80]] ^ lC2[R7[95:88]] ^ l10[R7[103:96]] ^ l85[R7[111:104]] ^ l20[R7[119:112]] ^ l94[R7[127:120]];
      R9[119:0] = R8[127:8];
      R9[127:120] = R8[7:0] ^ l94[R8[15:8]] ^ l20[R8[23:16]] ^ l85[R8[31:24]] ^ l10[R8[39:32]] ^ lC2[R8[47:40]] ^ lC0[R8[55:48]] ^ R8[63:56] ^ lFB[R8[71:64]] ^
                    R8[79:72] ^ lC0[R8[87:80]] ^ lC2[R8[95:88]] ^ l10[R8[103:96]] ^ l85[R8[111:104]] ^ l20[R8[119:112]] ^ l94[R8[127:120]];
      R10[119:0] = R9[127:8];
      R10[127:120] = R9[7:0] ^ l94[R9[15:8]] ^ l20[R9[23:16]] ^ l85[R9[31:24]] ^ l10[R9[39:32]] ^ lC2[R9[47:40]] ^ lC0[R9[55:48]] ^ R9[63:56] ^ lFB[R9[71:64]] ^
                    R9[79:72] ^ lC0[R9[87:80]] ^ lC2[R9[95:88]] ^ l10[R9[103:96]] ^ l85[R9[111:104]] ^ l20[R9[119:112]] ^ l94[R9[127:120]];
      R11[119:0] = R10[127:8];
      R11[127:120] = R10[7:0] ^ l94[R10[15:8]] ^ l20[R10[23:16]] ^ l85[R10[31:24]] ^ l10[R10[39:32]] ^ lC2[R10[47:40]] ^ lC0[R10[55:48]] ^ R10[63:56] ^ lFB[R10[71:64]] ^
                    R10[79:72] ^ lC0[R10[87:80]] ^ lC2[R10[95:88]] ^ l10[R10[103:96]] ^ l85[R10[111:104]] ^ l20[R10[119:112]] ^ l94[R10[127:120]];
      R12[119:0] = R11[127:8];
      R12[127:120] = R11[7:0] ^ l94[R11[15:8]] ^ l20[R11[23:16]] ^ l85[R11[31:24]] ^ l10[R11[39:32]] ^ lC2[R11[47:40]] ^ lC0[R11[55:48]] ^ R11[63:56] ^ lFB[R11[71:64]] ^
                    R11[79:72] ^ lC0[R11[87:80]] ^ lC2[R11[95:88]] ^ l10[R11[103:96]] ^ l85[R11[111:104]] ^ l20[R11[119:112]] ^ l94[R11[127:120]];
      R13[119:0] = R12[127:8];
      R13[127:120] = R12[7:0] ^ l94[R12[15:8]] ^ l20[R12[23:16]] ^ l85[R12[31:24]] ^ l10[R12[39:32]] ^ lC2[R12[47:40]] ^ lC0[R12[55:48]] ^ R12[63:56] ^ lFB[R12[71:64]] ^
                    R12[79:72] ^ lC0[R12[87:80]] ^ lC2[R12[95:88]] ^ l10[R12[103:96]] ^ l85[R12[111:104]] ^ l20[R12[119:112]] ^ l94[R12[127:120]];
      R14[119:0] = R13[127:8];
      R14[127:120] = R13[7:0] ^ l94[R13[15:8]] ^ l20[R13[23:16]] ^ l85[R13[31:24]] ^ l10[R13[39:32]] ^ lC2[R13[47:40]] ^ lC0[R13[55:48]] ^ R13[63:56] ^ lFB[R13[71:64]] ^
                    R13[79:72] ^ lC0[R13[87:80]] ^ lC2[R13[95:88]] ^ l10[R13[103:96]] ^ l85[R13[111:104]] ^ l20[R13[119:112]] ^ l94[R13[127:120]];
      R15[119:0] = R14[127:8];
      R15[127:120] = R14[7:0] ^ l94[R14[15:8]] ^ l20[R14[23:16]] ^ l85[R14[31:24]] ^ l10[R14[39:32]] ^ lC2[R14[47:40]] ^ lC0[R14[55:48]] ^ R14[63:56] ^ lFB[R14[71:64]] ^
                    R14[79:72] ^ lC0[R14[87:80]] ^ lC2[R14[95:88]] ^ l10[R14[103:96]] ^ l85[R14[111:104]] ^ l20[R14[119:112]] ^ l94[R14[127:120]];
      lBlock[119:0] = R15[127:8];
      lBlock[127:120] = R15[7:0] ^ l94[R15[15:8]] ^ l20[R15[23:16]] ^ l85[R15[31:24]] ^ l10[R15[39:32]] ^ lC2[R15[47:40]] ^ lC0[R15[55:48]] ^ R15[63:56] ^ lFB[R15[71:64]] ^
                    R15[79:72] ^ lC0[R15[87:80]] ^ lC2[R15[95:88]] ^ l10[R15[103:96]] ^ l85[R15[111:104]] ^ l20[R15[119:112]] ^ l94[R15[127:120]];
    end
  endfunction
  
  // CONSTS
  reg [4095:0] consts;
    assign consts[127:0]     = 128'h6ea276726c487ab85d27bd10dd849401;
    assign consts[255:128]   = 128'hdc87ece4d890f4b3ba4eb92079cbeb02;
    assign consts[383:256]   = 128'hb2259a96b4d88e0be7690430a44f7f03;
    assign consts[511:384]   = 128'h7bcd1b0b73e32ba5b79cb140f2551504;
    assign consts[639:512]   = 128'h156f6d791fab511deabb0c502fd18105;
    assign consts[767:640]   = 128'ha74af7efab73df160dd208608b9efe06;
    assign consts[895:768]   = 128'hc9e8819dc73ba5ae50f5b570561a6a07;
    assign consts[1023:896]  = 128'hf6593616e6055689adfba18027aa2a08;
    assign consts[1151:1024] = 128'h98fb40648a4d2c31f0dc1c90fa2ebe09;
    assign consts[1279:1152] = 128'h2adedaf23e95a23a17b518a05e61c10a;
    assign consts[1407:1280] = 128'h447cac8052ddd8824a92a5b083e5550b;
    assign consts[1535:1408] = 128'h8d942d1d95e67d2c1a6710c0d5ff3f0c;
    assign consts[1663:1536] = 128'he3365b6ff9ae07944740add0087bab0d;
    assign consts[1791:1664] = 128'h5113c1f94d76899fa029a9e0ac34d40e;
    assign consts[1919:1792] = 128'h3fb1b78b213ef327fd0e14f071b0400f;
    assign consts[2047:1920] = 128'h2fb26c2c0f0aacd1993581c34e975410;
    assign consts[2175:2048] = 128'h41101a5e6342d669c4123cd39313c011;
    assign consts[2303:2176] = 128'hf33580c8d79a5862237b38e3375cbf12;
    assign consts[2431:2304] = 128'h9d97f6babbd222da7e5c85f3ead82b13;
    assign consts[2559:2432] = 128'h547f77277ce987742ea93083bcc24114;
    assign consts[2687:2560] = 128'h3add015510a1fdcc738e8d936146d515;
    assign consts[2815:2688] = 128'h88f89bc3a47973c794e789a3c509aa16;
    assign consts[2943:2816] = 128'he65aedb1c831097fc9c034b3188d3e17;
    assign consts[3071:2944] = 128'hd9eb5a3ae90ffa5834ce2043693d7e18;
    assign consts[3199:3072] = 128'hb7492c48854780e069e99d53b4b9ea19;
    assign consts[3327:3200] = 128'h056cb6de319f0eeb8e80996310f6951a;
    assign consts[3455:3328] = 128'h6bcec0ac5dd77453d3a72473cd72011b;
    assign consts[3583:3456] = 128'ha22641319aecd1fd835291039b686b1c;
    assign consts[3711:3584] = 128'hcc843743f6a4ab45de752c1346ecff1d;
    assign consts[3839:3712] = 128'h7ea1add5427c254e391c2823e2a3801e;
    assign consts[3967:3840] = 128'h1003dba72e345ff6643b95333f27141f;
    assign consts[4095:3968] = 128'h5ea7d8581e149b61f16ac1459ceda820;

  //-------------------------------------------------------------------------------------------------------------------------------------------//
  // KEYS
  //-------------------------------------------------------------------------------------------------------------------------------------------//
  reg [127:0] xorK11; reg [127:0] sK11; reg [127:0] lK11; reg [127:0] k11;
  reg [127:0] xorK12; reg [127:0] sK12; reg [127:0] lK12; reg [127:0] k12;
  reg [127:0] xorK13; reg [127:0] sK13; reg [127:0] lK13; reg [127:0] k13;
  reg [127:0] xorK14; reg [127:0] sK14; reg [127:0] lK14; reg [127:0] k14;
  reg [127:0] xorK15; reg [127:0] sK15; reg [127:0] lK15; reg [127:0] k15;
  reg [127:0] xorK16; reg [127:0] sK16; reg [127:0] lK16; reg [127:0] k16;
  reg [127:0] xorK17; reg [127:0] sK17; reg [127:0] lK17; /*key4*/
  reg [127:0] xorK18; reg [127:0] sK18; reg [127:0] lK18; /*key3*/

  reg [127:0] xorK21; reg [127:0] sK21; reg [127:0] lK21; reg [127:0] k21;
  reg [127:0] xorK22; reg [127:0] sK22; reg [127:0] lK22; reg [127:0] k22;
  reg [127:0] xorK23; reg [127:0] sK23; reg [127:0] lK23; reg [127:0] k23;
  reg [127:0] xorK24; reg [127:0] sK24; reg [127:0] lK24; reg [127:0] k24;
  reg [127:0] xorK25; reg [127:0] sK25; reg [127:0] lK25; reg [127:0] k25;
  reg [127:0] xorK26; reg [127:0] sK26; reg [127:0] lK26; reg [127:0] k26;
  reg [127:0] xorK27; reg [127:0] sK27; reg [127:0] lK27; /*key6*/
  reg [127:0] xorK28; reg [127:0] sK28; reg [127:0] lK28; /*key5*/
  
  reg [127:0] xorK31; reg [127:0] sK31; reg [127:0] lK31; reg [127:0] k31;
  reg [127:0] xorK32; reg [127:0] sK32; reg [127:0] lK32; reg [127:0] k32;
  reg [127:0] xorK33; reg [127:0] sK33; reg [127:0] lK33; reg [127:0] k33;
  reg [127:0] xorK34; reg [127:0] sK34; reg [127:0] lK34; reg [127:0] k34;
  reg [127:0] xorK35; reg [127:0] sK35; reg [127:0] lK35; reg [127:0] k35;
  reg [127:0] xorK36; reg [127:0] sK36; reg [127:0] lK36; reg [127:0] k36;
  reg [127:0] xorK37; reg [127:0] sK37; reg [127:0] lK37; /*key8*/
  reg [127:0] xorK38; reg [127:0] sK38; reg [127:0] lK38; /*key7*/
  
  reg [127:0] xorK41; reg [127:0] sK41; reg [127:0] lK41; reg [127:0] k41;
  reg [127:0] xorK42; reg [127:0] sK42; reg [127:0] lK42; reg [127:0] k42;
  reg [127:0] xorK43; reg [127:0] sK43; reg [127:0] lK43; reg [127:0] k43;
  reg [127:0] xorK44; reg [127:0] sK44; reg [127:0] lK44; reg [127:0] k44;
  reg [127:0] xorK45; reg [127:0] sK45; reg [127:0] lK45; reg [127:0] k45;
  reg [127:0] xorK46; reg [127:0] sK46; reg [127:0] lK46; reg [127:0] k46;
  reg [127:0] xorK47; reg [127:0] sK47; reg [127:0] lK47; /*key10*/
  reg [127:0] xorK48; reg [127:0] sK48; reg [127:0] lK48; /*key9*/

  /// K_3 and K_4
  always @(posedge clk) begin
    xorK11 = key[255:128] ^ consts[127:0]; // X
    sK11 = sBlock(xorK11);                 // S
    lK11 = lBlock(sK11);                   // L
    k11 = lK11 ^ key[127:0];
  end
  always @(posedge clk) begin
    xorK12 = k11 ^ consts[255:128]; // X
    sK12 = sBlock(xorK12);          // S
    lK12 = lBlock(sK12);            // L
    k12 = lK12 ^ key[255:128];
  end
  always @(posedge clk) begin
    xorK13 = k12 ^ consts[383:256]; // X
    sK13 = sBlock(xorK13);          // S
    lK13 = lBlock(sK13);            // L
    k13 = lK13 ^ k11;
  end
  always @(posedge clk) begin
    xorK14 = k13 ^ consts[511:384]; // X
    sK14 = sBlock(xorK14);          // S
    lK14 = lBlock(sK14);            // L
    k14 = lK14 ^ k12;
  end
  always @(posedge clk) begin
    xorK15 = k14 ^ consts[639:512]; // X
    sK15 = sBlock(xorK15);          // S
    lK15 = lBlock(sK15);            // L
    k15 = lK15 ^ k13;
  end
  always @(posedge clk) begin
    xorK16 = k15 ^ consts[767:640]; // X
    sK16 = sBlock(xorK16);          // S
    lK16 = lBlock(sK16);            // L
    k16 = lK16 ^ k14;
  end
  always @(posedge clk) begin
    xorK17 = k16 ^ consts[895:768]; // X
    sK17 = sBlock(xorK17);          // S
    lK17 = lBlock(sK17);            // L
    key4 = lK17 ^ k15;
  end
  always @(posedge clk) begin
    xorK18 = key4 ^ consts[1023:896]; // X
    sK18 = sBlock(xorK18);            // S
    lK18 = lBlock(sK18);              // L
    key3 = lK18 ^ k16;
  end
  
  /// K_5 and K_6
  always @(posedge clk) begin
    xorK21 = key3 ^ consts[1151:1024]; // X
    sK21 = sBlock(xorK21);             // S
    lK21 = lBlock(sK21);               // L
    k21 = lK21 ^ key4;
  end
  always @(posedge clk) begin
    xorK22 = k21 ^ consts[1279:1152]; // X
    sK22 = sBlock(xorK22);            // S
    lK22 = lBlock(sK22);              // L
    k22 = lK22 ^ key3;
  end
  always @(posedge clk) begin
    xorK23 = k22 ^ consts[1407:1280]; // X
    sK23 = sBlock(xorK23);            // S
    lK23 = lBlock(sK23);              // L
    k23 = lK23 ^ k21;
  end
  always @(posedge clk) begin
    xorK24 = k23 ^ consts[1535:1408]; // X
    sK24 = sBlock(xorK24);            // S
    lK24 = lBlock(sK24);              // L
    k24 = lK24 ^ k22;
  end
  always @(posedge clk) begin
    xorK25 = k24 ^ consts[1663:1536]; // X
    sK25 = sBlock(xorK25);            // S
    lK25 = lBlock(sK25);              // L
    k25 = lK25 ^ k23;
  end
  always @(posedge clk) begin
    xorK26 = k25 ^ consts[1791:1664]; // X
    sK26 = sBlock(xorK26);            // S
    lK26 = lBlock(sK26);              // L
    k26 = lK26 ^ k24;
  end
  always @(posedge clk) begin
    xorK27 = k26 ^ consts[1919:1792]; // X
    sK27 = sBlock(xorK27);            // S
    lK27 = lBlock(sK27);              // L
    key6 = lK27 ^ k25;
  end
  always @(posedge clk) begin
    xorK28 = key6 ^ consts[2047:1920]; // X
    sK28 = sBlock(xorK28);             // S
    lK28 = lBlock(sK28);               // L
    key5 = lK28 ^ k26;
  end
  
  /// K_7 and K_8
  always @(posedge clk) begin
    xorK31 = key5 ^ consts[2175:2048]; // X
    sK31 = sBlock(xorK31);             // S
    lK31 = lBlock(sK31);               // L
    k31 = lK31 ^ key6;
  end
  always @(posedge clk) begin
    xorK32 = k31 ^ consts[2303:2176]; // X
    sK32 = sBlock(xorK32);            // S
    lK32 = lBlock(sK32);              // L
    k32 = lK32 ^ key5;
  end
  always @(posedge clk) begin
    xorK33 = k32 ^ consts[2431:2304]; // X
    sK33 = sBlock(xorK33);            // S
    lK33 = lBlock(sK33);              // L
    k33 = lK33 ^ k31;
  end
  always @(posedge clk) begin
    xorK34 = k33 ^ consts[2559:2432]; // X
    sK34 = sBlock(xorK34);            // S
    lK34 = lBlock(sK34);              // L
    k34 = lK34 ^ k32;
  end
  always @(posedge clk) begin
    xorK35 = k34 ^ consts[2687:2560]; // X
    sK35 = sBlock(xorK35);            // S
    lK35 = lBlock(sK35);              // L
    k35 = lK35 ^ k33;
  end
  always @(posedge clk) begin
    xorK36 = k35 ^ consts[2815:2688]; // X
    sK36 = sBlock(xorK36);            // S
    lK36 = lBlock(sK36);              // L
    k36 = lK36 ^ k34;
  end
  always @(posedge clk) begin
    xorK37 = k36 ^ consts[2943:2816]; // X
    sK37 = sBlock(xorK37);            // S
    lK37 = lBlock(sK37);              // L
    key8 = lK37 ^ k35;
  end
  always @(posedge clk) begin
    xorK38 = key8 ^ consts[3071:2944]; // X
    sK38 = sBlock(xorK38);             // S
    lK38 = lBlock(sK38);               // L
    key7 = lK38 ^ k36;
  end
  
  /// K_9 and K_10
  always @(posedge clk) begin
    xorK41 = key7 ^ consts[3199:3072]; // X
    sK41 = sBlock(xorK41);             // S
    lK41 = lBlock(sK41);               // L
    k41 = lK41 ^ key8;
  end
  always @(posedge clk) begin
    xorK42 = k41 ^ consts[3327:3200]; // X
    sK42 = sBlock(xorK42);            // S
    lK42 = lBlock(sK42);              // L
    k42 = lK42 ^ key7;
  end
  always @(posedge clk) begin
    xorK43 = k42 ^ consts[3455:3328]; // X
    sK43 = sBlock(xorK43);            // S
    lK43 = lBlock(sK43);              // L
    k43 = lK43 ^ k41;
  end
  always @(posedge clk) begin
    xorK44 = k43 ^ consts[3583:3456]; // X
    sK44 = sBlock(xorK44);            // S
    lK44 = lBlock(sK44);              // L
    k44 = lK44 ^ k42;
  end
  always @(posedge clk) begin
    xorK45 = k44 ^ consts[3711:3584]; // X
    sK45 = sBlock(xorK45);            // S
    lK45 = lBlock(sK45);              // L
    k45 = lK45 ^ k43;
  end
  always @(posedge clk) begin
    xorK46 = k45 ^ consts[3839:3712]; // X
    sK46 = sBlock(xorK46);            // S
    lK46 = lBlock(sK46);              // L
    k46 = lK46 ^ k44;
  end
  always @(posedge clk) begin
    xorK47 = k46 ^ consts[3967:3840]; // X
    sK47 = sBlock(xorK47);            // S
    lK47 = lBlock(sK47);              // L
    key10 = lK47 ^ k45;
  end
  always @(posedge clk) begin
    xorK48 = key10 ^ consts[4095:3968]; // X
    sK48 = sBlock(xorK48);              // S
    lK48 = lBlock(sK48);                // L
    key9 = lK48 ^ k46;
  end
  
  //-------------------------------------------------------------------------------------------------------------------------------------------//
  // ROUNDS
  //-------------------------------------------------------------------------------------------------------------------------------------------//
  
  reg [127:0] xR1; reg [127:0] sR1; reg [127:0] lR1;
  reg [127:0] xR2; reg [127:0] sR2; reg [127:0] lR2;
  reg [127:0] xR3; reg [127:0] sR3; reg [127:0] lR3;
  reg [127:0] xR4; reg [127:0] sR4; reg [127:0] lR4;
  reg [127:0] xR5; reg [127:0] sR5; reg [127:0] lR5;
  reg [127:0] xR6; reg [127:0] sR6; reg [127:0] lR6;
  reg [127:0] xR7; reg [127:0] sR7; reg [127:0] lR7;
  reg [127:0] xR8; reg [127:0] sR8; reg [127:0] lR8;
  reg [127:0] xR9; reg [127:0] sR9; reg [127:0] lR9;
  
  // ROUND 1
  always @(posedge clk) begin
    xR1 = block ^ key[255:128]; // X
    sR1 = sBlock(xR1);          // S
    lR1 = lBlock(sR1);          // L
  end
  // ROUND 2
  always @(posedge clk) begin
    xR2 = lR1 ^ key[127:0]; // X
    sR2 = sBlock(xR2);      // S
    lR2 = lBlock(sR2);      // L
  end
  // ROUND 3
  always @(posedge clk) begin
    xR3 = lR2 ^ key3;  // X
    sR3 = sBlock(xR3); // S
    lR3 = lBlock(sR3); // L
  end
  // ROUND 4
  always @(posedge clk) begin
    xR4 = lR3 ^ key4;  // X
    sR4 = sBlock(xR4); // S
    lR4 = lBlock(sR4); // L
  end
  // ROUND 5
  always @(posedge clk) begin
    xR5 = lR4 ^ key5;  // X
    sR5 = sBlock(xR5); // S
    lR5 = lBlock(sR5); // L
  end
  // ROUND 6
  always @(posedge clk) begin
    xR6 = lR5 ^ key6;  // X
    sR6 = sBlock(xR6); // S
    lR6 = lBlock(sR6); // L
  end
  // ROUND 7
  always @(posedge clk) begin
    xR7 = lR6 ^ key7;  // X
    sR7 = sBlock(xR7); // S
    lR7 = lBlock(sR7); // L
  end
  // ROUND 8
  always @(posedge clk) begin
    xR8 = lR7 ^ key8;  // X
    sR8 = sBlock(xR8); // S
    lR8 = lBlock(sR8); // L
  end
  // ROUND 9 and 10
  always @(posedge clk) begin
    xR9 = lR8 ^ key9;  // X
    sR9 = sBlock(xR9); // S
    lR9 = lBlock(sR9); // L
    enc = lR9 ^ key10;
  end
endmodule

