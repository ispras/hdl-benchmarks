//NOTE: no-implementation module stub

module GTECH_MUX4 (
    input wire D0,
    input wire D1,
    input wire D2,
    input wire D3,
    input wire A,
    input wire B,
    output wire Z
);

endmodule
