// IWLS benchmark module "i6" printed on Wed May 29 17:26:49 2002
module i6(\V138(0) , \V138(2) , \V32(27) , \V32(26) , \V32(25) , \V32(24) , \V32(23) , \V32(22) , \V32(21) , \V32(20) , \V32(19) , \V32(18) , \V32(17) , \V32(16) , \V32(15) , \V32(14) , \V32(13) , \V32(12) , \V32(11) , \V32(10) , \V32(9) , \V32(8) , \V32(7) , \V32(6) , \V32(5) , \V32(4) , \V32(3) , \V32(2) , \V32(1) , \V32(0) , \V64(27) , \V64(26) , \V64(25) , \V64(24) , \V64(23) , \V64(22) , \V64(21) , \V64(20) , \V64(19) , \V64(18) , \V64(17) , \V64(16) , \V64(15) , \V64(14) , \V64(13) , \V64(12) , \V64(11) , \V64(10) , \V64(9) , \V64(8) , \V64(7) , \V64(6) , \V64(5) , \V64(4) , \V64(3) , \V64(2) , \V64(1) , \V64(0) , \V96(27) , \V138(4) , \V96(26) , \V96(25) , \V96(24) , \V96(23) , \V96(22) , \V96(21) , \V96(20) , \V96(19) , \V96(18) , \V96(17) , \V96(16) , \V96(15) , \V96(14) , \V96(13) , \V96(12) , \V96(11) , \V96(10) , \V96(9) , \V96(8) , \V96(7) , \V96(6) , \V96(5) , \V96(4) , \V96(3) , \V96(2) , \V96(1) , \V96(0) , \V32(31) , \V32(30) , \V32(29) , \V32(28) , \V131(27) , \V131(26) , \V131(25) , \V131(24) , \V131(23) , \V131(22) , \V131(21) , \V131(20) , \V131(19) , \V131(18) , \V131(17) , \V131(16) , \V131(15) , \V131(14) , \V131(13) , \V131(12) , \V131(11) , \V131(10) , \V131(9) , \V131(8) , \V131(7) , \V131(6) , \V131(5) , \V131(4) , \V131(3) , \V131(2) , \V131(1) , \V131(0) , \V64(31) , \V64(30) , \V64(29) , \V64(28) , \V99(0) , \V138(3) , \V98(0) , \V97(0) , \V96(31) , \V96(30) , \V96(29) , \V96(28) , \V134(0) , \V133(1) , \V133(0) , \V131(31) , \V131(30) , \V131(29) , \V131(28) , \V166(27) , \V166(26) , \V166(25) , \V166(24) , \V166(23) , \V166(22) , \V166(21) , \V166(20) , \V166(19) , \V166(18) , \V166(17) , \V166(16) , \V166(15) , \V166(14) , \V166(13) , \V166(12) , \V166(11) , \V166(10) , \V166(9) , \V166(8) , \V166(7) , \V166(6) , \V166(5) , \V166(4) , \V166(3) , \V166(2) , \V166(1) , \V166(0) , \V198(31) , \V198(30) , \V198(29) , \V198(28) , \V198(27) , \V198(26) , \V198(25) , \V198(24) , \V198(23) , \V198(22) , \V198(21) , \V198(20) , \V198(19) , \V198(18) , \V198(17) , \V198(16) , \V198(15) , \V198(14) , \V198(13) , \V198(12) , \V198(11) , \V198(10) , \V198(9) , \V198(8) , \V198(7) , \V198(6) , \V198(5) , \V198(4) , \V198(3) , \V198(2) , \V198(1) , \V198(0) , \V205(6) , \V205(5) , \V205(4) , \V205(3) , \V205(2) , \V205(1) , \V205(0) );
input
  \V32(30) ,
  \V138(3) ,
  \V138(2) ,
  \V138(4) ,
  \V138(0) ,
  \V32(0) ,
  \V32(1) ,
  \V32(2) ,
  \V32(3) ,
  \V32(4) ,
  \V32(5) ,
  \V131(27) ,
  \V32(6) ,
  \V131(26) ,
  \V32(7) ,
  \V131(29) ,
  \V32(8) ,
  \V131(28) ,
  \V32(9) ,
  \V96(0) ,
  \V96(1) ,
  \V131(21) ,
  \V96(2) ,
  \V131(20) ,
  \V96(3) ,
  \V131(23) ,
  \V96(4) ,
  \V96(13) ,
  \V131(22) ,
  \V96(5) ,
  \V96(12) ,
  \V131(25) ,
  \V96(6) ,
  \V97(0) ,
  \V96(15) ,
  \V131(24) ,
  \V96(7) ,
  \V96(14) ,
  \V131(17) ,
  \V96(8) ,
  \V131(16) ,
  \V96(9) ,
  \V131(19) ,
  \V96(11) ,
  \V131(18) ,
  \V96(10) ,
  \V98(0) ,
  \V96(17) ,
  \V96(16) ,
  \V131(11) ,
  \V96(19) ,
  \V131(10) ,
  \V99(0) ,
  \V96(18) ,
  \V131(13) ,
  \V96(23) ,
  \V131(12) ,
  \V96(22) ,
  \V131(15) ,
  \V64(13) ,
  \V96(25) ,
  \V131(14) ,
  \V64(12) ,
  \V96(24) ,
  \V64(15) ,
  \V64(14) ,
  \V96(21) ,
  \V96(20) ,
  \V64(11) ,
  \V64(10) ,
  \V96(27) ,
  \V96(26) ,
  \V64(17) ,
  \V96(29) ,
  \V64(16) ,
  \V96(28) ,
  \V131(3) ,
  \V64(19) ,
  \V131(2) ,
  \V64(18) ,
  \V131(5) ,
  \V64(23) ,
  \V131(4) ,
  \V64(22) ,
  \V32(13) ,
  \V64(25) ,
  \V32(12) ,
  \V64(24) ,
  \V32(15) ,
  \V131(1) ,
  \V32(14) ,
  \V96(31) ,
  \V131(0) ,
  \V96(30) ,
  \V64(21) ,
  \V64(20) ,
  \V32(11) ,
  \V32(10) ,
  \V131(7) ,
  \V131(6) ,
  \V131(9) ,
  \V131(31) ,
  \V64(27) ,
  \V131(8) ,
  \V131(30) ,
  \V64(26) ,
  \V32(17) ,
  \V64(29) ,
  \V32(16) ,
  \V64(28) ,
  \V32(19) ,
  \V32(18) ,
  \V133(1) ,
  \V32(23) ,
  \V133(0) ,
  \V64(0) ,
  \V32(22) ,
  \V64(1) ,
  \V32(25) ,
  \V64(2) ,
  \V32(24) ,
  \V64(3) ,
  \V64(4) ,
  \V64(31) ,
  \V64(5) ,
  \V64(30) ,
  \V32(21) ,
  \V64(6) ,
  \V134(0) ,
  \V32(20) ,
  \V64(7) ,
  \V64(8) ,
  \V64(9) ,
  \V32(27) ,
  \V32(26) ,
  \V32(29) ,
  \V32(28) ,
  \V32(31) ;
output
  \V198(7) ,
  \V198(6) ,
  \V198(9) ,
  \V198(8) ,
  \V166(3) ,
  \V166(2) ,
  \V166(5) ,
  \V166(4) ,
  \V166(1) ,
  \V166(0) ,
  \V166(7) ,
  \V166(6) ,
  \V166(9) ,
  \V198(27) ,
  \V166(8) ,
  \V205(3) ,
  \V198(26) ,
  \V205(2) ,
  \V198(29) ,
  \V205(5) ,
  \V198(28) ,
  \V205(4) ,
  \V205(1) ,
  \V205(0) ,
  \V198(21) ,
  \V198(20) ,
  \V198(23) ,
  \V198(22) ,
  \V205(6) ,
  \V198(25) ,
  \V198(24) ,
  \V198(17) ,
  \V198(16) ,
  \V166(27) ,
  \V198(19) ,
  \V166(26) ,
  \V198(18) ,
  \V198(11) ,
  \V198(10) ,
  \V166(21) ,
  \V198(13) ,
  \V166(20) ,
  \V198(12) ,
  \V166(23) ,
  \V198(15) ,
  \V166(22) ,
  \V198(14) ,
  \V166(25) ,
  \V166(24) ,
  \V166(17) ,
  \V166(16) ,
  \V166(19) ,
  \V166(18) ,
  \V166(11) ,
  \V166(10) ,
  \V166(13) ,
  \V166(12) ,
  \V166(15) ,
  \V166(14) ,
  \V198(3) ,
  \V198(2) ,
  \V198(5) ,
  \V198(4) ,
  \V198(31) ,
  \V198(30) ,
  \V198(1) ,
  \V198(0) ;
wire
  \[60] ,
  \[61] ,
  \[62] ,
  \[63] ,
  \[64] ,
  \[65] ,
  \[66] ,
  \[67] ,
  \[68] ,
  \[69] ,
  \[0] ,
  \[1] ,
  \[2] ,
  \[3] ,
  \[4] ,
  \[70] ,
  \[5] ,
  \[71] ,
  \[6] ,
  \[72] ,
  \[7] ,
  \[73] ,
  \[8] ,
  \[74] ,
  \[9] ,
  \[10] ,
  \[11] ,
  \[12] ,
  \[13] ,
  \[14] ,
  \[15] ,
  \[16] ,
  \[17] ,
  \[18] ,
  \[19] ,
  \[20] ,
  \[21] ,
  \[22] ,
  V451,
  \[23] ,
  \[24] ,
  \[25] ,
  \[26] ,
  \[27] ,
  \[28] ,
  \[29] ,
  \[30] ,
  \[31] ,
  \[32] ,
  \[33] ,
  \[34] ,
  \[35] ,
  \[36] ,
  \[37] ,
  \[38] ,
  \[39] ,
  \[40] ,
  \[41] ,
  \[42] ,
  \[43] ,
  \[44] ,
  \[45] ,
  \[46] ,
  \[47] ,
  \[48] ,
  \[49] ,
  \[50] ,
  \[51] ,
  \[52] ,
  \[53] ,
  \[54] ,
  \[55] ,
  \[56] ,
  \[57] ,
  \[58] ,
  \[59] ;
assign
  \[60]  = (\V134(0)  & (\V138(3)  & \V138(0) )) | (\[72]  & \V99(0) ),
  \[61]  = (\[73]  & \V133(1) ) | ((\[72]  & \V98(0) ) | ((\[69]  & ~\V133(1) ) | \[74] )),
  \[62]  = (\[73]  & \V133(0) ) | ((\[72]  & \V97(0) ) | ((\[69]  & ~\V133(0) ) | \[74] )),
  \V198(7)  = \[52] ,
  \[63]  = (\[73]  & \V131(31) ) | ((\[72]  & \V96(31) ) | ((\[69]  & ~\V131(31) ) | \[74] )),
  \V198(6)  = \[53] ,
  \[64]  = (\[73]  & \V131(30) ) | ((\[72]  & \V96(30) ) | ((\[69]  & ~\V131(30) ) | \[74] )),
  \V198(9)  = \[50] ,
  \[65]  = (\[73]  & \V131(29) ) | ((\[72]  & \V96(29) ) | ((\[69]  & ~\V131(29) ) | \[74] )),
  \V198(8)  = \[51] ,
  \[66]  = (\[73]  & \V131(28) ) | ((\[72]  & \V96(28) ) | ((\[69]  & ~\V131(28) ) | \[74] )),
  \[67]  = ~\V138(2)  & ~\V138(0) ,
  \[68]  = ~\V138(2)  & \V138(0) ,
  \[69]  = \V138(2)  & \V138(0) ,
  \[0]  = (\[69]  & ~\V64(27) ) | ((\[68]  & \V64(27) ) | (\[67]  & \V32(27) )),
  \[1]  = (\[69]  & ~\V64(26) ) | ((\[68]  & \V64(26) ) | (\[67]  & \V32(26) )),
  \[2]  = (\[69]  & ~\V64(25) ) | ((\[68]  & \V64(25) ) | (\[67]  & \V32(25) )),
  \[3]  = (\[69]  & ~\V64(24) ) | ((\[68]  & \V64(24) ) | (\[67]  & \V32(24) )),
  \[4]  = (\[69]  & ~\V64(23) ) | ((\[68]  & \V64(23) ) | (\[67]  & \V32(23) )),
  \[70]  = \[68]  & \V138(4) ,
  \[5]  = (\[69]  & ~\V64(22) ) | ((\[68]  & \V64(22) ) | (\[67]  & \V32(22) )),
  \[71]  = \[67]  & \V138(4) ,
  \[6]  = (\[69]  & ~\V64(21) ) | ((\[68]  & \V64(21) ) | (\[67]  & \V32(21) )),
  \[72]  = \[67]  & \V138(3) ,
  \[7]  = (\[69]  & ~\V64(20) ) | ((\[68]  & \V64(20) ) | (\[67]  & \V32(20) )),
  \[73]  = \[68]  & \V138(3) ,
  \[8]  = (\[69]  & ~\V64(19) ) | ((\[68]  & \V64(19) ) | (\[67]  & \V32(19) )),
  \[74]  = ~\V138(3)  & \V138(2) ,
  \[9]  = (\[69]  & ~\V64(18) ) | ((\[68]  & \V64(18) ) | (\[67]  & \V32(18) )),
  \[10]  = (\[69]  & ~\V64(17) ) | ((\[68]  & \V64(17) ) | (\[67]  & \V32(17) )),
  \[11]  = (\[69]  & ~\V64(16) ) | ((\[68]  & \V64(16) ) | (\[67]  & \V32(16) )),
  \V166(3)  = \[24] ,
  \[12]  = (\[69]  & ~\V64(15) ) | ((\[68]  & \V64(15) ) | (\[67]  & \V32(15) )),
  \V166(2)  = \[25] ,
  \[13]  = (\[69]  & ~\V64(14) ) | ((\[68]  & \V64(14) ) | (\[67]  & \V32(14) )),
  \V166(5)  = \[22] ,
  \[14]  = (\[69]  & ~\V64(13) ) | ((\[68]  & \V64(13) ) | (\[67]  & \V32(13) )),
  \V166(4)  = \[23] ,
  \[15]  = (\[69]  & ~\V64(12) ) | ((\[68]  & \V64(12) ) | (\[67]  & \V32(12) )),
  \[16]  = (\[69]  & ~\V64(11) ) | ((\[68]  & \V64(11) ) | (\[67]  & \V32(11) )),
  \[17]  = (\[69]  & ~\V64(10) ) | ((\[68]  & \V64(10) ) | (\[67]  & \V32(10) )),
  \V166(1)  = \[26] ,
  \[18]  = (\[69]  & ~\V64(9) ) | ((\[68]  & \V64(9) ) | (\[67]  & \V32(9) )),
  \V166(0)  = \[27] ,
  \[19]  = (\[69]  & ~\V64(8) ) | ((\[68]  & \V64(8) ) | (\[67]  & \V32(8) )),
  \V166(7)  = \[20] ,
  \V166(6)  = \[21] ,
  \V166(9)  = \[18] ,
  \V198(27)  = \[32] ,
  \[20]  = (\[69]  & ~\V64(7) ) | ((\[68]  & \V64(7) ) | (\[67]  & \V32(7) )),
  \V166(8)  = \[19] ,
  \V205(3)  = \[63] ,
  \V198(26)  = \[33] ,
  \[21]  = (\[69]  & ~\V64(6) ) | ((\[68]  & \V64(6) ) | (\[67]  & \V32(6) )),
  \V205(2)  = \[64] ,
  \V198(29)  = \[30] ,
  \[22]  = (\[69]  & ~\V64(5) ) | ((\[68]  & \V64(5) ) | (\[67]  & \V32(5) )),
  \V205(5)  = \[61] ,
  V451 = ~\V138(4)  & \V138(2) ,
  \V198(28)  = \[31] ,
  \[23]  = (\[69]  & ~\V64(4) ) | ((\[68]  & \V64(4) ) | (\[67]  & \V32(4) )),
  \V205(4)  = \[62] ,
  \[24]  = (\[69]  & ~\V64(3) ) | ((\[68]  & \V64(3) ) | (\[67]  & \V32(3) )),
  \[25]  = (\[69]  & ~\V64(2) ) | ((\[68]  & \V64(2) ) | (\[67]  & \V32(2) )),
  \[26]  = (\[69]  & ~\V64(1) ) | ((\[68]  & \V64(1) ) | (\[67]  & \V32(1) )),
  \V205(1)  = \[65] ,
  \[27]  = (\[69]  & ~\V64(0) ) | ((\[68]  & \V64(0) ) | (\[67]  & \V32(0) )),
  \V205(0)  = \[66] ,
  \[28]  = (\[71]  & \V96(27) ) | ((\[70]  & \V131(27) ) | ((\[69]  & ~\V131(27) ) | V451)),
  \[29]  = (\[71]  & \V96(26) ) | ((\[70]  & \V131(26) ) | ((\[69]  & ~\V131(26) ) | V451)),
  \V198(21)  = \[38] ,
  \V198(20)  = \[39] ,
  \V198(23)  = \[36] ,
  \V198(22)  = \[37] ,
  \V205(6)  = \[60] ,
  \V198(25)  = \[34] ,
  \V198(24)  = \[35] ,
  \V198(17)  = \[42] ,
  \[30]  = (\[71]  & \V96(25) ) | ((\[70]  & \V131(25) ) | ((\[69]  & ~\V131(25) ) | V451)),
  \V198(16)  = \[43] ,
  \V166(27)  = \[0] ,
  \[31]  = (\[71]  & \V96(24) ) | ((\[70]  & \V131(24) ) | ((\[69]  & ~\V131(24) ) | V451)),
  \V198(19)  = \[40] ,
  \V166(26)  = \[1] ,
  \[32]  = (\[71]  & \V96(23) ) | ((\[70]  & \V131(23) ) | ((\[69]  & ~\V131(23) ) | V451)),
  \V198(18)  = \[41] ,
  \[33]  = (\[71]  & \V96(22) ) | ((\[70]  & \V131(22) ) | ((\[69]  & ~\V131(22) ) | V451)),
  \[34]  = (\[71]  & \V96(21) ) | ((\[70]  & \V131(21) ) | ((\[69]  & ~\V131(21) ) | V451)),
  \[35]  = (\[71]  & \V96(20) ) | ((\[70]  & \V131(20) ) | ((\[69]  & ~\V131(20) ) | V451)),
  \[36]  = (\[71]  & \V96(19) ) | ((\[70]  & \V131(19) ) | ((\[69]  & ~\V131(19) ) | V451)),
  \[37]  = (\[71]  & \V96(18) ) | ((\[70]  & \V131(18) ) | ((\[69]  & ~\V131(18) ) | V451)),
  \[38]  = (\[71]  & \V96(17) ) | ((\[70]  & \V131(17) ) | ((\[69]  & ~\V131(17) ) | V451)),
  \[39]  = (\[71]  & \V96(16) ) | ((\[70]  & \V131(16) ) | ((\[69]  & ~\V131(16) ) | V451)),
  \V198(11)  = \[48] ,
  \V198(10)  = \[49] ,
  \V166(21)  = \[6] ,
  \V198(13)  = \[46] ,
  \V166(20)  = \[7] ,
  \V198(12)  = \[47] ,
  \V166(23)  = \[4] ,
  \V198(15)  = \[44] ,
  \V166(22)  = \[5] ,
  \V198(14)  = \[45] ,
  \V166(25)  = \[2] ,
  \V166(24)  = \[3] ,
  \[40]  = (\[71]  & \V96(15) ) | ((\[70]  & \V131(15) ) | ((\[69]  & ~\V131(15) ) | V451)),
  \V166(17)  = \[10] ,
  \[41]  = (\[71]  & \V96(14) ) | ((\[70]  & \V131(14) ) | ((\[69]  & ~\V131(14) ) | V451)),
  \V166(16)  = \[11] ,
  \[42]  = (\[71]  & \V96(13) ) | ((\[70]  & \V131(13) ) | ((\[69]  & ~\V131(13) ) | V451)),
  \V166(19)  = \[8] ,
  \[43]  = (\[71]  & \V96(12) ) | ((\[70]  & \V131(12) ) | ((\[69]  & ~\V131(12) ) | V451)),
  \V166(18)  = \[9] ,
  \[44]  = (\[71]  & \V96(11) ) | ((\[70]  & \V131(11) ) | ((\[69]  & ~\V131(11) ) | V451)),
  \[45]  = (\[71]  & \V96(10) ) | ((\[70]  & \V131(10) ) | ((\[69]  & ~\V131(10) ) | V451)),
  \[46]  = (\[71]  & \V96(9) ) | ((\[70]  & \V131(9) ) | ((\[69]  & ~\V131(9) ) | V451)),
  \[47]  = (\[71]  & \V96(8) ) | ((\[70]  & \V131(8) ) | ((\[69]  & ~\V131(8) ) | V451)),
  \[48]  = (\[71]  & \V96(7) ) | ((\[70]  & \V131(7) ) | ((\[69]  & ~\V131(7) ) | V451)),
  \[49]  = (\[71]  & \V96(6) ) | ((\[70]  & \V131(6) ) | ((\[69]  & ~\V131(6) ) | V451)),
  \V166(11)  = \[16] ,
  \V166(10)  = \[17] ,
  \V166(13)  = \[14] ,
  \V166(12)  = \[15] ,
  \V166(15)  = \[12] ,
  \V166(14)  = \[13] ,
  \[50]  = (\[71]  & \V96(5) ) | ((\[70]  & \V131(5) ) | ((\[69]  & ~\V131(5) ) | V451)),
  \[51]  = (\[71]  & \V96(4) ) | ((\[70]  & \V131(4) ) | ((\[69]  & ~\V131(4) ) | V451)),
  \[52]  = (\[71]  & \V96(3) ) | ((\[70]  & \V131(3) ) | ((\[69]  & ~\V131(3) ) | V451)),
  \[53]  = (\[71]  & \V96(2) ) | ((\[70]  & \V131(2) ) | ((\[69]  & ~\V131(2) ) | V451)),
  \[54]  = (\[71]  & \V96(1) ) | ((\[70]  & \V131(1) ) | ((\[69]  & ~\V131(1) ) | V451)),
  \[55]  = (\[71]  & \V96(0) ) | ((\[70]  & \V131(0) ) | ((\[69]  & ~\V131(0) ) | V451)),
  \[56]  = (\[71]  & \V32(31) ) | ((\[70]  & \V64(31) ) | ((\[69]  & ~\V64(31) ) | V451)),
  \V198(3)  = \[56] ,
  \[57]  = (\[71]  & \V32(30) ) | ((\[70]  & \V64(30) ) | ((\[69]  & ~\V64(30) ) | V451)),
  \V198(2)  = \[57] ,
  \[58]  = (\[71]  & \V32(29) ) | ((\[70]  & \V64(29) ) | ((\[69]  & ~\V64(29) ) | V451)),
  \V198(5)  = \[54] ,
  \[59]  = (\[71]  & \V32(28) ) | ((\[70]  & \V64(28) ) | ((\[69]  & ~\V64(28) ) | V451)),
  \V198(4)  = \[55] ,
  \V198(31)  = \[28] ,
  \V198(30)  = \[29] ,
  \V198(1)  = \[58] ,
  \V198(0)  = \[59] ;
endmodule

