// IWLS benchmark module "sbc" printed on Wed May 29 21:45:20 2002
module sbc(ACKl, BUS_Inactive, GRANTi, LastRQSTi, SBCResetPCC, PCCReq, PCCReqCode0, PCCReqCode1, PCCReqCode2, PCCReqCode3, PCCConfirm, RQSTi, SingleStep, STARTi, TM0i, TM1i, VACKl, VTM0i, VSACKi, ACKi, RESETi, SlotSpace_Id_Match, PCCSawReset, CoherencyState1i, CoherencyState2i, NuBusActive, PCCAck, PCCsync, STARTo, Tag_Match, TM1l, VTM0l, VTM1l, PCCAckCode, VACKi, physrecXXXXstate0, physrecXXXXstate1, wdcntXXXXstate1, wdcntXXXXstate2, wdcntXXXXstate3, physrecXXXXNextState0, physrecXXXXNextState1, wdcntXXXXNextState1, wdcntXXXXNextState2, wdcntXXXXNextState3, masterXXXXArb_active, masterXXXXEn_ABufo, masterXXXXEn_PDBufi, masterXXXXL_PDBufi, masterXXXXEn_VDBufi, masterXXXXEn_PDBufo, masterXXXXL_DBufo_if_TM0, masterXXXXRQSTo, masterXXXXSBC_WriteCache, nubusXXXXNuBusActive, nubusXXXXL_PABufi, resetXXXXSBCResetPCC, resetXXXXReset, slaveXXXXL_VABufi, slaveXXXXSBCReq, slaveXXXXSBCReqCode0, slaveXXXXSBCReqCode1, slaveXXXXSBCReqCode2, slaveXXXXSnoopAddrFromProc, slaveXXXXSnoopVTag_W, slaveXXXXSnoopState_W, slaveXXXXGenerateNextState, slaveXXXXSnoopVTagState_R, virmachXXXXEn_VDBufo, virmachXXXXSBCsetDirty, virmachXXXXSBCCacheRelease, virmachXXXXSBCConfigure, wdcntXXXXwd_cnt0, wdcntXXXXwd_cnt1, wdcntXXXXwd_cnt2, encodemuxXXXXMX_AD_8, nextstateXXXXCoherencyState2o, orXXXXACKo, orXXXXEn_CNTL, orXXXXRESETo, orXXXXTM0o, orXXXXTM1o, orXXXXEn_START, orXXXXSBCAck, orXXXXSBCAckCodelatch, orXXXXSBCAckCode0, orXXXXSBCAckCode1, orXXXXSBCAckCode2, orXXXXSBCAckCode3, orXXXXSTARTo, orXXXXEn_VCNTL, orXXXXVSACKo, orXXXXVACKo, orXXXXVTM0o, orXXXXVTM1o, orXXXXL_DBufo);
input
  GRANTi,
  LastRQSTi,
  PCCSawReset,
  TM0i,
  TM1i,
  TM1l,
  STARTi,
  STARTo,
  SBCResetPCC,
  SlotSpace_Id_Match,
  wdcntXXXXstate1,
  wdcntXXXXstate2,
  wdcntXXXXstate3,
  NuBusActive,
  RESETi,
  PCCsync,
  RQSTi,
  VSACKi,
  BUS_Inactive,
  VACKi,
  VACKl,
  SingleStep,
  PCCReqCode0,
  PCCReqCode1,
  PCCReqCode2,
  PCCReqCode3,
  PCCAck,
  PCCConfirm,
  ACKi,
  ACKl,
  PCCAckCode,
  CoherencyState1i,
  CoherencyState2i,
  PCCReq,
  physrecXXXXstate0,
  physrecXXXXstate1,
  VTM0i,
  VTM0l,
  VTM1l,
  Tag_Match;
output
  masterXXXXArb_active,
  orXXXXVSACKo,
  slaveXXXXGenerateNextState,
  masterXXXXEn_VDBufi,
  slaveXXXXL_VABufi,
  resetXXXXSBCResetPCC,
  orXXXXRESETo,
  slaveXXXXSnoopVTag_W,
  masterXXXXEn_ABufo,
  orXXXXSBCAck,
  orXXXXEn_VCNTL,
  resetXXXXReset,
  encodemuxXXXXMX_AD_8,
  masterXXXXEn_PDBufi,
  masterXXXXEn_PDBufo,
  physrecXXXXNextState0,
  physrecXXXXNextState1,
  slaveXXXXSBCReq,
  orXXXXVTM1o,
  orXXXXVTM0o,
  orXXXXL_DBufo,
  nextstateXXXXCoherencyState2o,
  orXXXXSBCAckCodelatch,
  slaveXXXXSnoopVTagState_R,
  masterXXXXL_PDBufi,
  wdcntXXXXNextState1,
  wdcntXXXXNextState2,
  wdcntXXXXNextState3,
  virmachXXXXSBCCacheRelease,
  orXXXXEn_CNTL,
  slaveXXXXSBCReqCode0,
  slaveXXXXSBCReqCode1,
  slaveXXXXSBCReqCode2,
  wdcntXXXXwd_cnt0,
  wdcntXXXXwd_cnt1,
  wdcntXXXXwd_cnt2,
  orXXXXACKo,
  orXXXXSTARTo,
  virmachXXXXEn_VDBufo,
  slaveXXXXSnoopAddrFromProc,
  nubusXXXXNuBusActive,
  virmachXXXXSBCsetDirty,
  orXXXXTM1o,
  virmachXXXXSBCConfigure,
  masterXXXXRQSTo,
  orXXXXTM0o,
  slaveXXXXSnoopState_W,
  masterXXXXL_DBufo_if_TM0,
  orXXXXEn_START,
  orXXXXVACKo,
  orXXXXSBCAckCode0,
  orXXXXSBCAckCode1,
  orXXXXSBCAckCode2,
  orXXXXSBCAckCode3,
  nubusXXXXL_PABufi,
  masterXXXXSBC_WriteCache;
reg
  wd_cnt_test,
  nubusXXXXstate0,
  nubusXXXXstate1,
  Set_ex_wd_cnt1,
  Incr_wd_cnt,
  Intr_done,
  wdcntXXXXstate0,
  slaveXXXXstate0,
  slaveXXXXstate1,
  slaveXXXXstate2,
  Reset_wd_cnt,
  P_receive_cancel,
  resetXXXXstate0,
  resetXXXXstate1,
  resetXXXXstate2,
  Intr_req,
  V_transmit_begin,
  UpdateReq,
  virmachXXXXstate0,
  virmachXXXXstate1,
  masterXXXXstate0,
  masterXXXXstate1,
  masterXXXXstate2,
  masterXXXXstate3,
  UpdateDone,
  P_receive_begin,
  Gen_Reset;
wire
  \[10936]_inv ,
  \[15357] ,
  \[15446] ,
  \[15541] ,
  \[15079] ,
  \[10899]_inv ,
  \{physrecXXXXNextState1} ,
  \[15074] ,
  \[15637] ,
  \[10748]_inv ,
  I515,
  I516,
  I88,
  \[14627]* ,
  I91,
  \[15353] ,
  \{masterXXXXNextState1} ,
  \[15452] ,
  \[10307] ,
  I536,
  \{masterXXXXNextState2} ,
  I537,
  I543,
  \[15355] ,
  \{masterXXXXNextState3} ,
  \[14411] ,
  \[14508] ,
  \[15081] ,
  \[10573]_inv ,
  \[15362] ,
  \[15266] ,
  \{orXXXXSBCAckCodelatch} ,
  \{masterXXXXNextState0} ,
  I599,
  \[14503] ,
  \[15545] ,
  \{nubusXXXXNuBusActive} ,
  \[14417] ,
  \[84] ,
  \[15550] ,
  \[85] ,
  \{orXXXXVSACKo} ,
  \[14505] ,
  \[15176] ,
  \[14419] ,
  \[86] ,
  \[14797]* ,
  \[15367] ,
  \[87] ,
  \[15456] ,
  \[15089] ,
  \[88] ,
  \[14512] ,
  \[15369] ,
  \[89] ,
  \[15182] ,
  \[10126] ,
  \[15085] ,
  \[15558] ,
  \[15643] ,
  \[10696]_inv ,
  \[15646] ,
  \[14421] ,
  \[14603] ,
  \{orXXXXL_DBufo} ,
  \[14517] ,
  \[15091] ,
  \[90] ,
  \[15276] ,
  \[91] ,
  \[10749]_inv ,
  \[15553] ,
  \[92] ,
  \{slaveXXXXNextState1} ,
  \[15280] ,
  \[93] ,
  \[15184] ,
  \{slaveXXXXNextState2} ,
  \[94] ,
  \[10923]_inv ,
  \[15560] ,
  \[95] ,
  \[15097] ,
  \{slaveXXXXNextState0} ,
  \[96] ,
  \[15377] ,
  \[97] ,
  \[100] ,
  \[10921]_inv ,
  \[14709] ,
  \[15658] ,
  \[15190] ,
  \[98] ,
  \[101] ,
  \[15465] ,
  \[10458]_inv ,
  \[15379] ,
  \[99] ,
  \[102] ,
  \[14521] ,
  \[10823]_inv ,
  \[15192] ,
  \[14802] ,
  \[2536] ,
  \[103] ,
  \[14617] ,
  \[15288] ,
  \[2537] ,
  \[104] ,
  \[10327] ,
  \[105] ,
  \[15471] ,
  \[14619] ,
  \[10821]_inv ,
  \[15653] ,
  \[106] ,
  \[10721]_inv ,
  \[107] ,
  \[15655] ,
  \[15284] ,
  \[108] ,
  \[15569] ,
  \[10422] ,
  \[10817]_inv ,
  \[14711] ,
  \[10662]_inv ,
  \[15198] ,
  \[14808] ,
  \[15382] ,
  \[109] ,
  \[1] ,
  \[10483]_inv ,
  \[14529] ,
  \[2] ,
  masterXXXXACKo,
  \[15566] ,
  \[15661] ,
  \[3] ,
  \[10658]_inv ,
  \[10946]_inv ,
  \[15290] ,
  \[14900] ,
  \[14523] ,
  \[4] ,
  \[14804] ,
  \[5] ,
  \[15292] ,
  \[14902] ,
  \[14525] ,
  \[14717] ,
  \[6] ,
  \[15572] ,
  \[7] ,
  \[15668] ,
  \[8] ,
  \[111] ,
  \[14862]* ,
  \[9] ,
  \[15389] ,
  \[14531] ,
  \[14627] ,
  \[15298] ,
  \[10930]_inv ,
  \[15481] ,
  \[15663] ,
  \[10339] ,
  \[15577] ,
  \[14909] ,
  \[14441] ,
  \{resetXXXXNextState1} ,
  \[15665] ,
  \[15294] ,
  \[14537] ,
  \{resetXXXXNextState2} ,
  \[15670] ,
  \[15574] ,
  \[15296] ,
  \[15391] ,
  \[14539] ,
  \[10335] ,
  \[15487] ,
  \[14448] ,
  \[10877]_inv ,
  \[14533] ,
  \[10061] ,
  \[15489] ,
  \[10912]_inv ,
  \[14535] ,
  \[14816] ,
  \[1048] ,
  \[14911] ,
  \[15582] ,
  \[10718] ,
  \[10525] ,
  \[14443] ,
  \[10612]_inv ,
  \[10908]_inv ,
  \[15399] ,
  \[14541] ,
  \[14723] ,
  \[14726] ,
  \[14821] ,
  \[14450] ,
  \[15393] ,
  \[15492] ,
  \[10559]_inv ,
  \[2836] ,
  \[15674] ,
  \[14917] ,
  \[15396] ,
  \[14730] ,
  \[14634] ,
  \[15587] ,
  \[2838] ,
  \[15676] ,
  \{resetXXXXSBCResetPCC} ,
  \[14547] ,
  \[15680] ,
  \[10933]_inv ,
  \[14640] ,
  \[13378]_inv ,
  \[14915] ,
  \[14543] ,
  \[15499] ,
  \[10890]_inv ,
  \[14823] ,
  \[14922] ,
  \[14737] ,
  \[10533] ,
  \[10632] ,
  \[15591] ,
  \[14830] ,
  \[15495] ,
  \[14733] ,
  \[14928] ,
  \[15686] ,
  \{orXXXXIncr_wd_cnt} ,
  \[14924] ,
  \[15599] ,
  \{orXXXXSBCAckCode1} ,
  \[14838] ,
  \{orXXXXSBCAckCode2} ,
  \{nubusXXXXNextState0} ,
  \[15692] ,
  \{orXXXXSBCAckCode3} ,
  \[10640] ,
  \[14467] ,
  \{nubusXXXXNextState1} ,
  \[14747] ,
  \[14469] ,
  \{orXXXXSBCAckCode0} ,
  \[10940]_inv ,
  \[15697] ,
  \[10089] ,
  \[14659] ,
  \[14654] ,
  \[10924]_inv ,
  \[14567] ,
  \[10363] ,
  \[14751] ,
  \[10624]_inv ,
  \{orXXXXTM1o} ,
  \[14940] ,
  \[14478] ,
  \[10918]_inv ,
  \[14661] ,
  \[14942] ,
  \[14757] ,
  \[14846] ,
  \[10822]_inv ,
  \[14387] ,
  \[14571] ,
  \[14668] ,
  \[14852] ,
  \[14480] ,
  \[10506]_inv ,
  \[10190] ,
  \[10943]_inv ,
  \[14760] ,
  \[13753]_inv ,
  \[14944] ,
  \[14666] ,
  \[10643]_inv ,
  \[14857] ,
  \[10653] ,
  \[14946] ,
  \[10375] ,
  \[10937]_inv ,
  \[14950] ,
  \[14488] ,
  \[530] ,
  \{orXXXXEn_CNTL} ,
  \[14952] ,
  \[14575] ,
  \[14767] ,
  \[14484] ,
  \[14769] ,
  \[10682]_inv ,
  \[14860] ,
  \[14764] ,
  \[10882]_inv ,
  \[14862] ,
  \[14490] ,
  \[10878]_inv ,
  \{slaveXXXXL_VABufi} ,
  \[14492] ,
  \[14674] ,
  \[14959] ,
  \{orXXXXSBCAck} ,
  \[15003] ,
  \[14676] ,
  \[14771] ,
  \[10866]_inv ,
  \[10819]_inv ,
  \[14955] ,
  \[14676]* ,
  \{virmachXXXXNextState1} ,
  \[15011] ,
  \[14681] ,
  \[10] ,
  \[10296] ,
  \[14585] ,
  \[11] ,
  \[12] ,
  \[14494] ,
  \[15109] ,
  \{virmachXXXXNextState0} ,
  \[13] ,
  \[10580] ,
  \[14] ,
  \[14496] ,
  \[14688] ,
  \[15] ,
  \[10750]_inv ,
  \[10934]_inv ,
  \[15017] ,
  \[14871] ,
  \[16] ,
  \[10897]_inv ,
  \[15105] ,
  \[17] ,
  \{virmachXXXXSBCConfigure} ,
  \[10685]_inv ,
  \[18] ,
  \[14857]* ,
  \[10932]_inv ,
  \[10492] ,
  \[14781] ,
  \[14963] ,
  \[10928]_inv ,
  \{wdcntXXXXwd_cnt_test} ,
  \[14966] ,
  \{orXXXXEn_START} ,
  \[14879] ,
  \[15300] ,
  \[14970] ,
  \[14593] ,
  \[15021] ,
  \[15302] ,
  \[14972] ,
  \[14595] ,
  \[15206] ,
  \[10497] ,
  \[10586] ,
  \[14902]* ,
  \[10816]_inv ,
  \[14698] ,
  \[10493] ,
  \[15211] ,
  \[10591] ,
  \[15120] ,
  \[14984]* ,
  \[14693] ,
  \[10651]_inv ,
  \[15304] ,
  \[15026] ,
  \[14976] ,
  \[15030] ,
  \[10935]_inv ,
  \[15219] ,
  \[10894]_inv ,
  \[15310] ,
  \[14980] ,
  \[14883] ,
  \[14982] ,
  \[14797] ,
  \[15215] ,
  \[10688]_inv ,
  \[15407] ,
  \[15129] ,
  \[10929]_inv ,
  \[10888]_inv ,
  \[15123] ,
  \[15037] ,
  \[15403] ,
  \[14987] ,
  \[15039] ,
  \{orXXXXReset_wd_cnt_x} ,
  \[15405] ,
  I105,
  \[15319] ,
  I108,
  \[15410] ,
  I109,
  \[14984] ,
  \[15228] ,
  I126,
  I128,
  \[15412] ,
  \[15035] ,
  I130,
  I131,
  \[14897] ,
  I139,
  \[15508] ,
  I140,
  \[14990] ,
  I163,
  I164,
  I167,
  \[10901]_inv ,
  \[15041] ,
  I172,
  \[15223] ,
  I173,
  I177,
  I179,
  \[15137] ,
  I187,
  I188,
  \[15418] ,
  \[10944]_inv ,
  I192,
  \{orXXXXEn_VCNTL} ,
  I193,
  \[15030]* ,
  I199,
  \[10703]_inv ,
  \[15506] ,
  \[15230] ,
  \[15510] ,
  \[15133] ,
  \[15232] ,
  \[10544]_inv ,
  \{orXXXXRESETo} ,
  \[15512] ,
  \[15135] ,
  \[15327] ,
  \[14997] ,
  \[15416] ,
  \[10938]_inv ,
  I201,
  \[15329] ,
  I207,
  I208,
  I211,
  I214,
  I215,
  I219,
  \[15046] ,
  \{orXXXXACKo} ,
  \[15141] ,
  I220,
  I222,
  I223,
  \[14993] ,
  I229,
  \[15604] ,
  \[10889]_inv ,
  I231,
  I232,
  I235,
  I236,
  \[15050] ,
  \[15702] ,
  \{slaveXXXXSBCReq} ,
  \[15052] ,
  \[15148] ,
  \{nubusXXXXL_PABufi} ,
  I273,
  I276,
  I279,
  \{slaveXXXXSnoopState_W} ,
  I280,
  I282,
  I284,
  I285,
  I287,
  I288,
  I292,
  \[15235] ,
  I295,
  I296,
  \[15427] ,
  I299,
  \[15240] ,
  \[15707] ,
  \[15143] ,
  \[10863]_inv ,
  \[15338] ,
  \[15521] ,
  \[15425] ,
  \{orXXXXVTM0o} ,
  \[15054] ,
  I300,
  I304,
  \[10657]_inv ,
  I305,
  \[10945]_inv ,
  \[15334] ,
  \[15056] ,
  \[15710] ,
  I322,
  I323,
  \[15614] ,
  \[15247] ,
  \[15336] ,
  I340,
  I341,
  \[15712] ,
  I348,
  \{slaveXXXXSBCReqCode0} ,
  I354,
  \[10845]_inv ,
  I357,
  \{masterXXXXSBC_WriteCache} ,
  I361,
  I363,
  I364,
  I366,
  \[10939]_inv ,
  I368,
  I369,
  \[15529] ,
  I373,
  I374,
  I377,
  \[10686]_inv ,
  \{orXXXXVACKo} ,
  I398,
  I399,
  \[15526] ,
  \[15159] ,
  \[10886]_inv ,
  \[15439] ,
  \[15068] ,
  \[15252] ,
  \{slaveXXXXSBCReqCode1} ,
  \[15064] ,
  \[15349] ,
  \[15344] ,
  \[15066] ,
  \[15442] ,
  \[10911]_inv ,
  \[15624] ,
  \[10703]_inv* ,
  \[15538] ,
  \{masterXXXXUpdateReq} ,
  \[10813]_inv ,
  I450,
  I451,
  I453,
  \[10907]_inv ,
  I465,
  \[10511]_inv ,
  I475,
  I476,
  \[15536] ,
  \[10507]_inv ,
  \[10854]_inv ,
  \[15169] ,
  \[15444] ,
  masterXXXXVSACKo,
  \[14409] ;
assign
  \[10936]_inv  = RESETi | slaveXXXXstate0,
  \[15357]  = \[15712]  & ~\[15529] ,
  \[15446]  = ~\[10923]_inv  & nubusXXXXstate1,
  \[15541]  = ~Intr_done & nubusXXXXstate1,
  \[15079]  = ~\[15637]  & ~\[15319] ,
  \[10899]_inv  = RQSTi | SingleStep,
  \{physrecXXXXNextState1}  = I287 | I288,
  \[15074]  = ~\[15355]  & ~masterXXXXstate1,
  \[15637]  = STARTi & VSACKi,
  masterXXXXArb_active = \[14529] ,
  \[10748]_inv  = \[10813]_inv  | ~PCCReqCode3,
  I515 = STARTi & ACKi,
  I516 = ~\[10912]_inv  & slaveXXXXstate0,
  I88 = ~\[10483]_inv  & PCCReqCode2,
  \[14627]*  = ~\[14627] ,
  I91 = ~\[10889]_inv  & \[10089] ,
  \[15353]  = ~\[15712]  & CoherencyState1i,
  \{masterXXXXNextState1}  = ~\[14411]  | I91,
  \[15452]  = ~\[10946]_inv  & ~virmachXXXXstate1,
  \[10307]  = \[2536]  | I377,
  orXXXXVSACKo = \{orXXXXVSACKo} ,
  I536 = PCCReqCode2 & ~PCCReqCode0,
  \{masterXXXXNextState2}  = ~\[14769]  | ~\[14419] ,
  I537 = ~PCCReqCode2 & PCCReqCode0,
  I543 = VTM0l & ~STARTo,
  \[15355]  = ~\[15661]  & ~\[10894]_inv ,
  \{masterXXXXNextState3}  = I108 | I109,
  \[14411]  = ~\[14448]  & \[14902] ,
  \[14508]  = ~\[14917]  & (~\[2838]  & ~\[14723] ),
  \[15081]  = ~\[15298]  & ~\[15439] ,
  \[10573]_inv  = \[10929]_inv  | (\[15329]  | (masterXXXXstate1 | \[10882]_inv )),
  \[15362]  = ~\[15558]  & ~\[10901]_inv ,
  \[15266]  = ~\[2537]  & ~physrecXXXXstate0,
  \{orXXXXSBCAckCodelatch}  = \[2836]  | (\[15041]  | (\[14469]  | \[15336] )),
  \{masterXXXXNextState0}  = \[14541]  | (\[15247]  | \[10632] ),
  I599 = ~P_receive_cancel & ~TM0i,
  \[14503]  = ~\[14802]  & (~\[14640]  & (~\[2838]  & ~\[14717] )),
  \[15545]  = masterXXXXstate1 & masterXXXXstate3,
  \{nubusXXXXNuBusActive}  = \[14990]  | \[15240] ,
  \[14417]  = \[14443]  & PCCReqCode1,
  \[84]  = \{masterXXXXNextState0} ,
  \[15550]  = ~PCCReqCode2 & PCCReqCode1,
  \[85]  = \{masterXXXXNextState1} ,
  \{orXXXXVSACKo}  = ~\[14698]  | ~\[14387] ,
  \[14505]  = ~\[15550]  & \[10507]_inv ,
  \[15176]  = ~\[15412]  & ~\[15574] ,
  \[14419]  = ~\[15105]  & (~\[14492]  & ~\[14757] ),
  \[86]  = \{masterXXXXNextState2} ,
  \[14797]*  = ~\[14797] ,
  \[15367]  = ~\[15680]  & PCCsync,
  \[87]  = \{masterXXXXNextState3} ,
  \[15456]  = ~\[10890]_inv  & Incr_wd_cnt,
  \[15089]  = ~\[15353]  & ~CoherencyState2i,
  \[88]  = \{nubusXXXXNextState0} ,
  \[14512]  = ~\[10507]_inv  & ~PCCReqCode2,
  \[15369]  = ~\[15697]  & ~\[15550] ,
  \[89]  = \{nubusXXXXNextState1} ,
  \[15182]  = ~\[10918]_inv  & ~\[15349] ,
  \[10126]  = I536 | I537,
  \[15085]  = ~\[15288]  & \[15418] ,
  \[15558]  = ~VSACKi & STARTi,
  \[15643]  = PCCReqCode1 & ~PCCReqCode0,
  \[10696]_inv  = \[10335]  | \[15707] ,
  \[15646]  = ~masterXXXXstate2 & ~masterXXXXstate1,
  \[14421]  = ~\[14862]  & \[14450] ,
  \[14603]  = ~\[14711]  & ~VSACKi,
  \{orXXXXL_DBufo}  = \[14952]  | (\[15159]  | (\[14450]  | \[14441] )),
  \[14517]  = ~\[10586]  & ~\[14575] ,
  \[15091]  = ~\[15284]  & ~PCCReqCode3,
  \[90]  = \{slaveXXXXNextState0} ,
  \[15276]  = ~\[10888]_inv  & (~\[10939]_inv  & (~nubusXXXXstate1 & ACKi)),
  \[91]  = \{slaveXXXXNextState1} ,
  \[10749]_inv  = ~\[15344]  | SingleStep,
  \[15553]  = slaveXXXXstate0 & ~RESETi,
  \[92]  = \{slaveXXXXNextState2} ,
  \{slaveXXXXNextState1}  = ~\[14478]  | I105,
  \[15280]  = ~\[10912]_inv  & (~\[10908]_inv  & ~slaveXXXXstate2),
  \[93]  = \[14976] ,
  \[15184]  = \[15452]  & ~PCCAckCode,
  \{slaveXXXXNextState2}  = ~\[14484]  | I126,
  \[94]  = \{resetXXXXNextState1} ,
  \[10923]_inv  = nubusXXXXstate0 | ~SlotSpace_Id_Match,
  \[15560]  = resetXXXXstate1 & ~PCCSawReset,
  \[95]  = \{resetXXXXNextState2} ,
  slaveXXXXGenerateNextState = \[14676]* ,
  \[15097]  = ~\[10877]_inv  & ~\[15294] ,
  \{slaveXXXXNextState0}  = I130 | I131,
  \[96]  = \{virmachXXXXNextState0} ,
  \[15377]  = ~\[15541]  & \[10923]_inv ,
  \[97]  = \{virmachXXXXNextState1} ,
  \[100]  = \[14883] ,
  \[10921]_inv  = slaveXXXXstate2 | ~STARTi,
  \[14709]  = ~\[15452]  & ~\[14852] ,
  \[15658]  = ~resetXXXXstate1 & ~resetXXXXstate0,
  \[15190]  = ~\[15489]  & \[10936]_inv ,
  \[98]  = \[15030]* ,
  \[101]  = \[15190] ,
  \[15465]  = \[15686]  & PCCReqCode0,
  \[10458]_inv  = ~\[10483]_inv  | \[15614] ,
  \[15379]  = \[15646]  & ~\[15702] ,
  \[99]  = \[14627]* ,
  \[102]  = \{masterXXXXUpdateReq} ,
  \[14521]  = ~\[10822]_inv  & ~\[14603] ,
  \[10823]_inv  = masterXXXXstate3 | \[10932]_inv ,
  \[15192]  = ~\[15481]  & ~\[13753]_inv ,
  \[14802]  = ~\[10918]_inv  & ~\[10685]_inv ,
  \[2536]  = I450 | I451,
  \[103]  = \[14681] ,
  \[14617]  = ~\[14666]  & masterXXXXstate3,
  \[15288]  = ~\[15624]  & Incr_wd_cnt,
  \[2537]  = I599 | ~wd_cnt_test,
  \[104]  = \{orXXXXReset_wd_cnt_x} ,
  \[10327]  = I368 | I369,
  \[105]  = \[14467] ,
  \[15471]  = ~\[10921]_inv  & ~slaveXXXXstate1,
  \[14619]  = ~\[15021]  & ~\[14730] ,
  \[10821]_inv  = ~\[15646]  | ~masterXXXXstate3,
  \[15653]  = ~VSACKi & ~STARTi,
  \[106]  = \{orXXXXIncr_wd_cnt} ,
  \[10721]_inv  = I543 | ~STARTi,
  \[107]  = \{wdcntXXXXwd_cnt_test} ,
  \[15655]  = ~TM1l & CoherencyState2i,
  \[15284]  = ~\[15686]  & ~SingleStep,
  masterXXXXEn_VDBufi = \[14902]* ,
  \[108]  = \[14443] ,
  \[15569]  = ~PCCReqCode1 & PCCReqCode0,
  \[10422]  = I515 | I516,
  \[10817]_inv  = \[10889]_inv  | ~masterXXXXstate3,
  \[14711]  = ~\[14871]  & masterXXXXstate2,
  \[10662]_inv  = ~\[10888]_inv  | \[10307] ,
  \[15198]  = ~\[15569]  & (~PCCReqCode3 & ~PCCReqCode2),
  \[14808]  = ~\[14987]  & ~\[15159] ,
  \[15382]  = ~\[15574]  & VACKl,
  \[109]  = \[15017] ,
  \[1]  = ~\[10339]  | ~\[14537] ,
  \[10483]_inv  = PCCReqCode1 | \[10507]_inv ,
  \[14529]  = ~\[14595]  & ~SBCResetPCC,
  \[2]  = ~\[15465]  | ~\[14911] ,
  masterXXXXACKo = \[10506]_inv  | ~\[15041] ,
  \[15566]  = masterXXXXstate2 & ~VSACKi,
  \[15661]  = masterXXXXstate3 & ~SingleStep,
  \[3]  = ~\[15396]  | ~\[14823] ,
  \[10658]_inv  = ~\[10899]_inv  | \[15512] ,
  \[10946]_inv  = ~virmachXXXXstate0 | SBCResetPCC,
  \[15290]  = ~\[15521]  & VSACKi,
  \[14900]  = ~\[10422]  & \[7] ,
  slaveXXXXL_VABufi = \{slaveXXXXL_VABufi} ,
  \[14523]  = ~\[10749]_inv  & (~\[14668]  & ~SBCResetPCC),
  \[4]  = ~\[10924]_inv  | ~\[15074] ,
  \[14804]  = ~\[15120]  & ~\[10750]_inv ,
  \[5]  = ~\[10819]_inv  | \[15655] ,
  \[15292]  = ~\[15521]  & ~\[15591] ,
  \[14902]  = \[8]  & \[10889]_inv ,
  \[14525]  = ~\[15302]  & ~\[10533] ,
  \[14717]  = \[14897]  & PCCReqCode0,
  \[6]  = ~\[15109]  | ~\[15247] ,
  \[15572]  = P_receive_cancel & ~physrecXXXXstate0,
  \[7]  = ~\[15425]  | NuBusActive,
  \[15668]  = ~wdcntXXXXstate3 & ~wdcntXXXXstate2,
  \[8]  = ~\[15382]  | ~\[15017] ,
  \[111]  = \[14852] ,
  \[14862]*  = ~\[14862] ,
  \[9]  = ~\[15037]  | ~masterXXXXstate2,
  \[15389]  = ~\[15670]  & ~\[15541] ,
  \[14531]  = ~\[14593]  & ~SBCResetPCC,
  \[14627]  = ~\[14879]  & \[2] ,
  \[15298]  = ~\[15572]  & physrecXXXXstate1,
  \[10930]_inv  = ~PCCReqCode3 | ~PCCReq,
  \[15481]  = \[18]  & ~virmachXXXXstate1,
  \[15663]  = ~P_receive_cancel & ~TM1i,
  \[10339]  = I279 | I280,
  \[15577]  = slaveXXXXstate1 & slaveXXXXstate2,
  \[14909]  = \[9]  & UpdateDone,
  \[14441]  = ~\[14496]  & ~PCCReqCode2,
  \{resetXXXXNextState1}  = \[15676]  | I292,
  \[15665]  = P_receive_cancel & physrecXXXXstate1,
  \[15294]  = ~\[15526]  & STARTi,
  \[14537]  = \[10061]  & (\[15553]  & slaveXXXXstate2),
  \{resetXXXXNextState2}  = \[15676]  | I354,
  \[15670]  = ~nubusXXXXstate1 & nubusXXXXstate0,
  \[15574]  = ~masterXXXXstate3 & masterXXXXstate1,
  \[15296]  = ~\[10945]_inv  & ~\[15582] ,
  \[15391]  = ~\[15541]  & ~\[15692] ,
  \[14539]  = ~\[13378]_inv  & slaveXXXXstate2,
  \[10335]  = I284 | I285,
  \[15487]  = Incr_wd_cnt & (wdcntXXXXstate3 & ~wdcntXXXXstate1),
  \[14448]  = ~\[14488]  & ~SBCResetPCC,
  \[10877]_inv  = slaveXXXXstate1 | slaveXXXXstate2,
  \[14533]  = ~\[14760]  & ~\[14585] ,
  \[10061]  = I235 | I236,
  resetXXXXSBCResetPCC = \{resetXXXXSBCResetPCC} ,
  \[15489]  = ~slaveXXXXstate2 & (slaveXXXXstate1 & PCCAck),
  orXXXXRESETo = \{orXXXXRESETo} ,
  \[10912]_inv  = STARTi | ACKi,
  \[14535]  = ~\[10749]_inv  & (~\[14688]  & ~SBCResetPCC),
  \[14816]  = ~\[10685]_inv  & ~SBCResetPCC,
  \[1048]  = I299 | I300,
  \[14911]  = ~\[10935]_inv  & (~\[15230]  & (physrecXXXXstate1 & ~physrecXXXXstate0)),
  \[15582]  = physrecXXXXstate0 & physrecXXXXstate1,
  \[10718]  = I322 | I323,
  \[10525]  = ~\[14709]  | I167,
  \[14443]  = ~\[14512]  & PCCReqCode0,
  \[10612]_inv  = P_receive_cancel | (\[10945]_inv  | \[10911]_inv ),
  \[10908]_inv  = slaveXXXXstate0 | slaveXXXXstate1,
  \[15399]  = ~\[15653]  & ~\[15637] ,
  \[14541]  = ~\[10296]  & SBCResetPCC,
  \[14723]  = ~\[15232]  & ~\[10643]_inv ,
  \[14726]  = ~\[10544]_inv  & \[4] ,
  \[14821]  = ~\[15643]  & (~\[15091]  & (~\[15614]  & PCCReq)),
  \[14450]  = ~\[14505]  & ~PCCReqCode0,
  \[15393]  = \[15591]  & ~masterXXXXstate3,
  slaveXXXXSnoopVTag_W = \[14681] ,
  \[15492]  = P_receive_cancel & (~virmachXXXXstate1 & ~virmachXXXXstate0),
  \[10559]_inv  = \[10912]_inv  | I361,
  \[2836]  = \[14816]  | (\[15604]  | \[15052] ),
  \[15674]  = ~TM0i & ~STARTi,
  \[14917]  = ~\[10748]_inv  & PCCReqCode0,
  \[15396]  = \[15646]  & ~RQSTi,
  \[14730]  = ~\[15512]  & (~\[10657]_inv  & (~RQSTi & ~PCCReqCode3)),
  \[14634]  = ~\[10934]_inv  & (~\[14900]  & (~Intr_req & slaveXXXXstate2)),
  \[15587]  = VSACKi & ~STARTi,
  \[2838]  = \[1048]  | I201,
  \[15676]  = RESETi & resetXXXXstate2,
  \{resetXXXXSBCResetPCC}  = resetXXXXstate0 | (resetXXXXstate2 | (RESETi | \[15560] )),
  \[14547]  = ~\[14982]  & (~\[14917]  & (~\[1048]  & ~\[14897] )),
  \[15680]  = ~Intr_req & ~SlotSpace_Id_Match,
  \[10933]_inv  = ~NuBusActive | STARTi,
  \[14640]  = ~\[15344]  & (~\[10643]_inv  & PCCConfirm),
  \[13378]_inv  = \[10061]  | I177,
  \[14915]  = ~\[15056]  & ~\[15553] ,
  \[14543]  = \[10375]  & (\[15553]  & ~slaveXXXXstate1),
  masterXXXXEn_ABufo = \[14535] ,
  \[15499]  = virmachXXXXstate1 & (virmachXXXXstate0 & ~VACKi),
  \[10890]_inv  = ~Reset_wd_cnt | ~SBCResetPCC,
  \[14823]  = \[15021]  & PCCConfirm,
  \[14922]  = ~\[15074]  & ~RQSTi,
  \[14737]  = ~\[15026]  & (VTM0i & ~SBCResetPCC),
  \[10533]  = ~\[14661]  | I179,
  \[10632]  = I219 | I220,
  \[15591]  = masterXXXXstate2 & ~STARTi,
  \[14830]  = ~\[14980]  & ~physrecXXXXstate0,
  \[15495]  = ~\[10877]_inv  & ~PCCsync,
  \[14733]  = ~\[15382]  & (~\[15362]  & (~\[10640]  & ~\[10089] )),
  \[14928]  = ~\[10945]_inv  & \[10] ,
  \[15686]  = ~PCCReqCode2 & ~PCCReqCode1,
  \{orXXXXIncr_wd_cnt}  = \[15066]  | (\[15159]  | (\[14737]  | \[15054] )),
  orXXXXSBCAck = \{orXXXXSBCAck} ,
  orXXXXEn_VCNTL = \{orXXXXEn_VCNTL} ,
  \[14924]  = ~\[15079]  & ~ACKl,
  resetXXXXReset = \[15676] ,
  \[15599]  = ~VSACKi & VTM0i,
  \{orXXXXSBCAckCode1}  = I187 | I188,
  \[14838]  = ~\[14970]  & ~masterXXXXstate1,
  \{orXXXXSBCAckCode2}  = \[10492]  | \[10493] ,
  \{nubusXXXXNextState0}  = \[14990]  | I276,
  encodemuxXXXXMX_AD_8 = \[15198] ,
  \[15692]  = ~nubusXXXXstate1 & ~ACKi,
  \{orXXXXSBCAckCode3}  = ~\[14627]  | \[15604] ,
  \[10640]  = I340 | I341,
  \[14467]  = ~\[10126]  & \[10483]_inv ,
  \{nubusXXXXNextState1}  = \[15219]  | I211,
  masterXXXXEn_PDBufi = \[10703]_inv* ,
  masterXXXXEn_PDBufo = \[15247] ,
  \[14747]  = ~\[15182]  & ~\[10497] ,
  \[14469]  = ~\[14508]  & ~SBCResetPCC,
  \{orXXXXSBCAckCode0}  = \[14469]  | \[14911] ,
  \[10940]_inv  = nubusXXXXstate0 | ~STARTi,
  \[15697]  = ~PCCReqCode1 & ~PCCReqCode0,
  physrecXXXXNextState0 = \[14928] ,
  physrecXXXXNextState1 = \{physrecXXXXNextState1} ,
  \[10089]  = I475 | I476,
  \[14659]  = ~\[14771]  & ~\[15545] ,
  \[14654]  = ~\[10907]_inv  & (~\[14950]  & slaveXXXXstate2),
  \[10924]_inv  = masterXXXXstate0 | masterXXXXstate2,
  \[14567]  = ~\[14619]  & ~\[10937]_inv ,
  \[10363]  = I398 | I399,
  \[14751]  = ~\[10932]_inv  & (~\[15035]  & \[15143] ),
  \[10624]_inv  = \[10750]_inv  | ~TM1l,
  \{orXXXXTM1o}  = ~\[14421]  | I88,
  \[14940]  = ~\[10816]_inv  & (\[15344]  & PCCConfirm),
  \[14478]  = \[1]  & ~slaveXXXXstate1,
  slaveXXXXSBCReq = \{slaveXXXXSBCReq} ,
  \[10918]_inv  = TM1i | ~TM0i,
  \[14661]  = ~\[10653]  & (~\[15039]  & ~\[14966] ),
  \[14942]  = ~\[15097]  & ~\[15577] ,
  \[14757]  = ~\[10878]_inv  & ~\[14909] ,
  \[14846]  = ~\[14922]  & ~\[15545] ,
  \[10822]_inv  = ~\[15574]  | ~GRANTi,
  orXXXXVTM1o = \[14417] ,
  orXXXXVTM0o = \{orXXXXVTM0o} ,
  \[14387]  = ~\[15192]  & (~\[15159]  & (~masterXXXXVSACKo & ~\[14764] )),
  \[14571]  = ~\[15489]  & ~\[10718] ,
  \[14668]  = ~\[15137]  & ~\[14823] ,
  orXXXXL_DBufo = \{orXXXXL_DBufo} ,
  \[14852]  = \[15655]  & ~\[10750]_inv ,
  \[14480]  = ~\[14517]  & ~RQSTi,
  \[10506]_inv  = \[14723]  | ~SBCResetPCC,
  \[10190]  = I295 | I296,
  \[10943]_inv  = ~masterXXXXstate0 | ~ACKl,
  \[14760]  = ~\[10822]_inv  & (~\[15068]  & masterXXXXstate2),
  \[13753]_inv  = SBCResetPCC | virmachXXXXstate0,
  \[14944]  = ~\[15123]  & ~ACKl,
  \[14666]  = ~\[15338]  & (~\[15396]  & (~\[15379]  & ~\[14924] )),
  \[10643]_inv  = ~\[15021]  | SingleStep,
  \[14857]  = ~\[15442]  & ~\[15064] ,
  \[10653]  = I363 | I364,
  \[14946]  = ~\[15405]  & (~\[15471]  & ~\[15577] ),
  \[10375]  = I231 | I232,
  \[10937]_inv  = SBCResetPCC | SingleStep,
  \[14950]  = \[11]  & \[10908]_inv ,
  \[14488]  = ~\[14959]  & (~\[14726]  & ~\[14521] ),
  \[530]  = \[10894]_inv  | ~PCCConfirm,
  \{orXXXXEn_CNTL}  = I172 | I173,
  \[14952]  = ~\[15192]  & ~PCCAck,
  \[14575]  = ~\[14821]  & (~\[10882]_inv  & ~masterXXXXstate1),
  \[14767]  = ~\[15120]  & \[5] ,
  \[14484]  = ~\[14860]  & ~\[14543] ,
  \[14769]  = \[6]  & \[10889]_inv ,
  \[10682]_inv  = \[10907]_inv  | \[10921]_inv ,
  \[14860]  = ~\[10907]_inv  & (~\[15215]  & STARTi),
  \[14764]  = ~\[10877]_inv  & ~\[14915] ,
  \[10882]_inv  = ~masterXXXXstate3 | masterXXXXstate0,
  \[14862]  = ~\[15041]  & ~\[15219] ,
  \[14490]  = ~\[10591]  & ~\[14617] ,
  \[10878]_inv  = masterXXXXstate1 | (SBCResetPCC | masterXXXXstate0),
  \{slaveXXXXL_VABufi}  = \[14634]  | (\[15280]  | (RESETi | \[14674] )),
  \[14492]  = ~\[14533]  & ~SBCResetPCC,
  \[14674]  = ~\[14946]  & (~slaveXXXXstate0 & ACKi),
  \[14959]  = \[15223]  & STARTi,
  \{orXXXXSBCAck}  = \[2836]  | (masterXXXXACKo | (\[14494]  | \[14911] )),
  \[15003]  = \[15418]  & (Incr_wd_cnt & ~wdcntXXXXstate2),
  \[14676]  = ~\[14804]  & ~\[14852] ,
  \[14771]  = ~\[14955]  & ACKl,
  \[10866]_inv  = \[13753]_inv  | I465,
  \[10819]_inv  = \[10944]_inv  | (~\[15553]  | ~Tag_Match),
  \[14955]  = ~\[15290]  & (~\[15393]  & ~\[15566] ),
  \[14676]*  = ~\[14676] ,
  \{virmachXXXXNextState1}  = \[14987]  | I273,
  \[15011]  = ~\[10886]_inv  & (~\[10936]_inv  & (~\[10944]_inv  & ~slaveXXXXstate2)),
  \[14681]  = ~\[14942]  & (\[15707]  & (UpdateReq & ~RESETi)),
  \[10]  = ~\[15349]  | \[15439] ,
  \[10296]  = I214 | I215,
  \[14585]  = ~\[14838]  & (~\[10882]_inv  & ~masterXXXXstate2),
  \[11]  = ~\[15310]  | ~\[15252] ,
  \[12]  = ~\[15444]  | ~\[15329] ,
  \[14494]  = ~\[14547]  & ~SBCResetPCC,
  \[15109]  = ~\[15399]  & ~\[10901]_inv ,
  \{virmachXXXXNextState0}  = ~\[14808]  | I199,
  \[13]  = ~\[15710]  | ~\[15456] ,
  \[10580]  = ~\[10573]_inv  | I282,
  \[14]  = ~\[15499]  | ~\[15492] ,
  \[14496]  = ~\[15697]  & \[10507]_inv ,
  \[14688]  = \[3]  & \[10882]_inv ,
  \[15]  = ~\[15668]  | ~\[15410] ,
  \[10750]_inv  = \[10819]_inv  | ~slaveXXXXstate2,
  nextstateXXXXCoherencyState2o = \[15334] ,
  \[10934]_inv  = ~slaveXXXXstate1 | VSACKi,
  \[15017]  = \[15591]  & (~\[10817]_inv  & (VSACKi & VTM0i)),
  \[14871]  = ~\[15465]  & (\[15232]  & (~SingleStep & BUS_Inactive)),
  \[16]  = ~\[15637]  | ~\[15646] ,
  \[10897]_inv  = ~nubusXXXXstate1 | STARTi,
  \[15105]  = ~\[15338]  & \[10817]_inv ,
  \[17]  = ~\[15526]  | VTM0l,
  \{virmachXXXXSBCConfigure}  = \[14952]  | \[15452] ,
  \[10685]_inv  = \[10943]_inv  | I348,
  \[18]  = ~V_transmit_begin | P_receive_cancel,
  \[14857]*  = ~\[14857] ,
  \[10932]_inv  = ~masterXXXXstate2 | ~masterXXXXstate1,
  \[10492]  = I139 | I140,
  \[14781]  = ~\[14940]  & GRANTi,
  \[14963]  = ~\[15089]  & Tag_Match,
  \[10928]_inv  = ~masterXXXXstate3 | ~masterXXXXstate2,
  orXXXXSBCAckCodelatch = \{orXXXXSBCAckCodelatch} ,
  \{wdcntXXXXwd_cnt_test}  = ~\[10686]_inv  | ~\[15030] ,
  \[14966]  = ~\[10821]_inv  & \[12] ,
  \{orXXXXEn_START}  = ~\[15046]  | I128,
  slaveXXXXSnoopVTagState_R = \[14764] ,
  \[14879]  = ~\[10748]_inv  & ~SBCResetPCC,
  \[15300]  = ~\[15587]  & ~\[15599] ,
  \[14970]  = ~\[10899]_inv  & (~\[15369]  & ~\[10894]_inv ),
  \[14593]  = ~\[14993]  & (~\[15223]  & ~\[14693] ),
  \[15021]  = ~\[10822]_inv  & (\[15566]  & BUS_Inactive),
  \[15302]  = \[15582]  & P_receive_begin,
  \[14972]  = ~\[10938]_inv  & (~\[15391]  & STARTi),
  masterXXXXL_PDBufi = \[10703]_inv* ,
  \[14595]  = ~\[15235]  & (~\[14959]  & ~\[14693] ),
  \[15206]  = ~\[15536]  & (~\[15506]  & ~\[15707] ),
  \[10497]  = I373 | I374,
  \[10586]  = I304 | I305,
  wdcntXXXXNextState1 = \[14857]* ,
  wdcntXXXXNextState2 = \[14797]* ,
  wdcntXXXXNextState3 = \[14984]* ,
  \[14902]*  = ~\[14902] ,
  \[10816]_inv  = ~\[15702]  | ~BUS_Inactive,
  virmachXXXXSBCCacheRelease = \[15169] ,
  \[14698]  = ~\[15304]  & ~\[14767] ,
  \[10493]  = I222 | I223,
  \[15211]  = ~\[15499]  & ~\[15492] ,
  \[10591]  = I163 | I164,
  \[15120]  = ~\[15357]  & ~\[15529] ,
  \[14984]*  = ~\[14984] ,
  orXXXXEn_CNTL = \{orXXXXEn_CNTL} ,
  \[14693]  = ~\[10924]_inv  & ~\[14846] ,
  \[10651]_inv  = LastRQSTi | I453,
  \[15304]  = \[15553]  & (~slaveXXXXstate2 & ~PCCAck),
  \[15026]  = \[14]  & V_transmit_begin,
  \[14976]  = \[15407]  & (~resetXXXXstate2 & RESETi),
  slaveXXXXSBCReqCode0 = \{slaveXXXXSBCReqCode0} ,
  slaveXXXXSBCReqCode1 = \{slaveXXXXSBCReqCode1} ,
  slaveXXXXSBCReqCode2 = \[14654] ,
  \[15030]  = ~\[15508]  & \[15] ,
  \[10935]_inv  = ~ACKi | SBCResetPCC,
  wdcntXXXXwd_cnt0 = \[14984]* ,
  wdcntXXXXwd_cnt1 = \[14797]* ,
  \[15219]  = ~\[10938]_inv  & (\[15692]  & (Intr_done & ~STARTi)),
  wdcntXXXXwd_cnt2 = \[14857]* ,
  \[10894]_inv  = PCCReqCode3 | ~PCCReq,
  \[15310]  = ~\[15680]  & ~PCCsync,
  \[14980]  = ~\[15135]  & wd_cnt_test,
  \[14883]  = ~\[10888]_inv  & (~\[15141]  & ~\[10912]_inv ),
  \[14982]  = ~\[15292]  & (~\[10943]_inv  & ~VSACKi),
  \[14797]  = ~\[15133]  & ~\[15003] ,
  \[15215]  = ~\[15495]  & ~\[15577] ,
  \[10688]_inv  = \[10327]  | ~Intr_done,
  \[15407]  = Gen_Reset & \[15658] ,
  orXXXXACKo = \{orXXXXACKo} ,
  \[15129]  = ~\[15403]  & ~resetXXXXstate2,
  \[10929]_inv  = masterXXXXstate2 | \[10930]_inv ,
  \[10888]_inv  = RESETi | Intr_done,
  \[15123]  = ~\[15338]  & ~masterXXXXstate1,
  \[15037]  = \[15686]  & (~\[10929]_inv  & ~PCCReqCode0),
  \[15403]  = ~\[15658]  & ~RESETi,
  orXXXXSTARTo = \[14567] ,
  \[14987]  = ~\[15211]  & ~SBCResetPCC,
  \[15039]  = ~\[15235]  & ~BUS_Inactive,
  \{orXXXXReset_wd_cnt_x}  = \[14496]  | (\[14512]  | (\[15011]  | \[15017] )),
  \[15405]  = ~\[15680]  & ~slaveXXXXstate2,
  I105 = ~\[10696]_inv  & ~RESETi,
  \[15319]  = \[15566]  & ~STARTi,
  I108 = ~\[14409]  & ~SBCResetPCC,
  \[15410]  = ~\[10890]_inv  & wdcntXXXXstate0,
  I109 = ~\[10889]_inv  & ~\[14490] ,
  \[14984]  = ~\[15085]  & \[13] ,
  \[15228]  = ~\[10946]_inv  & (virmachXXXXstate1 & (VACKi & VTM0i)),
  I126 = ~\[14571]  & ~RESETi,
  I128 = ~\[14525]  & ~SBCResetPCC,
  \[15412]  = ~\[10894]_inv  & ~masterXXXXstate3,
  \[15035]  = ~\[15643]  & (~\[530]  & (~\[15686]  & ~\[15614] )),
  I130 = ~\[10682]_inv  & ~\[10944]_inv ,
  I131 = ~\[14539]  & \[15553] ,
  \[14897]  = ~\[10748]_inv  & PCCReqCode2,
  I139 = ~\[14503]  & ~SBCResetPCC,
  \[15508]  = Set_ex_wd_cnt1 & (Reset_wd_cnt & (~wdcntXXXXstate1 & ~SBCResetPCC)),
  I140 = \[15604]  & ~resetXXXXstate1,
  virmachXXXXEn_VDBufo = \[15452] ,
  \[14990]  = ~\[15389]  & (~\[10907]_inv  & ~STARTi),
  I163 = ~\[14659]  & ~LastRQSTi,
  I164 = \[15545]  & ~ACKl,
  I167 = ~\[15148]  & ~\[10817]_inv ,
  \[10901]_inv  = ~masterXXXXstate2 | ACKl,
  \[15041]  = ~\[10821]_inv  & (\[15702]  & ~\[10889]_inv ),
  I172 = ~\[14661]  & ~SBCResetPCC,
  \[15223]  = \[15646]  & (~masterXXXXstate3 & masterXXXXstate0),
  I173 = ~\[10559]_inv  & ~RESETi,
  I177 = VSACKi & slaveXXXXstate1,
  I179 = ~\[14830]  & ~LastRQSTi,
  \[15137]  = ~\[10821]_inv  & ~RQSTi,
  I187 = \[14816]  & ~TM0i,
  I188 = ~\[10935]_inv  & \[10190] ,
  \[15418]  = ~\[10890]_inv  & wdcntXXXXstate3,
  \[10944]_inv  = slaveXXXXstate1 | ~VTM0l,
  I192 = \[14852]  & VTM1l,
  \{orXXXXEn_VCNTL}  = \[14523]  | (\[15192]  | \[10525] ),
  I193 = ~\[10624]_inv  & \[15529] ,
  \[15030]*  = ~\[15030] ,
  I199 = ~\[10866]_inv  & PCCAck,
  \[10703]_inv  = \[10817]_inv  | I229,
  \[15506]  = ~Intr_req & (NuBusActive & ~ACKi),
  \[15230]  = ~\[15663]  & ~\[2537] ,
  \[15510]  = CoherencyState1i & (CoherencyState2i & TM1l),
  \[15133]  = ~\[15487]  & ~\[10854]_inv ,
  \[15232]  = ~\[15512]  & ~\[530] ,
  \[10544]_inv  = \[10894]_inv  | I357,
  \{orXXXXRESETo}  = ~\[14627]  | (\[14972]  | \[15276] ),
  \[15512]  = PCCReqCode1 & PCCReqCode2,
  \[15135]  = ~\[15665]  & ~\[15427] ,
  \[15327]  = \[17]  & TM1l,
  \[14997]  = ~\[15206]  & ~slaveXXXXstate2,
  \[15416]  = ~\[10918]_inv  & ~P_receive_cancel,
  \[10938]_inv  = ~nubusXXXXstate0 | RESETi,
  I201 = \[14897]  & masterXXXXstate3,
  \[15329]  = \[15569]  & ~PCCReqCode2,
  I207 = ~\[10750]_inv  & \[15357] ,
  I208 = ~\[10624]_inv  & \[15529] ,
  I211 = ~\[10662]_inv  & ~ACKi,
  I214 = ~\[10823]_inv  & ~\[14781] ,
  I215 = \[15223]  & ~STARTi,
  I219 = ~\[14733]  & ~\[10889]_inv ,
  \[15046]  = ~\[15296]  & ~\[15247] ,
  \{orXXXXACKo}  = masterXXXXACKo | \[15219] ,
  \[15141]  = ~\[15670]  & ~\[15446] ,
  I220 = \[14730]  & ~\[10937]_inv ,
  I222 = ~\[10935]_inv  & ~\[14747] ,
  I223 = \[14816]  & \[15538] ,
  \[14993]  = ~\[10823]_inv  & ~\[15143] ,
  I229 = ~\[15109]  & ~\[14944] ,
  \[15604]  = resetXXXXstate2 & ~RESETi,
  \[10889]_inv  = ~masterXXXXstate0 | SBCResetPCC,
  I231 = ~slaveXXXXstate2 & ~PCCsync,
  I232 = ~\[14963]  & slaveXXXXstate2,
  I235 = ~\[14963]  & ~slaveXXXXstate1,
  I236 = ~\[15510]  & ~\[10944]_inv ,
  \[15050]  = ~\[15416]  & (~\[15538]  & (wd_cnt_test & ~physrecXXXXstate0)),
  \[15702]  = ~VSACKi & ~SingleStep,
  \{slaveXXXXSBCReq}  = ~\[14676]  | \[14654] ,
  \[15052]  = ~\[10878]_inv  & (UpdateDone & masterXXXXstate2),
  \[15148]  = \[16]  & \[10901]_inv ,
  \{nubusXXXXL_PABufi}  = \[10688]_inv  | ~RESETi,
  I273 = ~\[10866]_inv  & ~PCCAck,
  I276 = ~\[10863]_inv  & ~TM1i,
  I279 = ~\[10933]_inv  & ~\[10907]_inv ,
  \{slaveXXXXSnoopState_W}  = ~\[14676]  | \[14681] ,
  slaveXXXXSnoopAddrFromProc = \[14681] ,
  I280 = ~\[14997]  & ~RESETi,
  I282 = ~\[10928]_inv  & masterXXXXstate1,
  I284 = ~\[10921]_inv  & ~\[15327] ,
  I285 = ~\[15367]  & slaveXXXXstate2,
  I287 = ~\[10945]_inv  & ~\[15081] ,
  I288 = ~\[10845]_inv  & \[15582] ,
  I292 = ~\[15129]  & ~PCCSawReset,
  \[15235]  = ~\[10823]_inv  & GRANTi,
  I295 = ~\[15349]  & ~TM0i,
  I296 = ~\[15050]  & physrecXXXXstate1,
  nubusXXXXNuBusActive = \{nubusXXXXNuBusActive} ,
  \[15427]  = ~\[10911]_inv  & TM1i,
  I299 = ~\[10658]_inv  & ~\[10657]_inv ,
  \[15240]  = ~\[10863]_inv  & (~Intr_done & ~nubusXXXXstate1),
  \[15707]  = ~slaveXXXXstate0 & ~ACKi,
  \[15143]  = ~\[10816]_inv  & GRANTi,
  \[10863]_inv  = \[10940]_inv  | \[10907]_inv ,
  \[15338]  = ~\[15599]  & ~masterXXXXstate2,
  \[15521]  = VACKl & masterXXXXstate1,
  \[15425]  = ~\[10933]_inv  & ACKi,
  \{orXXXXVTM0o}  = masterXXXXVSACKo | (\[15159]  | (\[14852]  | \[15184] )),
  \[15054]  = ~\[10612]_inv  & (~wd_cnt_test & ~physrecXXXXstate0),
  I300 = ~\[10748]_inv  & PCCReqCode1,
  I304 = ~\[10924]_inv  & ~\[15176] ,
  \[10657]_inv  = \[10813]_inv  | ~masterXXXXstate3,
  I305 = ~\[10928]_inv  & ~masterXXXXstate0,
  \[10945]_inv  = SBCResetPCC | ACKi,
  \[15334]  = \[15655]  & ~VTM1l,
  \[15056]  = ~\[10886]_inv  & (VTM0l & ~RESETi),
  \[15710]  = wdcntXXXXstate3 & wdcntXXXXstate0,
  I322 = ~\[15206]  & \[15577] ,
  I323 = \[10363]  & \[15707] ,
  \[15614]  = PCCReqCode0 & PCCReqCode2,
  \[15247]  = ~\[10901]_inv  & (~\[10889]_inv  & ~masterXXXXstate3),
  \[15336]  = ~\[10935]_inv  & ~\[15582] ,
  I340 = ~\[10928]_inv  & ~\[15300] ,
  I341 = \[15379]  & masterXXXXstate3,
  \[15712]  = ~VTM1l & ~TM1l,
  I348 = ~\[15393]  & ~\[15545] ,
  virmachXXXXSBCsetDirty = \[15228] ,
  \{slaveXXXXSBCReqCode0}  = I192 | I193,
  I354 = ~\[15407]  & RESETi,
  \[10845]_inv  = ~P_receive_begin | SBCResetPCC,
  I357 = ~\[15465]  & ~RQSTi,
  \{masterXXXXSBC_WriteCache}  = \[10511]_inv  | \[14902] ,
  I361 = ~\[15670]  & ~\[15377] ,
  I363 = ~\[10651]_inv  & ~\[10943]_inv ,
  I364 = ~\[10882]_inv  & masterXXXXstate2,
  I366 = ~\[15456]  & ~\[15418] ,
  \[10939]_inv  = STARTi | nubusXXXXstate0,
  I368 = ~\[10939]_inv  & \[15692] ,
  I369 = \[2536]  & ACKi,
  \[15529]  = ~CoherencyState2i & CoherencyState1i,
  I373 = ~\[15582]  & \[15538] ,
  I374 = ~\[15266]  & physrecXXXXstate1,
  I377 = ~\[10897]_inv  & ~SlotSpace_Id_Match,
  \[10686]_inv  = ~\[15624]  | I366,
  \{orXXXXVACKo}  = \[15041]  | \[15169] ,
  I398 = ~\[10877]_inv  & ~\[10721]_inv ,
  I399 = ~\[15310]  & slaveXXXXstate2,
  \[15526]  = STARTo & VTM0l,
  \[15159]  = \[15452]  & ~wd_cnt_test,
  \[10886]_inv  = STARTo | (ACKi | ~STARTi),
  orXXXXTM1o = \{orXXXXTM1o} ,
  \[15439]  = ~\[10911]_inv  & wd_cnt_test,
  virmachXXXXSBCConfigure = \{virmachXXXXSBCConfigure} ,
  masterXXXXRQSTo = \[14531] ,
  \[15068]  = ~\[530]  & (~\[10816]_inv  & \[15569] ),
  orXXXXTM0o = \[14862]* ,
  \[15252]  = ~\[10934]_inv  & (~\[10933]_inv  & (Intr_req & slaveXXXXstate0)),
  \{slaveXXXXSBCReqCode1}  = I207 | I208,
  slaveXXXXSnoopState_W = \{slaveXXXXSnoopState_W} ,
  \[15064]  = ~\[10854]_inv  & (Incr_wd_cnt & wdcntXXXXstate3),
  \[15349]  = ~\[15665]  & ~physrecXXXXstate0,
  \[15344]  = ~\[15512]  & ~\[10894]_inv ,
  \[15066]  = ~\[15674]  & \[15247] ,
  \[15442]  = ~\[10890]_inv  & wdcntXXXXstate1,
  \[10911]_inv  = ~physrecXXXXstate1 | ~TM0i,
  \[15624]  = wdcntXXXXstate1 & wdcntXXXXstate2,
  masterXXXXL_DBufo_if_TM0 = \[15247] ,
  \[10703]_inv*  = ~\[10703]_inv ,
  \[15538]  = TM1i & ~TM0i,
  orXXXXEn_START = \{orXXXXEn_START} ,
  \{masterXXXXUpdateReq}  = masterXXXXVSACKo | (\[14505]  | \[14757] ),
  \[10813]_inv  = ~\[15646]  | (masterXXXXstate0 | ~PCCReq),
  I450 = ~\[10940]_inv  & ~nubusXXXXstate1,
  I451 = ~\[10897]_inv  & nubusXXXXstate0,
  I453 = ~\[15591]  & ~masterXXXXstate1,
  orXXXXVACKo = \{orXXXXVACKo} ,
  \[10907]_inv  = ACKi | RESETi,
  I465 = ~V_transmit_begin & ~virmachXXXXstate1,
  \[10511]_inv  = \[15362]  | ~\[10817]_inv ,
  I475 = \[15574]  & VSACKi,
  I476 = masterXXXXstate1 & ~ACKl,
  \[15536]  = VSACKi & slaveXXXXstate0,
  \[10507]_inv  = \[10894]_inv  | (\[14688]  | \[10937]_inv ),
  \[10854]_inv  = \[10890]_inv  | ~wdcntXXXXstate2,
  \[15169]  = \[15452]  & wd_cnt_test,
  orXXXXSBCAckCode0 = \{orXXXXSBCAckCode0} ,
  orXXXXSBCAckCode1 = \{orXXXXSBCAckCode1} ,
  orXXXXSBCAckCode2 = \{orXXXXSBCAckCode2} ,
  orXXXXSBCAckCode3 = \{orXXXXSBCAckCode3} ,
  nubusXXXXL_PABufi = \{nubusXXXXL_PABufi} ,
  \[15444]  = ~\[10930]_inv  & ~masterXXXXstate0,
  masterXXXXSBC_WriteCache = \{masterXXXXSBC_WriteCache} ,
  masterXXXXVSACKo = \[10458]_inv  | ~\[14443] ,
  \[14409]  = ~\[14959]  & (~\[10580]  & (~\[14751]  & ~\[14480] ));
always begin
  wd_cnt_test = \[107] ;
  nubusXXXXstate0 = \[88] ;
  nubusXXXXstate1 = \[89] ;
  Set_ex_wd_cnt1 = \[105] ;
  Incr_wd_cnt = \[106] ;
  Intr_done = \[101] ;
  wdcntXXXXstate0 = \[98] ;
  slaveXXXXstate0 = \[90] ;
  slaveXXXXstate1 = \[91] ;
  slaveXXXXstate2 = \[92] ;
  Reset_wd_cnt = \[104] ;
  P_receive_cancel = \[109] ;
  resetXXXXstate0 = \[93] ;
  resetXXXXstate1 = \[94] ;
  resetXXXXstate2 = \[95] ;
  Intr_req = \[100] ;
  V_transmit_begin = \[111] ;
  UpdateReq = \[102] ;
  virmachXXXXstate0 = \[96] ;
  virmachXXXXstate1 = \[97] ;
  masterXXXXstate0 = \[84] ;
  masterXXXXstate1 = \[85] ;
  masterXXXXstate2 = \[86] ;
  masterXXXXstate3 = \[87] ;
  UpdateDone = \[103] ;
  P_receive_begin = \[108] ;
  Gen_Reset = \[99] ;
end
initial begin
  wd_cnt_test = 0;
  nubusXXXXstate0 = 0;
  nubusXXXXstate1 = 0;
  Set_ex_wd_cnt1 = 0;
  Incr_wd_cnt = 0;
  Intr_done = 0;
  wdcntXXXXstate0 = 0;
  slaveXXXXstate0 = 0;
  slaveXXXXstate1 = 0;
  slaveXXXXstate2 = 0;
  Reset_wd_cnt = 0;
  P_receive_cancel = 0;
  resetXXXXstate0 = 0;
  resetXXXXstate1 = 0;
  resetXXXXstate2 = 0;
  Intr_req = 0;
  V_transmit_begin = 0;
  UpdateReq = 0;
  virmachXXXXstate0 = 0;
  virmachXXXXstate1 = 0;
  masterXXXXstate0 = 0;
  masterXXXXstate1 = 0;
  masterXXXXstate2 = 0;
  masterXXXXstate3 = 0;
  UpdateDone = 0;
  P_receive_begin = 0;
  Gen_Reset = 0;
end
endmodule

